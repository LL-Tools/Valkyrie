

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756;

  INV_X4 U7146 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  OR2_X1 U7147 ( .A1(n10422), .A2(n7763), .ZN(n7762) );
  XNOR2_X1 U7148 ( .A(n9105), .B(SI_22_), .ZN(n9897) );
  CLKBUF_X3 U7149 ( .A(n6411), .Z(n9131) );
  CLKBUF_X2 U7150 ( .A(n10459), .Z(n6399) );
  OR2_X1 U7151 ( .A1(n8915), .A2(n10797), .ZN(n8916) );
  BUF_X2 U7152 ( .A(n6456), .Z(n11095) );
  INV_X2 U7153 ( .A(n8950), .ZN(n6407) );
  INV_X4 U7154 ( .A(n8070), .ZN(n8357) );
  BUF_X1 U7155 ( .A(n13953), .Z(n7158) );
  NAND2_X1 U7156 ( .A1(n8681), .A2(n8680), .ZN(n13951) );
  INV_X1 U7157 ( .A(n8615), .ZN(n14031) );
  OR2_X1 U7158 ( .A1(n11332), .A2(n6553), .ZN(n7135) );
  NAND4_X2 U7159 ( .A1(n6902), .A2(n6474), .A3(n6903), .A4(n6901), .ZN(n14626)
         );
  CLKBUF_X2 U7160 ( .A(n10032), .Z(n6403) );
  INV_X1 U7161 ( .A(n11239), .ZN(n11255) );
  AND2_X1 U7162 ( .A1(n8562), .A2(n8563), .ZN(n7184) );
  NOR2_X1 U7163 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7879) );
  NOR2_X2 U7164 ( .A1(n11408), .A2(n9494), .ZN(n15479) );
  NAND2_X1 U7165 ( .A1(n11896), .A2(n11690), .ZN(n11408) );
  AND2_X1 U7166 ( .A1(n8668), .A2(n8667), .ZN(n8695) );
  AND2_X1 U7167 ( .A1(n7496), .A2(n7495), .ZN(n11248) );
  AND2_X1 U7168 ( .A1(n6743), .A2(n6476), .ZN(n7757) );
  NAND2_X1 U7169 ( .A1(n11555), .A2(n13313), .ZN(n10448) );
  NOR2_X1 U7170 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7881) );
  NOR2_X1 U7171 ( .A1(n12913), .A2(n12912), .ZN(n12915) );
  NOR2_X1 U7172 ( .A1(n11422), .A2(n11427), .ZN(n11491) );
  NAND2_X1 U7173 ( .A1(n8038), .A2(n7913), .ZN(n7146) );
  INV_X2 U7174 ( .A(n9451), .ZN(n9454) );
  NOR3_X2 U7175 ( .A1(n14119), .A2(n7429), .A3(n14298), .ZN(n10440) );
  XNOR2_X1 U7176 ( .A(n6827), .B(n8578), .ZN(n9328) );
  INV_X1 U7177 ( .A(n12855), .ZN(n12877) );
  AND2_X1 U7178 ( .A1(n10921), .A2(n10920), .ZN(n12875) );
  INV_X1 U7179 ( .A(n10660), .ZN(n9848) );
  AND3_X1 U7180 ( .A1(n9550), .A2(n9522), .A3(n9521), .ZN(n9524) );
  INV_X2 U7181 ( .A(n10572), .ZN(n6776) );
  NAND2_X1 U7182 ( .A1(n9511), .A2(n9622), .ZN(n9551) );
  OAI21_X1 U7184 ( .B1(n12964), .B2(n6930), .A(n6928), .ZN(n12954) );
  INV_X2 U7185 ( .A(n8676), .ZN(n8948) );
  INV_X1 U7187 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14440) );
  AND2_X1 U7188 ( .A1(n14479), .A2(n6475), .ZN(n7725) );
  INV_X1 U7189 ( .A(n10029), .ZN(n9985) );
  INV_X1 U7190 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U7191 ( .A1(n8856), .A2(n8855), .ZN(n14382) );
  OR2_X1 U7192 ( .A1(n14755), .A2(n14760), .ZN(n14756) );
  INV_X1 U7193 ( .A(n15514), .ZN(n13128) );
  INV_X1 U7194 ( .A(n13321), .ZN(n13313) );
  NAND2_X1 U7195 ( .A1(n8684), .A2(n8726), .ZN(n10877) );
  INV_X2 U7196 ( .A(n14716), .ZN(n7274) );
  INV_X1 U7197 ( .A(n14940), .ZN(n14920) );
  INV_X1 U7198 ( .A(n14956), .ZN(n14937) );
  BUF_X1 U7199 ( .A(n9542), .Z(n15144) );
  INV_X1 U7200 ( .A(n9543), .ZN(n12896) );
  INV_X1 U7201 ( .A(n10923), .ZN(n10007) );
  INV_X1 U7202 ( .A(n10268), .ZN(n8398) );
  INV_X1 U7203 ( .A(n10459), .ZN(n10509) );
  OR2_X1 U7204 ( .A1(n8979), .A2(n8978), .ZN(n6398) );
  NAND2_X2 U7205 ( .A1(n11694), .A2(n10151), .ZN(n11792) );
  NAND2_X2 U7206 ( .A1(n11692), .A2(n11709), .ZN(n11694) );
  NAND2_X2 U7207 ( .A1(n8480), .A2(n8479), .ZN(n8752) );
  AND2_X2 U7208 ( .A1(n11662), .A2(n8614), .ZN(n9337) );
  NAND2_X1 U7209 ( .A1(n6734), .A2(n6732), .ZN(n7101) );
  NOR2_X1 U7210 ( .A1(n12384), .A2(n12139), .ZN(n10113) );
  NAND2_X2 U7211 ( .A1(n12686), .A2(n12685), .ZN(n14959) );
  NAND2_X2 U7212 ( .A1(n6906), .A2(n6904), .ZN(n12686) );
  XNOR2_X2 U7213 ( .A(n11133), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n15155) );
  NAND2_X2 U7214 ( .A1(n6824), .A2(n11127), .ZN(n11133) );
  AOI22_X2 U7215 ( .A1(n13267), .A2(n13266), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n13274), .ZN(n13294) );
  OAI22_X2 U7216 ( .A1(n13248), .A2(n13247), .B1(n13246), .B2(n13245), .ZN(
        n13267) );
  XNOR2_X2 U7217 ( .A(n14976), .B(n12707), .ZN(n14997) );
  NOR2_X2 U7218 ( .A1(n11248), .A2(n7494), .ZN(n11275) );
  OR2_X2 U7219 ( .A1(n8683), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8726) );
  NAND2_X2 U7220 ( .A1(n7460), .A2(n7459), .ZN(n8273) );
  XNOR2_X2 U7221 ( .A(n8939), .B(n8938), .ZN(n11060) );
  NAND4_X2 U7222 ( .A1(n7331), .A2(n7992), .A3(n7993), .A4(n7994), .ZN(n15536)
         );
  NAND2_X2 U7223 ( .A1(n8981), .A2(n8982), .ZN(n8520) );
  AOI211_X2 U7224 ( .C1(n10228), .C2(n13438), .A(n10227), .B(n10226), .ZN(
        n10230) );
  NAND2_X2 U7225 ( .A1(n11250), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n11315) );
  XNOR2_X2 U7226 ( .A(n7135), .B(n11263), .ZN(n11250) );
  OR2_X2 U7227 ( .A1(n14746), .A2(n14737), .ZN(n6413) );
  OAI211_X2 U7228 ( .C1(n11937), .C2(n6860), .A(n6541), .B(n6859), .ZN(n12035)
         );
  INV_X1 U7229 ( .A(n12755), .ZN(n11168) );
  BUF_X4 U7230 ( .A(n7991), .Z(n8375) );
  AND2_X2 U7231 ( .A1(n7896), .A2(n7897), .ZN(n7991) );
  CLKBUF_X1 U7232 ( .A(n10032), .Z(n6401) );
  BUF_X4 U7233 ( .A(n10032), .Z(n6402) );
  NAND2_X2 U7234 ( .A1(n9541), .A2(n12896), .ZN(n10032) );
  CLKBUF_X3 U7235 ( .A(n11096), .Z(n6404) );
  NAND2_X1 U7237 ( .A1(n8393), .A2(n8394), .ZN(n11096) );
  NAND2_X2 U7238 ( .A1(n9558), .A2(n9563), .ZN(n14716) );
  NAND2_X2 U7239 ( .A1(n9733), .A2(n9732), .ZN(n12295) );
  BUF_X1 U7240 ( .A(n11607), .Z(n6406) );
  XNOR2_X2 U7241 ( .A(n13200), .B(n13183), .ZN(n13202) );
  AOI21_X2 U7242 ( .B1(n13179), .B2(n13178), .A(n6599), .ZN(n13200) );
  AND2_X1 U7243 ( .A1(n12546), .A2(n10362), .ZN(n7118) );
  XNOR2_X2 U7244 ( .A(n13753), .B(n12422), .ZN(n12546) );
  NAND2_X2 U7245 ( .A1(n10115), .A2(n15146), .ZN(n10660) );
  XNOR2_X2 U7246 ( .A(n8715), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10896) );
  NAND2_X2 U7247 ( .A1(n7244), .A2(n7241), .ZN(n15322) );
  NAND2_X1 U7248 ( .A1(n6826), .A2(n15160), .ZN(n15170) );
  NAND2_X1 U7249 ( .A1(n14772), .A2(n12731), .ZN(n14755) );
  AND2_X1 U7250 ( .A1(n12688), .A2(n10089), .ZN(n14931) );
  INV_X1 U7251 ( .A(n10391), .ZN(n11414) );
  INV_X1 U7252 ( .A(n13129), .ZN(n15515) );
  INV_X2 U7253 ( .A(n11619), .ZN(n15472) );
  AND2_X1 U7254 ( .A1(n10104), .A2(n10103), .ZN(n10583) );
  INV_X1 U7255 ( .A(n14626), .ZN(n6900) );
  INV_X1 U7256 ( .A(n14621), .ZN(n6862) );
  XNOR2_X1 U7257 ( .A(n8384), .B(P3_IR_REG_22__SCAN_IN), .ZN(n10338) );
  INV_X1 U7258 ( .A(n11407), .ZN(n11345) );
  AND2_X2 U7259 ( .A1(n6408), .A2(n10567), .ZN(n9214) );
  INV_X2 U7260 ( .A(n8061), .ZN(n8085) );
  OR2_X1 U7261 ( .A1(n10029), .A2(n9578), .ZN(n9579) );
  INV_X2 U7262 ( .A(n9592), .ZN(n9849) );
  XNOR2_X1 U7264 ( .A(n8580), .B(n8576), .ZN(n14449) );
  INV_X2 U7265 ( .A(n11255), .ZN(n7497) );
  NAND4_X1 U7266 ( .A1(n7880), .A2(n7879), .A3(n8179), .A4(n8132), .ZN(n8205)
         );
  INV_X1 U7267 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8604) );
  INV_X1 U7268 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8600) );
  INV_X1 U7269 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8597) );
  NOR2_X1 U7270 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8586) );
  NOR2_X2 U7271 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8662) );
  INV_X1 U7272 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8591) );
  OAI21_X1 U7273 ( .B1(n13289), .B2(n13310), .A(n13311), .ZN(n6682) );
  AND3_X1 U7274 ( .A1(n13288), .A2(n13287), .A3(n13286), .ZN(n13289) );
  NAND2_X1 U7275 ( .A1(n6821), .A2(n7151), .ZN(n15209) );
  AND2_X1 U7276 ( .A1(n7190), .A2(n9333), .ZN(n7556) );
  INV_X1 U7277 ( .A(n13272), .ZN(n6654) );
  NAND2_X1 U7278 ( .A1(n6701), .A2(n13287), .ZN(n13272) );
  AND2_X1 U7279 ( .A1(n9457), .A2(n6676), .ZN(n13712) );
  NAND2_X1 U7280 ( .A1(n7663), .A2(n7664), .ZN(n13023) );
  NAND2_X1 U7281 ( .A1(n14296), .A2(n10385), .ZN(n10387) );
  AND2_X1 U7282 ( .A1(n13018), .A2(n13431), .ZN(n7663) );
  NAND2_X1 U7283 ( .A1(n13837), .A2(n7529), .ZN(n7020) );
  NOR2_X1 U7284 ( .A1(n14564), .A2(n6417), .ZN(n14471) );
  NOR2_X1 U7285 ( .A1(n10283), .A2(n7172), .ZN(n7171) );
  OAI21_X1 U7286 ( .B1(n7717), .B2(n7055), .A(n7054), .ZN(n12854) );
  AND2_X1 U7287 ( .A1(n7717), .A2(n7716), .ZN(n14564) );
  XNOR2_X1 U7288 ( .A(n9438), .B(n7165), .ZN(n13875) );
  NAND2_X1 U7289 ( .A1(n14112), .A2(n10427), .ZN(n7792) );
  NAND2_X1 U7290 ( .A1(n14134), .A2(n10379), .ZN(n14118) );
  NAND2_X1 U7291 ( .A1(n6696), .A2(n6695), .ZN(n15160) );
  NAND2_X1 U7292 ( .A1(n7767), .A2(n6666), .ZN(n14134) );
  NAND2_X1 U7293 ( .A1(n7101), .A2(n10426), .ZN(n14112) );
  NAND2_X1 U7294 ( .A1(n13777), .A2(n13776), .ZN(n13775) );
  NAND2_X1 U7295 ( .A1(n6641), .A2(n6494), .ZN(n7767) );
  NAND2_X1 U7296 ( .A1(n6734), .A2(n6736), .ZN(n14128) );
  OR2_X1 U7297 ( .A1(n14840), .A2(n14839), .ZN(n14788) );
  CLKBUF_X1 U7298 ( .A(n13758), .Z(n7163) );
  AOI21_X1 U7299 ( .B1(n7725), .B2(n7723), .A(n6534), .ZN(n7722) );
  AND2_X1 U7300 ( .A1(n13615), .A2(n13387), .ZN(n10236) );
  NAND2_X1 U7301 ( .A1(n14195), .A2(n10374), .ZN(n14172) );
  NAND2_X1 U7302 ( .A1(n6857), .A2(n7814), .ZN(n14851) );
  AND2_X1 U7303 ( .A1(n10428), .A2(n7791), .ZN(n7789) );
  NAND2_X1 U7304 ( .A1(n8349), .A2(n8348), .ZN(n13615) );
  OAI21_X1 U7305 ( .B1(n13477), .B2(n6546), .A(n7611), .ZN(n7610) );
  NOR2_X1 U7306 ( .A1(n6733), .A2(n14127), .ZN(n6732) );
  NAND2_X1 U7307 ( .A1(n13372), .A2(n10238), .ZN(n13386) );
  AOI21_X1 U7308 ( .B1(n12723), .B2(n7844), .A(n6527), .ZN(n6915) );
  AOI21_X1 U7309 ( .B1(n7612), .B2(n10225), .A(n10222), .ZN(n7611) );
  INV_X1 U7310 ( .A(n6736), .ZN(n6733) );
  NAND2_X1 U7311 ( .A1(n6858), .A2(n12717), .ZN(n14883) );
  CLKBUF_X1 U7312 ( .A(n14215), .Z(n7138) );
  AND2_X2 U7313 ( .A1(n9861), .A2(n12694), .ZN(n14853) );
  NAND2_X2 U7314 ( .A1(n9912), .A2(n9911), .ZN(n15025) );
  XOR2_X1 U7315 ( .A(n12820), .B(n12821), .Z(n14574) );
  NAND2_X1 U7316 ( .A1(n8338), .A2(n8337), .ZN(n12992) );
  NAND2_X1 U7317 ( .A1(n14861), .A2(n14866), .ZN(n12694) );
  NAND2_X1 U7318 ( .A1(n12715), .A2(n12714), .ZN(n14902) );
  NAND2_X1 U7319 ( .A1(n7485), .A2(n7486), .ZN(n8356) );
  NAND2_X1 U7320 ( .A1(n7520), .A2(n6504), .ZN(n13843) );
  NAND2_X1 U7321 ( .A1(n9145), .A2(n9144), .ZN(n14151) );
  NAND2_X1 U7322 ( .A1(n8279), .A2(n8278), .ZN(n13641) );
  NAND2_X1 U7323 ( .A1(n8256), .A2(n8255), .ZN(n13465) );
  NAND2_X1 U7324 ( .A1(n12722), .A2(n12720), .ZN(n14870) );
  NAND2_X1 U7325 ( .A1(n9127), .A2(n9126), .ZN(n14138) );
  XNOR2_X1 U7326 ( .A(n14336), .B(n13933), .ZN(n14159) );
  CLKBUF_X1 U7327 ( .A(n15058), .Z(n7159) );
  XNOR2_X1 U7328 ( .A(n9028), .B(n9027), .ZN(n11585) );
  NAND2_X1 U7329 ( .A1(n9535), .A2(n9534), .ZN(n15058) );
  CLKBUF_X1 U7330 ( .A(n12454), .Z(n6644) );
  AOI21_X1 U7331 ( .B1(n13161), .B2(n13145), .A(n13162), .ZN(n7511) );
  AOI21_X1 U7332 ( .B1(n7623), .B2(n7627), .A(n7621), .ZN(n7620) );
  NAND2_X1 U7333 ( .A1(n9092), .A2(n9091), .ZN(n14312) );
  NAND2_X1 U7334 ( .A1(n12297), .A2(n12296), .ZN(n12299) );
  AND2_X1 U7335 ( .A1(n13459), .A2(n10214), .ZN(n13484) );
  NAND2_X1 U7336 ( .A1(n13144), .A2(n13155), .ZN(n13161) );
  AND2_X1 U7337 ( .A1(n7626), .A2(n7624), .ZN(n7623) );
  NAND2_X1 U7338 ( .A1(n8987), .A2(n8986), .ZN(n14222) );
  NAND2_X1 U7339 ( .A1(n6923), .A2(n6925), .ZN(n13053) );
  XNOR2_X1 U7340 ( .A(n9039), .B(SI_20_), .ZN(n9137) );
  OR2_X1 U7341 ( .A1(n15085), .A2(n14555), .ZN(n12687) );
  NAND2_X1 U7342 ( .A1(n7024), .A2(n6418), .ZN(n9039) );
  XNOR2_X1 U7343 ( .A(n8536), .B(SI_24_), .ZN(n9089) );
  NAND2_X1 U7344 ( .A1(n9820), .A2(n9819), .ZN(n15073) );
  NAND2_X1 U7345 ( .A1(n7021), .A2(n7025), .ZN(n8536) );
  NAND2_X1 U7346 ( .A1(n11884), .A2(n6510), .ZN(n12092) );
  NAND2_X1 U7347 ( .A1(n12107), .A2(n11871), .ZN(n12090) );
  NAND2_X1 U7348 ( .A1(n8879), .A2(n8878), .ZN(n13793) );
  OAI21_X1 U7349 ( .B1(n8937), .B2(n8936), .A(n8935), .ZN(n8939) );
  NAND2_X1 U7350 ( .A1(n8900), .A2(n8899), .ZN(n12589) );
  NAND2_X1 U7351 ( .A1(n9749), .A2(n9748), .ZN(n12532) );
  AOI21_X1 U7352 ( .B1(n7643), .B2(n7646), .A(n7642), .ZN(n7641) );
  NAND2_X2 U7353 ( .A1(n8835), .A2(n8834), .ZN(n13753) );
  NAND2_X1 U7354 ( .A1(n8935), .A2(n8916), .ZN(n8937) );
  NAND2_X1 U7355 ( .A1(n11913), .A2(n6492), .ZN(n12070) );
  NAND2_X2 U7356 ( .A1(n8813), .A2(n8812), .ZN(n13851) );
  XNOR2_X1 U7357 ( .A(n8831), .B(n8830), .ZN(n10686) );
  NAND2_X2 U7358 ( .A1(n11716), .A2(n15509), .ZN(n15524) );
  XNOR2_X1 U7359 ( .A(n8173), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U7360 ( .A1(n8798), .A2(n8797), .ZN(n12159) );
  NAND2_X1 U7361 ( .A1(n11301), .A2(n11300), .ZN(n11302) );
  NAND2_X1 U7362 ( .A1(n7468), .A2(n7929), .ZN(n8173) );
  AOI21_X1 U7363 ( .B1(n15153), .B2(n15154), .A(n10645), .ZN(n10647) );
  INV_X1 U7364 ( .A(n11957), .ZN(n6860) );
  AND2_X1 U7365 ( .A1(n10126), .A2(n10139), .ZN(n11722) );
  INV_X1 U7366 ( .A(n15478), .ZN(n11656) );
  NAND4_X1 U7367 ( .A1(n8764), .A2(n8763), .A3(n8762), .A4(n8761), .ZN(n13948)
         );
  INV_X4 U7368 ( .A(n12857), .ZN(n11176) );
  NAND2_X1 U7369 ( .A1(n8638), .A2(n6517), .ZN(n13954) );
  BUF_X2 U7370 ( .A(n9344), .Z(n9451) );
  NAND4_X1 U7371 ( .A1(n8739), .A2(n8738), .A3(n8737), .A4(n8736), .ZN(n13949)
         );
  NAND2_X1 U7372 ( .A1(n8717), .A2(n8716), .ZN(n15478) );
  NAND4_X2 U7373 ( .A1(n8712), .A2(n8711), .A3(n8710), .A4(n8709), .ZN(n13950)
         );
  XNOR2_X1 U7374 ( .A(n13951), .B(n10391), .ZN(n7117) );
  CLKBUF_X1 U7375 ( .A(n10391), .Z(n11667) );
  NAND2_X1 U7376 ( .A1(n11207), .A2(n10920), .ZN(n12755) );
  XNOR2_X1 U7377 ( .A(n13126), .B(n10465), .ZN(n12167) );
  INV_X2 U7378 ( .A(n12875), .ZN(n12866) );
  NAND4_X2 U7379 ( .A1(n8657), .A2(n8656), .A3(n8655), .A4(n8654), .ZN(n13952)
         );
  AND4_X1 U7380 ( .A1(n8005), .A2(n8004), .A3(n8003), .A4(n8002), .ZN(n15514)
         );
  NAND4_X1 U7381 ( .A1(n7105), .A2(n8651), .A3(n8650), .A4(n8649), .ZN(n13953)
         );
  INV_X2 U7382 ( .A(n12747), .ZN(n14277) );
  CLKBUF_X1 U7383 ( .A(n8673), .Z(n8924) );
  OR2_X1 U7384 ( .A1(n8675), .A2(n8648), .ZN(n8649) );
  AND2_X1 U7386 ( .A1(n7684), .A2(n8499), .ZN(n7683) );
  OR2_X1 U7387 ( .A1(n11704), .A2(n11555), .ZN(n10451) );
  OR2_X1 U7388 ( .A1(n11225), .A2(n14623), .ZN(n9602) );
  NAND3_X1 U7389 ( .A1(n9585), .A2(n9586), .A3(n6872), .ZN(n14622) );
  NAND4_X1 U7390 ( .A1(n7215), .A2(n7214), .A3(n7216), .A4(n7977), .ZN(n13129)
         );
  CLKBUF_X1 U7391 ( .A(n8944), .Z(n9149) );
  CLKBUF_X3 U7392 ( .A(n8687), .Z(n9125) );
  NAND2_X1 U7393 ( .A1(n8391), .A2(n8390), .ZN(n11555) );
  INV_X1 U7394 ( .A(n9214), .ZN(n8666) );
  NAND2_X1 U7396 ( .A1(n8624), .A2(n12937), .ZN(n8673) );
  MUX2_X1 U7397 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10102), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n10104) );
  AOI21_X1 U7398 ( .B1(n8484), .B2(n6972), .A(n6530), .ZN(n6971) );
  MUX2_X1 U7399 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8388), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8391) );
  NAND2_X2 U7400 ( .A1(n8623), .A2(n8624), .ZN(n9234) );
  INV_X1 U7401 ( .A(n10920), .ZN(n10749) );
  INV_X1 U7402 ( .A(n10935), .ZN(n11909) );
  OR2_X1 U7403 ( .A1(n6401), .A2(n9571), .ZN(n6902) );
  NAND2_X1 U7404 ( .A1(n10107), .A2(n10108), .ZN(n12384) );
  INV_X1 U7405 ( .A(n8614), .ZN(n11690) );
  INV_X1 U7406 ( .A(n8623), .ZN(n12937) );
  CLKBUF_X2 U7407 ( .A(n10255), .Z(n10265) );
  MUX2_X1 U7408 ( .A(n8634), .B(n14452), .S(n8690), .Z(n11407) );
  NAND2_X2 U7409 ( .A1(n8606), .A2(n9324), .ZN(n11896) );
  MUX2_X1 U7410 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8602), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n8606) );
  NAND2_X1 U7411 ( .A1(n8605), .A2(n8604), .ZN(n9324) );
  XNOR2_X1 U7412 ( .A(n9555), .B(n9554), .ZN(n10006) );
  NAND2_X1 U7413 ( .A1(n6683), .A2(n8592), .ZN(n8594) );
  XNOR2_X1 U7414 ( .A(n7080), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U7415 ( .A1(n10007), .A2(n10011), .ZN(n10920) );
  XNOR2_X1 U7416 ( .A(n10112), .B(n10111), .ZN(n12139) );
  AND2_X1 U7417 ( .A1(n8386), .A2(n8382), .ZN(n8389) );
  NAND2_X1 U7418 ( .A1(n6636), .A2(n6633), .ZN(n13697) );
  OR2_X1 U7419 ( .A1(n6741), .A2(n10684), .ZN(n6740) );
  OAI21_X1 U7420 ( .B1(n9005), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U7421 ( .A1(n9590), .A2(n9619), .ZN(n14639) );
  AOI21_X1 U7422 ( .B1(n8590), .B2(P2_IR_REG_31__SCAN_IN), .A(n7535), .ZN(
        n6684) );
  XNOR2_X1 U7423 ( .A(n7213), .B(n7212), .ZN(n8394) );
  OR2_X1 U7424 ( .A1(n8601), .A2(n14440), .ZN(n8589) );
  XNOR2_X1 U7425 ( .A(n9564), .B(P1_IR_REG_20__SCAN_IN), .ZN(n10923) );
  XNOR2_X1 U7426 ( .A(n9561), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10011) );
  NAND2_X2 U7427 ( .A1(n10572), .A2(P3_U3151), .ZN(n13707) );
  AOI21_X1 U7428 ( .B1(n7476), .B2(n7474), .A(n7473), .ZN(n7472) );
  NAND2_X1 U7429 ( .A1(n15138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9539) );
  NAND2_X1 U7430 ( .A1(n10103), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9520) );
  NAND2_X1 U7431 ( .A1(n6755), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6754) );
  CLKBUF_X2 U7432 ( .A(n8579), .Z(n9321) );
  NAND2_X1 U7433 ( .A1(n8209), .A2(n7711), .ZN(n8381) );
  NOR2_X1 U7434 ( .A1(n10099), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U7435 ( .A1(n7965), .A2(n7894), .ZN(n13687) );
  NAND2_X2 U7436 ( .A1(n10567), .A2(P2_U3088), .ZN(n14447) );
  OAI21_X1 U7437 ( .B1(n10567), .B2(n10670), .A(n7715), .ZN(n8475) );
  NOR2_X2 U7438 ( .A1(n8429), .A2(n8205), .ZN(n8209) );
  AND2_X1 U7439 ( .A1(n7184), .A2(n8566), .ZN(n8574) );
  NAND2_X1 U7440 ( .A1(n6661), .A2(n7889), .ZN(n8429) );
  AND3_X1 U7441 ( .A1(n9550), .A2(n9549), .A3(n9521), .ZN(n7541) );
  AND2_X1 U7442 ( .A1(n9523), .A2(n9526), .ZN(n6756) );
  AND2_X1 U7443 ( .A1(n8659), .A2(n7242), .ZN(n7241) );
  AND3_X1 U7444 ( .A1(n9514), .A2(n9513), .A3(n9512), .ZN(n9550) );
  NAND2_X1 U7445 ( .A1(n10674), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7916) );
  AND2_X1 U7446 ( .A1(n9549), .A2(n9519), .ZN(n9523) );
  CLKBUF_X1 U7447 ( .A(n8597), .Z(n8598) );
  NAND3_X1 U7448 ( .A1(n8570), .A2(n8569), .A3(n8568), .ZN(n8595) );
  NAND3_X1 U7449 ( .A1(n8875), .A2(n8565), .A3(n8564), .ZN(n8584) );
  AND3_X1 U7450 ( .A1(n8662), .A2(n8586), .A3(n8585), .ZN(n9311) );
  NOR2_X2 U7451 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n11104) );
  INV_X4 U7452 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7453 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9675) );
  INV_X1 U7454 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10674) );
  INV_X1 U7455 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10654) );
  NOR2_X1 U7456 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n9508) );
  INV_X4 U7457 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7458 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9514) );
  NOR2_X1 U7459 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n9513) );
  NOR2_X1 U7460 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n9512) );
  NOR2_X1 U7461 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9549) );
  NOR2_X1 U7462 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9509) );
  NOR2_X1 U7463 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9510) );
  INV_X1 U7464 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8570) );
  INV_X1 U7465 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8569) );
  INV_X1 U7466 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8568) );
  INV_X1 U7467 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8132) );
  INV_X1 U7468 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8875) );
  INV_X1 U7469 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8565) );
  INV_X1 U7470 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8564) );
  BUF_X1 U7471 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n15321) );
  INV_X1 U7472 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8631) );
  INV_X1 U7473 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U7474 ( .A1(n9328), .A2(n14449), .ZN(n6408) );
  NAND2_X1 U7475 ( .A1(n9328), .A2(n14449), .ZN(n8690) );
  NAND2_X2 U7476 ( .A1(n12185), .A2(n12184), .ZN(n12188) );
  NAND2_X2 U7477 ( .A1(n7309), .A2(n7308), .ZN(n9105) );
  NAND2_X1 U7479 ( .A1(n10660), .A2(n10572), .ZN(n10015) );
  INV_X2 U7480 ( .A(n9542), .ZN(n9541) );
  XNOR2_X2 U7481 ( .A(n8589), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8614) );
  AOI21_X2 U7482 ( .B1(n11315), .B2(n6457), .A(n11314), .ZN(n11420) );
  NOR2_X1 U7483 ( .A1(n11108), .A2(n11109), .ZN(n11247) );
  INV_X2 U7484 ( .A(n6421), .ZN(n8965) );
  NAND2_X1 U7485 ( .A1(n12937), .A2(n12741), .ZN(n8675) );
  INV_X1 U7486 ( .A(n9269), .ZN(n6409) );
  INV_X1 U7487 ( .A(n6409), .ZN(n6410) );
  INV_X1 U7488 ( .A(n6409), .ZN(n6411) );
  INV_X2 U7489 ( .A(n6409), .ZN(n6412) );
  NAND2_X1 U7490 ( .A1(n9722), .A2(n9719), .ZN(n7587) );
  INV_X1 U7491 ( .A(n7789), .ZN(n7788) );
  INV_X1 U7492 ( .A(n9179), .ZN(n8542) );
  AND2_X1 U7493 ( .A1(n7890), .A2(n6580), .ZN(n7658) );
  INV_X1 U7494 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U7495 ( .A1(n7074), .A2(n6437), .ZN(n10369) );
  INV_X1 U7496 ( .A(n8595), .ZN(n8596) );
  NAND2_X1 U7497 ( .A1(n12092), .A2(n7842), .ZN(n12185) );
  NOR2_X1 U7498 ( .A1(n11888), .A2(n7843), .ZN(n7842) );
  INV_X1 U7499 ( .A(n11887), .ZN(n7843) );
  NAND2_X1 U7500 ( .A1(n6725), .A2(n10236), .ZN(n7036) );
  AND2_X2 U7501 ( .A1(n8623), .A2(n12741), .ZN(n8676) );
  AND2_X1 U7502 ( .A1(n7770), .A2(n14127), .ZN(n6666) );
  NAND2_X1 U7503 ( .A1(n12434), .A2(n7076), .ZN(n7074) );
  OR2_X1 U7504 ( .A1(n10545), .A2(n9498), .ZN(n10978) );
  AND2_X1 U7505 ( .A1(n6585), .A2(n7299), .ZN(n7270) );
  NOR2_X1 U7506 ( .A1(n10145), .A2(n10146), .ZN(n7336) );
  AND2_X1 U7507 ( .A1(n7586), .A2(n9736), .ZN(n7585) );
  NAND2_X1 U7508 ( .A1(n7588), .A2(n7587), .ZN(n7586) );
  AND2_X1 U7509 ( .A1(n13535), .A2(n6566), .ZN(n7346) );
  AOI21_X1 U7510 ( .B1(n6431), .B2(n7199), .A(n6551), .ZN(n7194) );
  AOI21_X1 U7511 ( .B1(n7209), .B2(n7208), .A(n7207), .ZN(n7206) );
  INV_X1 U7512 ( .A(n8933), .ZN(n7207) );
  NAND2_X1 U7513 ( .A1(n6952), .A2(n6945), .ZN(n6944) );
  NAND2_X1 U7514 ( .A1(n13482), .A2(n6946), .ZN(n6945) );
  NAND2_X1 U7515 ( .A1(n10213), .A2(n10204), .ZN(n6952) );
  NOR2_X1 U7516 ( .A1(n13585), .A2(n10197), .ZN(n6946) );
  INV_X1 U7517 ( .A(n10198), .ZN(n6949) );
  NAND2_X1 U7518 ( .A1(n7155), .A2(n7152), .ZN(n10193) );
  NOR2_X1 U7519 ( .A1(n13428), .A2(n7350), .ZN(n7349) );
  NAND2_X1 U7520 ( .A1(n13446), .A2(n6495), .ZN(n7350) );
  AOI21_X1 U7521 ( .B1(n6773), .B2(n6771), .A(n6769), .ZN(n6768) );
  NOR2_X1 U7522 ( .A1(n9124), .A2(SI_22_), .ZN(n7697) );
  INV_X1 U7523 ( .A(n8533), .ZN(n7698) );
  AOI21_X1 U7524 ( .B1(n14258), .B2(n10416), .A(n6496), .ZN(n7801) );
  OR2_X1 U7525 ( .A1(n13552), .A2(n12902), .ZN(n10244) );
  NAND2_X1 U7526 ( .A1(n11705), .A2(n8080), .ZN(n6721) );
  NAND2_X1 U7527 ( .A1(n8080), .A2(n8081), .ZN(n6720) );
  INV_X1 U7528 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7660) );
  AOI21_X1 U7529 ( .B1(n7564), .B2(n7561), .A(n7558), .ZN(n7557) );
  OR2_X1 U7530 ( .A1(n7565), .A2(n9053), .ZN(n7564) );
  AND2_X1 U7531 ( .A1(n7559), .A2(n7565), .ZN(n7558) );
  NOR2_X1 U7532 ( .A1(n7568), .A2(n7567), .ZN(n7565) );
  INV_X1 U7533 ( .A(n6912), .ZN(n6911) );
  OAI21_X1 U7534 ( .B1(n14958), .B2(n6913), .A(n14931), .ZN(n6912) );
  INV_X1 U7535 ( .A(n12687), .ZN(n6913) );
  AND2_X1 U7536 ( .A1(n8525), .A2(n9025), .ZN(n8526) );
  NAND2_X1 U7537 ( .A1(n8522), .A2(n7312), .ZN(n7311) );
  INV_X1 U7538 ( .A(n8522), .ZN(n7313) );
  NAND2_X1 U7539 ( .A1(n6415), .A2(n10495), .ZN(n6930) );
  AND2_X1 U7540 ( .A1(n10449), .A2(n10448), .ZN(n10450) );
  INV_X1 U7541 ( .A(n13697), .ZN(n7896) );
  NAND2_X1 U7542 ( .A1(n7395), .A2(n7394), .ZN(n7393) );
  AND2_X1 U7543 ( .A1(n7407), .A2(n7406), .ZN(n7405) );
  INV_X1 U7544 ( .A(n13136), .ZN(n7406) );
  OR2_X1 U7545 ( .A1(n12068), .A2(n12069), .ZN(n7407) );
  AOI21_X1 U7546 ( .B1(n7424), .B2(n8305), .A(n6515), .ZN(n7422) );
  INV_X1 U7547 ( .A(n12354), .ZN(n10452) );
  INV_X1 U7548 ( .A(n15511), .ZN(n10306) );
  NAND2_X1 U7549 ( .A1(n13128), .A2(n12354), .ZN(n10139) );
  NAND2_X1 U7550 ( .A1(n13129), .A2(n15526), .ZN(n10131) );
  OR2_X1 U7551 ( .A1(n13565), .A2(n13419), .ZN(n10231) );
  OR2_X1 U7552 ( .A1(n13635), .A2(n13418), .ZN(n10210) );
  AND2_X1 U7553 ( .A1(n13635), .A2(n13418), .ZN(n10208) );
  NOR2_X1 U7554 ( .A1(n7418), .A2(n8144), .ZN(n7417) );
  INV_X1 U7555 ( .A(n8128), .ZN(n7418) );
  OR2_X1 U7556 ( .A1(n11697), .A2(n10610), .ZN(n10347) );
  NOR2_X1 U7557 ( .A1(n8433), .A2(n12199), .ZN(n10530) );
  INV_X1 U7558 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7887) );
  NOR2_X1 U7559 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7888) );
  NAND2_X1 U7560 ( .A1(n6714), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7213) );
  INV_X1 U7561 ( .A(n7929), .ZN(n7471) );
  AND2_X1 U7562 ( .A1(n7918), .A2(n7477), .ZN(n7476) );
  AND2_X2 U7563 ( .A1(n11104), .A2(n7885), .ZN(n8008) );
  INV_X1 U7564 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7885) );
  NOR2_X1 U7565 ( .A1(n14387), .A2(n13928), .ZN(n9267) );
  NOR2_X1 U7566 ( .A1(n6532), .A2(n7100), .ZN(n7099) );
  INV_X1 U7567 ( .A(n10430), .ZN(n7100) );
  INV_X1 U7568 ( .A(n10426), .ZN(n7104) );
  INV_X1 U7569 ( .A(n14078), .ZN(n6753) );
  NOR2_X1 U7570 ( .A1(n14179), .A2(n14209), .ZN(n7438) );
  NAND2_X1 U7571 ( .A1(n8988), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9009) );
  INV_X1 U7572 ( .A(n10366), .ZN(n7077) );
  AND2_X1 U7573 ( .A1(n12430), .A2(n10405), .ZN(n10406) );
  AND2_X1 U7574 ( .A1(n12151), .A2(n10361), .ZN(n7181) );
  NAND2_X1 U7575 ( .A1(n11851), .A2(n10360), .ZN(n11770) );
  NAND2_X1 U7576 ( .A1(n9274), .A2(n14277), .ZN(n10389) );
  OR2_X1 U7577 ( .A1(n15058), .A2(n14889), .ZN(n12722) );
  NAND2_X1 U7578 ( .A1(n7116), .A2(n6606), .ZN(n8544) );
  AOI21_X1 U7579 ( .B1(n9075), .B2(n7015), .A(n7014), .ZN(n7013) );
  NOR2_X1 U7580 ( .A1(n9056), .A2(n12560), .ZN(n7014) );
  OAI21_X1 U7581 ( .B1(n9089), .B2(n7253), .A(n8537), .ZN(n9076) );
  INV_X1 U7582 ( .A(n9090), .ZN(n7253) );
  AND2_X1 U7583 ( .A1(n6740), .A2(n8496), .ZN(n8869) );
  NAND2_X1 U7584 ( .A1(n7314), .A2(n9569), .ZN(n8642) );
  INV_X1 U7585 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7661) );
  NAND2_X1 U7586 ( .A1(n10629), .A2(n10628), .ZN(n10627) );
  AOI21_X1 U7587 ( .B1(n7671), .B2(n7672), .A(n7670), .ZN(n7669) );
  NOR2_X1 U7588 ( .A1(n10486), .A2(n13525), .ZN(n7670) );
  AND2_X1 U7589 ( .A1(n7674), .A2(n6484), .ZN(n7671) );
  XNOR2_X1 U7590 ( .A(n11242), .B(n11281), .ZN(n11274) );
  NAND2_X1 U7591 ( .A1(n7393), .A2(n11425), .ZN(n7392) );
  INV_X1 U7592 ( .A(n7391), .ZN(n7390) );
  OAI21_X1 U7593 ( .B1(n7392), .B2(n6467), .A(n11430), .ZN(n7391) );
  NAND2_X1 U7594 ( .A1(n13271), .A2(n13299), .ZN(n13287) );
  NAND2_X1 U7595 ( .A1(n6654), .A2(n6625), .ZN(n7503) );
  NAND2_X1 U7596 ( .A1(n6654), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13288) );
  OAI21_X1 U7597 ( .B1(n13361), .B2(n7232), .A(n7231), .ZN(n7235) );
  AOI21_X1 U7598 ( .B1(n7233), .B2(n6725), .A(n7236), .ZN(n7231) );
  AND2_X1 U7599 ( .A1(n12633), .A2(n13548), .ZN(n7236) );
  AND2_X1 U7600 ( .A1(n8420), .A2(n10334), .ZN(n15521) );
  INV_X1 U7601 ( .A(n11095), .ZN(n10532) );
  OR2_X1 U7602 ( .A1(n13630), .A2(n13431), .ZN(n13398) );
  OR2_X1 U7603 ( .A1(n13429), .A2(n8305), .ZN(n7426) );
  NOR2_X1 U7604 ( .A1(n13416), .A2(n7425), .ZN(n7424) );
  INV_X1 U7605 ( .A(n8304), .ZN(n7425) );
  NAND2_X1 U7606 ( .A1(n13536), .A2(n10186), .ZN(n8190) );
  INV_X1 U7607 ( .A(n13535), .ZN(n10186) );
  OR2_X1 U7608 ( .A1(n10532), .A2(n10522), .ZN(n15513) );
  INV_X1 U7609 ( .A(n15535), .ZN(n15516) );
  AND2_X1 U7610 ( .A1(n11095), .A2(n10522), .ZN(n15535) );
  OR2_X1 U7611 ( .A1(n13683), .A2(n10530), .ZN(n11098) );
  NAND2_X1 U7612 ( .A1(n6969), .A2(n8440), .ZN(n8441) );
  NAND2_X1 U7613 ( .A1(n8435), .A2(n12452), .ZN(n6969) );
  XNOR2_X1 U7614 ( .A(n7895), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U7615 ( .A1(n13687), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7895) );
  NAND2_X1 U7616 ( .A1(n7967), .A2(n7968), .ZN(n8393) );
  MUX2_X1 U7617 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7966), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7968) );
  OR2_X1 U7618 ( .A1(n7965), .A2(n13686), .ZN(n7966) );
  OAI21_X1 U7619 ( .B1(n7949), .B2(n7449), .A(n7447), .ZN(n8309) );
  AND2_X1 U7620 ( .A1(n7448), .A2(n8306), .ZN(n7447) );
  OR2_X1 U7621 ( .A1(n6592), .A2(n7449), .ZN(n7448) );
  INV_X1 U7622 ( .A(n7951), .ZN(n7449) );
  NAND2_X1 U7623 ( .A1(n7949), .A2(n6592), .ZN(n8293) );
  NAND2_X1 U7624 ( .A1(n8381), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U7625 ( .A1(n7943), .A2(n7942), .ZN(n8232) );
  OAI21_X1 U7626 ( .B1(n9416), .B2(n6675), .A(n7007), .ZN(n13758) );
  INV_X1 U7627 ( .A(n6674), .ZN(n7007) );
  OAI21_X1 U7628 ( .B1(n6675), .B2(n9415), .A(n6543), .ZN(n6674) );
  OR2_X1 U7629 ( .A1(n9114), .A2(n13838), .ZN(n9094) );
  NAND2_X1 U7630 ( .A1(n13775), .A2(n9436), .ZN(n9438) );
  NAND2_X1 U7631 ( .A1(n7020), .A2(n7018), .ZN(n9457) );
  NOR2_X1 U7632 ( .A1(n7019), .A2(n13908), .ZN(n7018) );
  INV_X1 U7633 ( .A(n7531), .ZN(n7019) );
  NAND2_X1 U7634 ( .A1(n10435), .A2(n14048), .ZN(n7106) );
  AND4_X1 U7635 ( .A1(n8888), .A2(n8887), .A3(n8886), .A4(n8885), .ZN(n12583)
         );
  NAND2_X1 U7636 ( .A1(n7078), .A2(n10384), .ZN(n14072) );
  OAI21_X1 U7637 ( .B1(n14118), .B2(n7794), .A(n7795), .ZN(n7078) );
  NAND2_X1 U7638 ( .A1(n10382), .A2(n7800), .ZN(n7794) );
  INV_X1 U7639 ( .A(n7771), .ZN(n7770) );
  OR2_X1 U7640 ( .A1(n14151), .A2(n13932), .ZN(n7772) );
  NAND2_X1 U7641 ( .A1(n7775), .A2(n10378), .ZN(n7773) );
  AOI21_X1 U7642 ( .B1(n7759), .B2(n6476), .A(n7755), .ZN(n7754) );
  INV_X1 U7643 ( .A(n14159), .ZN(n7755) );
  AND2_X2 U7644 ( .A1(n7762), .A2(n7766), .ZN(n7761) );
  NAND2_X1 U7645 ( .A1(n10420), .A2(n10419), .ZN(n7763) );
  NAND2_X1 U7646 ( .A1(n7085), .A2(n10411), .ZN(n12635) );
  INV_X1 U7647 ( .A(n10412), .ZN(n7081) );
  OAI22_X2 U7648 ( .A1(n12429), .A2(n10365), .B1(n14382), .B2(n13942), .ZN(
        n12434) );
  AND2_X1 U7649 ( .A1(n9472), .A2(n9471), .ZN(n15458) );
  XNOR2_X1 U7650 ( .A(n9297), .B(n9296), .ZN(n10855) );
  NAND2_X1 U7651 ( .A1(n14439), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7080) );
  AND2_X1 U7652 ( .A1(n8577), .A2(n7782), .ZN(n8609) );
  XNOR2_X1 U7653 ( .A(n8599), .B(n8598), .ZN(n8615) );
  OAI211_X1 U7654 ( .C1(n11182), .C2(n11175), .A(n7049), .B(n11189), .ZN(
        n11193) );
  OR2_X1 U7655 ( .A1(n14639), .A2(n10704), .ZN(n6811) );
  NOR3_X1 U7656 ( .A1(n6413), .A2(n14986), .A3(n6791), .ZN(n6790) );
  NAND2_X1 U7657 ( .A1(n14974), .A2(n6792), .ZN(n6791) );
  OAI21_X1 U7658 ( .B1(n7822), .B2(n7320), .A(n7820), .ZN(n7319) );
  NAND2_X1 U7659 ( .A1(n14760), .A2(n12732), .ZN(n7320) );
  AOI21_X1 U7660 ( .B1(n7823), .B2(n7821), .A(n6535), .ZN(n7820) );
  NOR2_X1 U7661 ( .A1(n7822), .A2(n7322), .ZN(n7321) );
  INV_X1 U7662 ( .A(n12732), .ZN(n7322) );
  AND2_X1 U7663 ( .A1(n7318), .A2(n7317), .ZN(n14710) );
  NOR2_X1 U7664 ( .A1(n7319), .A2(n12735), .ZN(n7317) );
  AND2_X1 U7665 ( .A1(n9982), .A2(n9954), .ZN(n14747) );
  AND2_X1 U7666 ( .A1(n9953), .A2(n9935), .ZN(n14764) );
  NOR2_X1 U7667 ( .A1(n6468), .A2(n6877), .ZN(n6876) );
  INV_X1 U7668 ( .A(n12724), .ZN(n6877) );
  AOI21_X1 U7669 ( .B1(n7840), .B2(n7839), .A(n7838), .ZN(n7837) );
  INV_X1 U7670 ( .A(n12696), .ZN(n7838) );
  INV_X1 U7671 ( .A(n14824), .ZN(n7839) );
  NAND2_X2 U7672 ( .A1(n9851), .A2(n9850), .ZN(n14861) );
  NAND2_X1 U7673 ( .A1(n11585), .A2(n9591), .ZN(n9851) );
  NAND2_X1 U7674 ( .A1(n9538), .A2(n6845), .ZN(n9853) );
  AND2_X1 U7675 ( .A1(n7806), .A2(n12501), .ZN(n7805) );
  NAND2_X1 U7676 ( .A1(n7807), .A2(n12457), .ZN(n7806) );
  INV_X1 U7677 ( .A(n12453), .ZN(n7807) );
  XNOR2_X1 U7678 ( .A(n15097), .B(n12770), .ZN(n12457) );
  INV_X1 U7679 ( .A(n12095), .ZN(n11885) );
  OAI211_X1 U7680 ( .C1(n8553), .C2(n6993), .A(n6992), .B(n6988), .ZN(n14438)
         );
  INV_X1 U7681 ( .A(n6989), .ZN(n6988) );
  NAND2_X1 U7682 ( .A1(n8553), .A2(n6595), .ZN(n6992) );
  OAI21_X1 U7683 ( .B1(n6591), .B2(n6993), .A(n6990), .ZN(n6989) );
  NAND2_X1 U7684 ( .A1(n15249), .A2(n9575), .ZN(n9597) );
  NAND2_X1 U7685 ( .A1(n15159), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6826) );
  NAND2_X1 U7686 ( .A1(n15169), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7381) );
  NAND2_X1 U7687 ( .A1(n7383), .A2(n15442), .ZN(n7382) );
  OR2_X2 U7688 ( .A1(n13683), .A2(n10547), .ZN(n13130) );
  NOR2_X1 U7689 ( .A1(n6528), .A2(n6895), .ZN(n6894) );
  NOR2_X1 U7690 ( .A1(n6458), .A2(n11303), .ZN(n6895) );
  OAI22_X1 U7691 ( .A1(n13296), .A2(n15734), .B1(n13295), .B2(n13294), .ZN(
        n13319) );
  AOI21_X1 U7692 ( .B1(n7657), .B2(n7656), .A(n10236), .ZN(n13359) );
  AND2_X1 U7693 ( .A1(n9991), .A2(n9990), .ZN(n14732) );
  OR2_X1 U7694 ( .A1(n12703), .A2(n10026), .ZN(n9991) );
  INV_X1 U7695 ( .A(n14606), .ZN(n14798) );
  INV_X1 U7696 ( .A(n14604), .ZN(n14765) );
  AOI22_X1 U7697 ( .A1(n11072), .A2(n11071), .B1(n11070), .B2(n11069), .ZN(
        n11074) );
  AOI21_X1 U7698 ( .B1(n7291), .B2(P1_REG1_REG_18__SCAN_IN), .A(n14679), .ZN(
        n14680) );
  OAI21_X1 U7699 ( .B1(n14681), .B2(n14876), .A(n14684), .ZN(n14685) );
  NAND2_X1 U7700 ( .A1(n7825), .A2(n7823), .ZN(n14731) );
  NAND2_X1 U7701 ( .A1(n10650), .A2(n11127), .ZN(n10651) );
  INV_X1 U7702 ( .A(n12614), .ZN(n6695) );
  INV_X1 U7703 ( .A(n12615), .ZN(n6696) );
  OR2_X1 U7704 ( .A1(n15204), .A2(n15203), .ZN(n6821) );
  INV_X1 U7705 ( .A(n8637), .ZN(n8635) );
  OAI21_X1 U7706 ( .B1(n9610), .B2(n11596), .A(n11225), .ZN(n9608) );
  OAI21_X1 U7707 ( .B1(n8965), .B2(n12747), .A(n8652), .ZN(n8671) );
  NAND2_X1 U7708 ( .A1(n9649), .A2(n6767), .ZN(n6766) );
  NAND2_X1 U7709 ( .A1(n10142), .A2(n11095), .ZN(n7338) );
  AOI21_X1 U7710 ( .B1(n6432), .B2(n6781), .A(n6780), .ZN(n6779) );
  NAND2_X1 U7711 ( .A1(n7198), .A2(n7197), .ZN(n7196) );
  OAI21_X1 U7712 ( .B1(n8850), .B2(n8849), .A(n6498), .ZN(n6663) );
  NOR2_X1 U7713 ( .A1(n7583), .A2(n6464), .ZN(n7581) );
  OAI21_X1 U7714 ( .B1(n9720), .B2(n7588), .A(n7125), .ZN(n9738) );
  AND2_X1 U7715 ( .A1(n9784), .A2(n6540), .ZN(n6763) );
  AND2_X1 U7716 ( .A1(n14958), .A2(n9783), .ZN(n9784) );
  INV_X1 U7717 ( .A(n9750), .ZN(n7582) );
  NAND2_X1 U7718 ( .A1(n7346), .A2(n6514), .ZN(n7343) );
  INV_X1 U7719 ( .A(n7577), .ZN(n7203) );
  NAND2_X1 U7720 ( .A1(n7205), .A2(n6422), .ZN(n7204) );
  INV_X1 U7721 ( .A(n7206), .ZN(n7205) );
  NAND2_X1 U7722 ( .A1(n6460), .A2(n7577), .ZN(n7211) );
  OAI21_X1 U7723 ( .B1(n10199), .B2(n6943), .A(n6941), .ZN(n6950) );
  NAND2_X1 U7724 ( .A1(n6947), .A2(n10214), .ZN(n6943) );
  AND2_X1 U7725 ( .A1(n6951), .A2(n6942), .ZN(n6941) );
  AOI22_X1 U7726 ( .A1(n7600), .A2(n7595), .B1(n7592), .B2(n9887), .ZN(n7591)
         );
  NAND2_X1 U7727 ( .A1(n7608), .A2(n9932), .ZN(n7607) );
  INV_X1 U7728 ( .A(n9931), .ZN(n7608) );
  AOI21_X1 U7729 ( .B1(n7696), .B2(n7694), .A(n7693), .ZN(n7692) );
  INV_X1 U7730 ( .A(n8535), .ZN(n7693) );
  NAND2_X1 U7731 ( .A1(n7028), .A2(n6418), .ZN(n7027) );
  INV_X1 U7732 ( .A(n7030), .ZN(n7028) );
  NOR2_X1 U7733 ( .A1(n7029), .A2(n7023), .ZN(n7022) );
  INV_X1 U7734 ( .A(n8514), .ZN(n7023) );
  NAND2_X1 U7735 ( .A1(n7696), .A2(n6418), .ZN(n7029) );
  AND2_X1 U7736 ( .A1(n9026), .A2(n8521), .ZN(n8522) );
  AND2_X1 U7737 ( .A1(n7681), .A2(n7304), .ZN(n7303) );
  INV_X1 U7738 ( .A(n8896), .ZN(n7682) );
  INV_X1 U7739 ( .A(n7683), .ZN(n7306) );
  INV_X1 U7740 ( .A(n10290), .ZN(n7456) );
  AND2_X1 U7741 ( .A1(n9277), .A2(n6656), .ZN(n9278) );
  NOR2_X1 U7742 ( .A1(n6657), .A2(n11499), .ZN(n6656) );
  INV_X1 U7743 ( .A(n7562), .ZN(n7561) );
  INV_X1 U7744 ( .A(n9055), .ZN(n7566) );
  NAND2_X1 U7745 ( .A1(n7567), .A2(n9054), .ZN(n7563) );
  INV_X1 U7746 ( .A(n7560), .ZN(n7559) );
  OAI21_X1 U7747 ( .B1(n9037), .B2(n9036), .A(n9053), .ZN(n7560) );
  NAND2_X1 U7748 ( .A1(n7257), .A2(n6508), .ZN(n9164) );
  INV_X1 U7749 ( .A(n9167), .ZN(n7257) );
  NAND2_X1 U7750 ( .A1(n7438), .A2(n7437), .ZN(n7436) );
  INV_X1 U7751 ( .A(n14336), .ZN(n7437) );
  INV_X1 U7752 ( .A(n10395), .ZN(n7091) );
  INV_X1 U7753 ( .A(n10394), .ZN(n7088) );
  OAI21_X1 U7754 ( .B1(n7091), .B2(n11505), .A(n11859), .ZN(n7090) );
  INV_X1 U7755 ( .A(n8531), .ZN(n7310) );
  INV_X1 U7756 ( .A(n9040), .ZN(n9136) );
  NAND2_X1 U7757 ( .A1(n8981), .A2(n7030), .ZN(n7024) );
  NAND2_X1 U7758 ( .A1(n6741), .A2(n10684), .ZN(n8496) );
  OR2_X1 U7759 ( .A1(n8470), .A2(n10566), .ZN(n7715) );
  OAI21_X1 U7760 ( .B1(n8470), .B2(n7178), .A(n7177), .ZN(n8472) );
  NAND2_X1 U7761 ( .A1(n8470), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7177) );
  AOI21_X1 U7762 ( .B1(n12946), .B2(n7677), .A(n7676), .ZN(n7675) );
  NAND2_X1 U7763 ( .A1(n10476), .A2(n13122), .ZN(n7704) );
  NAND2_X1 U7764 ( .A1(n10131), .A2(n7609), .ZN(n10453) );
  AND2_X1 U7765 ( .A1(n11421), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U7766 ( .A1(n11914), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7134) );
  NAND2_X1 U7767 ( .A1(n7508), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U7768 ( .A1(n13141), .A2(n6604), .ZN(n13144) );
  INV_X1 U7769 ( .A(n13171), .ZN(n7402) );
  NAND2_X1 U7770 ( .A1(n13270), .A2(n13269), .ZN(n13271) );
  INV_X1 U7771 ( .A(n6491), .ZN(n7653) );
  OR2_X1 U7772 ( .A1(n8413), .A2(n10236), .ZN(n7652) );
  OAI21_X1 U7773 ( .B1(n7653), .B2(n7654), .A(n10123), .ZN(n7650) );
  NOR2_X1 U7774 ( .A1(n7655), .A2(n10319), .ZN(n7654) );
  NOR2_X1 U7775 ( .A1(n7656), .A2(n10236), .ZN(n7655) );
  NOR2_X1 U7776 ( .A1(n8213), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7176) );
  INV_X1 U7777 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7042) );
  INV_X1 U7778 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7872) );
  INV_X1 U7779 ( .A(n8163), .ZN(n7873) );
  OAI21_X1 U7780 ( .B1(n10165), .B2(n7637), .A(n7636), .ZN(n7635) );
  INV_X1 U7781 ( .A(n10170), .ZN(n7636) );
  INV_X1 U7782 ( .A(n7635), .ZN(n7631) );
  INV_X1 U7783 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7866) );
  AND3_X1 U7784 ( .A1(n8056), .A2(n8055), .A3(n8054), .ZN(n10465) );
  INV_X1 U7785 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U7786 ( .A1(n8246), .A2(n7329), .ZN(n7328) );
  OR2_X1 U7787 ( .A1(n13548), .A2(n13362), .ZN(n10123) );
  AOI21_X1 U7788 ( .B1(n7225), .B2(n7230), .A(n6524), .ZN(n6727) );
  AOI21_X1 U7789 ( .B1(n13386), .B2(n7229), .A(n6533), .ZN(n7228) );
  INV_X1 U7790 ( .A(n8333), .ZN(n7229) );
  INV_X1 U7791 ( .A(n13386), .ZN(n7230) );
  NAND2_X1 U7792 ( .A1(n13478), .A2(n13484), .ZN(n13477) );
  NOR2_X1 U7793 ( .A1(n8127), .A2(n6722), .ZN(n6719) );
  AND2_X1 U7794 ( .A1(n8126), .A2(n7637), .ZN(n7218) );
  INV_X1 U7795 ( .A(n7417), .ZN(n7415) );
  INV_X1 U7796 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7892) );
  INV_X1 U7797 ( .A(n7959), .ZN(n7488) );
  INV_X1 U7798 ( .A(n8290), .ZN(n7450) );
  NOR2_X1 U7799 ( .A1(n8381), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n8386) );
  INV_X1 U7800 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8208) );
  NOR2_X1 U7801 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7880) );
  INV_X1 U7802 ( .A(n7004), .ZN(n7002) );
  NAND2_X1 U7803 ( .A1(n7680), .A2(n7679), .ZN(n7678) );
  NOR2_X1 U7804 ( .A1(n9251), .A2(n9252), .ZN(n7679) );
  INV_X1 U7805 ( .A(n9253), .ZN(n7680) );
  NOR2_X1 U7806 ( .A1(n14292), .A2(n12678), .ZN(n6842) );
  OAI21_X1 U7807 ( .B1(n7788), .B2(n7103), .A(n7786), .ZN(n7102) );
  NAND2_X1 U7808 ( .A1(n14127), .A2(n10426), .ZN(n7103) );
  AOI21_X1 U7809 ( .B1(n7789), .B2(n7787), .A(n6445), .ZN(n7786) );
  NAND2_X1 U7810 ( .A1(n7430), .A2(n14070), .ZN(n7429) );
  INV_X1 U7811 ( .A(n7431), .ZN(n7430) );
  AND2_X1 U7812 ( .A1(n6749), .A2(n14063), .ZN(n6747) );
  NAND2_X1 U7813 ( .A1(n14404), .A2(n7432), .ZN(n7431) );
  NAND2_X1 U7814 ( .A1(n6735), .A2(n14148), .ZN(n6734) );
  AOI21_X1 U7815 ( .B1(n14148), .B2(n6737), .A(n6497), .ZN(n6736) );
  INV_X1 U7816 ( .A(n10424), .ZN(n6737) );
  OR2_X1 U7817 ( .A1(n9146), .A2(n13778), .ZN(n9148) );
  AND2_X1 U7818 ( .A1(n7094), .A2(n10418), .ZN(n7093) );
  AND2_X1 U7819 ( .A1(n8818), .A2(n8817), .ZN(n8836) );
  AND2_X1 U7820 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n8817) );
  NOR2_X1 U7821 ( .A1(n11651), .A2(n6836), .ZN(n6835) );
  NAND2_X1 U7822 ( .A1(n6837), .A2(n11656), .ZN(n6836) );
  NAND2_X1 U7823 ( .A1(n11081), .A2(n10357), .ZN(n11640) );
  OR2_X1 U7824 ( .A1(n7158), .A2(n14277), .ZN(n11079) );
  OR2_X1 U7825 ( .A1(n14250), .A2(n14258), .ZN(n14253) );
  NOR2_X1 U7826 ( .A1(n12151), .A2(n7784), .ZN(n7783) );
  INV_X1 U7827 ( .A(n10399), .ZN(n7784) );
  NAND2_X1 U7828 ( .A1(n11858), .A2(n10397), .ZN(n11772) );
  XNOR2_X1 U7829 ( .A(n13948), .B(n11856), .ZN(n11859) );
  OAI21_X1 U7830 ( .B1(n9485), .B2(n9484), .A(n15458), .ZN(n10442) );
  NOR2_X1 U7831 ( .A1(n8571), .A2(n8595), .ZN(n8572) );
  AND3_X1 U7832 ( .A1(n8662), .A2(n8567), .A3(n9316), .ZN(n8573) );
  NOR2_X1 U7833 ( .A1(n9864), .A2(n14546), .ZN(n7166) );
  BUF_X4 U7834 ( .A(n11168), .Z(n12871) );
  INV_X1 U7835 ( .A(n9963), .ZN(n6789) );
  NOR2_X1 U7836 ( .A1(n6522), .A2(n6786), .ZN(n6785) );
  AND2_X1 U7837 ( .A1(n6787), .A2(n9963), .ZN(n6786) );
  AND2_X1 U7838 ( .A1(n10092), .A2(n6852), .ZN(n6851) );
  NOR2_X1 U7839 ( .A1(n6853), .A2(n10095), .ZN(n6852) );
  AND4_X1 U7840 ( .A1(n14809), .A2(n10091), .A3(n14824), .A4(n14839), .ZN(
        n10092) );
  NAND2_X1 U7841 ( .A1(n7849), .A2(n6477), .ZN(n6853) );
  INV_X1 U7842 ( .A(n7823), .ZN(n7822) );
  NOR2_X1 U7843 ( .A1(n15043), .A2(n15036), .ZN(n6798) );
  OR2_X1 U7844 ( .A1(n7553), .A2(n7552), .ZN(n6799) );
  OR2_X1 U7845 ( .A1(n15012), .A2(n14781), .ZN(n7552) );
  NAND2_X1 U7846 ( .A1(n12756), .A2(n7554), .ZN(n7553) );
  NOR2_X1 U7847 ( .A1(n6846), .A2(n6848), .ZN(n6845) );
  INV_X1 U7848 ( .A(n6847), .ZN(n6846) );
  INV_X1 U7849 ( .A(n9795), .ZN(n9538) );
  NOR2_X1 U7850 ( .A1(n7159), .A2(n7544), .ZN(n7543) );
  INV_X1 U7851 ( .A(n7545), .ZN(n7544) );
  NOR2_X1 U7852 ( .A1(n14898), .A2(n15073), .ZN(n7545) );
  AOI21_X1 U7853 ( .B1(n7805), .B2(n7808), .A(n12507), .ZN(n7266) );
  NOR2_X1 U7854 ( .A1(n6425), .A2(n7828), .ZN(n6907) );
  NAND2_X1 U7855 ( .A1(n12299), .A2(n12298), .ZN(n12454) );
  INV_X1 U7856 ( .A(n7827), .ZN(n7826) );
  OAI21_X1 U7857 ( .B1(n12186), .B2(n7828), .A(n12286), .ZN(n7827) );
  INV_X1 U7858 ( .A(n14613), .ZN(n12770) );
  INV_X1 U7859 ( .A(n14615), .ZN(n12289) );
  NAND2_X1 U7860 ( .A1(n6909), .A2(n6910), .ZN(n14910) );
  AOI21_X1 U7861 ( .B1(n6911), .B2(n6913), .A(n6446), .ZN(n6910) );
  OAI21_X1 U7862 ( .B1(n14959), .B2(n6913), .A(n6911), .ZN(n14930) );
  NAND2_X1 U7863 ( .A1(n14959), .A2(n14958), .ZN(n14957) );
  OAI21_X1 U7864 ( .B1(n10963), .B2(P1_D_REG_1__SCAN_IN), .A(n10917), .ZN(
        n11736) );
  NAND2_X1 U7865 ( .A1(n6994), .A2(n9206), .ZN(n6993) );
  INV_X1 U7866 ( .A(n9209), .ZN(n6994) );
  AND2_X1 U7867 ( .A1(n9516), .A2(n9515), .ZN(n9521) );
  NAND2_X1 U7868 ( .A1(n8544), .A2(n6600), .ZN(n9227) );
  INV_X1 U7869 ( .A(n9224), .ZN(n8549) );
  AND2_X1 U7870 ( .A1(n9517), .A2(n9518), .ZN(n9522) );
  NAND2_X1 U7871 ( .A1(n9056), .A2(n12560), .ZN(n7016) );
  OR2_X1 U7872 ( .A1(n9076), .A2(n7011), .ZN(n7010) );
  NAND2_X1 U7873 ( .A1(n7017), .A2(n7012), .ZN(n7011) );
  INV_X1 U7874 ( .A(n7014), .ZN(n7012) );
  AND2_X1 U7875 ( .A1(n8519), .A2(n8518), .ZN(n8982) );
  INV_X1 U7876 ( .A(n6472), .ZN(n7685) );
  INV_X1 U7877 ( .A(n8867), .ZN(n7261) );
  AOI21_X1 U7878 ( .B1(n8493), .B2(n7305), .A(n7265), .ZN(n7264) );
  INV_X1 U7879 ( .A(n8851), .ZN(n7265) );
  NAND2_X1 U7880 ( .A1(n8492), .A2(n8491), .ZN(n8831) );
  AND2_X1 U7881 ( .A1(n9712), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9713) );
  OR2_X1 U7882 ( .A1(n9711), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9712) );
  XNOR2_X1 U7883 ( .A(n8472), .B(SI_3_), .ZN(n8685) );
  NAND2_X1 U7884 ( .A1(n10567), .A2(n10588), .ZN(n7249) );
  NAND2_X1 U7885 ( .A1(n10622), .A2(n10619), .ZN(n11129) );
  NAND2_X1 U7886 ( .A1(n11143), .A2(n11142), .ZN(n11149) );
  AOI21_X1 U7887 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n11453), .A(n11452), .ZN(
        n11580) );
  AND2_X1 U7888 ( .A1(n11575), .A2(n6820), .ZN(n6819) );
  OR2_X1 U7889 ( .A1(n15187), .A2(n15186), .ZN(n15189) );
  OAI21_X1 U7890 ( .B1(n10456), .B2(n6961), .A(n6960), .ZN(n11567) );
  OR2_X1 U7891 ( .A1(n10461), .A2(n15514), .ZN(n7691) );
  NOR2_X1 U7892 ( .A1(n15534), .A2(n12342), .ZN(n7609) );
  NAND2_X1 U7893 ( .A1(n7702), .A2(n6927), .ZN(n6926) );
  INV_X1 U7894 ( .A(n13030), .ZN(n6927) );
  INV_X1 U7895 ( .A(n6929), .ZN(n6928) );
  OAI21_X1 U7896 ( .B1(n6930), .B2(n12963), .A(n7706), .ZN(n6929) );
  AOI21_X1 U7897 ( .B1(n6415), .B2(n7708), .A(n7707), .ZN(n7706) );
  NAND2_X1 U7898 ( .A1(n10454), .A2(n10455), .ZN(n6961) );
  OR2_X1 U7899 ( .A1(n10459), .A2(n13129), .ZN(n10454) );
  OAI21_X1 U7900 ( .B1(n7668), .B2(n6958), .A(n13011), .ZN(n6957) );
  INV_X1 U7901 ( .A(n7669), .ZN(n6958) );
  NAND2_X1 U7902 ( .A1(n6921), .A2(n10322), .ZN(n6920) );
  NAND2_X1 U7903 ( .A1(n10300), .A2(n10299), .ZN(n6918) );
  OR2_X1 U7904 ( .A1(n11098), .A2(n11369), .ZN(n10538) );
  NAND2_X1 U7905 ( .A1(n10268), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7216) );
  OAI21_X1 U7906 ( .B1(n11297), .B2(n11105), .A(n11106), .ZN(n11291) );
  NOR2_X1 U7907 ( .A1(n11291), .A2(n15547), .ZN(n11290) );
  NOR2_X1 U7908 ( .A1(n7496), .A2(n7495), .ZN(n7494) );
  AOI21_X1 U7909 ( .B1(n11330), .B2(n11328), .A(n11329), .ZN(n11332) );
  NOR2_X1 U7910 ( .A1(n6893), .A2(n6897), .ZN(n6892) );
  INV_X1 U7911 ( .A(n11303), .ZN(n6893) );
  OR2_X1 U7912 ( .A1(n7507), .A2(n7506), .ZN(n12077) );
  INV_X1 U7913 ( .A(n12075), .ZN(n7506) );
  AOI21_X1 U7914 ( .B1(n7405), .B2(n12068), .A(n6544), .ZN(n7403) );
  NAND2_X1 U7915 ( .A1(n12070), .A2(n7405), .ZN(n7404) );
  NAND2_X1 U7916 ( .A1(n13201), .A2(n13226), .ZN(n6899) );
  OR2_X1 U7917 ( .A1(n8362), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n13336) );
  OR2_X1 U7918 ( .A1(n8350), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U7919 ( .A1(n7175), .A2(n7874), .ZN(n8296) );
  AND3_X1 U7920 ( .A1(n8254), .A2(n8253), .A3(n8252), .ZN(n13511) );
  INV_X1 U7921 ( .A(n8190), .ZN(n7222) );
  AOI21_X1 U7922 ( .B1(n7224), .B2(n13520), .A(n6519), .ZN(n7223) );
  INV_X1 U7923 ( .A(n8189), .ZN(n7224) );
  NAND2_X1 U7924 ( .A1(n6718), .A2(n7218), .ZN(n8129) );
  NAND2_X1 U7925 ( .A1(n7641), .A2(n8125), .ZN(n7639) );
  INV_X1 U7926 ( .A(n10156), .ZN(n7646) );
  AND2_X1 U7927 ( .A1(n10156), .A2(n10155), .ZN(n10466) );
  INV_X1 U7928 ( .A(SI_7_), .ZN(n7421) );
  NAND2_X1 U7929 ( .A1(n7868), .A2(n7867), .ZN(n8083) );
  INV_X1 U7930 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n7867) );
  INV_X1 U7931 ( .A(n8058), .ZN(n7868) );
  NAND2_X1 U7932 ( .A1(n7865), .A2(n12356), .ZN(n8041) );
  OAI211_X1 U7933 ( .C1(n10265), .C2(SI_3_), .A(n8010), .B(n8009), .ZN(n12354)
         );
  AND3_X2 U7934 ( .A1(n6470), .A2(n6426), .A3(n7982), .ZN(n15526) );
  AND2_X1 U7935 ( .A1(n7234), .A2(n6478), .ZN(n13351) );
  NAND2_X1 U7936 ( .A1(n8359), .A2(n8358), .ZN(n13552) );
  OR2_X1 U7937 ( .A1(n12992), .A2(n13404), .ZN(n13372) );
  NAND2_X1 U7938 ( .A1(n7426), .A2(n8304), .ZN(n13417) );
  AND2_X1 U7939 ( .A1(n8331), .A2(n8330), .ZN(n13419) );
  AND2_X1 U7940 ( .A1(n13398), .A2(n8319), .ZN(n13416) );
  NAND2_X1 U7941 ( .A1(n8289), .A2(n8288), .ZN(n13429) );
  INV_X1 U7942 ( .A(n10220), .ZN(n13438) );
  AOI21_X1 U7943 ( .B1(n7618), .B2(n7616), .A(n7615), .ZN(n7614) );
  INV_X1 U7944 ( .A(n10203), .ZN(n7616) );
  INV_X1 U7945 ( .A(n7618), .ZN(n7617) );
  OR2_X1 U7946 ( .A1(n13465), .A2(n13460), .ZN(n7413) );
  AND2_X1 U7947 ( .A1(n13446), .A2(n8230), .ZN(n7618) );
  OR2_X1 U7948 ( .A1(n13580), .A2(n13501), .ZN(n13459) );
  NAND2_X1 U7950 ( .A1(n8212), .A2(n8211), .ZN(n13585) );
  NAND2_X1 U7951 ( .A1(n7628), .A2(n10195), .ZN(n7626) );
  NAND2_X1 U7952 ( .A1(n10189), .A2(n10195), .ZN(n7627) );
  NAND2_X1 U7953 ( .A1(n8171), .A2(n8170), .ZN(n13536) );
  NAND2_X1 U7954 ( .A1(n7416), .A2(n8143), .ZN(n12469) );
  INV_X1 U7955 ( .A(n12468), .ZN(n7419) );
  NAND2_X1 U7956 ( .A1(n8129), .A2(n7417), .ZN(n7416) );
  AND4_X1 U7957 ( .A1(n8168), .A2(n8167), .A3(n8166), .A4(n8165), .ZN(n12948)
         );
  INV_X1 U7958 ( .A(n6405), .ZN(n8245) );
  OR2_X1 U7959 ( .A1(n10346), .A2(n8453), .ZN(n10525) );
  INV_X1 U7960 ( .A(n15513), .ZN(n15537) );
  INV_X1 U7961 ( .A(n15567), .ZN(n13586) );
  INV_X1 U7962 ( .A(n13687), .ZN(n6635) );
  NOR2_X1 U7963 ( .A1(P3_IR_REG_29__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6634) );
  NAND2_X1 U7964 ( .A1(n7963), .A2(n7962), .ZN(n8371) );
  OR2_X1 U7965 ( .A1(n8356), .A2(n7961), .ZN(n7963) );
  XNOR2_X1 U7966 ( .A(n8424), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U7967 ( .A1(n7957), .A2(n7956), .ZN(n8336) );
  OR2_X1 U7968 ( .A1(n7955), .A2(n12143), .ZN(n7956) );
  XNOR2_X1 U7969 ( .A(n7955), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n8320) );
  AND2_X1 U7970 ( .A1(n7954), .A2(n7953), .ZN(n8306) );
  AOI21_X1 U7971 ( .B1(n7462), .B2(n7464), .A(n6607), .ZN(n7459) );
  NAND2_X1 U7972 ( .A1(n8232), .A2(n7462), .ZN(n7460) );
  AND2_X1 U7973 ( .A1(n8208), .A2(n8220), .ZN(n7713) );
  INV_X1 U7974 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U7975 ( .A1(n7940), .A2(n7939), .ZN(n8243) );
  AOI21_X1 U7976 ( .B1(n7469), .B2(n7471), .A(n7466), .ZN(n7465) );
  INV_X1 U7977 ( .A(n7934), .ZN(n7466) );
  AND2_X1 U7978 ( .A1(n8008), .A2(n6662), .ZN(n6661) );
  AND2_X1 U7979 ( .A1(n7714), .A2(n8092), .ZN(n6662) );
  INV_X1 U7980 ( .A(n7916), .ZN(n7474) );
  INV_X1 U7981 ( .A(n7919), .ZN(n7473) );
  NOR2_X1 U7982 ( .A1(n7475), .A2(n6937), .ZN(n6936) );
  INV_X1 U7983 ( .A(n7914), .ZN(n6937) );
  AND2_X1 U7984 ( .A1(n7921), .A2(n7920), .ZN(n8099) );
  NAND2_X1 U7985 ( .A1(n7479), .A2(n7478), .ZN(n8069) );
  INV_X1 U7986 ( .A(n8066), .ZN(n7478) );
  INV_X1 U7987 ( .A(n8067), .ZN(n7479) );
  OR2_X1 U7988 ( .A1(n8052), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U7989 ( .A1(n7452), .A2(n7910), .ZN(n6964) );
  OAI21_X1 U7990 ( .B1(n8006), .B2(n7453), .A(n8017), .ZN(n7452) );
  NAND2_X1 U7991 ( .A1(n7995), .A2(n6434), .ZN(n6965) );
  AND2_X1 U7992 ( .A1(n7912), .A2(n7911), .ZN(n8048) );
  NAND3_X1 U7993 ( .A1(n6965), .A2(n6964), .A3(n8048), .ZN(n8051) );
  NAND2_X1 U7994 ( .A1(n7995), .A2(n7906), .ZN(n8007) );
  INV_X1 U7995 ( .A(n13854), .ZN(n7526) );
  NOR2_X1 U7996 ( .A1(n7526), .A2(n7523), .ZN(n7522) );
  INV_X1 U7997 ( .A(n13757), .ZN(n7523) );
  OR2_X1 U7998 ( .A1(n13768), .A2(n13767), .ZN(n13765) );
  NOR2_X1 U7999 ( .A1(n7540), .A2(n7539), .ZN(n7538) );
  INV_X1 U8000 ( .A(n13784), .ZN(n7540) );
  INV_X1 U8001 ( .A(n9394), .ZN(n7539) );
  INV_X1 U8002 ( .A(n13785), .ZN(n7537) );
  INV_X1 U8003 ( .A(n6997), .ZN(n7001) );
  OAI21_X1 U8004 ( .B1(n6469), .B2(n7002), .A(n7538), .ZN(n6997) );
  NAND2_X1 U8005 ( .A1(n7538), .A2(n7002), .ZN(n6998) );
  NAND2_X1 U8006 ( .A1(n6983), .A2(n6981), .ZN(n7520) );
  NAND2_X1 U8007 ( .A1(n13767), .A2(n9380), .ZN(n7519) );
  NAND2_X1 U8008 ( .A1(n9408), .A2(n9407), .ZN(n13805) );
  NOR2_X1 U8009 ( .A1(n11896), .A2(n11690), .ZN(n10856) );
  NOR2_X1 U8010 ( .A1(n9267), .A2(n6482), .ZN(n9294) );
  AND2_X1 U8011 ( .A1(n9120), .A2(n9119), .ZN(n13877) );
  AND3_X1 U8012 ( .A1(n9013), .A2(n9012), .A3(n9011), .ZN(n10421) );
  NAND2_X1 U8013 ( .A1(n8676), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9011) );
  AND4_X1 U8014 ( .A1(n8929), .A2(n8928), .A3(n8927), .A4(n8926), .ZN(n12584)
         );
  AND4_X1 U8015 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), .ZN(n12216)
         );
  AND4_X1 U8016 ( .A1(n8782), .A2(n8781), .A3(n8780), .A4(n8779), .ZN(n12152)
         );
  OR2_X1 U8017 ( .A1(n8673), .A2(n10865), .ZN(n8679) );
  OR2_X1 U8018 ( .A1(n8675), .A2(n8674), .ZN(n8678) );
  NAND2_X1 U8019 ( .A1(n15325), .A2(n10874), .ZN(n15338) );
  OAI21_X1 U8020 ( .B1(n15341), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6679), .ZN(
        n15339) );
  NAND2_X1 U8021 ( .A1(n15341), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U8022 ( .A1(n15379), .A2(n11033), .ZN(n15391) );
  NOR2_X1 U8023 ( .A1(n15443), .A2(n7240), .ZN(n7239) );
  AND2_X1 U8024 ( .A1(n15449), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7240) );
  NOR2_X1 U8025 ( .A1(n7239), .A2(n14012), .ZN(n14021) );
  OR2_X1 U8026 ( .A1(n14006), .A2(n14017), .ZN(n14025) );
  INV_X1 U8027 ( .A(n12911), .ZN(n7067) );
  NAND2_X1 U8028 ( .A1(n7792), .A2(n6751), .ZN(n6748) );
  NAND2_X1 U8029 ( .A1(n6753), .A2(n6750), .ZN(n6749) );
  AND3_X1 U8030 ( .A1(n14095), .A2(n14078), .A3(n14077), .ZN(n14079) );
  NOR2_X1 U8031 ( .A1(n14119), .A2(n7431), .ZN(n14086) );
  NOR2_X1 U8032 ( .A1(n14119), .A2(n14312), .ZN(n14103) );
  NOR2_X1 U8033 ( .A1(n14118), .A2(n10381), .ZN(n7793) );
  INV_X1 U8034 ( .A(n10377), .ZN(n6641) );
  INV_X1 U8035 ( .A(n10378), .ZN(n7774) );
  NOR2_X1 U8037 ( .A1(n10422), .A2(n7765), .ZN(n7764) );
  INV_X1 U8038 ( .A(n10419), .ZN(n7765) );
  AND3_X1 U8039 ( .A1(n14429), .A2(n12637), .A3(n6436), .ZN(n14221) );
  NAND2_X1 U8040 ( .A1(n11441), .A2(n9228), .ZN(n6731) );
  AND3_X1 U8041 ( .A1(n8994), .A2(n8993), .A3(n8992), .ZN(n14198) );
  NAND2_X1 U8042 ( .A1(n8676), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U8043 ( .A1(n7781), .A2(n13811), .ZN(n7780) );
  INV_X1 U8044 ( .A(n14433), .ZN(n7781) );
  NAND2_X1 U8045 ( .A1(n10369), .A2(n7778), .ZN(n7777) );
  NOR2_X1 U8046 ( .A1(n10370), .A2(n7779), .ZN(n7778) );
  INV_X1 U8047 ( .A(n10368), .ZN(n7779) );
  NAND2_X1 U8048 ( .A1(n7777), .A2(n7776), .ZN(n14189) );
  AND2_X1 U8049 ( .A1(n7780), .A2(n14233), .ZN(n7776) );
  NAND2_X1 U8050 ( .A1(n6839), .A2(n12637), .ZN(n14263) );
  NAND2_X1 U8051 ( .A1(n8901), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8946) );
  INV_X1 U8052 ( .A(n8903), .ZN(n8901) );
  AOI21_X1 U8053 ( .B1(n7076), .B2(n6424), .A(n6525), .ZN(n7075) );
  NAND2_X1 U8054 ( .A1(n12637), .A2(n12642), .ZN(n14260) );
  OR2_X1 U8055 ( .A1(n10407), .A2(n7803), .ZN(n7082) );
  INV_X1 U8056 ( .A(n7084), .ZN(n7083) );
  OAI21_X1 U8057 ( .B1(n10406), .B2(n7803), .A(n10410), .ZN(n7084) );
  OR2_X1 U8058 ( .A1(n10412), .A2(n9273), .ZN(n12582) );
  OR2_X1 U8059 ( .A1(n6488), .A2(n9279), .ZN(n7071) );
  NOR2_X1 U8060 ( .A1(n12222), .A2(n13851), .ZN(n12552) );
  NAND2_X1 U8061 ( .A1(n11769), .A2(n7181), .ZN(n12213) );
  CLKBUF_X1 U8062 ( .A(n11770), .Z(n6685) );
  NAND2_X1 U8063 ( .A1(n6685), .A2(n11771), .ZN(n11769) );
  NAND2_X1 U8064 ( .A1(n11501), .A2(n10359), .ZN(n11849) );
  OAI21_X1 U8065 ( .B1(n11620), .B2(n7753), .A(n7751), .ZN(n11643) );
  INV_X1 U8066 ( .A(n7117), .ZN(n7753) );
  NAND2_X1 U8067 ( .A1(n10389), .A2(n9275), .ZN(n10353) );
  NAND2_X1 U8068 ( .A1(n10434), .A2(n10433), .ZN(n14252) );
  NAND2_X1 U8069 ( .A1(n9078), .A2(n9077), .ZN(n14089) );
  AND2_X1 U8070 ( .A1(n10442), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10981) );
  OR2_X1 U8071 ( .A1(n12382), .A2(n12598), .ZN(n9326) );
  AND2_X1 U8072 ( .A1(n8576), .A2(n8578), .ZN(n7782) );
  AND2_X1 U8073 ( .A1(n9313), .A2(n9312), .ZN(n9317) );
  NAND2_X1 U8074 ( .A1(n9317), .A2(n9316), .ZN(n9319) );
  INV_X1 U8075 ( .A(n8603), .ZN(n8605) );
  NAND2_X1 U8076 ( .A1(n7315), .A2(n6531), .ZN(n7314) );
  INV_X1 U8077 ( .A(n7735), .ZN(n7734) );
  OAI21_X1 U8078 ( .B1(n14505), .B2(n7736), .A(n14583), .ZN(n7735) );
  INV_X1 U8079 ( .A(n12863), .ZN(n7736) );
  OR2_X1 U8080 ( .A1(n9773), .A2(n9766), .ZN(n9795) );
  INV_X1 U8081 ( .A(n14536), .ZN(n7057) );
  INV_X1 U8082 ( .A(n7058), .ZN(n7055) );
  INV_X1 U8083 ( .A(n7166), .ZN(n9876) );
  INV_X1 U8084 ( .A(n7725), .ZN(n7724) );
  NAND2_X1 U8085 ( .A1(n7166), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9890) );
  INV_X1 U8086 ( .A(n12267), .ZN(n7053) );
  NAND2_X1 U8087 ( .A1(n12267), .A2(n7052), .ZN(n7051) );
  OAI21_X1 U8088 ( .B1(n14463), .B2(n7739), .A(n7737), .ZN(n12812) );
  AOI21_X1 U8089 ( .B1(n7740), .B2(n7738), .A(n6542), .ZN(n7737) );
  INV_X1 U8090 ( .A(n7740), .ZN(n7739) );
  AOI21_X1 U8091 ( .B1(n15596), .B2(n10916), .A(n10915), .ZN(n11738) );
  INV_X1 U8092 ( .A(n10027), .ZN(n9988) );
  NAND2_X1 U8093 ( .A1(n14642), .A2(n7289), .ZN(n10777) );
  OR2_X1 U8094 ( .A1(n14639), .A2(n10694), .ZN(n7289) );
  NOR2_X1 U8095 ( .A1(n6801), .A2(n14647), .ZN(n6807) );
  INV_X1 U8096 ( .A(n14646), .ZN(n6802) );
  NAND2_X1 U8097 ( .A1(n6803), .A2(n6804), .ZN(n6808) );
  NAND2_X1 U8098 ( .A1(n14645), .A2(n10775), .ZN(n6803) );
  AOI21_X1 U8099 ( .B1(n10775), .B2(n6809), .A(n6805), .ZN(n6804) );
  INV_X1 U8100 ( .A(n6811), .ZN(n6809) );
  AOI21_X1 U8101 ( .B1(n11396), .B2(n11395), .A(n11394), .ZN(n11679) );
  OAI21_X1 U8102 ( .B1(n11064), .B2(n11063), .A(n11062), .ZN(n11396) );
  OR2_X1 U8103 ( .A1(n14692), .A2(n10038), .ZN(n7550) );
  AND2_X1 U8104 ( .A1(n14760), .A2(n6462), .ZN(n7850) );
  INV_X1 U8105 ( .A(n14806), .ZN(n14809) );
  NAND2_X1 U8106 ( .A1(n6914), .A2(n6915), .ZN(n14823) );
  NAND2_X1 U8107 ( .A1(n14823), .A2(n14824), .ZN(n14822) );
  NAND2_X1 U8108 ( .A1(n14854), .A2(n14853), .ZN(n14852) );
  AND2_X1 U8109 ( .A1(n7815), .A2(n12722), .ZN(n7814) );
  NAND2_X1 U8110 ( .A1(n14883), .A2(n7817), .ZN(n6857) );
  OR2_X1 U8111 ( .A1(n12721), .A2(n7816), .ZN(n7815) );
  INV_X1 U8112 ( .A(n12457), .ZN(n7808) );
  NAND2_X1 U8113 ( .A1(n9718), .A2(n9717), .ZN(n12183) );
  AND2_X1 U8114 ( .A1(n7811), .A2(n11888), .ZN(n7810) );
  OR2_X1 U8115 ( .A1(n12095), .A2(n7812), .ZN(n7811) );
  INV_X1 U8116 ( .A(n11872), .ZN(n7812) );
  NAND2_X1 U8117 ( .A1(n12090), .A2(n12095), .ZN(n12089) );
  NAND2_X1 U8118 ( .A1(n7833), .A2(n7836), .ZN(n7830) );
  NAND2_X1 U8119 ( .A1(n7804), .A2(n11590), .ZN(n11939) );
  OAI21_X2 U8120 ( .B1(n10015), .B2(n6871), .A(n6869), .ZN(n15234) );
  INV_X1 U8121 ( .A(n6870), .ZN(n6869) );
  OAI22_X1 U8122 ( .A1(n9592), .A2(n10568), .B1(n10660), .B2(n14639), .ZN(
        n6870) );
  OR2_X1 U8123 ( .A1(n10970), .A2(n15146), .ZN(n14918) );
  OR2_X1 U8124 ( .A1(n10970), .A2(n10928), .ZN(n14916) );
  INV_X1 U8125 ( .A(n14918), .ZN(n14962) );
  INV_X1 U8126 ( .A(n14949), .ZN(n14893) );
  AND2_X1 U8127 ( .A1(n10017), .A2(n10016), .ZN(n14974) );
  OR2_X1 U8128 ( .A1(n15143), .A2(n10015), .ZN(n10017) );
  OR2_X1 U8129 ( .A1(n7550), .A2(n7549), .ZN(n7548) );
  INV_X1 U8130 ( .A(n7551), .ZN(n7549) );
  AND2_X1 U8131 ( .A1(n14979), .A2(n6572), .ZN(n7112) );
  NAND2_X1 U8132 ( .A1(n10792), .A2(n9591), .ZN(n7269) );
  INV_X1 U8133 ( .A(n15302), .ZN(n15065) );
  INV_X1 U8134 ( .A(n15308), .ZN(n15007) );
  AND2_X1 U8135 ( .A1(n10954), .A2(n10953), .ZN(n15302) );
  OAI21_X1 U8136 ( .B1(n10963), .B2(P1_D_REG_0__SCAN_IN), .A(n10919), .ZN(
        n11748) );
  OR2_X1 U8137 ( .A1(n14873), .A2(n15282), .ZN(n15297) );
  AND2_X1 U8138 ( .A1(n11207), .A2(n10587), .ZN(n11740) );
  INV_X1 U8139 ( .A(n8557), .ZN(n6995) );
  INV_X1 U8140 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U8141 ( .A1(n9553), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U8142 ( .A1(n9588), .A2(n9587), .ZN(n9598) );
  INV_X1 U8143 ( .A(n7367), .ZN(n7366) );
  NAND2_X1 U8144 ( .A1(n10648), .A2(n10649), .ZN(n10650) );
  NAND2_X1 U8145 ( .A1(n11136), .A2(n11135), .ZN(n11146) );
  NAND2_X1 U8146 ( .A1(n12610), .A2(n12609), .ZN(n12615) );
  AND2_X1 U8147 ( .A1(n12352), .A2(n12353), .ZN(n6967) );
  NAND2_X1 U8148 ( .A1(n7689), .A2(n7688), .ZN(n7690) );
  AND3_X1 U8149 ( .A1(n8217), .A2(n8216), .A3(n8215), .ZN(n13525) );
  INV_X1 U8150 ( .A(n7690), .ZN(n12122) );
  AND4_X1 U8151 ( .A1(n8159), .A2(n8158), .A3(n8157), .A4(n8156), .ZN(n13076)
         );
  OR2_X1 U8152 ( .A1(n11703), .A2(n10519), .ZN(n13103) );
  INV_X1 U8153 ( .A(n13088), .ZN(n13111) );
  NAND2_X1 U8154 ( .A1(n8269), .A2(n8268), .ZN(n13470) );
  AND4_X1 U8155 ( .A1(n8142), .A2(n8141), .A3(n8140), .A4(n8139), .ZN(n13073)
         );
  NAND2_X1 U8156 ( .A1(n7991), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7331) );
  NAND2_X1 U8157 ( .A1(n11274), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11244) );
  INV_X1 U8158 ( .A(n11418), .ZN(n6896) );
  NAND2_X1 U8159 ( .A1(n11302), .A2(n6892), .ZN(n6887) );
  OAI21_X1 U8160 ( .B1(n6706), .B2(n7392), .A(n7390), .ZN(n11486) );
  NAND2_X1 U8161 ( .A1(n11488), .A2(n11487), .ZN(n11913) );
  XNOR2_X1 U8162 ( .A(n13244), .B(n7411), .ZN(n13248) );
  INV_X1 U8163 ( .A(n13303), .ZN(n13329) );
  INV_X1 U8164 ( .A(n7385), .ZN(n13298) );
  NAND2_X1 U8165 ( .A1(n13272), .A2(n13503), .ZN(n6640) );
  NAND2_X1 U8166 ( .A1(n13309), .A2(n7501), .ZN(n7500) );
  OR2_X1 U8167 ( .A1(n13272), .A2(n7499), .ZN(n7498) );
  NAND2_X1 U8168 ( .A1(n13319), .A2(n6454), .ZN(n6882) );
  AND2_X1 U8169 ( .A1(n11113), .A2(n13703), .ZN(n13322) );
  NAND2_X1 U8170 ( .A1(n6884), .A2(n6455), .ZN(n6883) );
  AOI21_X1 U8171 ( .B1(n8405), .B2(n15532), .A(n6609), .ZN(n13343) );
  XNOR2_X1 U8172 ( .A(n7235), .B(n10323), .ZN(n8405) );
  AND2_X1 U8173 ( .A1(n7039), .A2(n7038), .ZN(n13554) );
  AOI21_X1 U8174 ( .B1(n7427), .B2(n15532), .A(n13363), .ZN(n7038) );
  NAND2_X1 U8175 ( .A1(n13551), .A2(n15528), .ZN(n7039) );
  AND3_X1 U8176 ( .A1(n8027), .A2(n8026), .A3(n8025), .ZN(n12311) );
  NAND2_X1 U8177 ( .A1(n13343), .A2(n7647), .ZN(n10350) );
  OR2_X1 U8178 ( .A1(n13346), .A2(n12227), .ZN(n7647) );
  NAND2_X1 U8179 ( .A1(n8311), .A2(n8310), .ZN(n13630) );
  NAND2_X1 U8180 ( .A1(n8295), .A2(n8294), .ZN(n13635) );
  NAND2_X1 U8181 ( .A1(n7420), .A2(SI_22_), .ZN(n8294) );
  NAND2_X1 U8182 ( .A1(n8261), .A2(n8260), .ZN(n13646) );
  INV_X1 U8183 ( .A(n13708), .ZN(n6676) );
  AND2_X1 U8184 ( .A1(n9100), .A2(n9099), .ZN(n14114) );
  OAI21_X1 U8185 ( .B1(n11518), .B2(n6980), .A(n6979), .ZN(n13768) );
  AOI21_X1 U8186 ( .B1(n6986), .B2(n6985), .A(n6459), .ZN(n6979) );
  INV_X1 U8187 ( .A(n6986), .ZN(n6980) );
  NAND2_X1 U8188 ( .A1(n13798), .A2(n13797), .ZN(n13796) );
  NAND2_X1 U8189 ( .A1(n9416), .A2(n9415), .ZN(n13830) );
  NAND2_X1 U8190 ( .A1(n9442), .A2(n6671), .ZN(n13837) );
  NAND2_X1 U8191 ( .A1(n13875), .A2(n6672), .ZN(n6671) );
  OR2_X1 U8192 ( .A1(n13737), .A2(n13741), .ZN(n7856) );
  NAND2_X1 U8193 ( .A1(n9491), .A2(n14239), .ZN(n13926) );
  NOR2_X1 U8194 ( .A1(n9270), .A2(n6618), .ZN(n7187) );
  NAND2_X1 U8195 ( .A1(n9241), .A2(n9240), .ZN(n14050) );
  NAND2_X1 U8196 ( .A1(n9072), .A2(n9071), .ZN(n14083) );
  INV_X1 U8197 ( .A(n14114), .ZN(n14081) );
  INV_X1 U8198 ( .A(n13877), .ZN(n14098) );
  NAND2_X1 U8199 ( .A1(n9052), .A2(n9051), .ZN(n13933) );
  INV_X1 U8200 ( .A(n10417), .ZN(n13937) );
  INV_X1 U8201 ( .A(n12584), .ZN(n13939) );
  INV_X1 U8202 ( .A(n12152), .ZN(n13947) );
  NAND2_X1 U8203 ( .A1(n8676), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U8204 ( .A1(n6461), .A2(n6650), .ZN(n15375) );
  INV_X1 U8205 ( .A(n11046), .ZN(n6650) );
  OR2_X1 U8206 ( .A1(n15396), .A2(n15397), .ZN(n15398) );
  AOI21_X1 U8207 ( .B1(n14029), .B2(n15451), .A(n14031), .ZN(n6689) );
  AOI21_X1 U8208 ( .B1(n14030), .B2(n15402), .A(n6649), .ZN(n14032) );
  OAI21_X1 U8209 ( .B1(n14029), .B2(n15411), .A(n15405), .ZN(n6649) );
  OR2_X1 U8210 ( .A1(n12942), .A2(n14363), .ZN(n14039) );
  OR2_X1 U8211 ( .A1(n15143), .A2(n8666), .ZN(n8582) );
  OAI22_X1 U8212 ( .A1(n12914), .A2(n7067), .B1(n7065), .B2(n9293), .ZN(n7064)
         );
  NOR2_X1 U8213 ( .A1(n10386), .A2(n7067), .ZN(n7065) );
  NOR2_X1 U8214 ( .A1(n12914), .A2(n10435), .ZN(n7066) );
  NAND2_X1 U8215 ( .A1(n9182), .A2(n9181), .ZN(n14298) );
  NAND2_X1 U8216 ( .A1(n15466), .A2(n9490), .ZN(n14239) );
  INV_X1 U8217 ( .A(n10443), .ZN(n9490) );
  NAND2_X1 U8218 ( .A1(n9474), .A2(n9473), .ZN(n15462) );
  AND2_X1 U8219 ( .A1(n11527), .A2(n11192), .ZN(n7727) );
  INV_X1 U8220 ( .A(n11526), .ZN(n11527) );
  INV_X1 U8221 ( .A(n7859), .ZN(n7730) );
  NAND2_X1 U8222 ( .A1(n7729), .A2(n7728), .ZN(n11825) );
  AND2_X1 U8223 ( .A1(n11532), .A2(n7730), .ZN(n7728) );
  NAND2_X1 U8224 ( .A1(n12262), .A2(n12261), .ZN(n12268) );
  NAND2_X1 U8225 ( .A1(n7746), .A2(n7745), .ZN(n14494) );
  AND2_X1 U8226 ( .A1(n14495), .A2(n6444), .ZN(n7745) );
  INV_X1 U8227 ( .A(n14505), .ZN(n7131) );
  AND2_X1 U8228 ( .A1(n11208), .A2(n11740), .ZN(n15236) );
  INV_X1 U8229 ( .A(n14583), .ZN(n7179) );
  AND2_X1 U8230 ( .A1(n15236), .A2(n15302), .ZN(n14586) );
  NAND2_X1 U8231 ( .A1(n9972), .A2(n9971), .ZN(n14603) );
  NAND2_X1 U8232 ( .A1(n9960), .A2(n9959), .ZN(n14604) );
  NAND2_X1 U8233 ( .A1(n9941), .A2(n9940), .ZN(n14605) );
  NAND2_X1 U8234 ( .A1(n9928), .A2(n9927), .ZN(n14606) );
  OR2_X1 U8235 ( .A1(n14538), .A2(n10026), .ZN(n9928) );
  NAND2_X1 U8236 ( .A1(n9910), .A2(n9909), .ZN(n14607) );
  NAND2_X1 U8237 ( .A1(n9816), .A2(n9815), .ZN(n14610) );
  OR2_X1 U8238 ( .A1(n14891), .A2(n10026), .ZN(n9816) );
  INV_X1 U8239 ( .A(n6873), .ZN(n6872) );
  NAND2_X1 U8240 ( .A1(n6623), .A2(n14645), .ZN(n14649) );
  AOI21_X1 U8241 ( .B1(n7277), .B2(n7279), .A(n6608), .ZN(n7275) );
  INV_X1 U8242 ( .A(n6816), .ZN(n6815) );
  NOR2_X1 U8243 ( .A1(n14710), .A2(n14709), .ZN(n14711) );
  NAND2_X1 U8244 ( .A1(n9974), .A2(n9973), .ZN(n14737) );
  INV_X1 U8245 ( .A(n14733), .ZN(n7268) );
  NAND2_X1 U8246 ( .A1(n9962), .A2(n9961), .ZN(n14750) );
  NAND3_X1 U8247 ( .A1(n10660), .A2(n6775), .A3(n6518), .ZN(n6774) );
  MUX2_X1 U8248 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9557), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9558) );
  NAND2_X1 U8249 ( .A1(n10650), .A2(n7357), .ZN(n6824) );
  NAND2_X1 U8250 ( .A1(n10646), .A2(n10647), .ZN(n11127) );
  NAND2_X1 U8251 ( .A1(n7375), .A2(n7374), .ZN(n12405) );
  INV_X1 U8252 ( .A(n15170), .ZN(n7380) );
  NAND2_X1 U8253 ( .A1(n7376), .A2(n7114), .ZN(n15184) );
  NOR2_X1 U8254 ( .A1(n15180), .A2(n7115), .ZN(n7114) );
  INV_X1 U8255 ( .A(n7381), .ZN(n7115) );
  NAND2_X1 U8256 ( .A1(n15194), .A2(n15193), .ZN(n15199) );
  AND2_X1 U8257 ( .A1(n15208), .A2(n7364), .ZN(n7361) );
  INV_X1 U8258 ( .A(n15215), .ZN(n7364) );
  OAI21_X1 U8259 ( .B1(n8965), .B2(n15472), .A(n8669), .ZN(n8696) );
  NAND2_X1 U8260 ( .A1(n8635), .A2(n11345), .ZN(n8636) );
  NAND4_X1 U8261 ( .A1(n9618), .A2(n9617), .A3(n9616), .A4(n9615), .ZN(n9633)
         );
  OR2_X1 U8262 ( .A1(n9614), .A2(n9613), .ZN(n9617) );
  OAI21_X1 U8263 ( .B1(n10455), .B2(n10335), .A(n7144), .ZN(n10132) );
  NAND2_X1 U8264 ( .A1(n10335), .A2(n7145), .ZN(n7144) );
  INV_X1 U8265 ( .A(n10131), .ZN(n7145) );
  INV_X1 U8266 ( .A(n8721), .ZN(n7193) );
  NOR2_X1 U8267 ( .A1(n8724), .A2(n8721), .ZN(n7192) );
  INV_X1 U8268 ( .A(n9663), .ZN(n7602) );
  OR2_X1 U8269 ( .A1(n6782), .A2(n9682), .ZN(n6781) );
  INV_X1 U8270 ( .A(n9680), .ZN(n6782) );
  INV_X1 U8271 ( .A(n8805), .ZN(n7197) );
  INV_X1 U8272 ( .A(n8806), .ZN(n7198) );
  INV_X1 U8273 ( .A(n10154), .ZN(n7334) );
  INV_X1 U8274 ( .A(n8827), .ZN(n7569) );
  NOR2_X1 U8275 ( .A1(n7572), .A2(n7571), .ZN(n7570) );
  AND2_X1 U8276 ( .A1(n8805), .A2(n8806), .ZN(n7199) );
  NAND2_X1 U8277 ( .A1(n9703), .A2(n9702), .ZN(n9720) );
  NOR2_X1 U8278 ( .A1(n9722), .A2(n9719), .ZN(n7588) );
  AND2_X1 U8279 ( .A1(n9737), .A2(n7587), .ZN(n7125) );
  NOR2_X1 U8280 ( .A1(n9752), .A2(n9750), .ZN(n7583) );
  INV_X1 U8281 ( .A(n10182), .ZN(n7345) );
  NAND2_X1 U8282 ( .A1(n6536), .A2(n8865), .ZN(n7575) );
  INV_X1 U8283 ( .A(n8912), .ZN(n7576) );
  NOR2_X1 U8284 ( .A1(n7864), .A2(n9804), .ZN(n9805) );
  NAND2_X1 U8285 ( .A1(n6764), .A2(n6763), .ZN(n9806) );
  AND2_X1 U8286 ( .A1(n9832), .A2(n9831), .ZN(n7108) );
  NOR2_X1 U8287 ( .A1(n7154), .A2(n7153), .ZN(n7152) );
  INV_X1 U8288 ( .A(n10188), .ZN(n7153) );
  NOR2_X1 U8289 ( .A1(n13525), .A2(n13585), .ZN(n7154) );
  NAND2_X1 U8290 ( .A1(n6944), .A2(n10214), .ZN(n6942) );
  NOR2_X1 U8291 ( .A1(n7615), .A2(n10213), .ZN(n6951) );
  AOI21_X1 U8292 ( .B1(n7206), .B2(n7210), .A(n7202), .ZN(n7201) );
  NOR2_X1 U8293 ( .A1(n6422), .A2(n7203), .ZN(n7202) );
  NOR2_X1 U8294 ( .A1(n7596), .A2(n9886), .ZN(n7595) );
  NOR2_X1 U8295 ( .A1(n7596), .A2(n7594), .ZN(n7593) );
  INV_X1 U8296 ( .A(n9887), .ZN(n7594) );
  INV_X1 U8297 ( .A(n6944), .ZN(n6940) );
  INV_X1 U8298 ( .A(n13459), .ZN(n7352) );
  NAND2_X1 U8299 ( .A1(n6772), .A2(n9899), .ZN(n6771) );
  NOR2_X1 U8300 ( .A1(n6772), .A2(n9899), .ZN(n6773) );
  NAND2_X1 U8301 ( .A1(n11642), .A2(n6658), .ZN(n6657) );
  AND2_X1 U8302 ( .A1(n7117), .A2(n11622), .ZN(n6658) );
  AOI21_X1 U8303 ( .B1(n7254), .B2(n9131), .A(n6512), .ZN(n9173) );
  NAND2_X1 U8304 ( .A1(n9172), .A2(n9173), .ZN(n9177) );
  NAND2_X1 U8305 ( .A1(n7606), .A2(n9931), .ZN(n7605) );
  INV_X1 U8306 ( .A(n9932), .ZN(n7606) );
  INV_X1 U8307 ( .A(n8519), .ZN(n7312) );
  NOR2_X1 U8308 ( .A1(n7313), .A2(n7031), .ZN(n7030) );
  INV_X1 U8309 ( .A(n8982), .ZN(n7031) );
  OAI21_X1 U8310 ( .B1(n10572), .B2(P1_DATAO_REG_12__SCAN_IN), .A(n6739), .ZN(
        n6741) );
  OAI21_X1 U8311 ( .B1(n10572), .B2(P1_DATAO_REG_11__SCAN_IN), .A(n6699), .ZN(
        n8495) );
  NAND2_X1 U8312 ( .A1(n10572), .A2(n10731), .ZN(n6699) );
  INV_X1 U8313 ( .A(n11309), .ZN(n7395) );
  INV_X1 U8314 ( .A(SI_2_), .ZN(n7329) );
  INV_X1 U8315 ( .A(n13484), .ZN(n10315) );
  INV_X1 U8316 ( .A(n10427), .ZN(n7787) );
  OR2_X1 U8317 ( .A1(n7096), .A2(n10416), .ZN(n7094) );
  INV_X1 U8318 ( .A(n10353), .ZN(n10986) );
  XNOR2_X1 U8319 ( .A(n10006), .B(n7274), .ZN(n9562) );
  NAND2_X1 U8320 ( .A1(n6978), .A2(n9837), .ZN(n10068) );
  NOR2_X1 U8321 ( .A1(n9902), .A2(n9889), .ZN(n6844) );
  NOR2_X1 U8322 ( .A1(n12671), .A2(n9794), .ZN(n6847) );
  INV_X1 U8323 ( .A(n7026), .ZN(n7025) );
  OAI21_X1 U8324 ( .B1(n7695), .B2(n7027), .A(n7692), .ZN(n7026) );
  NAND2_X1 U8325 ( .A1(n8516), .A2(n15626), .ZN(n8519) );
  INV_X1 U8326 ( .A(n8503), .ZN(n7302) );
  INV_X1 U8327 ( .A(n8483), .ZN(n6972) );
  OAI21_X1 U8328 ( .B1(n10572), .B2(n10595), .A(n6713), .ZN(n8485) );
  NAND2_X1 U8329 ( .A1(n10572), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n6713) );
  OAI21_X1 U8330 ( .B1(n10572), .B2(n10571), .A(n6693), .ZN(n8482) );
  NAND2_X1 U8331 ( .A1(n10572), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6693) );
  INV_X1 U8332 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7971) );
  INV_X1 U8333 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U8334 ( .A1(n7353), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10613) );
  INV_X1 U8335 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7353) );
  AND2_X1 U8336 ( .A1(n10550), .A2(n10551), .ZN(n7705) );
  INV_X1 U8337 ( .A(n13043), .ZN(n7708) );
  INV_X1 U8338 ( .A(n10500), .ZN(n7707) );
  NAND2_X1 U8339 ( .A1(n10548), .A2(n7704), .ZN(n12978) );
  INV_X1 U8340 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n7035) );
  OAI211_X1 U8341 ( .C1(n10292), .C2(n10324), .A(n7457), .B(n7454), .ZN(n10293) );
  OAI21_X1 U8342 ( .B1(n10320), .B2(n13335), .A(n7458), .ZN(n7457) );
  NOR2_X1 U8343 ( .A1(n10291), .A2(n7455), .ZN(n7454) );
  NAND2_X1 U8344 ( .A1(n11255), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6680) );
  NAND2_X1 U8345 ( .A1(n13229), .A2(n7411), .ZN(n7493) );
  NAND2_X1 U8346 ( .A1(n13234), .A2(n13233), .ZN(n13258) );
  AND2_X1 U8347 ( .A1(n7385), .A2(n7384), .ZN(n13325) );
  NAND2_X1 U8348 ( .A1(n13300), .A2(n13299), .ZN(n7384) );
  NAND2_X1 U8349 ( .A1(n6723), .A2(n6727), .ZN(n13361) );
  NAND2_X1 U8350 ( .A1(n8334), .A2(n7225), .ZN(n6723) );
  NOR2_X1 U8351 ( .A1(n8324), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8323) );
  NOR2_X1 U8352 ( .A1(n8262), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7175) );
  AND2_X1 U8353 ( .A1(n15627), .A2(n7046), .ZN(n7045) );
  INV_X1 U8354 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7046) );
  AND2_X1 U8355 ( .A1(n6594), .A2(n7034), .ZN(n7033) );
  INV_X1 U8356 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n7034) );
  INV_X1 U8357 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7869) );
  INV_X1 U8358 ( .A(n8104), .ZN(n7870) );
  NAND2_X1 U8359 ( .A1(n7217), .A2(n15515), .ZN(n10455) );
  INV_X1 U8360 ( .A(n15526), .ZN(n7217) );
  NAND2_X1 U8361 ( .A1(n13350), .A2(n6478), .ZN(n7232) );
  NAND2_X1 U8362 ( .A1(n10243), .A2(n10237), .ZN(n10318) );
  INV_X1 U8363 ( .A(n10225), .ZN(n7613) );
  INV_X1 U8364 ( .A(n7614), .ZN(n7612) );
  AND2_X1 U8365 ( .A1(n10200), .A2(n8410), .ZN(n13482) );
  NAND2_X1 U8366 ( .A1(n13680), .A2(n13121), .ZN(n10187) );
  NAND2_X1 U8367 ( .A1(n6721), .A2(n6452), .ZN(n11839) );
  INV_X1 U8368 ( .A(n7463), .ZN(n7462) );
  OAI21_X1 U8369 ( .B1(n7944), .B2(n7464), .A(n8218), .ZN(n7463) );
  INV_X1 U8370 ( .A(n7945), .ZN(n7464) );
  AND2_X1 U8371 ( .A1(n7713), .A2(n7712), .ZN(n7711) );
  INV_X1 U8372 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7712) );
  INV_X1 U8373 ( .A(n7470), .ZN(n7469) );
  OAI21_X1 U8374 ( .B1(n7928), .B2(n7471), .A(n7930), .ZN(n7470) );
  INV_X1 U8375 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8092) );
  INV_X1 U8376 ( .A(n7326), .ZN(n7889) );
  OR2_X1 U8377 ( .A1(n8019), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8021) );
  NOR2_X1 U8378 ( .A1(n6985), .A2(n6459), .ZN(n6984) );
  INV_X1 U8379 ( .A(n6982), .ZN(n6981) );
  OAI21_X1 U8380 ( .B1(n6986), .B2(n6459), .A(n9380), .ZN(n6982) );
  OR4_X1 U8381 ( .A1(n14220), .A2(n14233), .A3(n14258), .A4(n9284), .ZN(n9286)
         );
  OR4_X1 U8382 ( .A1(n12546), .A2(n9280), .A3(n12151), .A4(n12215), .ZN(n9281)
         );
  AOI21_X1 U8383 ( .B1(n9038), .B2(n6509), .A(n7186), .ZN(n7185) );
  INV_X1 U8384 ( .A(n7557), .ZN(n7186) );
  NOR2_X1 U8385 ( .A1(n9164), .A2(n9135), .ZN(n9160) );
  NOR2_X1 U8386 ( .A1(n9158), .A2(n7862), .ZN(n7256) );
  NOR2_X1 U8387 ( .A1(n15432), .A2(n7247), .ZN(n13990) );
  AND2_X1 U8388 ( .A1(n15437), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7247) );
  INV_X1 U8389 ( .A(n7796), .ZN(n7795) );
  OAI21_X1 U8390 ( .B1(n7798), .B2(n7797), .A(n10383), .ZN(n7796) );
  OR2_X1 U8391 ( .A1(n14089), .A2(n14096), .ZN(n10383) );
  NOR2_X1 U8392 ( .A1(n14377), .A2(n14433), .ZN(n6839) );
  OR2_X1 U8393 ( .A1(n7181), .A2(n6488), .ZN(n7070) );
  XNOR2_X1 U8394 ( .A(n13950), .B(n11656), .ZN(n11639) );
  NOR2_X1 U8395 ( .A1(n7434), .A2(n7436), .ZN(n14150) );
  INV_X1 U8396 ( .A(n7090), .ZN(n7089) );
  NOR2_X1 U8397 ( .A1(n7091), .A2(n7088), .ZN(n7087) );
  NAND2_X1 U8398 ( .A1(n11504), .A2(n10395), .ZN(n11860) );
  NAND2_X1 U8399 ( .A1(n8597), .A2(n7119), .ZN(n8587) );
  INV_X1 U8400 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7119) );
  INV_X1 U8401 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7535) );
  OR2_X1 U8402 ( .A1(n8871), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U8403 ( .A1(n11172), .A2(n11173), .ZN(n11354) );
  INV_X1 U8404 ( .A(n9890), .ZN(n9888) );
  INV_X1 U8405 ( .A(n12261), .ZN(n7052) );
  AND2_X1 U8406 ( .A1(n12803), .A2(n7741), .ZN(n7740) );
  NAND2_X1 U8407 ( .A1(n14464), .A2(n12791), .ZN(n7741) );
  INV_X1 U8408 ( .A(n12791), .ZN(n7738) );
  OAI211_X1 U8409 ( .C1(n14697), .C2(n10068), .A(n6976), .B(n10062), .ZN(
        n10073) );
  NAND2_X1 U8410 ( .A1(n6977), .A2(n14697), .ZN(n6976) );
  INV_X1 U8411 ( .A(n10065), .ZN(n6977) );
  NAND2_X1 U8412 ( .A1(n10706), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6810) );
  INV_X1 U8413 ( .A(n6810), .ZN(n6805) );
  NOR2_X1 U8414 ( .A1(n7284), .A2(n11390), .ZN(n7280) );
  NOR2_X1 U8415 ( .A1(n14670), .A2(n6667), .ZN(n7292) );
  AND2_X1 U8416 ( .A1(n14671), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6667) );
  INV_X1 U8417 ( .A(n14745), .ZN(n7821) );
  OR2_X1 U8418 ( .A1(n9953), .A2(n9952), .ZN(n9982) );
  OR2_X1 U8419 ( .A1(n9934), .A2(n9933), .ZN(n9953) );
  NAND2_X1 U8420 ( .A1(n9888), .A2(n6844), .ZN(n9921) );
  NAND2_X1 U8421 ( .A1(n12719), .A2(n12718), .ZN(n7816) );
  NOR2_X1 U8422 ( .A1(n12721), .A2(n9829), .ZN(n7817) );
  NAND2_X1 U8423 ( .A1(n9538), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U8424 ( .A1(n6759), .A2(n6758), .ZN(n6757) );
  OR2_X1 U8425 ( .A1(n7266), .A2(n6480), .ZN(n6864) );
  INV_X1 U8426 ( .A(n7805), .ZN(n6867) );
  NOR2_X1 U8427 ( .A1(n12515), .A2(n15092), .ZN(n6759) );
  NOR2_X1 U8428 ( .A1(n11391), .A2(n9723), .ZN(n6843) );
  INV_X1 U8429 ( .A(n9724), .ZN(n9537) );
  NOR2_X1 U8430 ( .A1(n12183), .A2(n12101), .ZN(n6794) );
  INV_X1 U8431 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9704) );
  OR2_X1 U8432 ( .A1(n9705), .A2(n9704), .ZN(n9724) );
  NAND2_X1 U8433 ( .A1(n7835), .A2(n11601), .ZN(n7834) );
  INV_X1 U8434 ( .A(n11599), .ZN(n7835) );
  INV_X1 U8435 ( .A(n11601), .ZN(n7836) );
  NAND2_X1 U8436 ( .A1(n6900), .A2(n10935), .ZN(n10942) );
  AOI21_X1 U8437 ( .B1(n14986), .B2(n15302), .A(n14985), .ZN(n7551) );
  AND2_X1 U8438 ( .A1(n14983), .A2(n14977), .ZN(n14975) );
  NAND2_X1 U8439 ( .A1(n14855), .A2(n6798), .ZN(n14829) );
  NAND2_X1 U8440 ( .A1(n12725), .A2(n12724), .ZN(n14840) );
  NOR2_X1 U8441 ( .A1(n11949), .A2(n15234), .ZN(n11959) );
  NAND2_X1 U8442 ( .A1(n9209), .A2(n6991), .ZN(n6990) );
  INV_X1 U8443 ( .A(n9206), .ZN(n6991) );
  NAND2_X1 U8444 ( .A1(n7750), .A2(n7541), .ZN(n10099) );
  AOI21_X1 U8445 ( .B1(n6481), .B2(n7313), .A(n7694), .ZN(n7308) );
  NAND2_X1 U8446 ( .A1(n7589), .A2(n7750), .ZN(n9559) );
  AND2_X1 U8447 ( .A1(n6473), .A2(n7590), .ZN(n7589) );
  NOR2_X1 U8448 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n7590) );
  INV_X1 U8449 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U8450 ( .A1(n8520), .A2(n8519), .ZN(n9003) );
  OR2_X1 U8451 ( .A1(n9817), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n9807) );
  AND2_X1 U8452 ( .A1(n8509), .A2(n8506), .ZN(n8938) );
  OR2_X1 U8453 ( .A1(n9659), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9674) );
  NAND2_X1 U8454 ( .A1(n7161), .A2(n8476), .ZN(n6970) );
  NAND2_X1 U8455 ( .A1(n8685), .A2(n8473), .ZN(n7162) );
  NAND2_X1 U8456 ( .A1(n7315), .A2(n10593), .ZN(n6665) );
  INV_X1 U8457 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10559) );
  AND2_X1 U8458 ( .A1(n10617), .A2(n10616), .ZN(n10628) );
  INV_X1 U8459 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7147) );
  AOI21_X1 U8460 ( .B1(n11151), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n11150), .ZN(
        n11451) );
  OAI22_X1 U8461 ( .A1(n12612), .A2(n12611), .B1(P1_ADDR_REG_12__SCAN_IN), 
        .B2(n13160), .ZN(n15163) );
  OR2_X1 U8462 ( .A1(n15175), .A2(n15174), .ZN(n15178) );
  NAND2_X1 U8463 ( .A1(n10549), .A2(n7705), .ZN(n10548) );
  INV_X1 U8464 ( .A(n10498), .ZN(n7709) );
  NAND2_X1 U8465 ( .A1(n13044), .A2(n13043), .ZN(n7710) );
  AOI21_X1 U8466 ( .B1(n7675), .B2(n7673), .A(n6438), .ZN(n7672) );
  INV_X1 U8467 ( .A(n7677), .ZN(n7673) );
  AND2_X1 U8468 ( .A1(n7672), .A2(n6484), .ZN(n7668) );
  NAND2_X1 U8469 ( .A1(n7666), .A2(n7665), .ZN(n7664) );
  INV_X1 U8470 ( .A(n7667), .ZN(n7666) );
  NAND2_X1 U8471 ( .A1(n7667), .A2(n12956), .ZN(n13018) );
  INV_X1 U8472 ( .A(n6924), .ZN(n13029) );
  NAND2_X1 U8473 ( .A1(n12954), .A2(n12953), .ZN(n12955) );
  NAND2_X1 U8474 ( .A1(n7870), .A2(n6594), .ZN(n8137) );
  NAND2_X1 U8475 ( .A1(n11567), .A2(n6962), .ZN(n11566) );
  INV_X1 U8476 ( .A(n6963), .ZN(n6962) );
  OAI21_X1 U8477 ( .B1(n10509), .B2(n10457), .A(n15531), .ZN(n6963) );
  OR2_X1 U8478 ( .A1(n10484), .A2(n13121), .ZN(n7677) );
  INV_X1 U8479 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8383) );
  AND2_X1 U8480 ( .A1(n8369), .A2(n8368), .ZN(n12902) );
  OAI21_X1 U8481 ( .B1(n7497), .B2(P3_REG1_REG_2__SCAN_IN), .A(n6703), .ZN(
        n11119) );
  NAND2_X1 U8482 ( .A1(n7497), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8483 ( .A1(n11285), .A2(n7860), .ZN(n11118) );
  NAND2_X1 U8484 ( .A1(n11119), .A2(n11118), .ZN(n11241) );
  AND2_X1 U8485 ( .A1(n7410), .A2(n7409), .ZN(n11101) );
  NAND2_X1 U8486 ( .A1(n8394), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7409) );
  OR2_X1 U8487 ( .A1(n13703), .A2(n15547), .ZN(n7410) );
  XNOR2_X1 U8488 ( .A(n11101), .B(n7124), .ZN(n11287) );
  NAND2_X1 U8489 ( .A1(n11275), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U8490 ( .A1(n6706), .A2(n11266), .ZN(n11311) );
  INV_X1 U8491 ( .A(n7135), .ZN(n11249) );
  NAND2_X1 U8492 ( .A1(n6878), .A2(n11246), .ZN(n11299) );
  CLKBUF_X1 U8493 ( .A(n11265), .Z(n6706) );
  NAND2_X1 U8494 ( .A1(n7389), .A2(n7393), .ZN(n11432) );
  NAND2_X1 U8495 ( .A1(n6706), .A2(n6467), .ZN(n7389) );
  INV_X1 U8496 ( .A(n6892), .ZN(n6889) );
  AND2_X1 U8497 ( .A1(n11424), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U8498 ( .A1(n7141), .A2(n11912), .ZN(n12065) );
  NAND2_X1 U8499 ( .A1(n12073), .A2(n12074), .ZN(n13141) );
  NAND2_X1 U8500 ( .A1(n7512), .A2(n13161), .ZN(n13146) );
  NAND2_X1 U8501 ( .A1(n7514), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n13163) );
  INV_X1 U8502 ( .A(n13146), .ZN(n7514) );
  AND2_X1 U8503 ( .A1(n13212), .A2(n13213), .ZN(n7412) );
  XNOR2_X1 U8504 ( .A(n13258), .B(n7411), .ZN(n13236) );
  NOR2_X1 U8505 ( .A1(n13236), .A2(n13235), .ZN(n13257) );
  NOR2_X1 U8506 ( .A1(n13257), .A2(n6669), .ZN(n13261) );
  AND2_X1 U8507 ( .A1(n13258), .A2(n7411), .ZN(n6669) );
  NAND2_X1 U8508 ( .A1(n13261), .A2(n13260), .ZN(n13273) );
  OR2_X1 U8509 ( .A1(n13276), .A2(n13277), .ZN(n7385) );
  NAND2_X1 U8510 ( .A1(n6702), .A2(n13295), .ZN(n6701) );
  NAND2_X1 U8511 ( .A1(n6625), .A2(n7501), .ZN(n7499) );
  INV_X1 U8512 ( .A(n6624), .ZN(n7501) );
  OAI21_X1 U8513 ( .B1(n6886), .B2(n13318), .A(n6453), .ZN(n6885) );
  INV_X1 U8514 ( .A(n7650), .ZN(n7649) );
  NOR2_X1 U8515 ( .A1(n7653), .A2(n7652), .ZN(n7651) );
  NAND2_X1 U8516 ( .A1(n12633), .A2(n15535), .ZN(n8404) );
  AOI21_X1 U8517 ( .B1(n13349), .B2(n8375), .A(n7901), .ZN(n13362) );
  XNOR2_X1 U8518 ( .A(n13361), .B(n10319), .ZN(n7427) );
  NAND2_X1 U8519 ( .A1(n8334), .A2(n8333), .ZN(n13385) );
  AOI21_X1 U8520 ( .B1(n13375), .B2(n8375), .A(n8354), .ZN(n13387) );
  OR2_X1 U8521 ( .A1(n8312), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8324) );
  OR2_X1 U8522 ( .A1(n8296), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8312) );
  INV_X1 U8523 ( .A(n7175), .ZN(n8280) );
  NAND2_X1 U8524 ( .A1(n7176), .A2(n7043), .ZN(n8262) );
  AND2_X1 U8525 ( .A1(n7045), .A2(n7044), .ZN(n7043) );
  INV_X1 U8526 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7044) );
  INV_X1 U8527 ( .A(n7176), .ZN(n8249) );
  AND2_X1 U8528 ( .A1(n6450), .A2(n7041), .ZN(n7040) );
  INV_X1 U8529 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7041) );
  NAND2_X1 U8530 ( .A1(n7873), .A2(n6450), .ZN(n8197) );
  NAND2_X1 U8531 ( .A1(n7873), .A2(n7872), .ZN(n8183) );
  NAND2_X1 U8532 ( .A1(n7870), .A2(n7032), .ZN(n8163) );
  AND2_X1 U8533 ( .A1(n7033), .A2(n7871), .ZN(n7032) );
  INV_X1 U8534 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n7871) );
  NOR2_X1 U8535 ( .A1(n7635), .A2(n7644), .ZN(n7633) );
  NAND2_X1 U8536 ( .A1(n7870), .A2(n7869), .ZN(n8118) );
  OR2_X1 U8537 ( .A1(n8083), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8104) );
  AND4_X1 U8538 ( .A1(n8034), .A2(n8033), .A3(n8032), .A4(n8031), .ZN(n11790)
         );
  AND2_X1 U8539 ( .A1(n10151), .A2(n10152), .ZN(n11709) );
  INV_X1 U8540 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U8541 ( .A1(n11725), .A2(n8011), .ZN(n12307) );
  NAND2_X1 U8542 ( .A1(n15510), .A2(n6715), .ZN(n11725) );
  NOR2_X1 U8543 ( .A1(n11722), .A2(n6716), .ZN(n6715) );
  INV_X1 U8544 ( .A(n11727), .ZN(n6716) );
  INV_X1 U8545 ( .A(n11722), .ZN(n11726) );
  OR2_X1 U8546 ( .A1(n11098), .A2(n15567), .ZN(n11703) );
  INV_X1 U8547 ( .A(n15536), .ZN(n7330) );
  INV_X1 U8548 ( .A(n7609), .ZN(n15527) );
  NAND2_X1 U8549 ( .A1(n10455), .A2(n10131), .ZN(n15530) );
  NAND2_X1 U8550 ( .A1(n10267), .A2(n10266), .ZN(n10286) );
  NAND2_X1 U8551 ( .A1(n10123), .A2(n8415), .ZN(n13350) );
  INV_X1 U8552 ( .A(n6727), .ZN(n6726) );
  AOI21_X1 U8553 ( .B1(n6727), .B2(n7226), .A(n6725), .ZN(n6724) );
  INV_X1 U8554 ( .A(n7232), .ZN(n7233) );
  NAND2_X1 U8555 ( .A1(n7227), .A2(n7228), .ZN(n13377) );
  OR2_X1 U8556 ( .A1(n8334), .A2(n7230), .ZN(n7227) );
  NAND2_X1 U8557 ( .A1(n13379), .A2(n15537), .ZN(n6631) );
  INV_X1 U8558 ( .A(n10318), .ZN(n13376) );
  AND2_X1 U8559 ( .A1(n10231), .A2(n13383), .ZN(n13401) );
  NAND2_X1 U8560 ( .A1(n13414), .A2(n13416), .ZN(n13413) );
  OR2_X1 U8561 ( .A1(n10205), .A2(n10208), .ZN(n13428) );
  AND2_X1 U8562 ( .A1(n8286), .A2(n8285), .ZN(n13454) );
  AND2_X1 U8563 ( .A1(n8230), .A2(n10206), .ZN(n13460) );
  NAND2_X1 U8564 ( .A1(n7219), .A2(n7220), .ZN(n13463) );
  AOI21_X1 U8565 ( .B1(n6416), .B2(n10311), .A(n6526), .ZN(n7220) );
  NAND2_X1 U8566 ( .A1(n8190), .A2(n6416), .ZN(n7219) );
  INV_X1 U8567 ( .A(n13482), .ZN(n13496) );
  AOI21_X1 U8568 ( .B1(n6414), .B2(n7415), .A(n6485), .ZN(n7414) );
  OR2_X1 U8569 ( .A1(n10190), .A2(n10184), .ZN(n12564) );
  INV_X1 U8570 ( .A(n10466), .ZN(n11791) );
  NAND2_X1 U8571 ( .A1(n8418), .A2(n8417), .ZN(n10529) );
  NOR2_X1 U8572 ( .A1(n10347), .A2(n8453), .ZN(n10527) );
  INV_X1 U8573 ( .A(n8205), .ZN(n7323) );
  AND2_X1 U8574 ( .A1(n8008), .A2(n7212), .ZN(n7324) );
  AOI21_X1 U8575 ( .B1(n7482), .B2(n7481), .A(n6616), .ZN(n7480) );
  INV_X1 U8576 ( .A(n8372), .ZN(n7481) );
  AOI21_X1 U8577 ( .B1(n7487), .B2(n7958), .A(n6619), .ZN(n7486) );
  INV_X1 U8578 ( .A(n8394), .ZN(n13214) );
  NAND2_X1 U8579 ( .A1(n8431), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8425) );
  XNOR2_X1 U8580 ( .A(n8423), .B(n8422), .ZN(n11094) );
  INV_X1 U8581 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8422) );
  OAI21_X1 U8582 ( .B1(n8421), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8423) );
  XNOR2_X1 U8583 ( .A(n8385), .B(P3_IR_REG_21__SCAN_IN), .ZN(n11704) );
  OR2_X1 U8584 ( .A1(n8389), .A2(n13686), .ZN(n8385) );
  INV_X1 U8585 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8382) );
  INV_X1 U8586 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8179) );
  OR2_X1 U8587 ( .A1(n8178), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8193) );
  OR2_X1 U8588 ( .A1(n8147), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U8589 ( .A1(n7927), .A2(n7926), .ZN(n8146) );
  NAND2_X1 U8590 ( .A1(n6938), .A2(n7921), .ZN(n8112) );
  AND2_X1 U8591 ( .A1(n7923), .A2(n7922), .ZN(n8111) );
  AND2_X1 U8592 ( .A1(n8008), .A2(n7889), .ZN(n8093) );
  NAND2_X1 U8593 ( .A1(n7146), .A2(n7914), .ZN(n8067) );
  XNOR2_X1 U8594 ( .A(n7517), .B(n7981), .ZN(n11297) );
  AND2_X1 U8595 ( .A1(n9438), .A2(n9437), .ZN(n13736) );
  INV_X1 U8596 ( .A(n9371), .ZN(n6985) );
  AOI21_X1 U8597 ( .B1(n11517), .B2(n9371), .A(n6987), .ZN(n6986) );
  INV_X1 U8598 ( .A(n11796), .ZN(n6987) );
  NAND2_X1 U8599 ( .A1(n11864), .A2(n9338), .ZN(n9344) );
  INV_X1 U8600 ( .A(n6673), .ZN(n6672) );
  OAI21_X1 U8601 ( .B1(n9439), .B2(n14098), .A(n13874), .ZN(n6673) );
  NAND2_X1 U8602 ( .A1(n13736), .A2(n6975), .ZN(n9441) );
  OR2_X1 U8603 ( .A1(n9439), .A2(n9440), .ZN(n6975) );
  NAND2_X1 U8604 ( .A1(n8775), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8816) );
  INV_X1 U8605 ( .A(n10985), .ZN(n7164) );
  OR2_X1 U8606 ( .A1(n8883), .A2(n8882), .ZN(n8903) );
  NAND2_X1 U8607 ( .A1(n7006), .A2(n7005), .ZN(n7004) );
  INV_X1 U8608 ( .A(n9387), .ZN(n7005) );
  INV_X1 U8609 ( .A(n9388), .ZN(n7006) );
  INV_X1 U8610 ( .A(n9386), .ZN(n7003) );
  OR2_X1 U8611 ( .A1(n13886), .A2(n13885), .ZN(n13883) );
  XNOR2_X1 U8612 ( .A(n9344), .B(n14277), .ZN(n9340) );
  AOI21_X1 U8613 ( .B1(n13797), .B2(n9445), .A(n9450), .ZN(n7531) );
  NOR2_X1 U8614 ( .A1(n7532), .A2(n7530), .ZN(n7529) );
  INV_X1 U8615 ( .A(n13836), .ZN(n7530) );
  INV_X1 U8616 ( .A(n13797), .ZN(n7532) );
  INV_X1 U8617 ( .A(n13891), .ZN(n13917) );
  NAND2_X1 U8618 ( .A1(n6554), .A2(n7700), .ZN(n7188) );
  OR2_X1 U8619 ( .A1(n9294), .A2(n7678), .ZN(n7861) );
  AND3_X1 U8620 ( .A1(n8973), .A2(n8972), .A3(n8971), .ZN(n10417) );
  NAND2_X1 U8621 ( .A1(n8676), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8971) );
  AND4_X1 U8622 ( .A1(n8844), .A2(n8843), .A3(n8842), .A4(n8841), .ZN(n12422)
         );
  AND4_X1 U8623 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(n12547)
         );
  OAI21_X1 U8624 ( .B1(n15322), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6692), .ZN(
        n15327) );
  NAND2_X1 U8625 ( .A1(n15322), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U8626 ( .A1(n15327), .A2(n15326), .ZN(n15325) );
  NAND2_X1 U8627 ( .A1(n15337), .A2(n10876), .ZN(n15350) );
  INV_X1 U8628 ( .A(n15392), .ZN(n6686) );
  NOR2_X1 U8629 ( .A1(n15419), .A2(n7248), .ZN(n15434) );
  AND2_X1 U8630 ( .A1(n15424), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7248) );
  NAND2_X1 U8631 ( .A1(n6708), .A2(n6707), .ZN(n14026) );
  INV_X1 U8632 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6707) );
  XNOR2_X1 U8633 ( .A(n14024), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14030) );
  NAND2_X1 U8634 ( .A1(n10440), .A2(n6842), .ZN(n14042) );
  NAND2_X1 U8635 ( .A1(n10440), .A2(n6439), .ZN(n14040) );
  NAND2_X1 U8636 ( .A1(n10440), .A2(n14398), .ZN(n12923) );
  INV_X1 U8637 ( .A(n10440), .ZN(n14052) );
  AOI21_X1 U8638 ( .B1(n7102), .B2(n10430), .A(n6539), .ZN(n7097) );
  AND2_X1 U8639 ( .A1(n9184), .A2(n9066), .ZN(n14068) );
  NAND2_X1 U8640 ( .A1(n6752), .A2(n6747), .ZN(n6745) );
  AND2_X1 U8641 ( .A1(n6747), .A2(n10427), .ZN(n6746) );
  AND2_X1 U8642 ( .A1(n10429), .A2(n10380), .ZN(n7798) );
  OR2_X1 U8643 ( .A1(n9287), .A2(n10381), .ZN(n14117) );
  NAND2_X1 U8644 ( .A1(n9044), .A2(n9043), .ZN(n9146) );
  INV_X1 U8645 ( .A(n9046), .ZN(n9044) );
  OR2_X1 U8646 ( .A1(n9009), .A2(n9008), .ZN(n9046) );
  INV_X1 U8647 ( .A(n7764), .ZN(n7758) );
  NAND2_X1 U8648 ( .A1(n7761), .A2(n6479), .ZN(n7759) );
  NAND2_X1 U8649 ( .A1(n14221), .A2(n7438), .ZN(n14177) );
  NAND2_X1 U8650 ( .A1(n14221), .A2(n14352), .ZN(n14207) );
  OAI21_X1 U8651 ( .B1(n7138), .B2(n10420), .A(n10419), .ZN(n14187) );
  OR2_X1 U8652 ( .A1(n14222), .A2(n13936), .ZN(n10372) );
  INV_X1 U8653 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8945) );
  OR3_X1 U8654 ( .A1(n8946), .A2(n12252), .A3(n8945), .ZN(n8969) );
  NOR2_X1 U8655 ( .A1(n7445), .A2(n12554), .ZN(n12637) );
  NOR2_X1 U8656 ( .A1(n12440), .A2(n13793), .ZN(n12587) );
  NAND2_X1 U8657 ( .A1(n12420), .A2(n10409), .ZN(n12437) );
  NAND2_X1 U8658 ( .A1(n7446), .A2(n7443), .ZN(n12440) );
  INV_X1 U8659 ( .A(n12554), .ZN(n7446) );
  NAND2_X1 U8660 ( .A1(n10407), .A2(n10406), .ZN(n12420) );
  NAND2_X1 U8661 ( .A1(n8836), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8883) );
  NAND3_X1 U8662 ( .A1(n6834), .A2(n6835), .A3(n15488), .ZN(n12222) );
  NOR2_X1 U8663 ( .A1(n13821), .A2(n12159), .ZN(n6834) );
  INV_X1 U8664 ( .A(n11859), .ZN(n11848) );
  INV_X1 U8665 ( .A(n13821), .ZN(n7073) );
  INV_X1 U8666 ( .A(n11499), .ZN(n11505) );
  NAND2_X1 U8667 ( .A1(n11641), .A2(n10394), .ZN(n11506) );
  NAND2_X1 U8668 ( .A1(n11506), .A2(n11505), .ZN(n11504) );
  AND2_X1 U8669 ( .A1(n11654), .A2(n11632), .ZN(n11853) );
  NOR2_X1 U8670 ( .A1(n11651), .A2(n15478), .ZN(n11654) );
  INV_X1 U8671 ( .A(n11639), .ZN(n11642) );
  OR2_X1 U8672 ( .A1(n11615), .A2(n11667), .ZN(n11651) );
  NOR2_X1 U8673 ( .A1(n9338), .A2(n11587), .ZN(n11664) );
  NAND2_X1 U8674 ( .A1(n9336), .A2(n11587), .ZN(n11864) );
  XNOR2_X1 U8675 ( .A(n9337), .B(n11896), .ZN(n9336) );
  NOR2_X1 U8676 ( .A1(n14277), .A2(n11345), .ZN(n11616) );
  OR2_X1 U8677 ( .A1(n14055), .A2(n14054), .ZN(n14297) );
  NAND2_X1 U8678 ( .A1(n14253), .A2(n10416), .ZN(n14234) );
  AND2_X1 U8679 ( .A1(n14255), .A2(n14254), .ZN(n14371) );
  NAND2_X1 U8680 ( .A1(n10369), .A2(n10368), .ZN(n14259) );
  NAND2_X1 U8681 ( .A1(n7785), .A2(n10399), .ZN(n12150) );
  BUF_X1 U8682 ( .A(n9328), .Z(n10859) );
  OR2_X1 U8683 ( .A1(n8832), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U8684 ( .A1(n14440), .A2(n7243), .ZN(n7242) );
  INV_X1 U8685 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7243) );
  INV_X1 U8686 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9766) );
  NAND2_X1 U8687 ( .A1(n7743), .A2(n7742), .ZN(n14461) );
  INV_X1 U8688 ( .A(n14464), .ZN(n7742) );
  INV_X1 U8689 ( .A(n14463), .ZN(n7743) );
  XNOR2_X1 U8690 ( .A(n12826), .B(n12866), .ZN(n12828) );
  NAND2_X1 U8691 ( .A1(n12825), .A2(n12824), .ZN(n12826) );
  NAND2_X1 U8692 ( .A1(n14573), .A2(n14574), .ZN(n7726) );
  INV_X1 U8693 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9684) );
  OR2_X1 U8694 ( .A1(n9685), .A2(n9684), .ZN(n9705) );
  AOI21_X1 U8695 ( .B1(n7059), .B2(n6417), .A(n6471), .ZN(n7058) );
  NAND2_X1 U8696 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9640) );
  OAI21_X1 U8697 ( .B1(n6900), .B2(n12855), .A(n10750), .ZN(n10751) );
  AOI22_X1 U8698 ( .A1(n11176), .A2(n10935), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n10752), .ZN(n10750) );
  NAND2_X1 U8699 ( .A1(n9538), .A2(n6451), .ZN(n9864) );
  INV_X1 U8700 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14546) );
  INV_X1 U8701 ( .A(n14565), .ZN(n7716) );
  XNOR2_X1 U8702 ( .A(n7048), .B(n12875), .ZN(n11159) );
  OAI22_X1 U8703 ( .A1(n11218), .A2(n12755), .B1(n11152), .B2(n12857), .ZN(
        n7048) );
  OR2_X1 U8704 ( .A1(n10970), .A2(n10952), .ZN(n11206) );
  NAND2_X1 U8705 ( .A1(n11441), .A2(n9591), .ZN(n9535) );
  NAND2_X1 U8706 ( .A1(n14461), .A2(n12791), .ZN(n14513) );
  OR2_X1 U8707 ( .A1(n10073), .A2(n10056), .ZN(n10060) );
  NAND2_X1 U8708 ( .A1(n6784), .A2(n6783), .ZN(n9996) );
  AOI21_X1 U8709 ( .B1(n6785), .B2(n6788), .A(n6545), .ZN(n6783) );
  AND2_X1 U8710 ( .A1(n9964), .A2(n6789), .ZN(n6788) );
  OR2_X1 U8711 ( .A1(n10058), .A2(n10061), .ZN(n10054) );
  XNOR2_X1 U8712 ( .A(n6849), .B(n7274), .ZN(n10098) );
  NOR2_X1 U8713 ( .A1(n12707), .A2(n10093), .ZN(n6854) );
  AND2_X1 U8714 ( .A1(n9896), .A2(n9895), .ZN(n14797) );
  OR2_X1 U8715 ( .A1(n14813), .A2(n10026), .ZN(n9896) );
  OAI22_X1 U8716 ( .A1(n10704), .A2(n6403), .B1(n10026), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U8717 ( .A1(n11678), .A2(n11677), .ZN(n7281) );
  NAND2_X1 U8718 ( .A1(n11386), .A2(n7280), .ZN(n7282) );
  NOR2_X1 U8719 ( .A1(n11679), .A2(n6596), .ZN(n11681) );
  NAND2_X1 U8720 ( .A1(n11681), .A2(n11682), .ZN(n11974) );
  NOR2_X1 U8721 ( .A1(n7278), .A2(n11970), .ZN(n7277) );
  NOR2_X1 U8722 ( .A1(n7280), .A2(n7279), .ZN(n7278) );
  INV_X1 U8723 ( .A(n7281), .ZN(n7279) );
  NAND2_X1 U8724 ( .A1(n12656), .A2(n7285), .ZN(n12659) );
  OR2_X1 U8725 ( .A1(n12657), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7285) );
  NAND2_X1 U8726 ( .A1(n7292), .A2(n14672), .ZN(n7291) );
  NAND2_X1 U8727 ( .A1(n14668), .A2(n6615), .ZN(n14683) );
  XNOR2_X1 U8728 ( .A(n9982), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n14736) );
  XNOR2_X1 U8729 ( .A(n14603), .B(n14737), .ZN(n14728) );
  NOR2_X1 U8730 ( .A1(n14728), .A2(n7824), .ZN(n7823) );
  INV_X1 U8731 ( .A(n12733), .ZN(n7824) );
  NAND2_X1 U8732 ( .A1(n14744), .A2(n14745), .ZN(n7825) );
  NAND2_X1 U8733 ( .A1(n6797), .A2(n6796), .ZN(n14746) );
  AND2_X1 U8734 ( .A1(n14855), .A2(n6569), .ZN(n6796) );
  INV_X1 U8735 ( .A(n6799), .ZN(n6797) );
  NAND2_X1 U8736 ( .A1(n14756), .A2(n12732), .ZN(n14744) );
  NAND2_X1 U8737 ( .A1(n12700), .A2(n7849), .ZN(n7848) );
  OR2_X1 U8738 ( .A1(n7850), .A2(n7847), .ZN(n7846) );
  INV_X1 U8739 ( .A(n12700), .ZN(n7847) );
  NOR2_X1 U8740 ( .A1(n14829), .A2(n6799), .ZN(n14762) );
  NOR3_X1 U8741 ( .A1(n14829), .A2(n7553), .A3(n14781), .ZN(n14779) );
  NOR2_X1 U8742 ( .A1(n14829), .A2(n7553), .ZN(n14795) );
  XNOR2_X1 U8743 ( .A(n15025), .B(n14607), .ZN(n14793) );
  NOR2_X1 U8744 ( .A1(n14837), .A2(n7845), .ZN(n7844) );
  INV_X1 U8745 ( .A(n12694), .ZN(n7845) );
  NAND2_X1 U8746 ( .A1(n14855), .A2(n14846), .ZN(n14845) );
  AND3_X1 U8747 ( .A1(n14903), .A2(n7542), .A3(n7543), .ZN(n14855) );
  NAND2_X1 U8748 ( .A1(n14903), .A2(n7545), .ZN(n14894) );
  NOR2_X2 U8749 ( .A1(n6757), .A2(n15078), .ZN(n14903) );
  NAND2_X1 U8750 ( .A1(n14903), .A2(n14909), .ZN(n14904) );
  INV_X1 U8751 ( .A(n14931), .ZN(n14927) );
  OAI21_X1 U8752 ( .B1(n6644), .B2(n6868), .A(n6866), .ZN(n14945) );
  INV_X1 U8753 ( .A(n7266), .ZN(n6868) );
  INV_X1 U8754 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9770) );
  OR2_X1 U8755 ( .A1(n9771), .A2(n9770), .ZN(n9773) );
  INV_X1 U8756 ( .A(n6905), .ZN(n6904) );
  OAI21_X1 U8757 ( .B1(n7826), .B2(n6425), .A(n12508), .ZN(n6905) );
  NAND2_X1 U8758 ( .A1(n9537), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U8759 ( .A1(n9537), .A2(n6843), .ZN(n9753) );
  AND3_X1 U8760 ( .A1(n12112), .A2(n6793), .A3(n6420), .ZN(n12514) );
  NAND2_X1 U8761 ( .A1(n12188), .A2(n12287), .ZN(n6908) );
  NAND2_X1 U8762 ( .A1(n12112), .A2(n6420), .ZN(n12291) );
  NAND2_X1 U8763 ( .A1(n6863), .A2(n7809), .ZN(n12178) );
  AOI21_X1 U8764 ( .B1(n7810), .B2(n7812), .A(n6523), .ZN(n7809) );
  NAND2_X1 U8765 ( .A1(n12090), .A2(n7810), .ZN(n6863) );
  NAND2_X1 U8766 ( .A1(n12178), .A2(n12187), .ZN(n12297) );
  NAND2_X1 U8767 ( .A1(n12112), .A2(n12103), .ZN(n12098) );
  AND2_X1 U8768 ( .A1(n12111), .A2(n12115), .ZN(n12112) );
  NAND2_X1 U8769 ( .A1(n11870), .A2(n11869), .ZN(n12109) );
  NAND2_X1 U8770 ( .A1(n9536), .A2(n6430), .ZN(n9667) );
  NAND2_X1 U8771 ( .A1(n9536), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9653) );
  NOR2_X1 U8772 ( .A1(n12042), .A2(n12012), .ZN(n12111) );
  INV_X1 U8773 ( .A(n14620), .ZN(n11600) );
  INV_X1 U8774 ( .A(n11878), .ZN(n11602) );
  NAND2_X1 U8775 ( .A1(n7832), .A2(n11601), .ZN(n11879) );
  NAND2_X1 U8776 ( .A1(n12037), .A2(n11599), .ZN(n7832) );
  NAND2_X1 U8777 ( .A1(n11963), .A2(n11959), .ZN(n12044) );
  NAND2_X1 U8778 ( .A1(n6761), .A2(n6760), .ZN(n12042) );
  INV_X1 U8779 ( .A(n12044), .ZN(n6761) );
  NAND2_X1 U8780 ( .A1(n11957), .A2(n6861), .ZN(n6859) );
  INV_X1 U8781 ( .A(n11591), .ZN(n6861) );
  INV_X1 U8782 ( .A(n14916), .ZN(n14960) );
  OAI21_X1 U8783 ( .B1(n11014), .B2(n11152), .A(n11218), .ZN(n10937) );
  NAND2_X1 U8784 ( .A1(n6762), .A2(n11218), .ZN(n11949) );
  AND2_X1 U8785 ( .A1(n11909), .A2(n11225), .ZN(n6762) );
  NAND2_X1 U8786 ( .A1(n11909), .A2(n11218), .ZN(n11016) );
  INV_X1 U8787 ( .A(n14622), .ZN(n11596) );
  NAND2_X1 U8788 ( .A1(n6776), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U8789 ( .A1(n14930), .A2(n12688), .ZN(n14912) );
  NAND2_X1 U8790 ( .A1(n14957), .A2(n12687), .ZN(n14932) );
  NAND2_X1 U8791 ( .A1(n12092), .A2(n11887), .ZN(n11889) );
  AND2_X1 U8792 ( .A1(n11738), .A2(n10918), .ZN(n10959) );
  XNOR2_X1 U8793 ( .A(n9213), .B(n9212), .ZN(n12894) );
  NAND2_X1 U8794 ( .A1(n8544), .A2(n8543), .ZN(n9225) );
  OR2_X1 U8795 ( .A1(n7015), .A2(n7014), .ZN(n7009) );
  INV_X1 U8796 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10100) );
  XNOR2_X1 U8797 ( .A(n9143), .B(n9142), .ZN(n11689) );
  OR2_X1 U8798 ( .A1(n9762), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n9789) );
  OAI21_X1 U8799 ( .B1(n8831), .B2(n7685), .A(n7683), .ZN(n8897) );
  INV_X1 U8800 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9527) );
  OAI21_X1 U8801 ( .B1(n7263), .B2(n7260), .A(n7258), .ZN(n8870) );
  AOI21_X1 U8802 ( .B1(n7259), .B2(n8830), .A(n8498), .ZN(n7258) );
  NAND2_X1 U8803 ( .A1(n7262), .A2(n7264), .ZN(n8868) );
  OR2_X1 U8804 ( .A1(n8492), .A2(n8830), .ZN(n7262) );
  AND2_X1 U8805 ( .A1(n9716), .A2(n9730), .ZN(n11002) );
  NAND2_X1 U8806 ( .A1(n8686), .A2(n8471), .ZN(n7252) );
  NAND2_X1 U8807 ( .A1(n7249), .A2(n6513), .ZN(n8465) );
  OR2_X1 U8808 ( .A1(n7359), .A2(n10620), .ZN(n7358) );
  NAND2_X1 U8809 ( .A1(n11148), .A2(n11147), .ZN(n11448) );
  NAND2_X1 U8810 ( .A1(n11445), .A2(n13970), .ZN(n7356) );
  AOI21_X1 U8811 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n11582), .A(n11581), .ZN(
        n12024) );
  NAND2_X1 U8812 ( .A1(n6818), .A2(n12021), .ZN(n6817) );
  AND3_X1 U8813 ( .A1(n8241), .A2(n8240), .A3(n8239), .ZN(n13501) );
  AND4_X1 U8814 ( .A1(n8065), .A2(n8064), .A3(n8063), .A4(n8062), .ZN(n12483)
         );
  NAND2_X1 U8815 ( .A1(n7710), .A2(n10498), .ZN(n12970) );
  OAI21_X1 U8816 ( .B1(n12945), .B2(n7674), .A(n7672), .ZN(n13005) );
  NAND2_X1 U8817 ( .A1(n7669), .A2(n6955), .ZN(n13012) );
  NAND2_X1 U8818 ( .A1(n12945), .A2(n7668), .ZN(n6955) );
  AND2_X1 U8819 ( .A1(n8345), .A2(n8344), .ZN(n13404) );
  AOI21_X1 U8820 ( .B1(n10504), .B2(n10503), .A(n10502), .ZN(n13021) );
  OR2_X1 U8821 ( .A1(n10538), .A2(n10523), .ZN(n13098) );
  NAND2_X1 U8822 ( .A1(n6931), .A2(n10495), .ZN(n13044) );
  NAND2_X1 U8823 ( .A1(n12964), .A2(n12963), .ZN(n6931) );
  AND2_X1 U8824 ( .A1(n7701), .A2(n6926), .ZN(n6925) );
  AOI21_X1 U8825 ( .B1(n7702), .B2(n6429), .A(n6537), .ZN(n7701) );
  NAND2_X1 U8826 ( .A1(n6956), .A2(n6958), .ZN(n6954) );
  INV_X1 U8827 ( .A(n13115), .ZN(n13095) );
  INV_X1 U8828 ( .A(n13109), .ZN(n13100) );
  INV_X1 U8829 ( .A(n13103), .ZN(n13112) );
  AND2_X1 U8830 ( .A1(n10328), .A2(n6918), .ZN(n6917) );
  NAND2_X1 U8831 ( .A1(n6921), .A2(n10298), .ZN(n6916) );
  INV_X1 U8832 ( .A(n13362), .ZN(n12633) );
  INV_X1 U8833 ( .A(n12902), .ZN(n13379) );
  INV_X1 U8834 ( .A(n13387), .ZN(n13118) );
  INV_X1 U8835 ( .A(n13404), .ZN(n13378) );
  INV_X1 U8836 ( .A(n13419), .ZN(n13119) );
  INV_X1 U8837 ( .A(n13454), .ZN(n13065) );
  INV_X1 U8838 ( .A(n13511), .ZN(n13487) );
  INV_X1 U8839 ( .A(n13525), .ZN(n13498) );
  INV_X1 U8840 ( .A(n12948), .ZN(n13537) );
  INV_X1 U8841 ( .A(n12483), .ZN(n13124) );
  INV_X1 U8842 ( .A(n11790), .ZN(n13125) );
  NAND2_X1 U8843 ( .A1(n8060), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7215) );
  NAND2_X1 U8844 ( .A1(n8061), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7214) );
  NOR2_X1 U8845 ( .A1(n11235), .A2(n11115), .ZN(n11286) );
  NAND2_X1 U8846 ( .A1(n7123), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n11285) );
  AOI21_X1 U8847 ( .B1(n7390), .B2(n7392), .A(n7388), .ZN(n7387) );
  INV_X1 U8848 ( .A(n11485), .ZN(n7388) );
  XNOR2_X1 U8849 ( .A(n12065), .B(n12067), .ZN(n12066) );
  NAND2_X1 U8850 ( .A1(n7508), .A2(n12075), .ZN(n11924) );
  NAND2_X1 U8851 ( .A1(n6881), .A2(n6880), .ZN(n13132) );
  NAND2_X1 U8852 ( .A1(n12065), .A2(n11922), .ZN(n6880) );
  NAND2_X1 U8853 ( .A1(n12066), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n6881) );
  AOI21_X1 U8854 ( .B1(n12070), .B2(n12069), .A(n12068), .ZN(n13137) );
  NAND2_X1 U8855 ( .A1(n7404), .A2(n7403), .ZN(n13172) );
  INV_X1 U8856 ( .A(n7399), .ZN(n7398) );
  NAND2_X1 U8857 ( .A1(n12070), .A2(n6440), .ZN(n7396) );
  OAI21_X1 U8858 ( .B1(n6466), .B2(n7400), .A(n13173), .ZN(n7399) );
  INV_X1 U8859 ( .A(n7397), .ZN(n13174) );
  AOI21_X1 U8860 ( .B1(n7404), .B2(n6466), .A(n7400), .ZN(n7397) );
  OR2_X1 U8861 ( .A1(n13130), .A2(n11100), .ZN(n13303) );
  NAND2_X1 U8862 ( .A1(n7503), .A2(n6419), .ZN(n13310) );
  NAND2_X1 U8863 ( .A1(n7976), .A2(n7975), .ZN(n13548) );
  NAND2_X1 U8864 ( .A1(n8322), .A2(n8321), .ZN(n13565) );
  NAND2_X1 U8865 ( .A1(n7221), .A2(n7223), .ZN(n13508) );
  NAND2_X1 U8866 ( .A1(n7222), .A2(n13520), .ZN(n7221) );
  NAND2_X1 U8867 ( .A1(n8129), .A2(n8128), .ZN(n12488) );
  INV_X1 U8868 ( .A(n7634), .ZN(n12228) );
  AOI21_X1 U8869 ( .B1(n7640), .B2(n7638), .A(n10167), .ZN(n7634) );
  INV_X1 U8870 ( .A(n7639), .ZN(n7638) );
  AOI21_X1 U8871 ( .B1(n11792), .B2(n10466), .A(n7646), .ZN(n11837) );
  AND3_X1 U8872 ( .A1(n8075), .A2(n8074), .A3(n8073), .ZN(n12366) );
  NAND2_X1 U8873 ( .A1(n8246), .A2(n7421), .ZN(n8074) );
  INV_X1 U8874 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n12356) );
  INV_X1 U8875 ( .A(n12166), .ZN(n12084) );
  OR2_X1 U8876 ( .A1(n11703), .A2(n15543), .ZN(n15509) );
  INV_X1 U8877 ( .A(n15524), .ZN(n15549) );
  INV_X1 U8878 ( .A(n15509), .ZN(n15544) );
  INV_X1 U8879 ( .A(n12480), .ZN(n12338) );
  INV_X1 U8880 ( .A(n10286), .ZN(n13604) );
  OAI211_X1 U8881 ( .C1(n13556), .C2(n13555), .A(n13554), .B(n13553), .ZN(
        n13612) );
  AOI21_X1 U8882 ( .B1(n6632), .B2(n15532), .A(n6629), .ZN(n13613) );
  NAND2_X1 U8883 ( .A1(n6631), .A2(n6630), .ZN(n6629) );
  XNOR2_X1 U8884 ( .A(n13377), .B(n13376), .ZN(n6632) );
  NAND2_X1 U8885 ( .A1(n13378), .A2(n15535), .ZN(n6630) );
  INV_X1 U8886 ( .A(n12992), .ZN(n13622) );
  NAND2_X1 U8887 ( .A1(n7426), .A2(n7424), .ZN(n13421) );
  NAND2_X1 U8888 ( .A1(n7420), .A2(SI_21_), .ZN(n8278) );
  OAI21_X1 U8889 ( .B1(n6668), .B2(n7617), .A(n7614), .ZN(n13436) );
  NAND2_X1 U8890 ( .A1(n7619), .A2(n7618), .ZN(n13445) );
  AND2_X1 U8891 ( .A1(n7619), .A2(n8230), .ZN(n13447) );
  NAND2_X1 U8892 ( .A1(n6668), .A2(n10203), .ZN(n7619) );
  INV_X1 U8893 ( .A(n13462), .ZN(n13651) );
  NAND2_X1 U8894 ( .A1(n8248), .A2(n8247), .ZN(n13660) );
  NAND2_X1 U8895 ( .A1(n7625), .A2(n7626), .ZN(n13506) );
  OR2_X1 U8896 ( .A1(n13531), .A2(n7627), .ZN(n7625) );
  NAND2_X1 U8897 ( .A1(n8190), .A2(n8189), .ZN(n13521) );
  NAND2_X1 U8898 ( .A1(n8196), .A2(n8195), .ZN(n13669) );
  NAND2_X1 U8899 ( .A1(n13530), .A2(n10189), .ZN(n13517) );
  NAND2_X1 U8900 ( .A1(n8162), .A2(n8161), .ZN(n13058) );
  NAND2_X1 U8901 ( .A1(n7416), .A2(n6414), .ZN(n12471) );
  INV_X1 U8902 ( .A(n8124), .ZN(n13038) );
  NAND2_X1 U8903 ( .A1(n7640), .A2(n7641), .ZN(n11803) );
  OAI21_X1 U8904 ( .B1(n8441), .B2(P3_D_REG_0__SCAN_IN), .A(n6968), .ZN(n10610) );
  OR2_X1 U8905 ( .A1(n8439), .A2(n8440), .ZN(n6968) );
  NAND2_X1 U8906 ( .A1(n11094), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13683) );
  OR2_X1 U8907 ( .A1(n7893), .A2(n6637), .ZN(n6636) );
  NOR2_X1 U8908 ( .A1(n6635), .A2(n6634), .ZN(n6633) );
  INV_X1 U8909 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U8910 ( .A1(n7489), .A2(n7959), .ZN(n8347) );
  OR2_X1 U8911 ( .A1(n8336), .A2(n7958), .ZN(n7489) );
  INV_X1 U8912 ( .A(n8434), .ZN(n12452) );
  INV_X1 U8913 ( .A(SI_23_), .ZN(n11785) );
  NAND2_X1 U8914 ( .A1(n8293), .A2(n7951), .ZN(n8307) );
  NAND2_X1 U8915 ( .A1(n7949), .A2(n7948), .ZN(n8291) );
  INV_X1 U8916 ( .A(n10338), .ZN(n11459) );
  INV_X1 U8917 ( .A(n11704), .ZN(n11766) );
  INV_X1 U8918 ( .A(SI_19_), .ZN(n12934) );
  NAND2_X1 U8919 ( .A1(n7461), .A2(n7945), .ZN(n8219) );
  NAND2_X1 U8920 ( .A1(n8232), .A2(n7944), .ZN(n7461) );
  INV_X1 U8921 ( .A(SI_18_), .ZN(n11013) );
  NAND2_X1 U8922 ( .A1(n8209), .A2(n7713), .ZN(n8233) );
  INV_X1 U8923 ( .A(SI_17_), .ZN(n15626) );
  INV_X1 U8924 ( .A(SI_15_), .ZN(n10786) );
  INV_X1 U8925 ( .A(SI_13_), .ZN(n10800) );
  NAND2_X1 U8926 ( .A1(n6934), .A2(n7472), .ZN(n8100) );
  NAND2_X1 U8927 ( .A1(n7146), .A2(n6936), .ZN(n6934) );
  NAND2_X1 U8928 ( .A1(n8069), .A2(n7916), .ZN(n8096) );
  XNOR2_X1 U8929 ( .A(n8036), .B(n8035), .ZN(n11421) );
  AND2_X1 U8930 ( .A1(n6965), .A2(n6964), .ZN(n8049) );
  NAND2_X1 U8931 ( .A1(n7908), .A2(n7451), .ZN(n8018) );
  NAND2_X1 U8932 ( .A1(n8007), .A2(n8006), .ZN(n7451) );
  NAND2_X1 U8933 ( .A1(n8019), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6879) );
  INV_X1 U8934 ( .A(n7903), .ZN(n7978) );
  CLKBUF_X1 U8935 ( .A(n11297), .Z(n7124) );
  AND4_X1 U8936 ( .A1(n8908), .A2(n8907), .A3(n8906), .A4(n8905), .ZN(n13730)
         );
  NAND2_X1 U8937 ( .A1(n13843), .A2(n9386), .ZN(n13748) );
  NAND2_X1 U8938 ( .A1(n11463), .A2(n9348), .ZN(n11348) );
  XNOR2_X1 U8939 ( .A(n9350), .B(n9351), .ZN(n11347) );
  NOR3_X1 U8940 ( .A1(n9457), .A2(n13709), .A3(n9465), .ZN(n9489) );
  INV_X1 U8941 ( .A(n7525), .ZN(n7524) );
  OAI21_X1 U8942 ( .B1(n13756), .B2(n7526), .A(n13855), .ZN(n7525) );
  AND2_X1 U8943 ( .A1(n13883), .A2(n9394), .ZN(n13786) );
  NAND2_X1 U8944 ( .A1(n13835), .A2(n9446), .ZN(n13798) );
  NAND2_X1 U8945 ( .A1(n13837), .A2(n13836), .ZN(n13835) );
  NAND2_X1 U8946 ( .A1(n13765), .A2(n9380), .ZN(n13844) );
  NAND2_X1 U8947 ( .A1(n7527), .A2(n13756), .ZN(n13856) );
  NAND2_X1 U8948 ( .A1(n7163), .A2(n13757), .ZN(n7527) );
  AND2_X1 U8949 ( .A1(n7536), .A2(n6998), .ZN(n6999) );
  AOI21_X1 U8950 ( .B1(n7538), .B2(n13885), .A(n7537), .ZN(n7536) );
  INV_X1 U8951 ( .A(n9437), .ZN(n7165) );
  INV_X1 U8952 ( .A(n13919), .ZN(n13888) );
  NAND2_X1 U8953 ( .A1(n11339), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13891) );
  NAND2_X1 U8954 ( .A1(n7000), .A2(n7004), .ZN(n13886) );
  NAND2_X1 U8955 ( .A1(n13843), .A2(n6469), .ZN(n7000) );
  NAND2_X1 U8956 ( .A1(n11464), .A2(n11465), .ZN(n11463) );
  AND2_X1 U8957 ( .A1(n9348), .A2(n9347), .ZN(n11465) );
  OR2_X1 U8958 ( .A1(n9346), .A2(n9345), .ZN(n9347) );
  NAND2_X1 U8959 ( .A1(n13830), .A2(n9421), .ZN(n13896) );
  NAND2_X1 U8960 ( .A1(n13830), .A2(n7528), .ZN(n13897) );
  AND2_X1 U8961 ( .A1(n9084), .A2(n9083), .ZN(n13913) );
  NAND2_X1 U8962 ( .A1(n7020), .A2(n7531), .ZN(n13907) );
  NAND2_X1 U8963 ( .A1(n9495), .A2(n9494), .ZN(n13919) );
  AND3_X1 U8964 ( .A1(n7107), .A2(n9291), .A3(n6563), .ZN(n9295) );
  INV_X1 U8965 ( .A(n9294), .ZN(n7107) );
  NAND2_X1 U8966 ( .A1(n8676), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8612) );
  INV_X1 U8967 ( .A(n13913), .ZN(n14096) );
  INV_X1 U8968 ( .A(n13730), .ZN(n13940) );
  INV_X1 U8969 ( .A(n12422), .ZN(n13943) );
  INV_X1 U8970 ( .A(n12547), .ZN(n13944) );
  OR2_X1 U8971 ( .A1(n9234), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8680) );
  AND3_X1 U8972 ( .A1(n8678), .A2(n8679), .A3(n8677), .ZN(n8681) );
  OAI21_X1 U8973 ( .B1(n15322), .B2(P2_REG2_REG_1__SCAN_IN), .A(n6653), .ZN(
        n15331) );
  NAND2_X1 U8974 ( .A1(n15322), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U8975 ( .A1(n15358), .A2(n15359), .ZN(n15357) );
  NAND2_X1 U8976 ( .A1(n10887), .A2(n10886), .ZN(n13959) );
  NAND2_X1 U8977 ( .A1(n15371), .A2(n15372), .ZN(n15370) );
  NAND2_X1 U8978 ( .A1(n15375), .A2(n11047), .ZN(n15396) );
  NAND2_X1 U8979 ( .A1(n6652), .A2(n6651), .ZN(n15413) );
  INV_X1 U8980 ( .A(n15409), .ZN(n6651) );
  AND2_X1 U8981 ( .A1(n15404), .A2(n15403), .ZN(n15407) );
  NOR2_X1 U8982 ( .A1(n15407), .A2(n7245), .ZN(n11036) );
  AND2_X1 U8983 ( .A1(n11050), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7245) );
  AND2_X1 U8984 ( .A1(n12240), .A2(n12239), .ZN(n15427) );
  XNOR2_X1 U8985 ( .A(n12243), .B(n12242), .ZN(n15438) );
  NOR2_X1 U8986 ( .A1(n7237), .A2(n14021), .ZN(n14013) );
  NAND2_X1 U8987 ( .A1(n14013), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n14023) );
  XNOR2_X1 U8988 ( .A(n10387), .B(n10386), .ZN(n12684) );
  AOI21_X1 U8989 ( .B1(n7170), .B2(n14252), .A(n7167), .ZN(n14305) );
  NAND2_X1 U8990 ( .A1(n7169), .A2(n7168), .ZN(n7167) );
  XNOR2_X1 U8991 ( .A(n14064), .B(n14071), .ZN(n7170) );
  NAND2_X1 U8992 ( .A1(n14096), .A2(n14097), .ZN(n7168) );
  XNOR2_X1 U8993 ( .A(n14076), .B(n14078), .ZN(n14309) );
  NAND2_X1 U8994 ( .A1(n14314), .A2(n10382), .ZN(n14076) );
  AND2_X1 U8995 ( .A1(n14085), .A2(n14084), .ZN(n14308) );
  NAND2_X1 U8996 ( .A1(n6748), .A2(n6749), .ZN(n14080) );
  OR2_X1 U8997 ( .A1(n14087), .A2(n14086), .ZN(n14307) );
  NAND2_X1 U8998 ( .A1(n7799), .A2(n7798), .ZN(n14314) );
  NAND2_X1 U8999 ( .A1(n7799), .A2(n10380), .ZN(n14100) );
  NAND2_X1 U9000 ( .A1(n7767), .A2(n7770), .ZN(n14132) );
  INV_X1 U9001 ( .A(n7768), .ZN(n14149) );
  AOI21_X1 U9002 ( .B1(n7136), .B2(n7769), .A(n7774), .ZN(n7768) );
  INV_X1 U9003 ( .A(n7775), .ZN(n7769) );
  NAND2_X1 U9004 ( .A1(n7760), .A2(n7761), .ZN(n14174) );
  NAND2_X1 U9005 ( .A1(n7138), .A2(n7764), .ZN(n7760) );
  NAND2_X1 U9006 ( .A1(n7777), .A2(n7780), .ZN(n14231) );
  NAND2_X1 U9007 ( .A1(n8964), .A2(n8963), .ZN(n14245) );
  NAND2_X1 U9008 ( .A1(n7074), .A2(n7075), .ZN(n12644) );
  NAND2_X1 U9009 ( .A1(n7082), .A2(n7083), .ZN(n12581) );
  OAI21_X1 U9010 ( .B1(n12434), .B2(n6424), .A(n10366), .ZN(n12580) );
  NAND2_X1 U9011 ( .A1(n11769), .A2(n10361), .ZN(n12145) );
  NAND2_X1 U9012 ( .A1(n11620), .A2(n10390), .ZN(n11084) );
  INV_X1 U9013 ( .A(n14273), .ZN(n14266) );
  AND2_X1 U9014 ( .A1(n14242), .A2(n11613), .ZN(n14278) );
  AND2_X1 U9015 ( .A1(n14242), .A2(n11587), .ZN(n14273) );
  INV_X1 U9016 ( .A(n11662), .ZN(n11410) );
  INV_X1 U9017 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7441) );
  NAND2_X1 U9018 ( .A1(n9211), .A2(n9210), .ZN(n14387) );
  AND2_X2 U9019 ( .A1(n10981), .A2(n10445), .ZN(n15502) );
  INV_X1 U9020 ( .A(n15502), .ZN(n15500) );
  OR2_X1 U9021 ( .A1(n15494), .A2(n14389), .ZN(n6830) );
  NAND2_X1 U9022 ( .A1(n14039), .A2(n14035), .ZN(n14388) );
  AND2_X1 U9023 ( .A1(n14294), .A2(n14293), .ZN(n7068) );
  NAND2_X1 U9024 ( .A1(n6642), .A2(n14308), .ZN(n14401) );
  INV_X1 U9025 ( .A(n6643), .ZN(n6642) );
  OAI21_X1 U9026 ( .B1(n14309), .B2(n14386), .A(n14307), .ZN(n6643) );
  INV_X1 U9027 ( .A(n14138), .ZN(n14411) );
  INV_X1 U9028 ( .A(n12589), .ZN(n13870) );
  OR2_X1 U9029 ( .A1(n6408), .A2(n15322), .ZN(n8645) );
  INV_X1 U9030 ( .A(n15459), .ZN(n15460) );
  INV_X1 U9031 ( .A(n15463), .ZN(n15466) );
  AND2_X1 U9032 ( .A1(n7782), .A2(n8607), .ZN(n7079) );
  INV_X1 U9033 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8607) );
  INV_X1 U9034 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12383) );
  NAND2_X1 U9035 ( .A1(n9318), .A2(n9319), .ZN(n12382) );
  OAI21_X1 U9036 ( .B1(n9324), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9325) );
  INV_X1 U9037 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11663) );
  CLKBUF_X1 U9038 ( .A(n8615), .Z(n11587) );
  INV_X1 U9039 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11093) );
  INV_X1 U9040 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10994) );
  INV_X1 U9041 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11078) );
  INV_X1 U9042 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n15714) );
  INV_X1 U9043 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10791) );
  INV_X1 U9044 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10688) );
  INV_X1 U9045 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10679) );
  INV_X1 U9046 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10657) );
  AND2_X1 U9047 ( .A1(n8796), .A2(n8832), .ZN(n13975) );
  INV_X1 U9048 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10592) );
  AOI21_X1 U9049 ( .B1(n7734), .B2(n7736), .A(n6516), .ZN(n7732) );
  NAND2_X1 U9050 ( .A1(n12268), .A2(n12267), .ZN(n12529) );
  NAND2_X1 U9051 ( .A1(n7050), .A2(n11175), .ZN(n15242) );
  XNOR2_X1 U9052 ( .A(n12828), .B(n12829), .ZN(n14479) );
  AND2_X1 U9053 ( .A1(n7726), .A2(n6475), .ZN(n14480) );
  NAND2_X1 U9054 ( .A1(n7725), .A2(n7726), .ZN(n14478) );
  AND2_X1 U9055 ( .A1(n12885), .A2(n7127), .ZN(n7126) );
  NOR2_X1 U9056 ( .A1(n7128), .A2(n15237), .ZN(n7127) );
  INV_X1 U9057 ( .A(n12884), .ZN(n7128) );
  NAND2_X1 U9058 ( .A1(n11825), .A2(n11824), .ZN(n11828) );
  NAND2_X1 U9059 ( .A1(n7056), .A2(n7058), .ZN(n14535) );
  NAND2_X1 U9060 ( .A1(n7059), .A2(n7717), .ZN(n7056) );
  AND2_X1 U9061 ( .A1(n11990), .A2(n11984), .ZN(n7744) );
  AND2_X1 U9062 ( .A1(n11985), .A2(n11984), .ZN(n11991) );
  AOI21_X1 U9063 ( .B1(n7722), .B2(n7724), .A(n7720), .ZN(n7719) );
  INV_X1 U9064 ( .A(n14544), .ZN(n7720) );
  NAND2_X1 U9065 ( .A1(n7722), .A2(n7718), .ZN(n14545) );
  OR2_X1 U9066 ( .A1(n14573), .A2(n7724), .ZN(n7718) );
  INV_X1 U9067 ( .A(n7717), .ZN(n14566) );
  INV_X1 U9068 ( .A(n14732), .ZN(n14708) );
  INV_X1 U9069 ( .A(n14797), .ZN(n14826) );
  NAND2_X1 U9070 ( .A1(n9883), .A2(n9882), .ZN(n14608) );
  OAI21_X1 U9071 ( .B1(n14842), .B2(n10026), .A(n9869), .ZN(n14825) );
  NAND2_X1 U9072 ( .A1(n9548), .A2(n9547), .ZN(n14889) );
  NAND2_X1 U9073 ( .A1(n9827), .A2(n9826), .ZN(n14887) );
  OR2_X1 U9074 ( .A1(n11207), .A2(n10546), .ZN(n14611) );
  OR3_X1 U9075 ( .A1(n9757), .A2(n9756), .A3(n9755), .ZN(n14613) );
  NAND2_X1 U9076 ( .A1(n14649), .A2(n6811), .ZN(n10776) );
  AND2_X1 U9077 ( .A1(n6808), .A2(n6800), .ZN(n10723) );
  NAND2_X1 U9078 ( .A1(n6806), .A2(n6808), .ZN(n10725) );
  INV_X1 U9079 ( .A(n6807), .ZN(n6806) );
  NAND2_X1 U9080 ( .A1(n10706), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7287) );
  AND2_X1 U9081 ( .A1(n10738), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7294) );
  NOR2_X1 U9082 ( .A1(n10737), .A2(n10736), .ZN(n10837) );
  NOR2_X1 U9083 ( .A1(n10837), .A2(n7293), .ZN(n10839) );
  AND2_X1 U9084 ( .A1(n10838), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7293) );
  NAND2_X1 U9085 ( .A1(n10839), .A2(n10840), .ZN(n10999) );
  NAND2_X1 U9086 ( .A1(n11386), .A2(n7283), .ZN(n11389) );
  AND2_X1 U9087 ( .A1(n7282), .A2(n7281), .ZN(n11971) );
  AND2_X1 U9088 ( .A1(n12388), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7286) );
  NAND2_X1 U9089 ( .A1(n12389), .A2(n12390), .ZN(n12656) );
  OAI22_X1 U9090 ( .A1(n15262), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n15264), 
        .B2(n12660), .ZN(n12661) );
  INV_X1 U9091 ( .A(n12659), .ZN(n12660) );
  OR2_X1 U9092 ( .A1(n15258), .A2(n10928), .ZN(n14686) );
  XNOR2_X1 U9093 ( .A(n14683), .B(n14682), .ZN(n14681) );
  XNOR2_X1 U9094 ( .A(n6790), .B(n14699), .ZN(n14693) );
  INV_X1 U9095 ( .A(n6790), .ZN(n14701) );
  NAND2_X1 U9096 ( .A1(n7318), .A2(n7316), .ZN(n12734) );
  INV_X1 U9097 ( .A(n7319), .ZN(n7316) );
  NAND2_X1 U9098 ( .A1(n7851), .A2(n7850), .ZN(n14759) );
  AND2_X1 U9099 ( .A1(n7851), .A2(n6462), .ZN(n14761) );
  NAND2_X1 U9100 ( .A1(n7298), .A2(n7299), .ZN(n14774) );
  NAND2_X1 U9101 ( .A1(n14822), .A2(n7840), .ZN(n14808) );
  NAND2_X1 U9102 ( .A1(n14852), .A2(n12694), .ZN(n14838) );
  NAND2_X1 U9103 ( .A1(n14852), .A2(n7844), .ZN(n15040) );
  CLKBUF_X1 U9104 ( .A(n14861), .Z(n6628) );
  NAND2_X1 U9105 ( .A1(n7813), .A2(n12718), .ZN(n14867) );
  OR2_X1 U9106 ( .A1(n14883), .A2(n12719), .ZN(n7813) );
  NAND2_X1 U9107 ( .A1(n9810), .A2(n9809), .ZN(n14898) );
  OAI21_X1 U9108 ( .B1(n6644), .B2(n7808), .A(n7805), .ZN(n12709) );
  NAND2_X1 U9109 ( .A1(n12455), .A2(n12457), .ZN(n12502) );
  NAND2_X1 U9110 ( .A1(n6644), .A2(n12453), .ZN(n12455) );
  OAI21_X1 U9111 ( .B1(n12090), .B2(n7812), .A(n7810), .ZN(n12177) );
  NAND2_X1 U9112 ( .A1(n12089), .A2(n11872), .ZN(n11873) );
  NAND2_X1 U9113 ( .A1(n11884), .A2(n11883), .ZN(n12094) );
  NAND2_X1 U9114 ( .A1(n11958), .A2(n11957), .ZN(n11956) );
  NAND2_X1 U9115 ( .A1(n11937), .A2(n11591), .ZN(n11958) );
  OR2_X1 U9116 ( .A1(n11750), .A2(n11739), .ZN(n11741) );
  AND2_X1 U9117 ( .A1(n14940), .A2(n11747), .ZN(n14956) );
  INV_X1 U9118 ( .A(n14754), .ZN(n14864) );
  INV_X1 U9119 ( .A(n15316), .ZN(n15314) );
  NAND2_X1 U9120 ( .A1(n7548), .A2(n7547), .ZN(n14987) );
  NOR3_X1 U9121 ( .A1(n14976), .A2(n14983), .A3(n14982), .ZN(n14989) );
  AOI21_X1 U9122 ( .B1(n14998), .B2(n15282), .A(n6875), .ZN(n6874) );
  NAND2_X1 U9123 ( .A1(n14999), .A2(n6597), .ZN(n6875) );
  AND2_X2 U9124 ( .A1(n10959), .A2(n11748), .ZN(n15310) );
  NAND2_X1 U9125 ( .A1(n11740), .A2(n10963), .ZN(n15596) );
  INV_X1 U9126 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n15135) );
  AND2_X1 U9127 ( .A1(n9523), .A2(n7852), .ZN(n7137) );
  AND2_X1 U9128 ( .A1(n9526), .A2(n9540), .ZN(n7852) );
  NAND2_X1 U9129 ( .A1(n9207), .A2(n8559), .ZN(n15143) );
  NAND2_X1 U9130 ( .A1(n6856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6855) );
  INV_X1 U9131 ( .A(n10583), .ZN(n12740) );
  INV_X1 U9132 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12386) );
  NAND2_X1 U9133 ( .A1(n6660), .A2(n10572), .ZN(n9898) );
  INV_X1 U9134 ( .A(n10011), .ZN(n12939) );
  INV_X1 U9135 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12933) );
  INV_X1 U9136 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11442) );
  INV_X1 U9137 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n15692) );
  INV_X1 U9138 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11061) );
  INV_X1 U9139 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10998) );
  INV_X1 U9140 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10788) );
  INV_X1 U9141 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10795) );
  INV_X1 U9142 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10731) );
  INV_X1 U9143 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10690) );
  INV_X1 U9144 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10681) );
  INV_X1 U9145 ( .A(n11002), .ZN(n11070) );
  INV_X1 U9146 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10672) );
  INV_X1 U9147 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10676) );
  INV_X1 U9148 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10568) );
  NAND2_X1 U9149 ( .A1(n9598), .A2(n7295), .ZN(n10766) );
  AOI21_X1 U9150 ( .B1(n9597), .B2(n6506), .A(n7296), .ZN(n7295) );
  NOR2_X1 U9151 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n7296) );
  NAND2_X1 U9152 ( .A1(n9597), .A2(n6812), .ZN(n10700) );
  INV_X1 U9153 ( .A(n6813), .ZN(n6812) );
  OAI21_X1 U9154 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_1__SCAN_IN), .A(
        n6814), .ZN(n6813) );
  NAND2_X1 U9155 ( .A1(n7369), .A2(n7368), .ZN(n10624) );
  XNOR2_X1 U9156 ( .A(n11146), .B(n11137), .ZN(n15157) );
  XNOR2_X1 U9157 ( .A(n11448), .B(n11446), .ZN(n11445) );
  NAND2_X1 U9158 ( .A1(n7356), .A2(n7354), .ZN(n11575) );
  AND2_X1 U9159 ( .A1(n11449), .A2(n7355), .ZN(n7354) );
  INV_X1 U9160 ( .A(n11455), .ZN(n7355) );
  INV_X1 U9161 ( .A(n12411), .ZN(n7372) );
  AOI21_X1 U9162 ( .B1(n7379), .B2(n7381), .A(n7378), .ZN(n7377) );
  INV_X1 U9163 ( .A(n7382), .ZN(n7379) );
  INV_X1 U9164 ( .A(n15191), .ZN(n6697) );
  INV_X1 U9165 ( .A(n7689), .ZN(n12124) );
  OAI211_X1 U9166 ( .C1(n11302), .C2(n6458), .A(n6894), .B(n6887), .ZN(n11481)
         );
  AOI21_X1 U9167 ( .B1(n6639), .B2(n13311), .A(n6638), .ZN(n13282) );
  OR2_X1 U9168 ( .A1(n13281), .A2(n13280), .ZN(n6638) );
  AND2_X1 U9169 ( .A1(n13331), .A2(n13332), .ZN(n6704) );
  OAI211_X1 U9170 ( .C1(n13319), .C2(n6883), .A(n6882), .B(n13322), .ZN(n7142)
         );
  AOI21_X1 U9171 ( .B1(n10350), .B2(n15595), .A(n6605), .ZN(n7853) );
  NAND2_X1 U9172 ( .A1(n15583), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U9173 ( .A1(n13610), .A2(n15585), .ZN(n6729) );
  INV_X1 U9174 ( .A(n13611), .ZN(n6730) );
  AND2_X1 U9175 ( .A1(n13716), .A2(n13717), .ZN(n6670) );
  NOR2_X1 U9176 ( .A1(n6678), .A2(n14033), .ZN(n6677) );
  NAND2_X1 U9177 ( .A1(n7442), .A2(n7439), .ZN(P2_U3530) );
  AOI21_X1 U9178 ( .B1(n14387), .B2(n14374), .A(n7440), .ZN(n7439) );
  NAND2_X1 U9179 ( .A1(n14388), .A2(n15502), .ZN(n7442) );
  NOR2_X1 U9180 ( .A1(n15502), .A2(n7441), .ZN(n7440) );
  NAND2_X1 U9181 ( .A1(n6831), .A2(n6828), .ZN(P2_U3498) );
  INV_X1 U9182 ( .A(n6829), .ZN(n6828) );
  NAND2_X1 U9183 ( .A1(n14388), .A2(n15494), .ZN(n6831) );
  OAI21_X1 U9184 ( .B1(n14390), .B2(n14428), .A(n6830), .ZN(n6829) );
  AND2_X1 U9185 ( .A1(n7729), .A2(n7730), .ZN(n11533) );
  OAI21_X1 U9186 ( .B1(n7130), .B2(n15237), .A(n14509), .ZN(P1_U3225) );
  XNOR2_X1 U9187 ( .A(n14504), .B(n7131), .ZN(n7130) );
  XNOR2_X1 U9188 ( .A(n7180), .B(n7179), .ZN(n14588) );
  AOI21_X1 U9189 ( .B1(n7273), .B2(n7274), .A(n7272), .ZN(n7271) );
  OAI21_X1 U9190 ( .B1(n15271), .B2(n7969), .A(n14691), .ZN(n7272) );
  NAND2_X1 U9191 ( .A1(n6823), .A2(n11127), .ZN(n11128) );
  INV_X1 U9192 ( .A(n6824), .ZN(n6823) );
  NAND2_X1 U9193 ( .A1(n15170), .A2(n15169), .ZN(n15172) );
  NAND2_X1 U9194 ( .A1(n7383), .A2(n7380), .ZN(n15173) );
  INV_X1 U9195 ( .A(n6821), .ZN(n15205) );
  AND2_X1 U9196 ( .A1(n7362), .A2(n15218), .ZN(n15227) );
  OAI21_X1 U9197 ( .B1(n6886), .B2(n6453), .A(n6885), .ZN(n6884) );
  AND2_X1 U9198 ( .A1(n7419), .A2(n8143), .ZN(n6414) );
  NOR2_X1 U9199 ( .A1(n12971), .A2(n7709), .ZN(n6415) );
  AND2_X2 U9200 ( .A1(n9566), .A2(n10019), .ZN(n9837) );
  AND2_X1 U9201 ( .A1(n7223), .A2(n6507), .ZN(n6416) );
  AND2_X1 U9202 ( .A1(n12839), .A2(n12840), .ZN(n6417) );
  AND2_X1 U9203 ( .A1(n7311), .A2(n8526), .ZN(n6418) );
  INV_X1 U9204 ( .A(n7254), .ZN(n14070) );
  NAND2_X1 U9205 ( .A1(n9060), .A2(n9059), .ZN(n7254) );
  OR2_X2 U9206 ( .A1(n13287), .A2(n13286), .ZN(n6419) );
  INV_X1 U9207 ( .A(n8530), .ZN(n7694) );
  INV_X1 U9208 ( .A(n10319), .ZN(n6725) );
  INV_X1 U9209 ( .A(n12699), .ZN(n7849) );
  INV_X1 U9210 ( .A(n10429), .ZN(n7791) );
  AND2_X1 U9211 ( .A1(n12179), .A2(n6794), .ZN(n6420) );
  AND3_X2 U9212 ( .A1(n9337), .A2(n14031), .A3(n11896), .ZN(n6421) );
  OR2_X1 U9213 ( .A1(n7208), .A2(n8934), .ZN(n6422) );
  AND2_X1 U9214 ( .A1(n14903), .A2(n7543), .ZN(n6423) );
  NOR2_X1 U9215 ( .A1(n13793), .A2(n13941), .ZN(n6424) );
  NAND2_X1 U9216 ( .A1(n12504), .A2(n12503), .ZN(n6425) );
  OR2_X1 U9217 ( .A1(n8070), .A2(n10666), .ZN(n6426) );
  NAND2_X1 U9218 ( .A1(n14870), .A2(n12692), .ZN(n6427) );
  NOR2_X1 U9219 ( .A1(n7254), .A2(n14083), .ZN(n6428) );
  INV_X1 U9220 ( .A(n14699), .ZN(n6978) );
  NAND2_X1 U9221 ( .A1(n9930), .A2(n9929), .ZN(n14781) );
  NAND2_X1 U9222 ( .A1(n7704), .A2(n6490), .ZN(n6429) );
  AND2_X1 U9223 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_REG3_REG_6__SCAN_IN), 
        .ZN(n6430) );
  AND2_X1 U9224 ( .A1(n6521), .A2(n7196), .ZN(n6431) );
  INV_X1 U9225 ( .A(n12756), .ZN(n15030) );
  NAND2_X1 U9226 ( .A1(n15150), .A2(n10660), .ZN(n12756) );
  NOR2_X1 U9227 ( .A1(n9680), .A2(n9683), .ZN(n6432) );
  INV_X1 U9228 ( .A(n14077), .ZN(n6750) );
  AND3_X1 U9229 ( .A1(n7546), .A2(n7550), .A3(n14949), .ZN(n6433) );
  INV_X1 U9230 ( .A(n6460), .ZN(n7208) );
  AND3_X1 U9231 ( .A1(n7908), .A2(n7910), .A3(n7906), .ZN(n6434) );
  OR2_X1 U9232 ( .A1(n6419), .A2(n6624), .ZN(n6435) );
  INV_X1 U9233 ( .A(n9270), .ZN(n7699) );
  NAND2_X1 U9234 ( .A1(n9230), .A2(n9229), .ZN(n12678) );
  AND2_X1 U9235 ( .A1(n6839), .A2(n6838), .ZN(n6436) );
  AND2_X1 U9236 ( .A1(n7075), .A2(n6590), .ZN(n6437) );
  AND4_X1 U9237 ( .A1(n8123), .A2(n8122), .A3(n8121), .A4(n8120), .ZN(n13033)
         );
  INV_X1 U9238 ( .A(n13033), .ZN(n13122) );
  AND2_X1 U9239 ( .A1(n10485), .A2(n13510), .ZN(n6438) );
  INV_X1 U9240 ( .A(n14127), .ZN(n6738) );
  NAND2_X1 U9241 ( .A1(n9873), .A2(n9872), .ZN(n7599) );
  INV_X1 U9242 ( .A(n7599), .ZN(n7596) );
  AND2_X1 U9243 ( .A1(n6841), .A2(n6842), .ZN(n6439) );
  AND2_X1 U9244 ( .A1(n7405), .A2(n7401), .ZN(n6440) );
  AND2_X1 U9245 ( .A1(n7700), .A2(n9263), .ZN(n6441) );
  NAND3_X1 U9246 ( .A1(n7290), .A2(P1_REG1_REG_18__SCAN_IN), .A3(n7291), .ZN(
        n6442) );
  AND2_X1 U9247 ( .A1(n7064), .A2(n14366), .ZN(n6443) );
  NAND2_X1 U9248 ( .A1(n12765), .A2(n12764), .ZN(n6444) );
  OR2_X1 U9249 ( .A1(n7790), .A2(n6750), .ZN(n6445) );
  NAND2_X1 U9250 ( .A1(n12689), .A2(n12688), .ZN(n6446) );
  AND2_X1 U9251 ( .A1(n7551), .A2(n10038), .ZN(n6447) );
  INV_X1 U9252 ( .A(n10311), .ZN(n13520) );
  AND2_X1 U9253 ( .A1(n7747), .A2(n7051), .ZN(n6448) );
  AND2_X1 U9254 ( .A1(n9205), .A2(n9204), .ZN(n6449) );
  NAND2_X1 U9255 ( .A1(n11792), .A2(n7643), .ZN(n7640) );
  INV_X1 U9256 ( .A(n15169), .ZN(n7383) );
  INV_X1 U9257 ( .A(n11836), .ZN(n7645) );
  AND2_X1 U9258 ( .A1(n7872), .A2(n7042), .ZN(n6450) );
  AND2_X1 U9259 ( .A1(n6845), .A2(n6603), .ZN(n6451) );
  AND2_X1 U9260 ( .A1(n6720), .A2(n8082), .ZN(n6452) );
  OR2_X1 U9261 ( .A1(n13324), .A2(n7122), .ZN(n6453) );
  INV_X1 U9262 ( .A(n13793), .ZN(n7444) );
  AND2_X1 U9263 ( .A1(n6884), .A2(n6617), .ZN(n6454) );
  NAND2_X1 U9264 ( .A1(n6453), .A2(n13326), .ZN(n6455) );
  BUF_X1 U9265 ( .A(n6421), .Z(n9269) );
  INV_X1 U9266 ( .A(n11427), .ZN(n6897) );
  AND2_X1 U9267 ( .A1(n10338), .A2(n11704), .ZN(n6456) );
  INV_X1 U9268 ( .A(n10174), .ZN(n7637) );
  OR2_X1 U9269 ( .A1(n11249), .A2(n11263), .ZN(n6457) );
  OR2_X1 U9270 ( .A1(n6896), .A2(n11427), .ZN(n6458) );
  NAND2_X1 U9271 ( .A1(n8236), .A2(n8235), .ZN(n13580) );
  AND2_X1 U9272 ( .A1(n9374), .A2(n9373), .ZN(n6459) );
  OR2_X1 U9273 ( .A1(n7576), .A2(n8913), .ZN(n6460) );
  AND2_X1 U9274 ( .A1(n13979), .A2(n11045), .ZN(n6461) );
  NAND2_X1 U9275 ( .A1(n6908), .A2(n7826), .ZN(n12505) );
  AND2_X1 U9276 ( .A1(n10037), .A2(n10036), .ZN(n10038) );
  INV_X1 U9277 ( .A(n11281), .ZN(n7495) );
  NAND2_X1 U9278 ( .A1(n14527), .A2(n12816), .ZN(n14573) );
  INV_X1 U9279 ( .A(n10038), .ZN(n14986) );
  INV_X1 U9280 ( .A(n14209), .ZN(n14352) );
  NAND2_X1 U9281 ( .A1(n8182), .A2(n8181), .ZN(n13680) );
  OR2_X1 U9282 ( .A1(n14781), .A2(n14798), .ZN(n6462) );
  AND2_X1 U9283 ( .A1(n7037), .A2(n7036), .ZN(n6463) );
  NOR2_X1 U9284 ( .A1(n9782), .A2(n9781), .ZN(n6464) );
  AND2_X1 U9285 ( .A1(n7288), .A2(n7287), .ZN(n6465) );
  AND2_X1 U9286 ( .A1(n7403), .A2(n7408), .ZN(n6466) );
  AND2_X1 U9287 ( .A1(n7395), .A2(n11266), .ZN(n6467) );
  NAND2_X1 U9288 ( .A1(n12730), .A2(n7819), .ZN(n6468) );
  NOR2_X1 U9289 ( .A1(n13747), .A2(n7003), .ZN(n6469) );
  INV_X1 U9290 ( .A(n12159), .ZN(n10439) );
  INV_X1 U9291 ( .A(n7793), .ZN(n7799) );
  INV_X1 U9292 ( .A(n13507), .ZN(n7624) );
  INV_X1 U9293 ( .A(n11263), .ZN(n7505) );
  OR2_X1 U9294 ( .A1(n10255), .A2(n10665), .ZN(n6470) );
  NOR2_X1 U9295 ( .A1(n12846), .A2(n12845), .ZN(n6471) );
  AND4_X1 U9296 ( .A1(n8852), .A2(n6740), .A3(n8496), .A4(n8851), .ZN(n6472)
         );
  AND2_X1 U9297 ( .A1(n9550), .A2(n9549), .ZN(n6473) );
  OR2_X1 U9298 ( .A1(n10029), .A2(n15247), .ZN(n6474) );
  NAND2_X1 U9299 ( .A1(n12822), .A2(n12823), .ZN(n6475) );
  NAND2_X1 U9300 ( .A1(n14179), .A2(n14200), .ZN(n6476) );
  XNOR2_X1 U9301 ( .A(n14986), .B(n10079), .ZN(n14983) );
  AND2_X1 U9302 ( .A1(n14760), .A2(n14793), .ZN(n6477) );
  OR2_X1 U9303 ( .A1(n13552), .A2(n13379), .ZN(n6478) );
  OR2_X1 U9304 ( .A1(n14179), .A2(n14200), .ZN(n6479) );
  NAND2_X1 U9306 ( .A1(n7010), .A2(n7009), .ZN(n9178) );
  NOR2_X1 U9307 ( .A1(n15092), .A2(n14963), .ZN(n6480) );
  NAND2_X1 U9308 ( .A1(n10425), .A2(n10424), .ZN(n14145) );
  INV_X1 U9309 ( .A(n7803), .ZN(n7802) );
  NAND2_X1 U9310 ( .A1(n9282), .A2(n10409), .ZN(n7803) );
  AND2_X1 U9311 ( .A1(n6418), .A2(n7310), .ZN(n6481) );
  INV_X1 U9312 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U9313 ( .A1(n10244), .A2(n13347), .ZN(n10319) );
  NAND2_X1 U9314 ( .A1(n10001), .A2(n10000), .ZN(n14699) );
  INV_X1 U9315 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9560) );
  AND2_X1 U9316 ( .A1(n14387), .A2(n13928), .ZN(n6482) );
  NAND2_X1 U9317 ( .A1(n15025), .A2(n14607), .ZN(n6483) );
  INV_X1 U9318 ( .A(n10320), .ZN(n7174) );
  OR2_X1 U9319 ( .A1(n13003), .A2(n13498), .ZN(n6484) );
  AND2_X1 U9320 ( .A1(n12988), .A2(n10479), .ZN(n6485) );
  NOR4_X1 U9321 ( .A1(n10318), .A2(n13386), .A3(n10317), .A4(n10316), .ZN(
        n6486) );
  INV_X1 U9322 ( .A(n9650), .ZN(n6767) );
  INV_X1 U9323 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9526) );
  OR2_X1 U9324 ( .A1(n8965), .A2(n11407), .ZN(n6487) );
  NAND2_X1 U9325 ( .A1(n12540), .A2(n12212), .ZN(n6488) );
  OR2_X1 U9326 ( .A1(n10456), .A2(n6959), .ZN(n6489) );
  INV_X1 U9327 ( .A(n10217), .ZN(n7615) );
  OR2_X1 U9328 ( .A1(n12977), .A2(n13073), .ZN(n6490) );
  AND2_X1 U9329 ( .A1(n8415), .A2(n13347), .ZN(n6491) );
  OR2_X1 U9330 ( .A1(n11915), .A2(n11914), .ZN(n6492) );
  INV_X1 U9331 ( .A(n9900), .ZN(n6772) );
  INV_X1 U9332 ( .A(n15180), .ZN(n7378) );
  INV_X1 U9333 ( .A(n15043), .ZN(n14846) );
  INV_X1 U9334 ( .A(n7139), .ZN(n12676) );
  INV_X1 U9335 ( .A(n7696), .ZN(n7695) );
  NAND2_X1 U9336 ( .A1(n7254), .A2(n14083), .ZN(n6493) );
  NOR2_X1 U9337 ( .A1(n14148), .A2(n7774), .ZN(n6494) );
  NOR2_X1 U9338 ( .A1(n10222), .A2(n10207), .ZN(n6495) );
  INV_X1 U9339 ( .A(n13510), .ZN(n13538) );
  AND4_X1 U9340 ( .A1(n8202), .A2(n8201), .A3(n8200), .A4(n8199), .ZN(n13510)
         );
  INV_X1 U9341 ( .A(n9551), .ZN(n9525) );
  AND2_X1 U9342 ( .A1(n14245), .A2(n10417), .ZN(n6496) );
  INV_X1 U9343 ( .A(n9700), .ZN(n6780) );
  AND2_X1 U9344 ( .A1(n14151), .A2(n13876), .ZN(n6497) );
  INV_X1 U9345 ( .A(n7226), .ZN(n7225) );
  INV_X1 U9346 ( .A(n9916), .ZN(n6769) );
  OR2_X1 U9347 ( .A1(n8865), .A2(n6536), .ZN(n6498) );
  AND2_X1 U9348 ( .A1(n12676), .A2(n12681), .ZN(n6499) );
  AND2_X1 U9349 ( .A1(n7792), .A2(n10428), .ZN(n6500) );
  INV_X1 U9350 ( .A(n7284), .ZN(n7283) );
  AND2_X1 U9351 ( .A1(n7819), .A2(n7818), .ZN(n6501) );
  AND2_X1 U9352 ( .A1(n7664), .A2(n13018), .ZN(n6502) );
  NAND2_X1 U9353 ( .A1(n9216), .A2(n9215), .ZN(n14292) );
  AND2_X1 U9354 ( .A1(n6822), .A2(n7366), .ZN(n6503) );
  AND2_X1 U9355 ( .A1(n13845), .A2(n7519), .ZN(n6504) );
  NAND2_X1 U9356 ( .A1(n9344), .A2(n11407), .ZN(n6505) );
  AND2_X1 U9357 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6506) );
  INV_X1 U9358 ( .A(n9977), .ZN(n7603) );
  NAND2_X1 U9359 ( .A1(n13585), .A2(n13498), .ZN(n6507) );
  NAND2_X1 U9360 ( .A1(n9166), .A2(n9165), .ZN(n6508) );
  INV_X1 U9361 ( .A(n7428), .ZN(n14066) );
  NOR2_X1 U9362 ( .A1(n14119), .A2(n7429), .ZN(n7428) );
  OR2_X1 U9363 ( .A1(n7561), .A2(n7559), .ZN(n6509) );
  AND2_X1 U9364 ( .A1(n11885), .A2(n11883), .ZN(n6510) );
  INV_X1 U9365 ( .A(n7210), .ZN(n7209) );
  NAND2_X1 U9366 ( .A1(n7211), .A2(n8934), .ZN(n7210) );
  NAND2_X1 U9367 ( .A1(n7870), .A2(n7033), .ZN(n6511) );
  AND2_X1 U9368 ( .A1(n14083), .A2(n9244), .ZN(n6512) );
  AND2_X1 U9369 ( .A1(n8464), .A2(SI_1_), .ZN(n6513) );
  OR2_X1 U9370 ( .A1(n12564), .A2(n7347), .ZN(n6514) );
  AND2_X1 U9371 ( .A1(n13630), .A2(n13120), .ZN(n6515) );
  AND2_X1 U9372 ( .A1(n12870), .A2(n12869), .ZN(n6516) );
  OR2_X1 U9373 ( .A1(n14775), .A2(n12699), .ZN(n7851) );
  AND2_X1 U9374 ( .A1(n8629), .A2(n8628), .ZN(n6517) );
  INV_X1 U9375 ( .A(n7644), .ZN(n7643) );
  OAI21_X1 U9376 ( .B1(n10466), .B2(n7646), .A(n7645), .ZN(n7644) );
  INV_X1 U9377 ( .A(n7401), .ZN(n7400) );
  NAND2_X1 U9378 ( .A1(n7402), .A2(n7408), .ZN(n7401) );
  NAND2_X1 U9379 ( .A1(n6776), .A2(n6777), .ZN(n6518) );
  AND2_X1 U9380 ( .A1(n13669), .A2(n13538), .ZN(n6519) );
  AND2_X1 U9381 ( .A1(n7710), .A2(n6415), .ZN(n6520) );
  NAND2_X1 U9382 ( .A1(n13169), .A2(n13170), .ZN(n7408) );
  OR2_X1 U9383 ( .A1(n8827), .A2(n8829), .ZN(n6521) );
  NOR2_X1 U9384 ( .A1(n9976), .A2(n7603), .ZN(n6522) );
  NOR2_X1 U9385 ( .A1(n12183), .A2(n14616), .ZN(n6523) );
  NOR2_X1 U9386 ( .A1(n13615), .A2(n13118), .ZN(n6524) );
  NOR2_X1 U9387 ( .A1(n12589), .A2(n13940), .ZN(n6525) );
  NOR2_X1 U9388 ( .A1(n13585), .A2(n13498), .ZN(n6526) );
  NOR2_X1 U9389 ( .A1(n15043), .A2(n14490), .ZN(n6527) );
  NOR2_X1 U9390 ( .A1(n11418), .A2(n6897), .ZN(n6528) );
  AND2_X1 U9391 ( .A1(n9160), .A2(n7256), .ZN(n6529) );
  AND2_X1 U9392 ( .A1(n8485), .A2(SI_7_), .ZN(n6530) );
  AND2_X1 U9393 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n6531) );
  NOR2_X1 U9394 ( .A1(n8912), .A2(n8914), .ZN(n7577) );
  INV_X1 U9395 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10569) );
  INV_X1 U9396 ( .A(n10381), .ZN(n7800) );
  OR2_X1 U9397 ( .A1(n7788), .A2(n7104), .ZN(n6532) );
  AND2_X1 U9398 ( .A1(n12992), .A2(n13378), .ZN(n6533) );
  NOR2_X1 U9399 ( .A1(n12830), .A2(n12829), .ZN(n6534) );
  NOR2_X1 U9400 ( .A1(n14737), .A2(n14603), .ZN(n6535) );
  AND2_X1 U9401 ( .A1(n8863), .A2(n8862), .ZN(n6536) );
  AND2_X1 U9402 ( .A1(n10480), .A2(n10479), .ZN(n6537) );
  AND2_X1 U9403 ( .A1(n8959), .A2(n8958), .ZN(n6538) );
  INV_X1 U9404 ( .A(n12287), .ZN(n7828) );
  AND2_X1 U9405 ( .A1(n7254), .A2(n13800), .ZN(n6539) );
  MUX2_X1 U9406 ( .A(n14608), .B(n15036), .S(n10045), .Z(n9886) );
  OR3_X1 U9407 ( .A1(n7582), .A2(n9751), .A3(n6464), .ZN(n6540) );
  INV_X1 U9408 ( .A(n8491), .ZN(n7305) );
  AND2_X1 U9409 ( .A1(n13651), .A2(n13085), .ZN(n10215) );
  INV_X1 U9410 ( .A(n6675), .ZN(n7528) );
  NAND2_X1 U9411 ( .A1(n9422), .A2(n9421), .ZN(n6675) );
  INV_X1 U9412 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10571) );
  INV_X1 U9413 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10595) );
  OR2_X1 U9414 ( .A1(n14621), .A2(n6406), .ZN(n6541) );
  NAND2_X1 U9415 ( .A1(n12807), .A2(n14523), .ZN(n6542) );
  NAND2_X1 U9416 ( .A1(n9424), .A2(n9423), .ZN(n6543) );
  NOR2_X1 U9417 ( .A1(n13135), .A2(n13140), .ZN(n6544) );
  INV_X1 U9418 ( .A(n7260), .ZN(n7259) );
  NAND2_X1 U9419 ( .A1(n7264), .A2(n7261), .ZN(n7260) );
  AND2_X1 U9420 ( .A1(n7603), .A2(n9976), .ZN(n6545) );
  OR2_X1 U9421 ( .A1(n7617), .A2(n7613), .ZN(n6546) );
  INV_X1 U9422 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10793) );
  OR2_X1 U9423 ( .A1(n9349), .A2(n11407), .ZN(n6547) );
  OR2_X1 U9424 ( .A1(n14829), .A2(n15030), .ZN(n6548) );
  INV_X1 U9425 ( .A(n10382), .ZN(n7797) );
  OR2_X1 U9426 ( .A1(n13680), .A2(n13121), .ZN(n10189) );
  AND2_X1 U9427 ( .A1(n7290), .A2(n7291), .ZN(n6549) );
  AND2_X1 U9428 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n15321), .ZN(n6550) );
  NOR2_X1 U9429 ( .A1(n7569), .A2(n8828), .ZN(n6551) );
  OAI21_X1 U9430 ( .B1(n11355), .B2(n11377), .A(n11354), .ZN(n11182) );
  AND2_X1 U9431 ( .A1(n14927), .A2(n12710), .ZN(n6552) );
  AND2_X1 U9432 ( .A1(n11327), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6553) );
  OAI21_X1 U9433 ( .B1(n13535), .B2(n7629), .A(n10311), .ZN(n7628) );
  INV_X1 U9434 ( .A(n9036), .ZN(n7567) );
  INV_X1 U9435 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7178) );
  INV_X1 U9436 ( .A(n6752), .ZN(n6751) );
  NAND2_X1 U9437 ( .A1(n7789), .A2(n6753), .ZN(n6752) );
  NAND2_X1 U9438 ( .A1(n7861), .A2(n9262), .ZN(n6554) );
  NAND2_X1 U9439 ( .A1(n9265), .A2(n9264), .ZN(n7700) );
  INV_X1 U9440 ( .A(n9964), .ZN(n6787) );
  NAND2_X1 U9441 ( .A1(n9538), .A2(n6847), .ZN(n6555) );
  AND2_X1 U9442 ( .A1(n10617), .A2(n7370), .ZN(n6556) );
  OR2_X1 U9443 ( .A1(n12832), .A2(n12833), .ZN(n6557) );
  AND2_X1 U9444 ( .A1(n7551), .A2(n14906), .ZN(n6558) );
  OR2_X1 U9445 ( .A1(n14336), .A2(n13933), .ZN(n6559) );
  NAND2_X1 U9446 ( .A1(n9943), .A2(n9942), .ZN(n15012) );
  INV_X1 U9447 ( .A(n10630), .ZN(n7182) );
  NAND2_X1 U9448 ( .A1(n9576), .A2(n6774), .ZN(n12007) );
  INV_X1 U9449 ( .A(n12007), .ZN(n11218) );
  AND2_X1 U9450 ( .A1(n12835), .A2(n12836), .ZN(n6560) );
  OR2_X1 U9451 ( .A1(n9293), .A2(n7067), .ZN(n6561) );
  OR2_X1 U9452 ( .A1(n9293), .A2(n7106), .ZN(n6562) );
  NOR2_X1 U9453 ( .A1(n9292), .A2(n6562), .ZN(n6563) );
  NOR2_X1 U9454 ( .A1(n10280), .A2(n10320), .ZN(n6564) );
  NOR2_X1 U9455 ( .A1(n7096), .A2(n7095), .ZN(n6565) );
  OR2_X1 U9456 ( .A1(n10185), .A2(n11095), .ZN(n6566) );
  INV_X1 U9457 ( .A(n7365), .ZN(n7368) );
  AND2_X1 U9458 ( .A1(n13416), .A2(n10211), .ZN(n6567) );
  NOR2_X1 U9459 ( .A1(n10054), .A2(n10043), .ZN(n6568) );
  AND2_X1 U9460 ( .A1(n15003), .A2(n6798), .ZN(n6569) );
  AND2_X1 U9461 ( .A1(n10188), .A2(n10195), .ZN(n10311) );
  NOR2_X1 U9462 ( .A1(n7595), .A2(n7593), .ZN(n6570) );
  AND2_X1 U9463 ( .A1(n13202), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n6571) );
  OR2_X1 U9464 ( .A1(n14980), .A2(n14981), .ZN(n6572) );
  INV_X1 U9465 ( .A(n14063), .ZN(n7790) );
  AND2_X1 U9466 ( .A1(n10153), .A2(n10466), .ZN(n6573) );
  AND2_X1 U9467 ( .A1(n13376), .A2(n10239), .ZN(n6574) );
  OR2_X1 U9468 ( .A1(n10289), .A2(n10288), .ZN(n6575) );
  NAND2_X1 U9469 ( .A1(n13615), .A2(n13118), .ZN(n6576) );
  AND2_X1 U9470 ( .A1(n11826), .A2(n11824), .ZN(n6577) );
  AND2_X1 U9471 ( .A1(n8938), .A2(n8507), .ZN(n6578) );
  OR2_X1 U9472 ( .A1(n9665), .A2(n9663), .ZN(n6579) );
  AND2_X1 U9473 ( .A1(n7660), .A2(n7659), .ZN(n6580) );
  NOR2_X1 U9474 ( .A1(n9873), .A2(n9872), .ZN(n7600) );
  AND2_X1 U9475 ( .A1(n7188), .A2(n7187), .ZN(n6581) );
  AND2_X1 U9476 ( .A1(n7188), .A2(n7699), .ZN(n6582) );
  AND2_X1 U9477 ( .A1(n14822), .A2(n12695), .ZN(n6583) );
  INV_X1 U9478 ( .A(n7060), .ZN(n7059) );
  OR2_X1 U9479 ( .A1(n14472), .A2(n7061), .ZN(n7060) );
  OR2_X1 U9480 ( .A1(n6767), .A2(n9649), .ZN(n6584) );
  AND2_X1 U9481 ( .A1(n6483), .A2(n12699), .ZN(n6585) );
  OR2_X1 U9482 ( .A1(n9664), .A2(n7602), .ZN(n6586) );
  INV_X1 U9483 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7212) );
  AND2_X1 U9484 ( .A1(n6552), .A2(n6864), .ZN(n6587) );
  INV_X1 U9485 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8578) );
  INV_X1 U9486 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9519) );
  INV_X1 U9487 ( .A(n8414), .ZN(n7656) );
  INV_X1 U9488 ( .A(n7703), .ZN(n7702) );
  OAI21_X1 U9489 ( .B1(n7705), .B2(n6429), .A(n10478), .ZN(n7703) );
  INV_X1 U9490 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7370) );
  INV_X1 U9491 ( .A(n7908), .ZN(n7453) );
  NAND2_X1 U9492 ( .A1(n7178), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7908) );
  OR2_X1 U9493 ( .A1(n7698), .A2(n7697), .ZN(n6588) );
  NAND2_X1 U9494 ( .A1(n9160), .A2(n9159), .ZN(n6589) );
  INV_X1 U9495 ( .A(SI_12_), .ZN(n10684) );
  INV_X1 U9496 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10566) );
  INV_X1 U9497 ( .A(n7841), .ZN(n7840) );
  NAND2_X1 U9498 ( .A1(n14809), .A2(n12695), .ZN(n7841) );
  OR2_X1 U9499 ( .A1(n14377), .A2(n13939), .ZN(n6590) );
  INV_X1 U9500 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10744) );
  INV_X1 U9501 ( .A(n6948), .ZN(n6947) );
  NAND2_X1 U9502 ( .A1(n13482), .A2(n6949), .ZN(n6948) );
  INV_X2 U9503 ( .A(n15583), .ZN(n15585) );
  INV_X1 U9504 ( .A(n14151), .ZN(n7435) );
  AND2_X1 U9505 ( .A1(n12351), .A2(n7691), .ZN(n7689) );
  NAND2_X1 U9506 ( .A1(n7829), .A2(n12186), .ZN(n12285) );
  AND2_X1 U9507 ( .A1(n6995), .A2(n8552), .ZN(n6591) );
  INV_X1 U9508 ( .A(n14245), .ZN(n6838) );
  NAND2_X1 U9509 ( .A1(n13029), .A2(n13030), .ZN(n10549) );
  NAND2_X1 U9510 ( .A1(n8582), .A2(n8581), .ZN(n14286) );
  INV_X1 U9511 ( .A(n14286), .ZN(n6841) );
  INV_X1 U9512 ( .A(n15237), .ZN(n14589) );
  NAND2_X1 U9513 ( .A1(n12112), .A2(n6794), .ZN(n6795) );
  AOI21_X1 U9514 ( .B1(n7266), .B2(n6867), .A(n6480), .ZN(n6866) );
  INV_X1 U9515 ( .A(n8085), .ZN(n8364) );
  NAND2_X1 U9516 ( .A1(n8029), .A2(n8028), .ZN(n11705) );
  AND2_X1 U9517 ( .A1(n7948), .A2(n7450), .ZN(n6592) );
  NAND2_X1 U9518 ( .A1(n8209), .A2(n8208), .ZN(n6593) );
  NAND2_X1 U9519 ( .A1(n9993), .A2(n9992), .ZN(n14991) );
  INV_X1 U9520 ( .A(n14991), .ZN(n6792) );
  AND2_X1 U9521 ( .A1(n7869), .A2(n7035), .ZN(n6594) );
  INV_X1 U9522 ( .A(n14312), .ZN(n7432) );
  INV_X1 U9523 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7714) );
  INV_X1 U9524 ( .A(n10196), .ZN(n7621) );
  AND2_X1 U9525 ( .A1(n6591), .A2(n9209), .ZN(n6595) );
  INV_X1 U9526 ( .A(n15025), .ZN(n7554) );
  AND2_X1 U9527 ( .A1(n11680), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U9528 ( .A1(n12420), .A2(n7802), .ZN(n12435) );
  OR2_X1 U9529 ( .A1(n15000), .A2(n15065), .ZN(n6597) );
  NAND2_X1 U9530 ( .A1(n6436), .A2(n12637), .ZN(n6840) );
  INV_X1 U9531 ( .A(n6628), .ZN(n7542) );
  AND2_X1 U9532 ( .A1(n8458), .A2(n8457), .ZN(n6598) );
  AND2_X1 U9533 ( .A1(n13180), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6599) );
  AND2_X1 U9534 ( .A1(n8549), .A2(n8543), .ZN(n6600) );
  OR2_X1 U9535 ( .A1(n14404), .A2(n14428), .ZN(n6601) );
  AND2_X1 U9536 ( .A1(n7690), .A2(n10463), .ZN(n6602) );
  AND2_X1 U9537 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6603) );
  INV_X1 U9538 ( .A(n8106), .ZN(n10270) );
  INV_X1 U9539 ( .A(n8060), .ZN(n8106) );
  OR2_X1 U9540 ( .A1(n13143), .A2(n13142), .ZN(n6604) );
  INV_X1 U9541 ( .A(n8082), .ZN(n6722) );
  NOR2_X1 U9542 ( .A1(n15595), .A2(n10351), .ZN(n6605) );
  OR2_X1 U9543 ( .A1(n8542), .A2(SI_27_), .ZN(n6606) );
  AND2_X1 U9544 ( .A1(n10275), .A2(n10274), .ZN(n13335) );
  AND2_X1 U9545 ( .A1(n11586), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n6607) );
  AND2_X1 U9546 ( .A1(n11684), .A2(n11675), .ZN(n6608) );
  NAND2_X1 U9547 ( .A1(n8404), .A2(n8403), .ZN(n6609) );
  OR2_X1 U9548 ( .A1(n13622), .A2(n13597), .ZN(n6610) );
  AND2_X1 U9549 ( .A1(n6843), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6611) );
  AND2_X1 U9550 ( .A1(n13226), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n6612) );
  INV_X1 U9551 ( .A(n9075), .ZN(n7017) );
  AND2_X1 U9552 ( .A1(n7746), .A2(n6444), .ZN(n6613) );
  AND2_X1 U9553 ( .A1(n8541), .A2(n7016), .ZN(n7015) );
  INV_X1 U9554 ( .A(n13246), .ZN(n7411) );
  INV_X1 U9555 ( .A(n12045), .ZN(n6760) );
  INV_X2 U9556 ( .A(n8470), .ZN(n10567) );
  INV_X1 U9557 ( .A(n11310), .ZN(n7394) );
  INV_X1 U9558 ( .A(n14382), .ZN(n7443) );
  OR2_X1 U9559 ( .A1(n6833), .A2(n6832), .ZN(n6614) );
  INV_X1 U9560 ( .A(n11844), .ZN(n6837) );
  NAND2_X1 U9561 ( .A1(n11193), .A2(n11192), .ZN(n11525) );
  INV_X1 U9562 ( .A(n12532), .ZN(n6793) );
  INV_X1 U9564 ( .A(n13418), .ZN(n13440) );
  AND2_X1 U9565 ( .A1(n8303), .A2(n8302), .ZN(n13418) );
  AND2_X1 U9566 ( .A1(n11864), .A2(n15484), .ZN(n14386) );
  INV_X1 U9567 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6848) );
  OR2_X1 U9568 ( .A1(n14669), .A2(n14892), .ZN(n6615) );
  AND2_X1 U9569 ( .A1(n12895), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U9570 ( .A1(n6886), .A2(n13318), .ZN(n6617) );
  NAND2_X1 U9571 ( .A1(n11932), .A2(n9307), .ZN(n6618) );
  INV_X1 U9572 ( .A(n13286), .ZN(n7504) );
  AND2_X1 U9573 ( .A1(n12738), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6619) );
  AND2_X1 U9574 ( .A1(n8941), .A2(n8983), .ZN(n13993) );
  INV_X1 U9575 ( .A(n13993), .ZN(n7246) );
  OR2_X1 U9576 ( .A1(n11746), .A2(n10923), .ZN(n14906) );
  INV_X1 U9577 ( .A(n14906), .ZN(n14949) );
  INV_X1 U9578 ( .A(n13431), .ZN(n13120) );
  AND2_X1 U9579 ( .A1(n8318), .A2(n8317), .ZN(n13431) );
  AND2_X1 U9580 ( .A1(n6844), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6620) );
  OR2_X1 U9581 ( .A1(n13275), .A2(n13274), .ZN(n6621) );
  NOR2_X1 U9582 ( .A1(n7960), .A2(n7488), .ZN(n7487) );
  INV_X1 U9583 ( .A(n7483), .ZN(n7482) );
  NAND2_X1 U9584 ( .A1(n10253), .A2(n7484), .ZN(n7483) );
  AND2_X1 U9585 ( .A1(n10567), .A2(P3_U3151), .ZN(n6622) );
  INV_X1 U9586 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8608) );
  XNOR2_X1 U9587 ( .A(n8686), .B(n8685), .ZN(n10564) );
  OR2_X1 U9588 ( .A1(n14647), .A2(n14646), .ZN(n6623) );
  INV_X1 U9589 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7357) );
  XOR2_X1 U9590 ( .A(n13321), .B(P3_REG2_REG_19__SCAN_IN), .Z(n6624) );
  NAND2_X1 U9591 ( .A1(n8577), .A2(n7079), .ZN(n14439) );
  AND2_X1 U9592 ( .A1(n7504), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U9593 ( .A1(n10777), .A2(n10778), .ZN(n7288) );
  INV_X1 U9594 ( .A(n13326), .ZN(n6886) );
  AND2_X1 U9595 ( .A1(n6624), .A2(n13308), .ZN(n6626) );
  INV_X1 U9596 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n7509) );
  INV_X1 U9597 ( .A(n11284), .ZN(n7123) );
  INV_X1 U9598 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n6655) );
  INV_X1 U9599 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6820) );
  INV_X1 U9600 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n7122) );
  NAND2_X1 U9601 ( .A1(n14065), .A2(n14082), .ZN(n7169) );
  AND2_X1 U9602 ( .A1(n13888), .A2(n14082), .ZN(n13909) );
  AOI22_X1 U9603 ( .A1(n13753), .A2(n9131), .B1(n13943), .B2(n9194), .ZN(n8847) );
  NAND2_X1 U9604 ( .A1(n7307), .A2(n8658), .ZN(n8469) );
  NAND2_X1 U9605 ( .A1(n6659), .A2(n8465), .ZN(n7307) );
  NAND2_X1 U9606 ( .A1(n6974), .A2(n8483), .ZN(n8771) );
  NAND2_X1 U9607 ( .A1(n7731), .A2(n7732), .ZN(n14455) );
  NAND2_X1 U9608 ( .A1(n7719), .A2(n7721), .ZN(n14543) );
  NAND2_X1 U9609 ( .A1(n7510), .A2(n12067), .ZN(n7508) );
  NAND2_X1 U9610 ( .A1(n13230), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n13250) );
  NAND2_X1 U9611 ( .A1(n6627), .A2(n13161), .ZN(n7133) );
  INV_X1 U9612 ( .A(n7512), .ZN(n6627) );
  NAND2_X1 U9613 ( .A1(n7513), .A2(n13170), .ZN(n7512) );
  NAND2_X1 U9614 ( .A1(n13288), .A2(n6640), .ZN(n6639) );
  NAND2_X1 U9615 ( .A1(n13182), .A2(n13181), .ZN(n13184) );
  NAND2_X1 U9616 ( .A1(n7133), .A2(n7511), .ZN(n13182) );
  NAND2_X1 U9617 ( .A1(n13250), .A2(n7493), .ZN(n13251) );
  INV_X1 U9618 ( .A(n11491), .ZN(n7516) );
  INV_X1 U9619 ( .A(n11923), .ZN(n7510) );
  NAND2_X1 U9620 ( .A1(n14543), .A2(n6557), .ZN(n14486) );
  NAND2_X1 U9621 ( .A1(n6681), .A2(n6680), .ZN(n7496) );
  NAND2_X1 U9622 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7517) );
  AOI21_X1 U9623 ( .B1(n14743), .B2(n12702), .A(n12701), .ZN(n14726) );
  NAND2_X1 U9624 ( .A1(n9024), .A2(n9023), .ZN(n9028) );
  NAND3_X1 U9626 ( .A1(n6721), .A2(n6719), .A3(n6720), .ZN(n6718) );
  NAND2_X1 U9627 ( .A1(n13451), .A2(n13450), .ZN(n13449) );
  NAND2_X1 U9628 ( .A1(n7098), .A2(n7097), .ZN(n14049) );
  NAND2_X1 U9629 ( .A1(n6698), .A2(n6697), .ZN(n15194) );
  OAI21_X1 U9630 ( .B1(n12024), .B2(n12025), .A(n12026), .ZN(n12407) );
  AOI21_X2 U9631 ( .B1(n13993), .B2(n13992), .A(n13991), .ZN(n13995) );
  NAND2_X1 U9632 ( .A1(n13961), .A2(n10899), .ZN(n10900) );
  NAND2_X1 U9633 ( .A1(n14028), .A2(n15402), .ZN(n6690) );
  NAND2_X1 U9634 ( .A1(n13973), .A2(n13974), .ZN(n15378) );
  NAND2_X1 U9635 ( .A1(n6690), .A2(n6689), .ZN(n6688) );
  NAND2_X1 U9636 ( .A1(n6687), .A2(n6686), .ZN(n15389) );
  NOR2_X1 U9637 ( .A1(n7238), .A2(n14017), .ZN(n7237) );
  AOI21_X1 U9638 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n14011), .A(n14010), .ZN(
        n15446) );
  INV_X1 U9639 ( .A(n15192), .ZN(n6698) );
  NAND2_X1 U9640 ( .A1(n7369), .A2(n6503), .ZN(n10626) );
  NAND2_X1 U9641 ( .A1(n8309), .A2(n7954), .ZN(n7955) );
  NAND2_X1 U9642 ( .A1(n7228), .A2(n6576), .ZN(n7226) );
  INV_X1 U9643 ( .A(n7476), .ZN(n7475) );
  NOR2_X1 U9644 ( .A1(n10367), .A2(n7077), .ZN(n7076) );
  NAND2_X1 U9645 ( .A1(n8320), .A2(n12140), .ZN(n7957) );
  OAI21_X1 U9646 ( .B1(n7146), .B2(n6935), .A(n6932), .ZN(n6938) );
  OAI21_X1 U9647 ( .B1(n8334), .B2(n6726), .A(n6724), .ZN(n7234) );
  OAI21_X1 U9648 ( .B1(n13353), .B2(n13352), .A(n13355), .ZN(n13610) );
  OAI21_X1 U9649 ( .B1(n14395), .B2(n15500), .A(n10446), .ZN(n10447) );
  NAND2_X1 U9650 ( .A1(n11593), .A2(n11602), .ZN(n11870) );
  NAND2_X1 U9651 ( .A1(n14403), .A2(n6601), .ZN(P2_U3492) );
  NAND2_X1 U9652 ( .A1(n14902), .A2(n12716), .ZN(n6858) );
  NAND2_X1 U9653 ( .A1(n14731), .A2(n14730), .ZN(n14998) );
  NAND2_X1 U9654 ( .A1(n6865), .A2(n6587), .ZN(n12715) );
  OR2_X1 U9655 ( .A1(n10169), .A2(n10168), .ZN(n10175) );
  NAND2_X1 U9656 ( .A1(n6645), .A2(n10289), .ZN(n7157) );
  NAND3_X1 U9657 ( .A1(n10249), .A2(n6646), .A3(n10248), .ZN(n6645) );
  NAND2_X1 U9658 ( .A1(n6647), .A2(n10246), .ZN(n6646) );
  INV_X1 U9659 ( .A(n10250), .ZN(n6647) );
  NAND2_X1 U9660 ( .A1(n7965), .A2(n7892), .ZN(n7967) );
  NOR2_X1 U9661 ( .A1(n7327), .A2(n7326), .ZN(n7325) );
  NAND2_X1 U9662 ( .A1(n6648), .A2(n10229), .ZN(n10235) );
  NAND3_X1 U9663 ( .A1(n7348), .A2(n6700), .A3(n6567), .ZN(n6648) );
  OR2_X1 U9664 ( .A1(n10183), .A2(n7344), .ZN(n7342) );
  NAND2_X1 U9665 ( .A1(n6922), .A2(n10324), .ZN(n6921) );
  NAND2_X1 U9666 ( .A1(n6920), .A2(n15507), .ZN(n6919) );
  NAND2_X1 U9667 ( .A1(n14025), .A2(n14007), .ZN(n14009) );
  NAND2_X1 U9668 ( .A1(n15427), .A2(n15426), .ZN(n15425) );
  NAND2_X1 U9669 ( .A1(n10867), .A2(n10866), .ZN(n13957) );
  INV_X1 U9670 ( .A(n15410), .ZN(n6652) );
  INV_X1 U9671 ( .A(n14009), .ZN(n6708) );
  NAND3_X1 U9672 ( .A1(n7503), .A2(n6419), .A3(n6626), .ZN(n7502) );
  XNOR2_X1 U9673 ( .A(n11239), .B(n6655), .ZN(n11109) );
  NOR2_X1 U9674 ( .A1(n13954), .A2(n11407), .ZN(n10985) );
  OAI21_X1 U9675 ( .B1(n9305), .B2(n11410), .A(n9299), .ZN(n9335) );
  NAND2_X1 U9676 ( .A1(n8642), .A2(n8463), .ZN(n6659) );
  INV_X1 U9677 ( .A(n7675), .ZN(n7674) );
  INV_X1 U9678 ( .A(n9897), .ZN(n6660) );
  INV_X1 U9679 ( .A(n13106), .ZN(n7676) );
  INV_X1 U9680 ( .A(n6957), .ZN(n6956) );
  NOR2_X1 U9681 ( .A1(n7716), .A2(n6417), .ZN(n7061) );
  NAND3_X1 U9682 ( .A1(n9335), .A2(n7556), .A3(n9334), .ZN(P2_U3328) );
  OAI21_X1 U9683 ( .B1(n9017), .B2(n9016), .A(n9015), .ZN(n9018) );
  OR2_X2 U9684 ( .A1(n8848), .A2(n6663), .ZN(n7574) );
  OAI21_X2 U9685 ( .B1(n7255), .B2(n6529), .A(n6441), .ZN(n7189) );
  OR2_X1 U9686 ( .A1(n9234), .A2(n11614), .ZN(n8655) );
  AOI21_X1 U9687 ( .B1(n9002), .B2(n9001), .A(n9000), .ZN(n9017) );
  OAI21_X1 U9688 ( .B1(n8699), .B2(n8698), .A(n8697), .ZN(n8705) );
  OAI21_X2 U9689 ( .B1(n6538), .B2(n8957), .A(n6664), .ZN(n8979) );
  OR2_X1 U9690 ( .A1(n8959), .A2(n8958), .ZN(n6664) );
  NAND2_X1 U9691 ( .A1(n8750), .A2(n8749), .ZN(n8769) );
  OAI22_X1 U9692 ( .A1(n7573), .A2(n7570), .B1(n8786), .B2(n8785), .ZN(n8807)
         );
  INV_X1 U9693 ( .A(n8767), .ZN(n6711) );
  OAI21_X1 U9694 ( .B1(n14823), .B2(n7841), .A(n7837), .ZN(n14794) );
  XNOR2_X2 U9695 ( .A(n8466), .B(SI_2_), .ZN(n8658) );
  NAND2_X2 U9696 ( .A1(n6665), .A2(n8460), .ZN(n8466) );
  OAI22_X1 U9697 ( .A1(n8722), .A2(n7192), .B1(n8723), .B2(n7193), .ZN(n8745)
         );
  OAI21_X2 U9698 ( .B1(n14775), .B2(n7848), .A(n7846), .ZN(n14743) );
  OAI21_X1 U9699 ( .B1(n14689), .B2(n14687), .A(n14686), .ZN(n6816) );
  OAI21_X1 U9700 ( .B1(n14688), .B2(n14677), .A(n6815), .ZN(n7273) );
  NAND2_X1 U9701 ( .A1(n6559), .A2(n10376), .ZN(n7775) );
  NAND2_X1 U9702 ( .A1(n15184), .A2(n15185), .ZN(n15192) );
  NAND2_X1 U9703 ( .A1(n14643), .A2(n14644), .ZN(n14642) );
  NAND2_X1 U9704 ( .A1(n7276), .A2(n7275), .ZN(n11972) );
  NOR2_X1 U9705 ( .A1(n10734), .A2(n7294), .ZN(n10737) );
  OAI21_X1 U9706 ( .B1(n14690), .B2(n7274), .A(n7271), .ZN(P1_U3262) );
  NOR2_X1 U9707 ( .A1(n12387), .A2(n7286), .ZN(n12389) );
  OAI21_X1 U9708 ( .B1(n14148), .B2(n7773), .A(n7772), .ZN(n7771) );
  XNOR2_X2 U9709 ( .A(n7330), .B(n10458), .ZN(n15511) );
  AOI21_X2 U9710 ( .B1(n12563), .B2(n10185), .A(n10190), .ZN(n13531) );
  INV_X1 U9711 ( .A(n7472), .ZN(n6935) );
  NAND2_X1 U9712 ( .A1(n7924), .A2(n7923), .ZN(n8131) );
  NAND2_X1 U9713 ( .A1(n7467), .A2(n7465), .ZN(n8192) );
  NAND2_X1 U9714 ( .A1(n7423), .A2(n7422), .ZN(n13402) );
  NAND2_X1 U9715 ( .A1(n7937), .A2(n7936), .ZN(n8204) );
  OAI21_X1 U9716 ( .B1(n13463), .B2(n7413), .A(n8259), .ZN(n13451) );
  NAND2_X1 U9717 ( .A1(n8066), .A2(n7916), .ZN(n7477) );
  INV_X1 U9718 ( .A(n6933), .ZN(n6932) );
  NOR2_X1 U9719 ( .A1(n13190), .A2(n13191), .ZN(n13211) );
  NOR2_X1 U9720 ( .A1(n13301), .A2(n13302), .ZN(n13323) );
  NAND2_X1 U9721 ( .A1(n13217), .A2(n13216), .ZN(n13234) );
  OAI22_X1 U9722 ( .A1(n11323), .A2(n11324), .B1(n11261), .B2(n11327), .ZN(
        n11265) );
  OAI21_X1 U9723 ( .B1(n13718), .B2(n13921), .A(n6670), .ZN(P2_U3186) );
  NAND2_X1 U9724 ( .A1(n7521), .A2(n7524), .ZN(n13777) );
  NAND2_X1 U9725 ( .A1(n14034), .A2(n6677), .ZN(P2_U3233) );
  NOR2_X1 U9726 ( .A1(n15457), .A2(n7970), .ZN(n6678) );
  INV_X1 U9727 ( .A(n15391), .ZN(n6687) );
  INV_X1 U9728 ( .A(n7239), .ZN(n7238) );
  INV_X1 U9729 ( .A(n11247), .ZN(n6681) );
  NAND4_X1 U9730 ( .A1(n6682), .A2(n13306), .A3(n13305), .A4(n13307), .ZN(
        P3_U3200) );
  NAND2_X1 U9731 ( .A1(n10355), .A2(n10356), .ZN(n11081) );
  INV_X1 U9732 ( .A(n6684), .ZN(n6683) );
  OR2_X1 U9733 ( .A1(n8895), .A2(n8894), .ZN(n7578) );
  NAND2_X2 U9734 ( .A1(n14055), .A2(n14054), .ZN(n14296) );
  OAI21_X1 U9735 ( .B1(n14395), .B2(n15492), .A(n14396), .ZN(n14397) );
  NAND2_X1 U9736 ( .A1(n6691), .A2(n6688), .ZN(n14034) );
  NAND2_X1 U9737 ( .A1(n14032), .A2(n14031), .ZN(n6691) );
  NAND2_X1 U9738 ( .A1(n15350), .A2(n15351), .ZN(n15349) );
  NAND2_X1 U9739 ( .A1(n14789), .A2(n14839), .ZN(n7819) );
  NAND2_X1 U9740 ( .A1(n15389), .A2(n11034), .ZN(n15404) );
  XNOR2_X1 U9741 ( .A(n13990), .B(n7246), .ZN(n12249) );
  NOR2_X1 U9742 ( .A1(n15434), .A2(n15433), .ZN(n15432) );
  NAND2_X1 U9743 ( .A1(n6694), .A2(n10622), .ZN(n10644) );
  NAND2_X1 U9744 ( .A1(n10621), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6694) );
  NAND2_X1 U9745 ( .A1(n15199), .A2(n15198), .ZN(n15204) );
  NAND2_X1 U9746 ( .A1(n12032), .A2(n12031), .ZN(n12404) );
  NAND2_X1 U9747 ( .A1(n11920), .A2(n7134), .ZN(n11923) );
  NAND2_X1 U9748 ( .A1(n13312), .A2(n13311), .ZN(n6705) );
  OAI21_X1 U9749 ( .B1(n9020), .B2(n9019), .A(n9018), .ZN(n9038) );
  NAND2_X1 U9750 ( .A1(n9321), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8580) );
  NOR2_X1 U9751 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  NAND2_X1 U9752 ( .A1(n7339), .A2(n7340), .ZN(n7155) );
  INV_X1 U9753 ( .A(n6950), .ZN(n10228) );
  AOI22_X1 U9754 ( .A1(n10140), .A2(n10139), .B1(n11095), .B2(n10138), .ZN(
        n10141) );
  NOR2_X1 U9755 ( .A1(n10194), .A2(n7621), .ZN(n10199) );
  INV_X1 U9756 ( .A(n10230), .ZN(n6700) );
  NOR3_X4 U9757 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .A3(
        P3_IR_REG_24__SCAN_IN), .ZN(n7890) );
  OAI21_X1 U9758 ( .B1(n10130), .B2(n10335), .A(n10455), .ZN(n10134) );
  AOI21_X1 U9759 ( .B1(n10212), .B2(n10214), .A(n7352), .ZN(n7351) );
  INV_X1 U9760 ( .A(n13271), .ZN(n6702) );
  NAND3_X1 U9761 ( .A1(n6705), .A2(n7142), .A3(n6704), .ZN(P3_U3201) );
  OAI21_X2 U9762 ( .B1(n14885), .B2(n6427), .A(n12693), .ZN(n7160) );
  NAND2_X1 U9763 ( .A1(n12698), .A2(n12697), .ZN(n14775) );
  NAND2_X1 U9764 ( .A1(n14742), .A2(n6874), .ZN(n15117) );
  AOI21_X2 U9765 ( .B1(n7121), .B2(n6493), .A(n6428), .ZN(n14055) );
  NAND2_X1 U9766 ( .A1(n8663), .A2(n8683), .ZN(n15341) );
  NAND2_X1 U9767 ( .A1(n13563), .A2(n6610), .ZN(P3_U3484) );
  AND3_X2 U9768 ( .A1(n7328), .A2(n8001), .A3(n8000), .ZN(n10458) );
  OAI21_X2 U9769 ( .B1(n13391), .B2(n15521), .A(n13390), .ZN(n13560) );
  NAND2_X1 U9770 ( .A1(n6709), .A2(n10125), .ZN(n11723) );
  NAND2_X1 U9771 ( .A1(n10306), .A2(n15504), .ZN(n6709) );
  AOI21_X2 U9772 ( .B1(n13493), .B2(n13482), .A(n10204), .ZN(n13478) );
  AND2_X1 U9773 ( .A1(n7342), .A2(n7343), .ZN(n10191) );
  NAND2_X1 U9774 ( .A1(n12306), .A2(n7338), .ZN(n7337) );
  AOI211_X2 U9775 ( .C1(n10175), .C2(n10174), .A(n10173), .B(n10172), .ZN(
        n10183) );
  NAND2_X1 U9776 ( .A1(n7157), .A2(n6564), .ZN(n6922) );
  AOI21_X1 U9777 ( .B1(n7332), .B2(n10164), .A(n10163), .ZN(n10169) );
  INV_X1 U9778 ( .A(n6939), .ZN(n10212) );
  NAND2_X1 U9779 ( .A1(n7335), .A2(n7334), .ZN(n7333) );
  OAI21_X1 U9780 ( .B1(n7351), .B2(n10215), .A(n7349), .ZN(n7348) );
  NOR2_X1 U9781 ( .A1(n11420), .A2(n7132), .ZN(n11422) );
  XNOR2_X2 U9782 ( .A(n8610), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8623) );
  OAI21_X1 U9783 ( .B1(n7185), .B2(n6589), .A(n6449), .ZN(n7255) );
  OAI21_X1 U9784 ( .B1(n8769), .B2(n8768), .A(n6710), .ZN(n7573) );
  NAND2_X1 U9785 ( .A1(n6712), .A2(n6711), .ZN(n6710) );
  NAND2_X1 U9786 ( .A1(n8769), .A2(n8768), .ZN(n6712) );
  OAI21_X2 U9787 ( .B1(n9321), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U9788 ( .A1(n11500), .A2(n11499), .ZN(n11501) );
  INV_X1 U9789 ( .A(n11770), .ZN(n7072) );
  INV_X4 U9790 ( .A(n8666), .ZN(n9228) );
  NAND2_X1 U9791 ( .A1(n7195), .A2(n7194), .ZN(n8850) );
  NAND2_X1 U9792 ( .A1(n9140), .A2(n9139), .ZN(n9143) );
  NAND2_X1 U9793 ( .A1(n8788), .A2(n8486), .ZN(n7129) );
  XNOR2_X2 U9794 ( .A(n14151), .B(n13932), .ZN(n14148) );
  NAND3_X1 U9795 ( .A1(n7658), .A2(n8093), .A3(n7891), .ZN(n6714) );
  NOR2_X2 U9796 ( .A1(n8205), .A2(n7327), .ZN(n7891) );
  NAND2_X1 U9797 ( .A1(n6717), .A2(n7414), .ZN(n12565) );
  NAND3_X1 U9798 ( .A1(n6718), .A2(n6414), .A3(n7218), .ZN(n6717) );
  NAND3_X1 U9799 ( .A1(n6730), .A2(n6729), .A3(n6728), .ZN(P3_U3455) );
  NAND2_X2 U9800 ( .A1(n8515), .A2(n8514), .ZN(n8981) );
  NAND2_X2 U9801 ( .A1(n8961), .A2(n8960), .ZN(n8515) );
  AND2_X2 U9802 ( .A1(n14209), .A2(n10421), .ZN(n10422) );
  NAND2_X2 U9803 ( .A1(n6731), .A2(n9007), .ZN(n14209) );
  XNOR2_X2 U9804 ( .A(n9022), .B(n9004), .ZN(n11441) );
  INV_X1 U9805 ( .A(n10425), .ZN(n6735) );
  INV_X1 U9806 ( .A(n8495), .ZN(n6742) );
  NAND2_X1 U9807 ( .A1(n10572), .A2(n10795), .ZN(n6739) );
  NAND2_X1 U9808 ( .A1(n6742), .A2(SI_11_), .ZN(n8852) );
  NAND3_X1 U9809 ( .A1(n7761), .A2(n7758), .A3(n6479), .ZN(n6743) );
  NAND2_X1 U9810 ( .A1(n14112), .A2(n6746), .ZN(n6744) );
  NAND2_X1 U9811 ( .A1(n6744), .A2(n6745), .ZN(n14064) );
  NAND2_X1 U9812 ( .A1(n7792), .A2(n7789), .ZN(n14095) );
  XNOR2_X2 U9813 ( .A(n6754), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9543) );
  NAND3_X1 U9814 ( .A1(n9525), .A2(n9524), .A3(n6756), .ZN(n6755) );
  INV_X1 U9815 ( .A(n6759), .ZN(n14948) );
  INV_X1 U9816 ( .A(n6757), .ZN(n14951) );
  INV_X1 U9817 ( .A(n15085), .ZN(n6758) );
  NAND3_X1 U9818 ( .A1(n9739), .A2(n9738), .A3(n7581), .ZN(n6764) );
  NAND3_X1 U9819 ( .A1(n9638), .A2(n6584), .A3(n9637), .ZN(n6765) );
  NAND3_X1 U9820 ( .A1(n6765), .A2(n6766), .A3(n6579), .ZN(n7601) );
  OAI21_X1 U9821 ( .B1(n9901), .B2(n6773), .A(n6771), .ZN(n9915) );
  NAND2_X1 U9822 ( .A1(n6770), .A2(n6768), .ZN(n9914) );
  NAND2_X1 U9823 ( .A1(n9901), .A2(n6771), .ZN(n6770) );
  NAND2_X1 U9824 ( .A1(n10589), .A2(n6777), .ZN(n6775) );
  NAND2_X2 U9825 ( .A1(n10660), .A2(n6776), .ZN(n9592) );
  NAND2_X1 U9826 ( .A1(n9681), .A2(n6781), .ZN(n6778) );
  OAI21_X1 U9827 ( .B1(n9681), .B2(n6432), .A(n6781), .ZN(n9699) );
  NAND2_X1 U9828 ( .A1(n6778), .A2(n6779), .ZN(n9698) );
  NAND2_X1 U9829 ( .A1(n9965), .A2(n6785), .ZN(n6784) );
  NOR3_X1 U9830 ( .A1(n6413), .A2(n14991), .A3(n14986), .ZN(n14712) );
  NOR2_X2 U9831 ( .A1(n6413), .A2(n14991), .ZN(n14692) );
  NOR2_X1 U9832 ( .A1(n6807), .A2(n10724), .ZN(n6800) );
  NAND3_X1 U9833 ( .A1(n6811), .A2(n6810), .A3(n6802), .ZN(n6801) );
  NAND3_X1 U9834 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U9835 ( .A1(n12023), .A2(n6817), .ZN(n12032) );
  NAND2_X1 U9836 ( .A1(n11576), .A2(n6819), .ZN(n6818) );
  NAND2_X1 U9837 ( .A1(n11576), .A2(n11575), .ZN(n12022) );
  NAND3_X1 U9838 ( .A1(n10629), .A2(n10628), .A3(P3_ADDR_REG_3__SCAN_IN), .ZN(
        n6822) );
  NAND2_X1 U9839 ( .A1(n10633), .A2(n10613), .ZN(n10629) );
  NAND2_X1 U9840 ( .A1(n7183), .A2(n7182), .ZN(n10633) );
  NAND2_X1 U9841 ( .A1(n6825), .A2(n7377), .ZN(n15183) );
  NAND3_X1 U9842 ( .A1(n6826), .A2(n7381), .A3(n15160), .ZN(n6825) );
  NAND2_X1 U9843 ( .A1(n12615), .A2(n12614), .ZN(n15159) );
  NAND3_X1 U9844 ( .A1(n7148), .A2(n10619), .A3(n7147), .ZN(n10622) );
  NAND2_X1 U9845 ( .A1(n7148), .A2(n10619), .ZN(n10621) );
  INV_X1 U9846 ( .A(n8579), .ZN(n8577) );
  NAND2_X1 U9847 ( .A1(n15488), .A2(n11632), .ZN(n6832) );
  INV_X1 U9848 ( .A(n6835), .ZN(n6833) );
  NAND3_X1 U9849 ( .A1(n15488), .A2(n11632), .A3(n11654), .ZN(n11852) );
  INV_X1 U9850 ( .A(n6840), .ZN(n14237) );
  NAND3_X1 U9851 ( .A1(n9536), .A2(n6430), .A3(P1_REG3_REG_7__SCAN_IN), .ZN(
        n9685) );
  NAND2_X1 U9852 ( .A1(n9537), .A2(n6611), .ZN(n9771) );
  NAND2_X1 U9853 ( .A1(n9888), .A2(n6620), .ZN(n9934) );
  NAND2_X1 U9854 ( .A1(n9888), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9903) );
  NAND4_X1 U9855 ( .A1(n6854), .A2(n6851), .A3(n6850), .A4(n14980), .ZN(n6849)
         );
  NOR2_X1 U9856 ( .A1(n14745), .A2(n10094), .ZN(n6850) );
  XNOR2_X2 U9857 ( .A(n6855), .B(n9526), .ZN(n15146) );
  NAND3_X1 U9858 ( .A1(n7750), .A2(n9524), .A3(n9523), .ZN(n6856) );
  NAND2_X1 U9859 ( .A1(n11939), .A2(n11938), .ZN(n11937) );
  XNOR2_X2 U9860 ( .A(n6862), .B(n11607), .ZN(n11957) );
  NAND2_X1 U9861 ( .A1(n12454), .A2(n6866), .ZN(n6865) );
  XNOR2_X1 U9862 ( .A(n14622), .B(n15234), .ZN(n11941) );
  INV_X1 U9863 ( .A(n10564), .ZN(n6871) );
  NAND2_X4 U9864 ( .A1(n9541), .A2(n9543), .ZN(n10026) );
  AOI21_X2 U9865 ( .B1(n14998), .B2(n14873), .A(n7267), .ZN(n14742) );
  NAND2_X1 U9866 ( .A1(n7270), .A2(n7297), .ZN(n14772) );
  NAND2_X1 U9867 ( .A1(n12725), .A2(n6876), .ZN(n7297) );
  OAI21_X1 U9868 ( .B1(n11325), .B2(n11326), .A(n6878), .ZN(n11336) );
  NAND2_X1 U9869 ( .A1(n11325), .A2(n11326), .ZN(n6878) );
  XNOR2_X2 U9870 ( .A(n6879), .B(P3_IR_REG_3__SCAN_IN), .ZN(n11281) );
  NAND2_X1 U9871 ( .A1(n11241), .A2(n11240), .ZN(n11242) );
  INV_X1 U9872 ( .A(n11302), .ZN(n6891) );
  NAND2_X1 U9873 ( .A1(n11302), .A2(n11303), .ZN(n11419) );
  NAND3_X1 U9874 ( .A1(n6890), .A2(P3_REG1_REG_7__SCAN_IN), .A3(n6888), .ZN(
        n11484) );
  NAND3_X1 U9875 ( .A1(n6894), .A2(n11302), .A3(n6889), .ZN(n6888) );
  NAND3_X1 U9876 ( .A1(n6891), .A2(n6894), .A3(n6458), .ZN(n6890) );
  NAND2_X1 U9877 ( .A1(n11419), .A2(n11418), .ZN(n11482) );
  NAND3_X1 U9878 ( .A1(n6899), .A2(n13231), .A3(n6898), .ZN(n13244) );
  NAND2_X1 U9879 ( .A1(n13202), .A2(n6612), .ZN(n6898) );
  NOR2_X1 U9880 ( .A1(n6571), .A2(n13201), .ZN(n13227) );
  OR2_X1 U9881 ( .A1(n10026), .A2(n11902), .ZN(n6901) );
  NAND2_X1 U9882 ( .A1(n10027), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6903) );
  NAND3_X1 U9883 ( .A1(n7137), .A2(n9525), .A3(n9524), .ZN(n15138) );
  NAND2_X1 U9884 ( .A1(n12188), .A2(n6907), .ZN(n6906) );
  NAND2_X1 U9885 ( .A1(n14959), .A2(n6911), .ZN(n6909) );
  NAND2_X1 U9886 ( .A1(n7160), .A2(n7844), .ZN(n6914) );
  INV_X1 U9887 ( .A(n7160), .ZN(n14854) );
  NAND3_X1 U9888 ( .A1(n6919), .A2(n6917), .A3(n6916), .ZN(n7143) );
  NAND2_X1 U9889 ( .A1(n6924), .A2(n7702), .ZN(n6923) );
  OR2_X1 U9890 ( .A1(n10475), .A2(n10474), .ZN(n6924) );
  OAI21_X1 U9891 ( .B1(n6935), .B2(n6936), .A(n8099), .ZN(n6933) );
  OAI21_X1 U9892 ( .B1(n10199), .B2(n6948), .A(n6940), .ZN(n6939) );
  NAND3_X1 U9893 ( .A1(n6954), .A2(n6953), .A3(n10489), .ZN(n13083) );
  NAND2_X1 U9894 ( .A1(n6956), .A2(n12945), .ZN(n6953) );
  INV_X1 U9895 ( .A(n6961), .ZN(n6959) );
  NAND2_X1 U9896 ( .A1(n10456), .A2(n15515), .ZN(n6960) );
  NAND2_X1 U9897 ( .A1(n11566), .A2(n6489), .ZN(n11559) );
  NAND4_X1 U9898 ( .A1(n7687), .A2(n7688), .A3(n7691), .A4(n12351), .ZN(n6966)
         );
  NAND2_X1 U9899 ( .A1(n11558), .A2(n6967), .ZN(n12351) );
  NAND2_X1 U9900 ( .A1(n7686), .A2(n6966), .ZN(n11758) );
  AND2_X2 U9901 ( .A1(n10187), .A2(n10189), .ZN(n13535) );
  OAI21_X2 U9902 ( .B1(n10451), .B2(n10610), .A(n10450), .ZN(n10459) );
  NAND3_X1 U9903 ( .A1(n7891), .A2(n8093), .A3(n7890), .ZN(n8431) );
  NAND2_X1 U9904 ( .A1(n6970), .A2(n8477), .ZN(n8480) );
  XNOR2_X1 U9905 ( .A(n6970), .B(n8725), .ZN(n10590) );
  INV_X1 U9906 ( .A(n8484), .ZN(n6973) );
  OAI21_X2 U9907 ( .B1(n6974), .B2(n6973), .A(n6971), .ZN(n8788) );
  NAND2_X1 U9908 ( .A1(n8752), .A2(n8481), .ZN(n6974) );
  NAND2_X2 U9909 ( .A1(n8594), .A2(n8593), .ZN(n11662) );
  NAND2_X1 U9910 ( .A1(n11518), .A2(n6984), .ZN(n6983) );
  OAI21_X1 U9911 ( .B1(n11518), .B2(n11517), .A(n9371), .ZN(n11795) );
  NAND2_X1 U9912 ( .A1(n8553), .A2(n6591), .ZN(n9207) );
  NAND2_X1 U9913 ( .A1(n8553), .A2(n8552), .ZN(n8558) );
  NAND2_X1 U9914 ( .A1(n13843), .A2(n7001), .ZN(n6996) );
  NAND2_X1 U9915 ( .A1(n6996), .A2(n6999), .ZN(n13719) );
  NAND2_X1 U9916 ( .A1(n13758), .A2(n7522), .ZN(n7521) );
  NAND2_X1 U9917 ( .A1(n9076), .A2(n7015), .ZN(n7008) );
  NAND2_X1 U9918 ( .A1(n7008), .A2(n7013), .ZN(n7116) );
  OAI21_X1 U9919 ( .B1(n9076), .B2(n9075), .A(n8541), .ZN(n9058) );
  INV_X1 U9920 ( .A(n9457), .ZN(n13906) );
  NAND2_X1 U9921 ( .A1(n8515), .A2(n7022), .ZN(n7021) );
  NAND3_X1 U9922 ( .A1(n7657), .A2(n6725), .A3(n7656), .ZN(n7037) );
  NAND2_X1 U9923 ( .A1(n7873), .A2(n7040), .ZN(n8213) );
  NAND2_X1 U9924 ( .A1(n7176), .A2(n7045), .ZN(n8238) );
  NAND2_X1 U9925 ( .A1(n7176), .A2(n15627), .ZN(n8251) );
  NAND3_X1 U9926 ( .A1(n7866), .A2(n7865), .A3(n12356), .ZN(n8043) );
  NAND4_X1 U9927 ( .A1(n12356), .A2(n7866), .A3(n7865), .A4(n7047), .ZN(n8058)
         );
  XNOR2_X1 U9928 ( .A(n11157), .B(n11159), .ZN(n11216) );
  XNOR2_X2 U9929 ( .A(n9520), .B(n9519), .ZN(n10115) );
  INV_X1 U9930 ( .A(n15239), .ZN(n7050) );
  NAND2_X1 U9931 ( .A1(n15239), .A2(n11183), .ZN(n7049) );
  OAI21_X1 U9932 ( .B1(n12262), .B2(n7053), .A(n6448), .ZN(n7746) );
  NAND2_X1 U9933 ( .A1(n11825), .A2(n6577), .ZN(n11985) );
  AOI21_X1 U9934 ( .B1(n7058), .B2(n7060), .A(n7057), .ZN(n7054) );
  NAND2_X1 U9935 ( .A1(n10387), .A2(n7066), .ZN(n7062) );
  NAND3_X1 U9936 ( .A1(n7063), .A2(n7062), .A3(n7064), .ZN(n14295) );
  NAND3_X1 U9937 ( .A1(n7063), .A2(n7062), .A3(n6443), .ZN(n7069) );
  OR2_X2 U9938 ( .A1(n10387), .A2(n6561), .ZN(n7063) );
  NAND2_X1 U9939 ( .A1(n7069), .A2(n7068), .ZN(n14394) );
  OAI211_X1 U9940 ( .C1(n7072), .C2(n7071), .A(n7118), .B(n7070), .ZN(n10364)
         );
  XNOR2_X1 U9941 ( .A(n13949), .B(n7073), .ZN(n11499) );
  NAND2_X1 U9942 ( .A1(n8676), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U9943 ( .A1(n10986), .A2(n10985), .ZN(n10984) );
  NAND3_X1 U9944 ( .A1(n7083), .A2(n7082), .A3(n7081), .ZN(n7085) );
  NAND2_X1 U9945 ( .A1(n11641), .A2(n7087), .ZN(n7086) );
  NAND2_X1 U9946 ( .A1(n7089), .A2(n7086), .ZN(n11858) );
  NAND2_X1 U9947 ( .A1(n10415), .A2(n6565), .ZN(n7092) );
  NAND2_X1 U9948 ( .A1(n7092), .A2(n7093), .ZN(n14215) );
  NAND2_X1 U9949 ( .A1(n10415), .A2(n10414), .ZN(n14250) );
  INV_X1 U9950 ( .A(n10414), .ZN(n7095) );
  INV_X1 U9951 ( .A(n7801), .ZN(n7096) );
  NAND2_X1 U9952 ( .A1(n14128), .A2(n7099), .ZN(n7098) );
  AOI21_X2 U9953 ( .B1(n14049), .B2(n14048), .A(n10432), .ZN(n10436) );
  NAND2_X1 U9954 ( .A1(n11640), .A2(n11639), .ZN(n11638) );
  NAND2_X1 U9955 ( .A1(n7120), .A2(n14186), .ZN(n14195) );
  NOR2_X1 U9956 ( .A1(n7117), .A2(n10354), .ZN(n10355) );
  NAND2_X1 U9957 ( .A1(n10364), .A2(n10363), .ZN(n12429) );
  INV_X1 U9958 ( .A(n13953), .ZN(n9274) );
  OR2_X1 U9959 ( .A1(n8673), .A2(n14281), .ZN(n8650) );
  NAND2_X1 U9960 ( .A1(n8944), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7105) );
  OR4_X2 U9961 ( .A1(n14127), .A2(n14186), .A3(n9286), .A4(n9285), .ZN(n9289)
         );
  NAND2_X1 U9962 ( .A1(n11772), .A2(n10398), .ZN(n7785) );
  NAND2_X1 U9963 ( .A1(n7109), .A2(n7108), .ZN(n9842) );
  NAND2_X1 U9964 ( .A1(n9806), .A2(n9805), .ZN(n7109) );
  INV_X4 U9965 ( .A(n9837), .ZN(n10045) );
  NAND2_X1 U9966 ( .A1(n9603), .A2(n7110), .ZN(n9604) );
  NAND2_X1 U9967 ( .A1(n9837), .A2(n11218), .ZN(n7110) );
  NAND3_X1 U9968 ( .A1(n7111), .A2(n10122), .A3(n10121), .ZN(P1_U3242) );
  NAND2_X1 U9969 ( .A1(n10044), .A2(n10053), .ZN(n7111) );
  NAND2_X1 U9970 ( .A1(n7113), .A2(n7112), .ZN(n14990) );
  NAND2_X1 U9971 ( .A1(n14976), .A2(n14975), .ZN(n7113) );
  NAND2_X2 U9972 ( .A1(n14910), .A2(n12691), .ZN(n14885) );
  NAND2_X1 U9973 ( .A1(n11964), .A2(n11598), .ZN(n12037) );
  NAND2_X1 U9974 ( .A1(n11595), .A2(n11594), .ZN(n11942) );
  INV_X1 U9975 ( .A(n7752), .ZN(n7751) );
  NAND2_X1 U9976 ( .A1(n7785), .A2(n7783), .ZN(n12148) );
  NAND2_X1 U9977 ( .A1(n7733), .A2(n12863), .ZN(n7180) );
  NOR2_X1 U9978 ( .A1(n14486), .A2(n14487), .ZN(n14485) );
  NAND2_X1 U9979 ( .A1(n14455), .A2(n12879), .ZN(n12890) );
  NAND2_X1 U9980 ( .A1(n12890), .A2(n7126), .ZN(n12889) );
  NAND2_X1 U9981 ( .A1(n7358), .A2(n11131), .ZN(n10649) );
  OAI21_X1 U9982 ( .B1(n8915), .B2(n8508), .A(n6578), .ZN(n8510) );
  NAND2_X1 U9983 ( .A1(n7300), .A2(n7301), .ZN(n8915) );
  XNOR2_X1 U9984 ( .A(n8475), .B(SI_4_), .ZN(n8713) );
  NAND2_X1 U9985 ( .A1(n9951), .A2(n9950), .ZN(n9965) );
  OAI21_X1 U9986 ( .B1(n9874), .B2(n6570), .A(n7591), .ZN(n9901) );
  INV_X1 U9987 ( .A(n7597), .ZN(n7592) );
  INV_X1 U9988 ( .A(n14072), .ZN(n7121) );
  NAND2_X1 U9989 ( .A1(n11638), .A2(n10358), .ZN(n11500) );
  NAND2_X1 U9990 ( .A1(n12404), .A2(n15607), .ZN(n7373) );
  NAND2_X1 U9991 ( .A1(n7360), .A2(n15215), .ZN(n15218) );
  NAND2_X1 U9992 ( .A1(n11456), .A2(n11455), .ZN(n11574) );
  NAND2_X1 U9993 ( .A1(n14172), .A2(n10375), .ZN(n10377) );
  NAND2_X1 U9994 ( .A1(n11849), .A2(n11848), .ZN(n11851) );
  NAND2_X1 U9995 ( .A1(n10373), .A2(n10372), .ZN(n7120) );
  XNOR2_X1 U9996 ( .A(n11129), .B(n11253), .ZN(n7359) );
  INV_X1 U9997 ( .A(n10751), .ZN(n10755) );
  NAND2_X1 U9998 ( .A1(n7750), .A2(n6473), .ZN(n9556) );
  AOI21_X1 U9999 ( .B1(n7683), .B2(n7685), .A(n7682), .ZN(n7681) );
  XNOR2_X1 U10000 ( .A(n8644), .B(n8643), .ZN(n9574) );
  NAND2_X2 U10001 ( .A1(n7129), .A2(n8488), .ZN(n8810) );
  XNOR2_X1 U10002 ( .A(n11181), .B(n12875), .ZN(n11377) );
  INV_X1 U10003 ( .A(n11182), .ZN(n11183) );
  NAND2_X1 U10004 ( .A1(n11985), .A2(n7744), .ZN(n12262) );
  NAND2_X1 U10005 ( .A1(n10101), .A2(n10100), .ZN(n10107) );
  NAND2_X1 U10006 ( .A1(n10107), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10102) );
  AND3_X2 U10007 ( .A1(n8646), .A2(n8647), .A3(n8645), .ZN(n12747) );
  INV_X1 U10008 ( .A(n9234), .ZN(n8944) );
  NAND2_X1 U10009 ( .A1(n7516), .A2(n12365), .ZN(n7515) );
  AND4_X2 U10010 ( .A1(n7324), .A2(n7323), .A3(n7325), .A4(n7658), .ZN(n7965)
         );
  AOI21_X2 U10011 ( .B1(n12467), .B2(n12468), .A(n8409), .ZN(n12563) );
  INV_X1 U10012 ( .A(n7610), .ZN(n13426) );
  NAND2_X1 U10013 ( .A1(n11643), .A2(n11642), .ZN(n11641) );
  NAND2_X1 U10014 ( .A1(n7622), .A2(n7620), .ZN(n13493) );
  NAND2_X1 U10015 ( .A1(n7632), .A2(n7630), .ZN(n12492) );
  OAI21_X1 U10016 ( .B1(n10437), .B2(n12913), .A(n10438), .ZN(n7139) );
  NAND2_X1 U10017 ( .A1(n13273), .A2(n6621), .ZN(n13276) );
  NOR2_X1 U10018 ( .A1(n13323), .A2(n7140), .ZN(n13328) );
  AND2_X1 U10019 ( .A1(n13325), .A2(n13324), .ZN(n7140) );
  NOR2_X1 U10020 ( .A1(n13211), .A2(n7412), .ZN(n13217) );
  AOI22_X1 U10021 ( .A1(n11287), .A2(n11286), .B1(n11102), .B2(n11101), .ZN(
        n11258) );
  INV_X1 U10022 ( .A(n14712), .ZN(n7546) );
  AND2_X1 U10023 ( .A1(n8626), .A2(n8625), .ZN(n8638) );
  INV_X8 U10024 ( .A(n7315), .ZN(n10572) );
  NAND2_X1 U10025 ( .A1(n7683), .A2(n7305), .ZN(n7304) );
  NAND2_X1 U10026 ( .A1(n11911), .A2(n11910), .ZN(n7141) );
  NAND2_X1 U10027 ( .A1(n14851), .A2(n12723), .ZN(n12725) );
  NAND2_X1 U10028 ( .A1(n7825), .A2(n12733), .ZN(n14729) );
  AND2_X1 U10029 ( .A1(n7156), .A2(n6725), .ZN(n10250) );
  NAND2_X1 U10030 ( .A1(n7143), .A2(n10329), .ZN(n10333) );
  NAND2_X1 U10031 ( .A1(n7333), .A2(n6573), .ZN(n7332) );
  OAI21_X1 U10032 ( .B1(n10141), .B2(n7337), .A(n7336), .ZN(n7335) );
  NAND2_X1 U10033 ( .A1(n7150), .A2(n7149), .ZN(n7148) );
  INV_X1 U10034 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7149) );
  INV_X1 U10035 ( .A(n10618), .ZN(n7150) );
  INV_X1 U10036 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U10037 ( .A1(n7359), .A2(n10620), .ZN(n11131) );
  OAI21_X1 U10038 ( .B1(n10240), .B2(n13386), .A(n6574), .ZN(n7156) );
  NAND2_X1 U10039 ( .A1(n7997), .A2(n7996), .ZN(n7995) );
  NAND2_X1 U10040 ( .A1(n12405), .A2(n7373), .ZN(n12412) );
  AND2_X1 U10041 ( .A1(n10187), .A2(n7343), .ZN(n7341) );
  NAND2_X1 U10042 ( .A1(n7346), .A2(n7345), .ZN(n7344) );
  NAND2_X1 U10043 ( .A1(n8146), .A2(n7928), .ZN(n7468) );
  NAND2_X1 U10044 ( .A1(n8469), .A2(n8468), .ZN(n8686) );
  NAND2_X1 U10045 ( .A1(n7252), .A2(n8473), .ZN(n8714) );
  AOI21_X1 U10046 ( .B1(n7341), .B2(n7344), .A(n13520), .ZN(n7339) );
  INV_X1 U10047 ( .A(n14574), .ZN(n7723) );
  NAND2_X1 U10048 ( .A1(n11940), .A2(n11597), .ZN(n11965) );
  NAND2_X1 U10049 ( .A1(n14734), .A2(n7268), .ZN(n7267) );
  NAND2_X1 U10050 ( .A1(n11942), .A2(n11941), .ZN(n11940) );
  NAND2_X2 U10051 ( .A1(n14725), .A2(n7855), .ZN(n14976) );
  NAND2_X1 U10052 ( .A1(n10947), .A2(n10946), .ZN(n11595) );
  NAND3_X1 U10053 ( .A1(n7251), .A2(n8474), .A3(n7162), .ZN(n7161) );
  XNOR2_X2 U10054 ( .A(n9003), .B(SI_18_), .ZN(n9022) );
  NAND2_X1 U10055 ( .A1(n11470), .A2(n9343), .ZN(n11464) );
  NAND2_X1 U10056 ( .A1(n8944), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U10057 ( .A1(n9339), .A2(n6505), .ZN(n11471) );
  NAND2_X1 U10058 ( .A1(n6547), .A2(n7164), .ZN(n11340) );
  INV_X1 U10059 ( .A(n7518), .ZN(n11547) );
  INV_X1 U10060 ( .A(n10120), .ZN(n10121) );
  NAND2_X1 U10061 ( .A1(n8323), .A2(n7875), .ZN(n8350) );
  NAND2_X1 U10062 ( .A1(n6486), .A2(n7171), .ZN(n10325) );
  OR2_X2 U10063 ( .A1(n7173), .A2(n13350), .ZN(n7172) );
  NAND4_X1 U10064 ( .A1(n10323), .A2(n10322), .A3(n7174), .A4(n6725), .ZN(
        n7173) );
  AOI22_X1 U10065 ( .A1(n10192), .A2(n10311), .B1(n10193), .B2(n10532), .ZN(
        n10194) );
  INV_X2 U10066 ( .A(n8470), .ZN(n7315) );
  INV_X1 U10067 ( .A(n10631), .ZN(n7183) );
  NAND2_X1 U10068 ( .A1(n15155), .A2(n15156), .ZN(n11136) );
  NAND2_X1 U10069 ( .A1(n12608), .A2(n12607), .ZN(n12610) );
  INV_X1 U10070 ( .A(n10649), .ZN(n10646) );
  NAND2_X1 U10071 ( .A1(n7356), .A2(n11449), .ZN(n11456) );
  NAND2_X1 U10072 ( .A1(n15218), .A2(n7363), .ZN(n15216) );
  NAND2_X1 U10073 ( .A1(n11965), .A2(n6860), .ZN(n11964) );
  AOI21_X1 U10074 ( .B1(n7303), .B2(n7306), .A(n7302), .ZN(n7301) );
  OR4_X2 U10075 ( .A1(n9289), .A2(n10429), .A3(n14078), .A4(n9288), .ZN(n9290)
         );
  NAND2_X1 U10076 ( .A1(n6472), .A2(n8830), .ZN(n7684) );
  NAND2_X1 U10077 ( .A1(n7184), .A2(n8583), .ZN(n8872) );
  NAND2_X1 U10078 ( .A1(n7189), .A2(n6581), .ZN(n7190) );
  NAND2_X1 U10079 ( .A1(n7189), .A2(n6582), .ZN(n9305) );
  INV_X1 U10080 ( .A(n9338), .ZN(n7191) );
  NAND2_X1 U10081 ( .A1(n8745), .A2(n8746), .ZN(n8744) );
  NAND2_X1 U10082 ( .A1(n8807), .A2(n6431), .ZN(n7195) );
  NAND2_X1 U10083 ( .A1(n7578), .A2(n7204), .ZN(n7200) );
  NAND2_X1 U10084 ( .A1(n7200), .A2(n7201), .ZN(n8959) );
  AND2_X1 U10085 ( .A1(n7234), .A2(n7233), .ZN(n13352) );
  NAND2_X1 U10086 ( .A1(n6550), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n7244) );
  MUX2_X1 U10087 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n10567), .Z(n8643) );
  NAND2_X2 U10088 ( .A1(n8810), .A2(n8808), .ZN(n8492) );
  NAND2_X1 U10089 ( .A1(n8469), .A2(n7250), .ZN(n7251) );
  AND2_X1 U10090 ( .A1(n8473), .A2(n8468), .ZN(n7250) );
  INV_X1 U10091 ( .A(n8492), .ZN(n7263) );
  MUX2_X1 U10092 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10567), .Z(n8478) );
  MUX2_X1 U10093 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10567), .Z(n8494) );
  MUX2_X1 U10094 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6776), .Z(n8487) );
  MUX2_X1 U10095 ( .A(n11061), .B(n11078), .S(n6776), .Z(n8504) );
  MUX2_X1 U10096 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6776), .Z(n8936) );
  MUX2_X1 U10097 ( .A(n12933), .B(n11663), .S(n6776), .Z(n9040) );
  MUX2_X1 U10098 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6776), .Z(n9108) );
  MUX2_X1 U10099 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6776), .Z(n8523) );
  MUX2_X1 U10100 ( .A(n11090), .B(n11093), .S(n6776), .Z(n8516) );
  MUX2_X1 U10101 ( .A(n12386), .B(n12383), .S(n6776), .Z(n8538) );
  MUX2_X1 U10102 ( .A(n12738), .B(n12597), .S(n10567), .Z(n9056) );
  MUX2_X1 U10103 ( .A(n15148), .B(n8545), .S(n10567), .Z(n8546) );
  MUX2_X1 U10104 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6776), .Z(n8554) );
  NAND2_X2 U10105 ( .A1(P1_U3086), .A2(n10572), .ZN(n15141) );
  NAND2_X2 U10106 ( .A1(n7269), .A2(n9761), .ZN(n15097) );
  NAND2_X1 U10107 ( .A1(n11386), .A2(n7277), .ZN(n7276) );
  INV_X1 U10108 ( .A(n7282), .ZN(n11676) );
  NOR2_X1 U10109 ( .A1(n11388), .A2(n11387), .ZN(n7284) );
  INV_X1 U10110 ( .A(n14679), .ZN(n7290) );
  AND2_X1 U10111 ( .A1(n7297), .A2(n6483), .ZN(n7298) );
  NAND2_X1 U10112 ( .A1(n12730), .A2(n6501), .ZN(n7299) );
  NAND2_X1 U10113 ( .A1(n8492), .A2(n7303), .ZN(n7300) );
  XNOR2_X1 U10114 ( .A(n7307), .B(n8658), .ZN(n10667) );
  NAND2_X1 U10115 ( .A1(n8520), .A2(n6481), .ZN(n7309) );
  NAND2_X1 U10116 ( .A1(n8633), .A2(n7314), .ZN(n14452) );
  NAND2_X1 U10117 ( .A1(n14755), .A2(n7321), .ZN(n7318) );
  NAND2_X2 U10118 ( .A1(n10080), .A2(n12696), .ZN(n14806) );
  OR2_X2 U10119 ( .A1(n12756), .A2(n14826), .ZN(n12696) );
  NAND4_X1 U10120 ( .A1(n7888), .A2(n7886), .A3(n7887), .A4(n8035), .ZN(n7326)
         );
  INV_X1 U10121 ( .A(n7891), .ZN(n8428) );
  NAND4_X1 U10122 ( .A1(n7882), .A2(n7883), .A3(n7884), .A4(n7881), .ZN(n7327)
         );
  NAND2_X1 U10123 ( .A1(n10183), .A2(n7341), .ZN(n7340) );
  INV_X1 U10124 ( .A(n10181), .ZN(n7347) );
  NAND2_X1 U10125 ( .A1(n15209), .A2(n15208), .ZN(n7360) );
  NAND2_X1 U10126 ( .A1(n15209), .A2(n7361), .ZN(n7363) );
  NAND3_X1 U10127 ( .A1(n7363), .A2(n14015), .A3(n15218), .ZN(n7362) );
  INV_X1 U10128 ( .A(n7362), .ZN(n15219) );
  AOI21_X1 U10129 ( .B1(n10627), .B2(n10617), .A(n7370), .ZN(n7365) );
  OAI21_X1 U10130 ( .B1(n10617), .B2(n7370), .A(n7371), .ZN(n7367) );
  NAND2_X1 U10131 ( .A1(n10627), .A2(n6556), .ZN(n7369) );
  INV_X1 U10132 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7371) );
  NAND3_X1 U10133 ( .A1(n7373), .A2(n12405), .A3(n7372), .ZN(n12608) );
  INV_X1 U10134 ( .A(n12031), .ZN(n7374) );
  INV_X1 U10135 ( .A(n12032), .ZN(n7375) );
  NAND2_X1 U10136 ( .A1(n15170), .A2(n7382), .ZN(n7376) );
  NAND2_X1 U10137 ( .A1(n7386), .A2(n7387), .ZN(n11488) );
  NAND2_X1 U10138 ( .A1(n11265), .A2(n7390), .ZN(n7386) );
  NAND2_X1 U10139 ( .A1(n7396), .A2(n7398), .ZN(n13187) );
  CLKBUF_X1 U10140 ( .A(n8246), .Z(n7420) );
  NAND2_X1 U10141 ( .A1(n7420), .A2(SI_24_), .ZN(n8321) );
  INV_X2 U10142 ( .A(n10255), .ZN(n8246) );
  NAND2_X1 U10143 ( .A1(n13429), .A2(n7424), .ZN(n7423) );
  NAND2_X1 U10144 ( .A1(n13402), .A2(n8332), .ZN(n8334) );
  NAND2_X1 U10145 ( .A1(n14221), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U10146 ( .A1(n7433), .A2(n14221), .ZN(n14166) );
  INV_X1 U10147 ( .A(n7436), .ZN(n7433) );
  NAND3_X1 U10148 ( .A1(n7444), .A2(n13870), .A3(n7443), .ZN(n7445) );
  NAND2_X1 U10149 ( .A1(n12552), .A2(n12555), .ZN(n12554) );
  XNOR2_X1 U10150 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n7903) );
  OAI21_X1 U10151 ( .B1(n10320), .B2(n6575), .A(n7456), .ZN(n7455) );
  NOR2_X1 U10152 ( .A1(n13604), .A2(n13321), .ZN(n7458) );
  NAND2_X1 U10153 ( .A1(n8146), .A2(n7469), .ZN(n7467) );
  OAI21_X1 U10154 ( .B1(n8371), .B2(n7483), .A(n7480), .ZN(n10261) );
  OAI21_X1 U10155 ( .B1(n8371), .B2(n8370), .A(n8372), .ZN(n10254) );
  NAND2_X1 U10156 ( .A1(n8370), .A2(n8372), .ZN(n7484) );
  NAND2_X1 U10157 ( .A1(n8336), .A2(n7487), .ZN(n7485) );
  NAND2_X2 U10158 ( .A1(n13185), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n13208) );
  AND2_X2 U10159 ( .A1(n7490), .A2(n13206), .ZN(n13185) );
  NAND2_X1 U10160 ( .A1(n13184), .A2(n13183), .ZN(n13206) );
  NAND2_X1 U10161 ( .A1(n7491), .A2(n13213), .ZN(n7490) );
  INV_X1 U10162 ( .A(n13184), .ZN(n7491) );
  AND2_X2 U10163 ( .A1(n7493), .A2(n7492), .ZN(n13230) );
  NAND3_X1 U10164 ( .A1(n13228), .A2(n13232), .A3(n13246), .ZN(n7492) );
  NAND4_X1 U10165 ( .A1(n7502), .A2(n6435), .A3(n7500), .A4(n7498), .ZN(n13312) );
  NAND2_X1 U10166 ( .A1(n7507), .A2(n12075), .ZN(n12073) );
  INV_X1 U10167 ( .A(n13144), .ZN(n7513) );
  OAI211_X1 U10168 ( .C1(n11424), .C2(n11491), .A(n7515), .B(n11490), .ZN(
        n11920) );
  XNOR2_X1 U10169 ( .A(n11422), .B(n6897), .ZN(n11424) );
  OAI21_X1 U10170 ( .B1(n11348), .B2(n11347), .A(n9354), .ZN(n7518) );
  NAND2_X1 U10171 ( .A1(n11547), .A2(n11546), .ZN(n11545) );
  INV_X1 U10172 ( .A(n8588), .ZN(n7533) );
  NAND2_X1 U10173 ( .A1(n8588), .A2(n7535), .ZN(n7534) );
  OR2_X2 U10174 ( .A1(n8919), .A2(n7533), .ZN(n8590) );
  NOR2_X2 U10175 ( .A1(n8919), .A2(n7534), .ZN(n8601) );
  OAI211_X2 U10176 ( .C1(n8666), .C2(n10667), .A(n8665), .B(n8664), .ZN(n11619) );
  INV_X1 U10177 ( .A(n11340), .ZN(n9339) );
  NAND2_X2 U10178 ( .A1(n14262), .A2(n11587), .ZN(n9349) );
  NAND3_X1 U10179 ( .A1(n9525), .A2(n7541), .A3(n9522), .ZN(n10103) );
  INV_X1 U10180 ( .A(n11225), .ZN(n11754) );
  AOI21_X1 U10181 ( .B1(n14692), .B2(n6447), .A(n6558), .ZN(n7547) );
  NAND2_X1 U10182 ( .A1(n7555), .A2(n9311), .ZN(n8919) );
  AND2_X1 U10183 ( .A1(n7555), .A2(n8596), .ZN(n9313) );
  NOR2_X2 U10184 ( .A1(n8872), .A2(n8584), .ZN(n7555) );
  OAI21_X1 U10185 ( .B1(n9037), .B2(n7563), .A(n7566), .ZN(n7562) );
  INV_X1 U10186 ( .A(n9037), .ZN(n7568) );
  INV_X1 U10187 ( .A(n8786), .ZN(n7571) );
  INV_X1 U10188 ( .A(n8785), .ZN(n7572) );
  NAND2_X1 U10189 ( .A1(n7574), .A2(n7575), .ZN(n8893) );
  NAND2_X1 U10190 ( .A1(n7580), .A2(n7579), .ZN(n10044) );
  NAND2_X1 U10191 ( .A1(n9999), .A2(n9998), .ZN(n7579) );
  NAND2_X1 U10192 ( .A1(n9995), .A2(n9994), .ZN(n7580) );
  NAND3_X1 U10193 ( .A1(n7580), .A2(n7579), .A3(n6568), .ZN(n10122) );
  NAND2_X1 U10194 ( .A1(n7584), .A2(n7585), .ZN(n9735) );
  NAND2_X1 U10195 ( .A1(n9720), .A2(n7587), .ZN(n7584) );
  INV_X1 U10196 ( .A(n9559), .ZN(n9552) );
  NAND3_X1 U10197 ( .A1(n7750), .A2(n6473), .A3(n7749), .ZN(n9563) );
  AOI21_X1 U10198 ( .B1(n7600), .B2(n7599), .A(n7598), .ZN(n7597) );
  INV_X1 U10199 ( .A(n9886), .ZN(n7598) );
  NAND2_X1 U10200 ( .A1(n7601), .A2(n6586), .ZN(n9681) );
  NAND3_X1 U10201 ( .A1(n9919), .A2(n9918), .A3(n7607), .ZN(n7604) );
  NAND2_X1 U10202 ( .A1(n7604), .A2(n7605), .ZN(n9946) );
  NOR2_X1 U10203 ( .A1(n10302), .A2(n7609), .ZN(n11540) );
  NAND2_X1 U10204 ( .A1(n13531), .A2(n7623), .ZN(n7622) );
  INV_X1 U10205 ( .A(n10189), .ZN(n7629) );
  NAND2_X1 U10206 ( .A1(n13531), .A2(n13535), .ZN(n13530) );
  NAND2_X1 U10207 ( .A1(n11792), .A2(n7633), .ZN(n7632) );
  OAI21_X1 U10208 ( .B1(n7639), .B2(n7637), .A(n7631), .ZN(n7630) );
  INV_X1 U10209 ( .A(n10159), .ZN(n7642) );
  NAND2_X1 U10210 ( .A1(n13414), .A2(n7651), .ZN(n7648) );
  NAND2_X1 U10211 ( .A1(n7649), .A2(n7648), .ZN(n10281) );
  NAND2_X1 U10212 ( .A1(n13414), .A2(n13370), .ZN(n7657) );
  NAND4_X1 U10213 ( .A1(n7891), .A2(n8093), .A3(n7890), .A4(n7660), .ZN(n8426)
         );
  NAND4_X2 U10214 ( .A1(n7969), .A2(n7970), .A3(n7661), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7974) );
  INV_X2 U10215 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7970) );
  INV_X1 U10216 ( .A(n13064), .ZN(n7662) );
  NAND2_X1 U10217 ( .A1(n7662), .A2(n13418), .ZN(n13062) );
  NAND2_X1 U10218 ( .A1(n13062), .A2(n12955), .ZN(n7667) );
  INV_X1 U10219 ( .A(n12956), .ZN(n7665) );
  OAI21_X1 U10220 ( .B1(n12945), .B2(n12946), .A(n7677), .ZN(n13105) );
  NAND2_X1 U10221 ( .A1(n10464), .A2(n7687), .ZN(n7686) );
  INV_X1 U10222 ( .A(n11759), .ZN(n7687) );
  INV_X1 U10223 ( .A(n12123), .ZN(n7688) );
  AOI21_X1 U10224 ( .B1(n8530), .B2(n8531), .A(n6588), .ZN(n7696) );
  NAND2_X1 U10225 ( .A1(n9227), .A2(n8550), .ZN(n9213) );
  NAND3_X1 U10226 ( .A1(n7889), .A2(n8008), .A3(n8092), .ZN(n8113) );
  INV_X1 U10227 ( .A(n8429), .ZN(n8114) );
  OR2_X2 U10228 ( .A1(n14485), .A2(n6560), .ZN(n7717) );
  NAND2_X1 U10229 ( .A1(n14573), .A2(n7722), .ZN(n7721) );
  NAND2_X1 U10230 ( .A1(n11193), .A2(n7727), .ZN(n7729) );
  NAND2_X1 U10231 ( .A1(n14504), .A2(n7734), .ZN(n7731) );
  NAND2_X1 U10232 ( .A1(n14504), .A2(n14505), .ZN(n7733) );
  NAND2_X1 U10233 ( .A1(n12529), .A2(n12528), .ZN(n12530) );
  INV_X1 U10234 ( .A(n7746), .ZN(n12766) );
  NOR2_X1 U10235 ( .A1(n12531), .A2(n7748), .ZN(n7747) );
  INV_X1 U10236 ( .A(n12528), .ZN(n7748) );
  NAND2_X1 U10237 ( .A1(n9563), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9564) );
  INV_X1 U10238 ( .A(n9551), .ZN(n7750) );
  OAI21_X1 U10239 ( .B1(n7753), .B2(n10390), .A(n10392), .ZN(n7752) );
  NAND2_X1 U10240 ( .A1(n7756), .A2(n7754), .ZN(n10425) );
  NAND2_X1 U10241 ( .A1(n14215), .A2(n7757), .ZN(n7756) );
  OAI21_X1 U10242 ( .B1(n7138), .B2(n7759), .A(n7757), .ZN(n14160) );
  OR2_X1 U10243 ( .A1(n14209), .A2(n10421), .ZN(n7766) );
  NAND2_X1 U10244 ( .A1(n7136), .A2(n10376), .ZN(n14158) );
  AND2_X1 U10245 ( .A1(n7804), .A2(n10941), .ZN(n11757) );
  NAND2_X1 U10246 ( .A1(n10939), .A2(n10940), .ZN(n7804) );
  INV_X1 U10247 ( .A(n14789), .ZN(n7818) );
  INV_X1 U10248 ( .A(n12188), .ZN(n7829) );
  NAND2_X1 U10249 ( .A1(n12037), .A2(n7833), .ZN(n7831) );
  AND2_X1 U10250 ( .A1(n7834), .A2(n11878), .ZN(n7833) );
  NAND3_X1 U10251 ( .A1(n7831), .A2(n7830), .A3(n11881), .ZN(n12118) );
  NAND2_X1 U10252 ( .A1(n8980), .A2(n6398), .ZN(n8999) );
  INV_X1 U10253 ( .A(n14262), .ZN(n14363) );
  NAND2_X1 U10254 ( .A1(n14262), .A2(n14031), .ZN(n10443) );
  CLKBUF_X1 U10255 ( .A(n8393), .Z(n13701) );
  NAND2_X1 U10256 ( .A1(n15151), .A2(n10011), .ZN(n10970) );
  AND2_X4 U10257 ( .A1(n7896), .A2(n13694), .ZN(n10268) );
  INV_X1 U10258 ( .A(n7897), .ZN(n13694) );
  INV_X1 U10259 ( .A(n10105), .ZN(n10101) );
  NAND2_X1 U10260 ( .A1(n9949), .A2(n9948), .ZN(n9950) );
  NAND2_X1 U10262 ( .A1(n7998), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U10263 ( .A1(n10350), .A2(n15585), .ZN(n8459) );
  NAND2_X1 U10264 ( .A1(n8641), .A2(n8640), .ZN(n8672) );
  AND2_X1 U10265 ( .A1(n11103), .A2(n6405), .ZN(n10522) );
  NAND2_X1 U10266 ( .A1(n8470), .A2(n10668), .ZN(n8460) );
  INV_X1 U10267 ( .A(n10448), .ZN(n10531) );
  AND2_X1 U10268 ( .A1(n11555), .A2(n13321), .ZN(n15507) );
  XNOR2_X1 U10269 ( .A(n9058), .B(n9057), .ZN(n12596) );
  NOR2_X1 U10270 ( .A1(n8595), .A2(n8587), .ZN(n8588) );
  XNOR2_X1 U10271 ( .A(n9323), .B(n9325), .ZN(n12141) );
  NAND2_X1 U10272 ( .A1(n12939), .A2(n10006), .ZN(n11746) );
  INV_X1 U10273 ( .A(n10006), .ZN(n15151) );
  NAND2_X4 U10274 ( .A1(n11207), .A2(n10749), .ZN(n12857) );
  NAND2_X4 U10275 ( .A1(n10583), .A2(n10113), .ZN(n11207) );
  AND4_X4 U10276 ( .A1(n9582), .A2(n9581), .A3(n9580), .A4(n9579), .ZN(n11152)
         );
  OR2_X1 U10277 ( .A1(n15583), .A2(n15567), .ZN(n13681) );
  INV_X1 U10278 ( .A(n15595), .ZN(n15593) );
  AND2_X2 U10279 ( .A1(n10349), .A2(n11702), .ZN(n15595) );
  INV_X1 U10280 ( .A(n10259), .ZN(n13340) );
  INV_X1 U10281 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10593) );
  OR2_X1 U10282 ( .A1(n14398), .A2(n14362), .ZN(n7854) );
  OR2_X1 U10283 ( .A1(n15000), .A2(n14603), .ZN(n7855) );
  NOR4_X1 U10284 ( .A1(n13428), .A2(n10315), .A3(n13467), .A4(n10314), .ZN(
        n7857) );
  AND2_X1 U10285 ( .A1(n9304), .A2(n11932), .ZN(n7858) );
  INV_X1 U10286 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13686) );
  NAND2_X1 U10287 ( .A1(n15595), .A2(n13586), .ZN(n13597) );
  INV_X1 U10288 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9540) );
  AND2_X1 U10289 ( .A1(n11200), .A2(n11199), .ZN(n7859) );
  OR2_X1 U10290 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n11232), .ZN(n7860) );
  NAND2_X2 U10291 ( .A1(n11741), .A2(n14946), .ZN(n14940) );
  INV_X2 U10292 ( .A(P2_U3947), .ZN(n13945) );
  INV_X1 U10293 ( .A(n12295), .ZN(n12179) );
  AND2_X1 U10294 ( .A1(n9156), .A2(n9155), .ZN(n7862) );
  NOR4_X1 U10295 ( .A1(n14886), .A2(n10090), .A3(n12711), .A4(n14927), .ZN(
        n7863) );
  INV_X1 U10296 ( .A(n14242), .ZN(n14264) );
  NAND2_X2 U10297 ( .A1(n14239), .A2(n11406), .ZN(n14242) );
  AND2_X2 U10298 ( .A1(n10981), .A2(n10980), .ZN(n15494) );
  INV_X1 U10299 ( .A(n15494), .ZN(n15492) );
  INV_X1 U10300 ( .A(n14082), .ZN(n14199) );
  NAND2_X1 U10301 ( .A1(n9467), .A2(n9466), .ZN(n9468) );
  AND4_X1 U10302 ( .A1(n14958), .A2(n9788), .A3(n9787), .A4(n9786), .ZN(n7864)
         );
  AOI22_X1 U10303 ( .A1(n8701), .A2(n8700), .B1(n8696), .B2(n8695), .ZN(n8697)
         );
  INV_X1 U10304 ( .A(n9751), .ZN(n9752) );
  NOR2_X1 U10305 ( .A1(n10132), .A2(n15511), .ZN(n10133) );
  NAND2_X1 U10306 ( .A1(n10162), .A2(n10161), .ZN(n10163) );
  NAND2_X1 U10307 ( .A1(n9917), .A2(n6769), .ZN(n9918) );
  INV_X1 U10308 ( .A(n9161), .ZN(n9158) );
  INV_X1 U10309 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7886) );
  INV_X1 U10310 ( .A(n9261), .ZN(n9262) );
  INV_X1 U10311 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9008) );
  INV_X1 U10312 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8545) );
  AND2_X1 U10313 ( .A1(n9136), .A2(SI_20_), .ZN(n8529) );
  INV_X1 U10314 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10614) );
  OR2_X1 U10315 ( .A1(n10532), .A2(n10531), .ZN(n11696) );
  NAND2_X1 U10316 ( .A1(n9062), .A2(n9061), .ZN(n9114) );
  AND2_X1 U10317 ( .A1(n13952), .A2(n11619), .ZN(n10354) );
  XNOR2_X1 U10318 ( .A(n11171), .B(n12866), .ZN(n11172) );
  OR2_X1 U10319 ( .A1(n10055), .A2(n11210), .ZN(n10043) );
  INV_X1 U10320 ( .A(n14913), .ZN(n12689) );
  OR2_X1 U10321 ( .A1(n12007), .A2(n11152), .ZN(n10944) );
  INV_X1 U10322 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n15674) );
  NOR2_X1 U10323 ( .A1(n11451), .A2(n11450), .ZN(n11452) );
  INV_X1 U10324 ( .A(n13076), .ZN(n10479) );
  OR2_X1 U10325 ( .A1(n10532), .A2(n10448), .ZN(n11369) );
  NAND2_X1 U10326 ( .A1(n12619), .A2(n13333), .ZN(n8403) );
  NAND2_X1 U10327 ( .A1(n7877), .A2(n7876), .ZN(n8362) );
  OR3_X1 U10328 ( .A1(n11459), .A2(n13321), .A3(n11555), .ZN(n10334) );
  NAND2_X1 U10329 ( .A1(n8389), .A2(n8383), .ZN(n8421) );
  NAND2_X1 U10330 ( .A1(n8243), .A2(n7941), .ZN(n7943) );
  OR2_X1 U10331 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  OR2_X1 U10332 ( .A1(n9094), .A2(n9063), .ZN(n9184) );
  INV_X1 U10333 ( .A(n8673), .ZN(n8706) );
  NAND2_X1 U10334 ( .A1(n8968), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8990) );
  OR2_X1 U10335 ( .A1(n13952), .A2(n11619), .ZN(n11080) );
  NAND2_X1 U10336 ( .A1(n8600), .A2(n8601), .ZN(n8603) );
  OR2_X1 U10337 ( .A1(n11173), .A2(n11172), .ZN(n11174) );
  OR2_X1 U10338 ( .A1(n12852), .A2(n12851), .ZN(n12853) );
  INV_X1 U10339 ( .A(n11829), .ZN(n11826) );
  INV_X1 U10340 ( .A(n11210), .ZN(n10050) );
  INV_X1 U10341 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12671) );
  AND2_X1 U10342 ( .A1(n14991), .A2(n14708), .ZN(n14709) );
  OR2_X1 U10343 ( .A1(n12875), .A2(n10922), .ZN(n11904) );
  INV_X1 U10344 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15627) );
  INV_X1 U10345 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11453) );
  OAI21_X1 U10346 ( .B1(n13021), .B2(n12995), .A(n12994), .ZN(n12993) );
  INV_X1 U10347 ( .A(n13488), .ZN(n13085) );
  INV_X1 U10348 ( .A(n10525), .ZN(n10537) );
  OR2_X1 U10349 ( .A1(n10451), .A2(n10336), .ZN(n10524) );
  INV_X1 U10350 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n11253) );
  INV_X1 U10351 ( .A(n13311), .ZN(n13164) );
  INV_X1 U10352 ( .A(n15503), .ZN(n13291) );
  OR2_X1 U10353 ( .A1(n13701), .A2(n13703), .ZN(n11103) );
  OR2_X1 U10354 ( .A1(n15585), .A2(n15671), .ZN(n8457) );
  INV_X1 U10355 ( .A(n15532), .ZN(n13522) );
  INV_X1 U10356 ( .A(n8441), .ZN(n10801) );
  AND2_X1 U10357 ( .A1(n7908), .A2(n7907), .ZN(n8006) );
  INV_X1 U10358 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9296) );
  AND2_X1 U10359 ( .A1(n9441), .A2(n7856), .ZN(n9442) );
  AND2_X1 U10360 ( .A1(n10856), .A2(n10859), .ZN(n14082) );
  OR2_X1 U10361 ( .A1(n13919), .A2(n14197), .ZN(n13912) );
  OR2_X1 U10362 ( .A1(n15462), .A2(n11402), .ZN(n9499) );
  INV_X1 U10363 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n12252) );
  AOI21_X1 U10364 ( .B1(n14291), .B2(n14273), .A(n12928), .ZN(n12929) );
  NAND2_X1 U10365 ( .A1(n10856), .A2(n9329), .ZN(n14197) );
  INV_X1 U10366 ( .A(n13753), .ZN(n12555) );
  INV_X1 U10367 ( .A(n14278), .ZN(n14226) );
  OR2_X1 U10368 ( .A1(n10976), .A2(n15462), .ZN(n10444) );
  AND2_X1 U10369 ( .A1(n12213), .A2(n12212), .ZN(n12542) );
  AND2_X1 U10370 ( .A1(n11851), .A2(n11850), .ZN(n15485) );
  INV_X1 U10371 ( .A(n14252), .ZN(n14217) );
  INV_X1 U10372 ( .A(n9497), .ZN(n9494) );
  OR2_X1 U10373 ( .A1(n10977), .A2(n10976), .ZN(n10979) );
  INV_X1 U10374 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9316) );
  NAND2_X1 U10375 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n8591), .ZN(n8592) );
  INV_X1 U10376 ( .A(n15238), .ZN(n11175) );
  INV_X1 U10377 ( .A(n14610), .ZN(n14915) );
  OR2_X1 U10378 ( .A1(n14595), .A2(n14916), .ZN(n14556) );
  INV_X1 U10379 ( .A(n10026), .ZN(n9966) );
  INV_X1 U10380 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11391) );
  OR2_X1 U10381 ( .A1(n14868), .A2(n10081), .ZN(n14886) );
  INV_X1 U10382 ( .A(n12286), .ZN(n12298) );
  NAND3_X1 U10383 ( .A1(n11740), .A2(n7274), .A3(n14949), .ZN(n14946) );
  NOR2_X1 U10384 ( .A1(n11904), .A2(n7274), .ZN(n14873) );
  AND2_X1 U10385 ( .A1(n11736), .A2(n10967), .ZN(n10918) );
  INV_X1 U10386 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10041) );
  AND2_X1 U10387 ( .A1(n8514), .A2(n8513), .ZN(n8960) );
  AND2_X1 U10388 ( .A1(n8503), .A2(n8502), .ZN(n8896) );
  OAI21_X1 U10389 ( .B1(n13366), .B2(n13103), .A(n10541), .ZN(n10542) );
  OR2_X1 U10390 ( .A1(n10538), .A2(n10521), .ZN(n13109) );
  INV_X1 U10391 ( .A(n13098), .ZN(n13107) );
  OAI211_X1 U10392 ( .C1(n10538), .C2(n10537), .A(n10536), .B(n11783), .ZN(
        n13045) );
  INV_X1 U10393 ( .A(n13314), .ZN(n13293) );
  OAI21_X1 U10394 ( .B1(n6725), .B2(n13360), .A(n6463), .ZN(n13551) );
  NAND2_X1 U10395 ( .A1(n10336), .A2(n10290), .ZN(n15532) );
  AND2_X1 U10396 ( .A1(n15524), .A2(n15523), .ZN(n15545) );
  INV_X1 U10397 ( .A(n13534), .ZN(n13519) );
  INV_X1 U10398 ( .A(n13597), .ZN(n13590) );
  NOR2_X1 U10399 ( .A1(n11098), .A2(n10348), .ZN(n11702) );
  NOR2_X1 U10400 ( .A1(n13335), .A2(n13334), .ZN(n13602) );
  AND2_X1 U10401 ( .A1(n10179), .A2(n10180), .ZN(n12468) );
  INV_X1 U10402 ( .A(n13681), .ZN(n13670) );
  INV_X1 U10403 ( .A(n12227), .ZN(n15569) );
  NAND2_X1 U10404 ( .A1(n11459), .A2(n11766), .ZN(n15567) );
  NAND2_X1 U10405 ( .A1(n8438), .A2(n8437), .ZN(n11697) );
  INV_X1 U10406 ( .A(n8389), .ZN(n8390) );
  AND2_X1 U10407 ( .A1(n8210), .A2(n6593), .ZN(n13259) );
  INV_X1 U10408 ( .A(n13921), .ZN(n13872) );
  NOR2_X1 U10409 ( .A1(n15463), .A2(n9499), .ZN(n9495) );
  AND2_X1 U10410 ( .A1(n9035), .A2(n9034), .ZN(n14200) );
  INV_X1 U10411 ( .A(n15411), .ZN(n15451) );
  OAI21_X1 U10412 ( .B1(n14294), .B2(n14280), .A(n12929), .ZN(n12930) );
  INV_X1 U10413 ( .A(n14197), .ZN(n14097) );
  INV_X1 U10414 ( .A(n14248), .ZN(n14268) );
  INV_X1 U10415 ( .A(n14239), .ZN(n14276) );
  NOR2_X1 U10416 ( .A1(n10444), .A2(n10978), .ZN(n10445) );
  OR2_X1 U10417 ( .A1(n15494), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n14396) );
  INV_X1 U10418 ( .A(n14386), .ZN(n14366) );
  NOR2_X1 U10419 ( .A1(n10979), .A2(n10978), .ZN(n10980) );
  NOR2_X1 U10420 ( .A1(n9326), .A2(n12141), .ZN(n10545) );
  INV_X1 U10421 ( .A(n9315), .ZN(n9318) );
  INV_X1 U10422 ( .A(n15246), .ZN(n14597) );
  AND3_X1 U10423 ( .A1(n10005), .A2(n10004), .A3(n10003), .ZN(n14697) );
  INV_X1 U10424 ( .A(n12658), .ZN(n15264) );
  INV_X1 U10425 ( .A(n14677), .ZN(n15267) );
  INV_X1 U10426 ( .A(n14687), .ZN(n15266) );
  INV_X1 U10427 ( .A(n14983), .ZN(n14980) );
  INV_X1 U10428 ( .A(n14953), .ZN(n14924) );
  AND2_X1 U10429 ( .A1(n14940), .A2(n11905), .ZN(n14841) );
  INV_X1 U10430 ( .A(n15297), .ZN(n15304) );
  NAND2_X1 U10431 ( .A1(n10926), .A2(n10925), .ZN(n15308) );
  AND2_X1 U10432 ( .A1(n10006), .A2(n10924), .ZN(n15282) );
  NAND2_X1 U10433 ( .A1(n10582), .A2(n10583), .ZN(n10963) );
  INV_X1 U10434 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10111) );
  AND2_X1 U10435 ( .A1(n9747), .A2(n9758), .ZN(n11680) );
  AND2_X1 U10436 ( .A1(n11111), .A2(n11110), .ZN(n15503) );
  INV_X1 U10437 ( .A(n13045), .ZN(n13088) );
  NAND2_X1 U10438 ( .A1(n10517), .A2(n10516), .ZN(n13115) );
  INV_X1 U10439 ( .A(n13501), .ZN(n13469) );
  MUX2_X1 U10440 ( .A(n13130), .B(n11112), .S(n13701), .Z(n13314) );
  INV_X1 U10441 ( .A(n13322), .ZN(n13283) );
  NAND2_X1 U10442 ( .A1(n12084), .A2(n13586), .ZN(n13534) );
  NAND2_X1 U10443 ( .A1(n15524), .A2(n12303), .ZN(n13529) );
  NAND2_X1 U10444 ( .A1(n15569), .A2(n15595), .ZN(n13592) );
  OR2_X1 U10445 ( .A1(n15583), .A2(n12227), .ZN(n13673) );
  AND2_X1 U10446 ( .A1(n8456), .A2(n8455), .ZN(n15583) );
  INV_X1 U10447 ( .A(SI_26_), .ZN(n12560) );
  INV_X1 U10448 ( .A(SI_21_), .ZN(n11767) );
  INV_X1 U10449 ( .A(SI_16_), .ZN(n10835) );
  INV_X1 U10450 ( .A(SI_11_), .ZN(n10608) );
  NOR2_X1 U10451 ( .A1(n10860), .A2(P2_U3088), .ZN(n15336) );
  INV_X1 U10452 ( .A(n13909), .ZN(n13900) );
  INV_X1 U10453 ( .A(n13926), .ZN(n13905) );
  NAND2_X1 U10454 ( .A1(n9495), .A2(n9487), .ZN(n13921) );
  NAND2_X1 U10455 ( .A1(n9191), .A2(n9190), .ZN(n14065) );
  INV_X1 U10456 ( .A(n14200), .ZN(n13934) );
  INV_X1 U10457 ( .A(n12583), .ZN(n13941) );
  NAND2_X1 U10458 ( .A1(n10861), .A2(n12916), .ZN(n15411) );
  INV_X1 U10459 ( .A(n12930), .ZN(n12931) );
  NAND2_X1 U10460 ( .A1(n14242), .A2(n11666), .ZN(n14248) );
  AND2_X1 U10461 ( .A1(n11501), .A2(n11502), .ZN(n11637) );
  NAND2_X1 U10462 ( .A1(n15502), .A2(n15479), .ZN(n14362) );
  INV_X1 U10463 ( .A(n14089), .ZN(n14404) );
  INV_X1 U10464 ( .A(n14222), .ZN(n14429) );
  NAND2_X1 U10465 ( .A1(n15494), .A2(n15479), .ZN(n14428) );
  NOR2_X1 U10466 ( .A1(n15458), .A2(n15463), .ZN(n15459) );
  OR2_X1 U10467 ( .A1(n10545), .A2(n9327), .ZN(n15463) );
  INV_X1 U10468 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12597) );
  INV_X1 U10469 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11443) );
  INV_X1 U10470 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10733) );
  AND2_X1 U10471 ( .A1(n10697), .A2(n10662), .ZN(n15255) );
  AND2_X1 U10472 ( .A1(n11211), .A2(n11210), .ZN(n15246) );
  NAND2_X1 U10473 ( .A1(n10972), .A2(n10971), .ZN(n15237) );
  INV_X1 U10474 ( .A(n14586), .ZN(n14600) );
  OR2_X1 U10475 ( .A1(n15258), .A2(n10756), .ZN(n14687) );
  OR2_X1 U10476 ( .A1(n15258), .A2(n10708), .ZN(n14677) );
  OR2_X1 U10477 ( .A1(n11750), .A2(n11749), .ZN(n14953) );
  INV_X1 U10478 ( .A(n14841), .ZN(n14969) );
  AND2_X2 U10479 ( .A1(n10959), .A2(n11739), .ZN(n15316) );
  INV_X1 U10480 ( .A(n15310), .ZN(n15309) );
  AND2_X1 U10481 ( .A1(n10114), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10587) );
  INV_X1 U10482 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15148) );
  INV_X1 U10483 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11090) );
  INV_X1 U10484 ( .A(n13130), .ZN(P3_U3897) );
  NAND2_X1 U10485 ( .A1(n8459), .A2(n6598), .ZN(P3_U3456) );
  AND2_X1 U10486 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10858), .ZN(P2_U3947) );
  INV_X2 U10487 ( .A(n14611), .ZN(P1_U4016) );
  INV_X1 U10488 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7874) );
  INV_X1 U10489 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n7875) );
  INV_X1 U10490 ( .A(n8360), .ZN(n7877) );
  INV_X1 U10491 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U10492 ( .A1(n8362), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n7878) );
  NAND2_X1 U10493 ( .A1(n13336), .A2(n7878), .ZN(n13349) );
  NOR2_X1 U10494 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n7883) );
  NOR2_X1 U10495 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), 
        .ZN(n7882) );
  NAND2_X1 U10496 ( .A1(n7967), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7893) );
  NOR2_X1 U10497 ( .A1(P3_IR_REG_29__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), 
        .ZN(n7894) );
  INV_X1 U10498 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n7900) );
  AND2_X2 U10499 ( .A1(n13694), .A2(n13697), .ZN(n8061) );
  INV_X2 U10500 ( .A(n8085), .ZN(n10269) );
  NAND2_X1 U10501 ( .A1(n10269), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7899) );
  AND2_X2 U10502 ( .A1(n7897), .A2(n13697), .ZN(n8060) );
  NAND2_X1 U10503 ( .A1(n8060), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n7898) );
  OAI211_X1 U10504 ( .C1(n8398), .C2(n7900), .A(n7899), .B(n7898), .ZN(n7901)
         );
  NAND2_X1 U10505 ( .A1(n8631), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7988) );
  INV_X1 U10506 ( .A(n7988), .ZN(n7902) );
  NAND2_X1 U10507 ( .A1(n7903), .A2(n7902), .ZN(n7979) );
  INV_X1 U10508 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U10509 ( .A1(n10588), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U10510 ( .A1(n7979), .A2(n7904), .ZN(n7997) );
  NAND2_X1 U10511 ( .A1(n10593), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7906) );
  INV_X1 U10512 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U10513 ( .A1(n10668), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7905) );
  AND2_X1 U10514 ( .A1(n7906), .A2(n7905), .ZN(n7996) );
  NAND2_X1 U10515 ( .A1(n10568), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7907) );
  NAND2_X1 U10516 ( .A1(n10566), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7910) );
  INV_X1 U10517 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10670) );
  NAND2_X1 U10518 ( .A1(n10670), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7909) );
  AND2_X1 U10519 ( .A1(n7910), .A2(n7909), .ZN(n8017) );
  NAND2_X1 U10520 ( .A1(n10592), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7912) );
  NAND2_X1 U10521 ( .A1(n10676), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U10522 ( .A1(n8051), .A2(n7912), .ZN(n8038) );
  NAND2_X1 U10523 ( .A1(n10672), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10524 ( .A1(n10571), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U10525 ( .A1(n10595), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U10526 ( .A1(n7916), .A2(n7915), .ZN(n8066) );
  NAND2_X1 U10527 ( .A1(n10654), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U10528 ( .A1(n10657), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U10529 ( .A1(n7919), .A2(n7917), .ZN(n8095) );
  INV_X1 U10530 ( .A(n8095), .ZN(n7918) );
  NAND2_X1 U10531 ( .A1(n10681), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10532 ( .A1(n10679), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U10533 ( .A1(n10690), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U10534 ( .A1(n10688), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7922) );
  NAND2_X1 U10535 ( .A1(n8112), .A2(n8111), .ZN(n7924) );
  NAND2_X1 U10536 ( .A1(n10733), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U10537 ( .A1(n8131), .A2(n7925), .ZN(n7927) );
  NAND2_X1 U10538 ( .A1(n10731), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7926) );
  XNOR2_X1 U10539 ( .A(n10795), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n8145) );
  INV_X1 U10540 ( .A(n8145), .ZN(n7928) );
  NAND2_X1 U10541 ( .A1(n10795), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7929) );
  AOI22_X1 U10542 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n10791), .B1(n15714), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10543 ( .A1(n10788), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U10544 ( .A1(n7931), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7933) );
  INV_X1 U10545 ( .A(n7931), .ZN(n7932) );
  AOI22_X1 U10546 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n7933), .B1(n7932), 
        .B2(n10998), .ZN(n7934) );
  XNOR2_X1 U10547 ( .A(n11061), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n8191) );
  INV_X1 U10548 ( .A(n8191), .ZN(n7935) );
  NAND2_X1 U10549 ( .A1(n8192), .A2(n7935), .ZN(n7937) );
  NAND2_X1 U10550 ( .A1(n11061), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7936) );
  XNOR2_X1 U10551 ( .A(n15692), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n8203) );
  INV_X1 U10552 ( .A(n8203), .ZN(n7938) );
  NAND2_X1 U10553 ( .A1(n8204), .A2(n7938), .ZN(n7940) );
  NAND2_X1 U10554 ( .A1(n15692), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7939) );
  XNOR2_X1 U10555 ( .A(n11090), .B(P1_DATAO_REG_17__SCAN_IN), .ZN(n8242) );
  INV_X1 U10556 ( .A(n8242), .ZN(n7941) );
  NAND2_X1 U10557 ( .A1(n11090), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7942) );
  XNOR2_X1 U10558 ( .A(n11442), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n8231) );
  INV_X1 U10559 ( .A(n8231), .ZN(n7944) );
  NAND2_X1 U10560 ( .A1(n11442), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7945) );
  XNOR2_X1 U10561 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .ZN(n8218) );
  INV_X1 U10562 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11586) );
  INV_X1 U10563 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11691) );
  NAND2_X1 U10564 ( .A1(n11691), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7946) );
  OAI211_X1 U10565 ( .C1(P1_DATAO_REG_20__SCAN_IN), .C2(n12933), .A(n8273), 
        .B(n7946), .ZN(n7949) );
  AND2_X1 U10566 ( .A1(n12933), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7947) );
  INV_X1 U10567 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U10568 ( .A1(n7947), .A2(n7946), .B1(P1_DATAO_REG_21__SCAN_IN), 
        .B2(n12941), .ZN(n7948) );
  INV_X1 U10569 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11898) );
  NAND2_X1 U10570 ( .A1(n11898), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U10571 ( .A1(n15674), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10572 ( .A1(n7951), .A2(n7950), .ZN(n8290) );
  INV_X1 U10573 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U10574 ( .A1(n7952), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7954) );
  INV_X1 U10575 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n15719) );
  NAND2_X1 U10576 ( .A1(n15719), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7953) );
  INV_X1 U10577 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12140) );
  INV_X1 U10578 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12143) );
  AND2_X1 U10579 ( .A1(n12386), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U10580 ( .A1(n12383), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7959) );
  AND2_X1 U10581 ( .A1(n12597), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7960) );
  INV_X1 U10582 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12738) );
  INV_X1 U10583 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n12893) );
  AND2_X1 U10584 ( .A1(n12893), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7961) );
  INV_X1 U10585 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14451) );
  NAND2_X1 U10586 ( .A1(n14451), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7962) );
  XNOR2_X1 U10587 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .ZN(n7964) );
  XNOR2_X1 U10588 ( .A(n8371), .B(n7964), .ZN(n13698) );
  NAND4_X2 U10589 ( .A1(n7972), .A2(n7971), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7973) );
  NAND2_X4 U10590 ( .A1(n7974), .A2(n7973), .ZN(n8470) );
  NAND2_X1 U10591 ( .A1(n13698), .A2(n8357), .ZN(n7976) );
  NAND2_X1 U10592 ( .A1(n6404), .A2(n10567), .ZN(n10255) );
  INV_X1 U10593 ( .A(SI_28_), .ZN(n13699) );
  OR2_X1 U10594 ( .A1(n10265), .A2(n13699), .ZN(n7975) );
  NAND2_X1 U10595 ( .A1(n7991), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7977) );
  INV_X1 U10596 ( .A(SI_1_), .ZN(n10665) );
  NAND2_X1 U10597 ( .A1(n7978), .A2(n7988), .ZN(n7980) );
  AND2_X1 U10598 ( .A1(n7980), .A2(n7979), .ZN(n10666) );
  INV_X1 U10599 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7981) );
  OR2_X1 U10600 ( .A1(n6404), .A2(n7124), .ZN(n7982) );
  NAND2_X1 U10601 ( .A1(n8363), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10602 ( .A1(n10268), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U10603 ( .A1(n8060), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U10604 ( .A1(n8061), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7983) );
  NAND4_X2 U10605 ( .A1(n7986), .A2(n7985), .A3(n7984), .A4(n7983), .ZN(n15534) );
  INV_X1 U10606 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11115) );
  INV_X1 U10607 ( .A(SI_0_), .ZN(n8632) );
  INV_X1 U10608 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U10609 ( .A1(n9567), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7987) );
  AND2_X1 U10610 ( .A1(n7988), .A2(n7987), .ZN(n7989) );
  MUX2_X1 U10611 ( .A(n8632), .B(n7989), .S(n10572), .Z(n10563) );
  MUX2_X1 U10612 ( .A(n11115), .B(n10563), .S(n6404), .Z(n12342) );
  INV_X1 U10613 ( .A(n12342), .ZN(n12085) );
  NAND2_X1 U10614 ( .A1(n15534), .A2(n12085), .ZN(n15531) );
  NAND2_X1 U10615 ( .A1(n15530), .A2(n15531), .ZN(n15529) );
  NAND2_X1 U10616 ( .A1(n15515), .A2(n15526), .ZN(n7990) );
  NAND2_X1 U10617 ( .A1(n15529), .A2(n7990), .ZN(n15512) );
  NAND2_X1 U10618 ( .A1(n10268), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10619 ( .A1(n8060), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U10620 ( .A1(n8061), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7992) );
  OAI21_X1 U10621 ( .B1(n7997), .B2(n7996), .A(n7995), .ZN(n10601) );
  OR2_X1 U10622 ( .A1(n8070), .A2(n10601), .ZN(n8001) );
  INV_X1 U10623 ( .A(n11104), .ZN(n7998) );
  OR2_X1 U10624 ( .A1(n6404), .A2(n7497), .ZN(n8000) );
  NAND2_X1 U10625 ( .A1(n15512), .A2(n15511), .ZN(n15510) );
  NAND2_X1 U10626 ( .A1(n8375), .A2(n12356), .ZN(n8005) );
  NAND2_X1 U10627 ( .A1(n10268), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8004) );
  NAND2_X1 U10628 ( .A1(n8060), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U10629 ( .A1(n8061), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8002) );
  XNOR2_X1 U10630 ( .A(n8007), .B(n8006), .ZN(n10605) );
  OR2_X1 U10631 ( .A1(n8070), .A2(n10605), .ZN(n8010) );
  INV_X1 U10632 ( .A(n8008), .ZN(n8019) );
  OR2_X1 U10633 ( .A1(n6405), .A2(n11281), .ZN(n8009) );
  NAND2_X1 U10634 ( .A1(n15514), .A2(n10452), .ZN(n10126) );
  INV_X1 U10635 ( .A(n15536), .ZN(n11724) );
  INV_X1 U10636 ( .A(n10458), .ZN(n15505) );
  NAND2_X1 U10637 ( .A1(n11724), .A2(n15505), .ZN(n11727) );
  NAND2_X1 U10638 ( .A1(n13128), .A2(n10452), .ZN(n8011) );
  NAND2_X1 U10639 ( .A1(n10268), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U10640 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8012) );
  NAND2_X1 U10641 ( .A1(n8041), .A2(n8012), .ZN(n12310) );
  NAND2_X1 U10642 ( .A1(n8375), .A2(n12310), .ZN(n8015) );
  NAND2_X1 U10643 ( .A1(n8060), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10644 ( .A1(n8061), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8013) );
  NAND4_X1 U10645 ( .A1(n8016), .A2(n8015), .A3(n8014), .A4(n8013), .ZN(n13127) );
  OR2_X1 U10646 ( .A1(n10265), .A2(SI_4_), .ZN(n8027) );
  XNOR2_X1 U10647 ( .A(n8018), .B(n8017), .ZN(n10597) );
  OR2_X1 U10648 ( .A1(n8070), .A2(n10597), .ZN(n8026) );
  NAND2_X1 U10649 ( .A1(n8021), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8020) );
  MUX2_X1 U10650 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8020), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8024) );
  INV_X1 U10651 ( .A(n8021), .ZN(n8023) );
  INV_X1 U10652 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8022) );
  NAND2_X1 U10653 ( .A1(n8023), .A2(n8022), .ZN(n8052) );
  NAND2_X1 U10654 ( .A1(n8024), .A2(n8052), .ZN(n11327) );
  INV_X1 U10655 ( .A(n11327), .ZN(n10596) );
  OR2_X1 U10656 ( .A1(n6405), .A2(n10596), .ZN(n8025) );
  XNOR2_X1 U10657 ( .A(n13127), .B(n12311), .ZN(n12306) );
  INV_X1 U10658 ( .A(n12306), .ZN(n12304) );
  NAND2_X1 U10659 ( .A1(n12307), .A2(n12304), .ZN(n8029) );
  NAND2_X1 U10660 ( .A1(n13127), .A2(n12311), .ZN(n8028) );
  NAND2_X1 U10661 ( .A1(n10268), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8034) );
  NAND2_X1 U10662 ( .A1(n8043), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8030) );
  NAND2_X1 U10663 ( .A1(n8058), .A2(n8030), .ZN(n12323) );
  NAND2_X1 U10664 ( .A1(n8375), .A2(n12323), .ZN(n8033) );
  NAND2_X1 U10665 ( .A1(n8060), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10666 ( .A1(n8061), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U10667 ( .A1(n8071), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8036) );
  INV_X1 U10668 ( .A(SI_6_), .ZN(n10573) );
  OR2_X1 U10669 ( .A1(n10265), .A2(n10573), .ZN(n8040) );
  XNOR2_X1 U10670 ( .A(n10672), .B(P1_DATAO_REG_6__SCAN_IN), .ZN(n8037) );
  XNOR2_X1 U10671 ( .A(n8038), .B(n8037), .ZN(n10574) );
  OR2_X1 U10672 ( .A1(n8070), .A2(n10574), .ZN(n8039) );
  OAI211_X1 U10673 ( .C1(n6405), .C2(n11421), .A(n8040), .B(n8039), .ZN(n12331) );
  NAND2_X1 U10674 ( .A1(n13125), .A2(n12331), .ZN(n11786) );
  NAND2_X1 U10675 ( .A1(n10268), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U10676 ( .A1(n8041), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8042) );
  NAND2_X1 U10677 ( .A1(n8043), .A2(n8042), .ZN(n12164) );
  NAND2_X1 U10678 ( .A1(n8375), .A2(n12164), .ZN(n8046) );
  NAND2_X1 U10679 ( .A1(n8060), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U10680 ( .A1(n10269), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8044) );
  NAND4_X1 U10681 ( .A1(n8047), .A2(n8046), .A3(n8045), .A4(n8044), .ZN(n13126) );
  OR2_X1 U10682 ( .A1(n8049), .A2(n8048), .ZN(n8050) );
  NAND2_X1 U10683 ( .A1(n8051), .A2(n8050), .ZN(n10599) );
  OR2_X1 U10684 ( .A1(n8070), .A2(n10599), .ZN(n8056) );
  OR2_X1 U10685 ( .A1(n10265), .A2(SI_5_), .ZN(n8055) );
  NAND2_X1 U10686 ( .A1(n8052), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8053) );
  XNOR2_X1 U10687 ( .A(n8053), .B(P3_IR_REG_5__SCAN_IN), .ZN(n11263) );
  OR2_X1 U10688 ( .A1(n6404), .A2(n11263), .ZN(n8054) );
  NAND2_X1 U10689 ( .A1(n13126), .A2(n10465), .ZN(n8057) );
  NAND2_X1 U10690 ( .A1(n11786), .A2(n8057), .ZN(n8081) );
  NAND2_X1 U10691 ( .A1(n11790), .A2(n12331), .ZN(n10151) );
  INV_X1 U10692 ( .A(n12331), .ZN(n11717) );
  NAND2_X1 U10693 ( .A1(n13125), .A2(n11717), .ZN(n10152) );
  INV_X1 U10694 ( .A(n11709), .ZN(n8078) );
  INV_X1 U10695 ( .A(n11786), .ZN(n8077) );
  NAND2_X1 U10696 ( .A1(n10268), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U10697 ( .A1(n8058), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U10698 ( .A1(n8083), .A2(n8059), .ZN(n12363) );
  NAND2_X1 U10699 ( .A1(n8363), .A2(n12363), .ZN(n8064) );
  NAND2_X1 U10700 ( .A1(n8060), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U10701 ( .A1(n8061), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8062) );
  NAND2_X1 U10702 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  AND2_X1 U10703 ( .A1(n8069), .A2(n8068), .ZN(n10603) );
  OR2_X1 U10704 ( .A1(n8070), .A2(n10603), .ZN(n8075) );
  OAI21_X1 U10705 ( .B1(n8071), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8072) );
  XNOR2_X1 U10706 ( .A(n8072), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11427) );
  OR2_X1 U10707 ( .A1(n6404), .A2(n11427), .ZN(n8073) );
  NAND2_X1 U10708 ( .A1(n12483), .A2(n12366), .ZN(n10156) );
  INV_X1 U10709 ( .A(n12366), .ZN(n12208) );
  NAND2_X1 U10710 ( .A1(n13124), .A2(n12208), .ZN(n10155) );
  NOR2_X1 U10711 ( .A1(n13126), .A2(n10465), .ZN(n11708) );
  NAND2_X1 U10712 ( .A1(n11708), .A2(n11786), .ZN(n8076) );
  OAI211_X1 U10713 ( .C1(n8078), .C2(n8077), .A(n11791), .B(n8076), .ZN(n8079)
         );
  INV_X1 U10714 ( .A(n8079), .ZN(n8080) );
  NAND2_X1 U10715 ( .A1(n13124), .A2(n12366), .ZN(n8082) );
  NAND2_X1 U10716 ( .A1(n10268), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10717 ( .A1(n8083), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8084) );
  NAND2_X1 U10718 ( .A1(n8104), .A2(n8084), .ZN(n12485) );
  NAND2_X1 U10719 ( .A1(n8375), .A2(n12485), .ZN(n8088) );
  NAND2_X1 U10720 ( .A1(n8060), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10721 ( .A1(n8364), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8086) );
  AND4_X2 U10722 ( .A1(n8089), .A2(n8088), .A3(n8087), .A4(n8086), .ZN(n13034)
         );
  INV_X1 U10723 ( .A(n8093), .ZN(n8090) );
  NAND2_X1 U10724 ( .A1(n8090), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8091) );
  MUX2_X1 U10725 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8091), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8094) );
  NAND2_X1 U10726 ( .A1(n8094), .A2(n8113), .ZN(n11914) );
  INV_X1 U10727 ( .A(n11914), .ZN(n11921) );
  AOI22_X1 U10728 ( .A1(n8246), .A2(SI_8_), .B1(n8245), .B2(n11921), .ZN(n8098) );
  XNOR2_X1 U10729 ( .A(n8096), .B(n8095), .ZN(n10575) );
  NAND2_X1 U10730 ( .A1(n10575), .A2(n8357), .ZN(n8097) );
  NAND2_X1 U10731 ( .A1(n8098), .A2(n8097), .ZN(n12480) );
  NAND2_X1 U10732 ( .A1(n13034), .A2(n12480), .ZN(n10159) );
  INV_X2 U10733 ( .A(n13034), .ZN(n12205) );
  NAND2_X1 U10734 ( .A1(n12205), .A2(n12338), .ZN(n10160) );
  NAND2_X1 U10735 ( .A1(n10159), .A2(n10160), .ZN(n11836) );
  XNOR2_X1 U10736 ( .A(n8100), .B(n8099), .ZN(n10664) );
  NAND2_X1 U10737 ( .A1(n10664), .A2(n8357), .ZN(n8103) );
  INV_X1 U10738 ( .A(SI_9_), .ZN(n10663) );
  NAND2_X1 U10739 ( .A1(n8113), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8101) );
  XNOR2_X1 U10740 ( .A(n8101), .B(n7714), .ZN(n11922) );
  AOI22_X1 U10741 ( .A1(n7420), .A2(n10663), .B1(n8245), .B2(n11922), .ZN(
        n8102) );
  NAND2_X1 U10742 ( .A1(n8103), .A2(n8102), .ZN(n8124) );
  NAND2_X1 U10743 ( .A1(n10268), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U10744 ( .A1(n8104), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U10745 ( .A1(n8118), .A2(n8105), .ZN(n13037) );
  NAND2_X1 U10746 ( .A1(n8363), .A2(n13037), .ZN(n8109) );
  NAND2_X1 U10747 ( .A1(n10270), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U10748 ( .A1(n8061), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8107) );
  NAND4_X1 U10749 ( .A1(n8110), .A2(n8109), .A3(n8108), .A4(n8107), .ZN(n13123) );
  NAND2_X1 U10750 ( .A1(n13038), .A2(n13123), .ZN(n12229) );
  NAND2_X1 U10751 ( .A1(n11836), .A2(n12229), .ZN(n8127) );
  XNOR2_X1 U10752 ( .A(n8112), .B(n8111), .ZN(n10579) );
  NAND2_X1 U10753 ( .A1(n10579), .A2(n8357), .ZN(n8117) );
  INV_X1 U10754 ( .A(SI_10_), .ZN(n10578) );
  NAND2_X1 U10755 ( .A1(n8429), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8115) );
  XNOR2_X1 U10756 ( .A(n8115), .B(n8132), .ZN(n13140) );
  AOI22_X1 U10757 ( .A1(n7420), .A2(n10578), .B1(n8245), .B2(n13140), .ZN(
        n8116) );
  NAND2_X1 U10758 ( .A1(n8117), .A2(n8116), .ZN(n12346) );
  NAND2_X1 U10759 ( .A1(n10268), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10760 ( .A1(n8118), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10761 ( .A1(n8137), .A2(n8119), .ZN(n12344) );
  NAND2_X1 U10762 ( .A1(n8363), .A2(n12344), .ZN(n8122) );
  NAND2_X1 U10763 ( .A1(n10270), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U10764 ( .A1(n10269), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8120) );
  XNOR2_X1 U10765 ( .A(n12346), .B(n13033), .ZN(n10174) );
  NOR2_X1 U10766 ( .A1(n8124), .A2(n13123), .ZN(n10166) );
  INV_X1 U10767 ( .A(n10166), .ZN(n8125) );
  NAND2_X1 U10768 ( .A1(n8124), .A2(n13123), .ZN(n10165) );
  NAND2_X1 U10769 ( .A1(n8125), .A2(n10165), .ZN(n11804) );
  NAND2_X1 U10770 ( .A1(n13034), .A2(n12338), .ZN(n11805) );
  NAND2_X1 U10771 ( .A1(n11804), .A2(n11805), .ZN(n11807) );
  NAND2_X1 U10772 ( .A1(n11807), .A2(n12229), .ZN(n8126) );
  OR2_X1 U10773 ( .A1(n12346), .A2(n13033), .ZN(n8128) );
  XNOR2_X1 U10774 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .ZN(n8130) );
  XNOR2_X1 U10775 ( .A(n8131), .B(n8130), .ZN(n10607) );
  NAND2_X1 U10776 ( .A1(n10607), .A2(n8357), .ZN(n8136) );
  NAND2_X1 U10777 ( .A1(n8114), .A2(n8132), .ZN(n8147) );
  NAND2_X1 U10778 ( .A1(n8147), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8134) );
  INV_X1 U10779 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8133) );
  XNOR2_X1 U10780 ( .A(n8134), .B(n8133), .ZN(n13155) );
  AOI22_X1 U10781 ( .A1(n8246), .A2(n10608), .B1(n8245), .B2(n13155), .ZN(
        n8135) );
  NAND2_X1 U10782 ( .A1(n8136), .A2(n8135), .ZN(n13601) );
  NAND2_X1 U10783 ( .A1(n10268), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U10784 ( .A1(n8137), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U10785 ( .A1(n6511), .A2(n8138), .ZN(n13078) );
  NAND2_X1 U10786 ( .A1(n8375), .A2(n13078), .ZN(n8141) );
  NAND2_X1 U10787 ( .A1(n10270), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U10788 ( .A1(n10269), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8139) );
  NOR2_X1 U10789 ( .A1(n13601), .A2(n13073), .ZN(n8144) );
  NAND2_X1 U10790 ( .A1(n13601), .A2(n13073), .ZN(n8143) );
  XNOR2_X1 U10791 ( .A(n8146), .B(n8145), .ZN(n10682) );
  NAND2_X1 U10792 ( .A1(n10682), .A2(n8357), .ZN(n8154) );
  NAND2_X1 U10793 ( .A1(n8149), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8148) );
  MUX2_X1 U10794 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8148), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8152) );
  INV_X1 U10795 ( .A(n8149), .ZN(n8151) );
  INV_X1 U10796 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U10797 ( .A1(n8151), .A2(n8150), .ZN(n8178) );
  NAND2_X1 U10798 ( .A1(n8152), .A2(n8178), .ZN(n13180) );
  INV_X1 U10799 ( .A(n13180), .ZN(n13189) );
  AOI22_X1 U10800 ( .A1(n8246), .A2(SI_12_), .B1(n8245), .B2(n13189), .ZN(
        n8153) );
  NAND2_X1 U10801 ( .A1(n8154), .A2(n8153), .ZN(n12988) );
  NAND2_X1 U10802 ( .A1(n10268), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10803 ( .A1(n6511), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U10804 ( .A1(n8163), .A2(n8155), .ZN(n12987) );
  NAND2_X1 U10805 ( .A1(n8363), .A2(n12987), .ZN(n8158) );
  NAND2_X1 U10806 ( .A1(n10270), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U10807 ( .A1(n10269), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8156) );
  OR2_X1 U10808 ( .A1(n12988), .A2(n13076), .ZN(n10179) );
  NAND2_X1 U10809 ( .A1(n12988), .A2(n13076), .ZN(n10180) );
  XNOR2_X1 U10810 ( .A(n8172), .B(n10791), .ZN(n10798) );
  NAND2_X1 U10811 ( .A1(n10798), .A2(n8357), .ZN(n8162) );
  NAND2_X1 U10812 ( .A1(n8178), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8160) );
  XNOR2_X1 U10813 ( .A(n8160), .B(P3_IR_REG_13__SCAN_IN), .ZN(n13213) );
  AOI22_X1 U10814 ( .A1(n8246), .A2(SI_13_), .B1(n8245), .B2(n13213), .ZN(
        n8161) );
  NAND2_X1 U10815 ( .A1(n8163), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10816 ( .A1(n8183), .A2(n8164), .ZN(n13057) );
  NAND2_X1 U10817 ( .A1(n8375), .A2(n13057), .ZN(n8168) );
  NAND2_X1 U10818 ( .A1(n10268), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U10819 ( .A1(n10270), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10820 ( .A1(n10269), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8165) );
  OR2_X1 U10821 ( .A1(n13058), .A2(n13537), .ZN(n8169) );
  NAND2_X1 U10822 ( .A1(n12565), .A2(n8169), .ZN(n8171) );
  NAND2_X1 U10823 ( .A1(n13058), .A2(n13537), .ZN(n8170) );
  NAND2_X1 U10824 ( .A1(n8172), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U10825 ( .A1(n8173), .A2(n10788), .ZN(n8174) );
  NAND2_X1 U10826 ( .A1(n8175), .A2(n8174), .ZN(n8177) );
  XNOR2_X1 U10827 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .ZN(n8176) );
  XNOR2_X1 U10828 ( .A(n8177), .B(n8176), .ZN(n10796) );
  NAND2_X1 U10829 ( .A1(n10796), .A2(n8357), .ZN(n8182) );
  INV_X1 U10830 ( .A(SI_14_), .ZN(n10797) );
  NAND2_X1 U10831 ( .A1(n8193), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8180) );
  XNOR2_X1 U10832 ( .A(n8180), .B(n8179), .ZN(n13221) );
  AOI22_X1 U10833 ( .A1(n8246), .A2(n10797), .B1(n13221), .B2(n8245), .ZN(
        n8181) );
  NAND2_X1 U10834 ( .A1(n10268), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U10835 ( .A1(n8183), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U10836 ( .A1(n8197), .A2(n8184), .ZN(n13532) );
  NAND2_X1 U10837 ( .A1(n8375), .A2(n13532), .ZN(n8187) );
  NAND2_X1 U10838 ( .A1(n10270), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U10839 ( .A1(n10269), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8185) );
  NAND4_X1 U10840 ( .A1(n8188), .A2(n8187), .A3(n8186), .A4(n8185), .ZN(n13121) );
  INV_X1 U10841 ( .A(n13121), .ZN(n13524) );
  OR2_X1 U10842 ( .A1(n13680), .A2(n13524), .ZN(n8189) );
  XNOR2_X1 U10843 ( .A(n8192), .B(n8191), .ZN(n10784) );
  NAND2_X1 U10844 ( .A1(n10784), .A2(n8357), .ZN(n8196) );
  OAI21_X1 U10845 ( .B1(n8193), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8194) );
  XNOR2_X1 U10846 ( .A(n8194), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U10847 ( .A1(n13246), .A2(n8245), .B1(n8246), .B2(SI_15_), .ZN(
        n8195) );
  NAND2_X1 U10848 ( .A1(n8197), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10849 ( .A1(n8213), .A2(n8198), .ZN(n13518) );
  NAND2_X1 U10850 ( .A1(n13518), .A2(n8375), .ZN(n8202) );
  NAND2_X1 U10851 ( .A1(n10268), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8201) );
  NAND2_X1 U10852 ( .A1(n10270), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10853 ( .A1(n10269), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8199) );
  OR2_X1 U10854 ( .A1(n13669), .A2(n13510), .ZN(n10188) );
  NAND2_X1 U10855 ( .A1(n13669), .A2(n13510), .ZN(n10195) );
  XNOR2_X1 U10856 ( .A(n8204), .B(n8203), .ZN(n10833) );
  NAND2_X1 U10857 ( .A1(n10833), .A2(n8357), .ZN(n8212) );
  INV_X1 U10858 ( .A(n8209), .ZN(n8206) );
  NAND2_X1 U10859 ( .A1(n8206), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8207) );
  MUX2_X1 U10860 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8207), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8210) );
  AOI22_X1 U10861 ( .A1(n8246), .A2(SI_16_), .B1(n8245), .B2(n13259), .ZN(
        n8211) );
  NAND2_X1 U10862 ( .A1(n8213), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U10863 ( .A1(n8249), .A2(n8214), .ZN(n13512) );
  NAND2_X1 U10864 ( .A1(n13512), .A2(n8363), .ZN(n8217) );
  AOI22_X1 U10865 ( .A1(n10268), .A2(P3_REG1_REG_16__SCAN_IN), .B1(n10270), 
        .B2(P3_REG2_REG_16__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U10866 ( .A1(n10269), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8215) );
  XNOR2_X1 U10867 ( .A(n8219), .B(n8218), .ZN(n12935) );
  NAND2_X1 U10868 ( .A1(n12935), .A2(n8357), .ZN(n8223) );
  XNOR2_X2 U10869 ( .A(n8221), .B(P3_IR_REG_19__SCAN_IN), .ZN(n13321) );
  AOI22_X1 U10870 ( .A1(n8246), .A2(n12934), .B1(n13313), .B2(n8245), .ZN(
        n8222) );
  NAND2_X1 U10871 ( .A1(n8223), .A2(n8222), .ZN(n13462) );
  NAND2_X1 U10872 ( .A1(n8238), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U10873 ( .A1(n8262), .A2(n8224), .ZN(n13475) );
  NAND2_X1 U10874 ( .A1(n13475), .A2(n8375), .ZN(n8229) );
  INV_X1 U10875 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U10876 ( .A1(n10269), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U10877 ( .A1(n10270), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8225) );
  OAI211_X1 U10878 ( .C1(n8398), .C2(n13320), .A(n8226), .B(n8225), .ZN(n8227)
         );
  INV_X1 U10879 ( .A(n8227), .ZN(n8228) );
  NAND2_X1 U10880 ( .A1(n8229), .A2(n8228), .ZN(n13488) );
  INV_X1 U10881 ( .A(n10215), .ZN(n8230) );
  NAND2_X1 U10882 ( .A1(n13462), .A2(n13488), .ZN(n10206) );
  XNOR2_X1 U10883 ( .A(n8232), .B(n8231), .ZN(n11011) );
  NAND2_X1 U10884 ( .A1(n11011), .A2(n8357), .ZN(n8236) );
  NAND2_X1 U10885 ( .A1(n8233), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8234) );
  XNOR2_X1 U10886 ( .A(n8234), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U10887 ( .A1(n8246), .A2(SI_18_), .B1(n8245), .B2(n13324), .ZN(
        n8235) );
  NAND2_X1 U10888 ( .A1(n8251), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8237) );
  NAND2_X1 U10889 ( .A1(n8238), .A2(n8237), .ZN(n13084) );
  NAND2_X1 U10890 ( .A1(n13084), .A2(n8363), .ZN(n8241) );
  AOI22_X1 U10891 ( .A1(n10268), .A2(P3_REG1_REG_18__SCAN_IN), .B1(n10270), 
        .B2(P3_REG2_REG_18__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U10892 ( .A1(n8364), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U10893 ( .A1(n13580), .A2(n13501), .ZN(n10214) );
  XNOR2_X1 U10894 ( .A(n8243), .B(n8242), .ZN(n10933) );
  NAND2_X1 U10895 ( .A1(n10933), .A2(n8357), .ZN(n8248) );
  NAND2_X1 U10896 ( .A1(n6593), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8244) );
  XNOR2_X1 U10897 ( .A(n8244), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13295) );
  AOI22_X1 U10898 ( .A1(n8246), .A2(SI_17_), .B1(n8245), .B2(n13295), .ZN(
        n8247) );
  NAND2_X1 U10899 ( .A1(n8249), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U10900 ( .A1(n8251), .A2(n8250), .ZN(n13494) );
  NAND2_X1 U10901 ( .A1(n13494), .A2(n8375), .ZN(n8254) );
  AOI22_X1 U10902 ( .A1(n10268), .A2(P3_REG1_REG_17__SCAN_IN), .B1(n10270), 
        .B2(P3_REG2_REG_17__SCAN_IN), .ZN(n8253) );
  NAND2_X1 U10903 ( .A1(n8364), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U10904 ( .A1(n13660), .A2(n13487), .ZN(n13483) );
  NAND2_X1 U10905 ( .A1(n10315), .A2(n13483), .ZN(n13464) );
  OR2_X1 U10906 ( .A1(n13660), .A2(n13511), .ZN(n10200) );
  NAND2_X1 U10907 ( .A1(n13660), .A2(n13511), .ZN(n8410) );
  OR2_X1 U10908 ( .A1(n13464), .A2(n13496), .ZN(n8256) );
  OR2_X1 U10909 ( .A1(n13580), .A2(n13469), .ZN(n8255) );
  INV_X1 U10910 ( .A(n13460), .ZN(n13467) );
  NAND2_X1 U10911 ( .A1(n13467), .A2(n13464), .ZN(n8257) );
  OAI22_X1 U10912 ( .A1(n13465), .A2(n8257), .B1(n13085), .B2(n13462), .ZN(
        n8258) );
  INV_X1 U10913 ( .A(n8258), .ZN(n8259) );
  XNOR2_X1 U10914 ( .A(n8273), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n8271) );
  XNOR2_X1 U10915 ( .A(n8271), .B(n12933), .ZN(n11554) );
  NAND2_X1 U10916 ( .A1(n11554), .A2(n8357), .ZN(n8261) );
  INV_X1 U10917 ( .A(SI_20_), .ZN(n11556) );
  OR2_X1 U10918 ( .A1(n10265), .A2(n11556), .ZN(n8260) );
  NAND2_X1 U10919 ( .A1(n8262), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10920 ( .A1(n8280), .A2(n8263), .ZN(n13448) );
  NAND2_X1 U10921 ( .A1(n13448), .A2(n8375), .ZN(n8269) );
  INV_X1 U10922 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U10923 ( .A1(n8364), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U10924 ( .A1(n8060), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8264) );
  OAI211_X1 U10925 ( .C1(n8398), .C2(n8266), .A(n8265), .B(n8264), .ZN(n8267)
         );
  INV_X1 U10926 ( .A(n8267), .ZN(n8268) );
  XNOR2_X1 U10927 ( .A(n13646), .B(n13470), .ZN(n13446) );
  INV_X1 U10928 ( .A(n13446), .ZN(n13450) );
  NAND2_X1 U10929 ( .A1(n13646), .A2(n13470), .ZN(n8270) );
  NAND2_X1 U10930 ( .A1(n13449), .A2(n8270), .ZN(n13439) );
  INV_X1 U10931 ( .A(n8271), .ZN(n8272) );
  NAND2_X1 U10932 ( .A1(n8272), .A2(n12933), .ZN(n8275) );
  NAND2_X1 U10933 ( .A1(n8273), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U10934 ( .A1(n8275), .A2(n8274), .ZN(n8277) );
  XNOR2_X1 U10935 ( .A(n12941), .B(P1_DATAO_REG_21__SCAN_IN), .ZN(n8276) );
  XNOR2_X1 U10936 ( .A(n8277), .B(n8276), .ZN(n11765) );
  NAND2_X1 U10937 ( .A1(n11765), .A2(n8357), .ZN(n8279) );
  NAND2_X1 U10938 ( .A1(n8280), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U10939 ( .A1(n8296), .A2(n8281), .ZN(n13437) );
  NAND2_X1 U10940 ( .A1(n13437), .A2(n8375), .ZN(n8286) );
  INV_X1 U10941 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13572) );
  NAND2_X1 U10942 ( .A1(n10269), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10943 ( .A1(n8060), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8282) );
  OAI211_X1 U10944 ( .C1(n8398), .C2(n13572), .A(n8283), .B(n8282), .ZN(n8284)
         );
  INV_X1 U10945 ( .A(n8284), .ZN(n8285) );
  OR2_X1 U10946 ( .A1(n13641), .A2(n13065), .ZN(n8287) );
  NAND2_X1 U10947 ( .A1(n13439), .A2(n8287), .ZN(n8289) );
  NAND2_X1 U10948 ( .A1(n13641), .A2(n13065), .ZN(n8288) );
  NAND2_X1 U10949 ( .A1(n8291), .A2(n8290), .ZN(n8292) );
  NAND2_X1 U10950 ( .A1(n8293), .A2(n8292), .ZN(n11461) );
  NAND2_X1 U10951 ( .A1(n11461), .A2(n8357), .ZN(n8295) );
  NAND2_X1 U10952 ( .A1(n8296), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U10953 ( .A1(n8312), .A2(n8297), .ZN(n13427) );
  NAND2_X1 U10954 ( .A1(n13427), .A2(n8363), .ZN(n8303) );
  INV_X1 U10955 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U10956 ( .A1(n8364), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U10957 ( .A1(n10270), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8298) );
  OAI211_X1 U10958 ( .C1(n8398), .C2(n8300), .A(n8299), .B(n8298), .ZN(n8301)
         );
  INV_X1 U10959 ( .A(n8301), .ZN(n8302) );
  AND2_X1 U10960 ( .A1(n13635), .A2(n13440), .ZN(n8305) );
  OR2_X1 U10961 ( .A1(n13635), .A2(n13440), .ZN(n8304) );
  OR2_X1 U10962 ( .A1(n8307), .A2(n8306), .ZN(n8308) );
  NAND2_X1 U10963 ( .A1(n8309), .A2(n8308), .ZN(n11782) );
  NAND2_X1 U10964 ( .A1(n11782), .A2(n8357), .ZN(n8311) );
  OR2_X1 U10965 ( .A1(n10265), .A2(n11785), .ZN(n8310) );
  NAND2_X1 U10966 ( .A1(n8312), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U10967 ( .A1(n8324), .A2(n8313), .ZN(n13415) );
  NAND2_X1 U10968 ( .A1(n13415), .A2(n8363), .ZN(n8318) );
  INV_X1 U10969 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13567) );
  NAND2_X1 U10970 ( .A1(n10269), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10971 ( .A1(n10270), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8314) );
  OAI211_X1 U10972 ( .C1(n8398), .C2(n13567), .A(n8315), .B(n8314), .ZN(n8316)
         );
  INV_X1 U10973 ( .A(n8316), .ZN(n8317) );
  AND2_X1 U10974 ( .A1(n13630), .A2(n13431), .ZN(n8411) );
  INV_X1 U10975 ( .A(n8411), .ZN(n8319) );
  XNOR2_X1 U10976 ( .A(n8320), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n12196) );
  NAND2_X1 U10977 ( .A1(n12196), .A2(n8357), .ZN(n8322) );
  INV_X1 U10978 ( .A(SI_24_), .ZN(n12197) );
  INV_X1 U10979 ( .A(n8323), .ZN(n8339) );
  NAND2_X1 U10980 ( .A1(n8324), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8325) );
  NAND2_X1 U10981 ( .A1(n8339), .A2(n8325), .ZN(n13408) );
  NAND2_X1 U10982 ( .A1(n13408), .A2(n8375), .ZN(n8331) );
  INV_X1 U10983 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U10984 ( .A1(n10268), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U10985 ( .A1(n8364), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8326) );
  OAI211_X1 U10986 ( .C1(n8106), .C2(n8328), .A(n8327), .B(n8326), .ZN(n8329)
         );
  INV_X1 U10987 ( .A(n8329), .ZN(n8330) );
  OR2_X1 U10988 ( .A1(n13565), .A2(n13119), .ZN(n8332) );
  NAND2_X1 U10989 ( .A1(n13565), .A2(n13119), .ZN(n8333) );
  XNOR2_X1 U10990 ( .A(n12386), .B(P1_DATAO_REG_25__SCAN_IN), .ZN(n8335) );
  XNOR2_X1 U10991 ( .A(n8336), .B(n8335), .ZN(n12449) );
  NAND2_X1 U10992 ( .A1(n12449), .A2(n8357), .ZN(n8338) );
  INV_X1 U10993 ( .A(SI_25_), .ZN(n12451) );
  OR2_X1 U10994 ( .A1(n10265), .A2(n12451), .ZN(n8337) );
  NAND2_X1 U10995 ( .A1(n8339), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U10996 ( .A1(n8350), .A2(n8340), .ZN(n13392) );
  NAND2_X1 U10997 ( .A1(n13392), .A2(n8375), .ZN(n8345) );
  INV_X1 U10998 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13562) );
  NAND2_X1 U10999 ( .A1(n8364), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U11000 ( .A1(n8060), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8341) );
  OAI211_X1 U11001 ( .C1(n8398), .C2(n13562), .A(n8342), .B(n8341), .ZN(n8343)
         );
  INV_X1 U11002 ( .A(n8343), .ZN(n8344) );
  NAND2_X1 U11003 ( .A1(n12992), .A2(n13404), .ZN(n10238) );
  XNOR2_X1 U11004 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .ZN(n8346) );
  XNOR2_X1 U11005 ( .A(n8347), .B(n8346), .ZN(n12559) );
  NAND2_X1 U11006 ( .A1(n12559), .A2(n8357), .ZN(n8349) );
  OR2_X1 U11007 ( .A1(n10265), .A2(n12560), .ZN(n8348) );
  NAND2_X1 U11008 ( .A1(n8350), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8351) );
  NAND2_X1 U11009 ( .A1(n8360), .A2(n8351), .ZN(n13375) );
  INV_X1 U11010 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13557) );
  NAND2_X1 U11011 ( .A1(n10269), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U11012 ( .A1(n8060), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8352) );
  OAI211_X1 U11013 ( .C1(n8398), .C2(n13557), .A(n8353), .B(n8352), .ZN(n8354)
         );
  XNOR2_X1 U11014 ( .A(n12893), .B(P1_DATAO_REG_27__SCAN_IN), .ZN(n8355) );
  XNOR2_X1 U11015 ( .A(n8356), .B(n8355), .ZN(n13702) );
  NAND2_X1 U11016 ( .A1(n13702), .A2(n8357), .ZN(n8359) );
  INV_X1 U11017 ( .A(SI_27_), .ZN(n13704) );
  OR2_X1 U11018 ( .A1(n10265), .A2(n13704), .ZN(n8358) );
  NAND2_X1 U11019 ( .A1(n8360), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U11020 ( .A1(n8362), .A2(n8361), .ZN(n13364) );
  NAND2_X1 U11021 ( .A1(n13364), .A2(n8363), .ZN(n8369) );
  INV_X1 U11022 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n15733) );
  NAND2_X1 U11023 ( .A1(n10268), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U11024 ( .A1(n8060), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8365) );
  OAI211_X1 U11025 ( .C1(n15733), .C2(n8085), .A(n8366), .B(n8365), .ZN(n8367)
         );
  INV_X1 U11026 ( .A(n8367), .ZN(n8368) );
  NAND2_X1 U11027 ( .A1(n13552), .A2(n12902), .ZN(n13347) );
  NAND2_X1 U11028 ( .A1(n13548), .A2(n13362), .ZN(n8415) );
  AND2_X1 U11029 ( .A1(n8545), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U11030 ( .A1(n15148), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8372) );
  INV_X1 U11031 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12895) );
  XNOR2_X1 U11032 ( .A(n12895), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n10252) );
  XNOR2_X1 U11033 ( .A(n10254), .B(n10252), .ZN(n13695) );
  NAND2_X1 U11034 ( .A1(n13695), .A2(n8357), .ZN(n8374) );
  INV_X1 U11035 ( .A(SI_29_), .ZN(n15690) );
  OR2_X1 U11036 ( .A1(n10265), .A2(n15690), .ZN(n8373) );
  NAND2_X2 U11037 ( .A1(n8374), .A2(n8373), .ZN(n10259) );
  INV_X1 U11038 ( .A(n13336), .ZN(n8376) );
  NAND2_X1 U11039 ( .A1(n8376), .A2(n8375), .ZN(n10275) );
  INV_X1 U11040 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n15671) );
  NAND2_X1 U11041 ( .A1(n10268), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U11042 ( .A1(n8060), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8377) );
  OAI211_X1 U11043 ( .C1(n8085), .C2(n15671), .A(n8378), .B(n8377), .ZN(n8379)
         );
  INV_X1 U11044 ( .A(n8379), .ZN(n8380) );
  NAND2_X1 U11045 ( .A1(n10275), .A2(n8380), .ZN(n13354) );
  XNOR2_X1 U11046 ( .A(n10259), .B(n13354), .ZN(n10323) );
  NAND2_X1 U11047 ( .A1(n8421), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U11048 ( .A1(n10338), .A2(n13321), .ZN(n10336) );
  INV_X1 U11049 ( .A(n8386), .ZN(n8387) );
  NAND2_X1 U11050 ( .A1(n8387), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8388) );
  INV_X1 U11051 ( .A(n11555), .ZN(n8392) );
  NAND2_X1 U11052 ( .A1(n11704), .A2(n8392), .ZN(n10290) );
  INV_X4 U11053 ( .A(n13214), .ZN(n13703) );
  INV_X1 U11054 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U11055 ( .A1(n10269), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U11056 ( .A1(n10270), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8395) );
  OAI211_X1 U11057 ( .C1(n8398), .C2(n8397), .A(n8396), .B(n8395), .ZN(n8399)
         );
  INV_X1 U11058 ( .A(n8399), .ZN(n8400) );
  NAND2_X1 U11059 ( .A1(n10275), .A2(n8400), .ZN(n12619) );
  INV_X1 U11060 ( .A(P3_B_REG_SCAN_IN), .ZN(n8401) );
  NOR2_X1 U11061 ( .A1(n13701), .A2(n8401), .ZN(n8402) );
  NOR2_X1 U11062 ( .A1(n15513), .A2(n8402), .ZN(n13333) );
  NAND2_X1 U11063 ( .A1(n10453), .A2(n10455), .ZN(n15504) );
  NAND2_X1 U11064 ( .A1(n11724), .A2(n10458), .ZN(n10125) );
  NAND2_X1 U11065 ( .A1(n11723), .A2(n11722), .ZN(n11721) );
  NAND2_X1 U11066 ( .A1(n11721), .A2(n10126), .ZN(n12305) );
  NAND2_X1 U11067 ( .A1(n12305), .A2(n12306), .ZN(n8407) );
  INV_X1 U11068 ( .A(n13127), .ZN(n12355) );
  NAND2_X1 U11069 ( .A1(n12355), .A2(n12311), .ZN(n8406) );
  NAND2_X1 U11070 ( .A1(n8407), .A2(n8406), .ZN(n12162) );
  NAND2_X1 U11071 ( .A1(n12162), .A2(n12167), .ZN(n8408) );
  INV_X1 U11072 ( .A(n13126), .ZN(n12328) );
  NAND2_X1 U11073 ( .A1(n12328), .A2(n10465), .ZN(n10147) );
  NAND2_X1 U11074 ( .A1(n8408), .A2(n10147), .ZN(n11692) );
  AND2_X1 U11075 ( .A1(n12346), .A2(n13122), .ZN(n10170) );
  XNOR2_X1 U11076 ( .A(n13601), .B(n13073), .ZN(n12491) );
  NAND2_X1 U11077 ( .A1(n12492), .A2(n12491), .ZN(n12490) );
  INV_X1 U11078 ( .A(n13601), .ZN(n12495) );
  NAND2_X1 U11079 ( .A1(n12495), .A2(n13073), .ZN(n10176) );
  NAND2_X1 U11080 ( .A1(n12490), .A2(n10176), .ZN(n12467) );
  INV_X1 U11081 ( .A(n10180), .ZN(n8409) );
  NAND2_X1 U11082 ( .A1(n13058), .A2(n12948), .ZN(n10185) );
  NOR2_X1 U11083 ( .A1(n13058), .A2(n12948), .ZN(n10190) );
  XNOR2_X1 U11084 ( .A(n13585), .B(n13525), .ZN(n13507) );
  NAND2_X1 U11085 ( .A1(n13585), .A2(n13525), .ZN(n10196) );
  INV_X1 U11086 ( .A(n8410), .ZN(n10204) );
  AND2_X1 U11087 ( .A1(n10206), .A2(n13459), .ZN(n10203) );
  INV_X1 U11088 ( .A(n13646), .ZN(n10216) );
  NAND2_X1 U11089 ( .A1(n10216), .A2(n13470), .ZN(n10217) );
  NAND2_X1 U11090 ( .A1(n13641), .A2(n13454), .ZN(n10225) );
  NOR2_X1 U11091 ( .A1(n13641), .A2(n13454), .ZN(n10222) );
  AOI21_X2 U11092 ( .B1(n13426), .B2(n10210), .A(n10208), .ZN(n13414) );
  NAND2_X1 U11093 ( .A1(n13565), .A2(n13419), .ZN(n13383) );
  NAND2_X1 U11094 ( .A1(n10231), .A2(n8411), .ZN(n8412) );
  NAND3_X1 U11095 ( .A1(n10238), .A2(n13383), .A3(n8412), .ZN(n8413) );
  INV_X1 U11096 ( .A(n8413), .ZN(n13370) );
  AND2_X1 U11097 ( .A1(n10231), .A2(n13398), .ZN(n13369) );
  OR2_X1 U11098 ( .A1(n13615), .A2(n13387), .ZN(n10237) );
  OAI211_X1 U11099 ( .C1(n8413), .C2(n13369), .A(n10237), .B(n13372), .ZN(
        n8414) );
  XNOR2_X1 U11100 ( .A(n10281), .B(n10323), .ZN(n13346) );
  AND2_X1 U11101 ( .A1(n11766), .A2(n11555), .ZN(n10337) );
  INV_X1 U11102 ( .A(n10337), .ZN(n8416) );
  XNOR2_X1 U11103 ( .A(n10338), .B(n8416), .ZN(n8418) );
  NAND2_X1 U11104 ( .A1(n11766), .A2(n13313), .ZN(n8417) );
  AND2_X1 U11105 ( .A1(n15567), .A2(n10531), .ZN(n8419) );
  NAND2_X1 U11106 ( .A1(n10529), .A2(n8419), .ZN(n8420) );
  NAND2_X1 U11107 ( .A1(n11459), .A2(n15507), .ZN(n13555) );
  AND2_X1 U11108 ( .A1(n15521), .A2(n13555), .ZN(n12227) );
  NAND2_X1 U11109 ( .A1(n8426), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8424) );
  MUX2_X1 U11110 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8425), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8427) );
  AND2_X1 U11111 ( .A1(n8427), .A2(n8426), .ZN(n8434) );
  NAND2_X1 U11112 ( .A1(n8440), .A2(n8434), .ZN(n8433) );
  OAI21_X1 U11113 ( .B1(n8429), .B2(n8428), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8430) );
  MUX2_X1 U11114 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8430), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8432) );
  NAND2_X1 U11115 ( .A1(n8432), .A2(n8431), .ZN(n12199) );
  OAI21_X1 U11116 ( .B1(n11098), .B2(n10524), .A(n10538), .ZN(n8452) );
  XNOR2_X1 U11117 ( .A(n12199), .B(P3_B_REG_SCAN_IN), .ZN(n8435) );
  INV_X1 U11118 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U11119 ( .A1(n10801), .A2(n8436), .ZN(n8438) );
  INV_X1 U11120 ( .A(n8440), .ZN(n12562) );
  NAND2_X1 U11121 ( .A1(n12562), .A2(n12452), .ZN(n8437) );
  INV_X1 U11122 ( .A(n12199), .ZN(n8439) );
  NOR2_X1 U11123 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .ZN(
        n8445) );
  NOR4_X1 U11124 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n8444) );
  NOR4_X1 U11125 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n8443) );
  NOR4_X1 U11126 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8442) );
  NAND4_X1 U11127 ( .A1(n8445), .A2(n8444), .A3(n8443), .A4(n8442), .ZN(n8451)
         );
  NOR4_X1 U11128 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8449) );
  NOR4_X1 U11129 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8448) );
  NOR4_X1 U11130 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8447) );
  NOR4_X1 U11131 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8446) );
  NAND4_X1 U11132 ( .A1(n8449), .A2(n8448), .A3(n8447), .A4(n8446), .ZN(n8450)
         );
  OAI21_X1 U11133 ( .B1(n8451), .B2(n8450), .A(n10801), .ZN(n10345) );
  INV_X1 U11134 ( .A(n10345), .ZN(n8453) );
  NAND2_X1 U11135 ( .A1(n8452), .A2(n10527), .ZN(n8456) );
  INV_X1 U11136 ( .A(n10529), .ZN(n8454) );
  NAND2_X1 U11137 ( .A1(n10610), .A2(n11697), .ZN(n10346) );
  OR3_X1 U11138 ( .A1(n8454), .A2(n11098), .A3(n10525), .ZN(n8455) );
  NAND2_X1 U11139 ( .A1(n10259), .A2(n13670), .ZN(n8458) );
  MUX2_X1 U11140 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n10572), .Z(n9124) );
  AND2_X1 U11141 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8461) );
  NAND2_X1 U11142 ( .A1(n8470), .A2(n8461), .ZN(n9569) );
  NAND2_X1 U11143 ( .A1(n8470), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8462) );
  OAI211_X1 U11144 ( .C1(n8470), .C2(n10588), .A(n8462), .B(n10665), .ZN(n8463) );
  NAND2_X1 U11145 ( .A1(n8470), .A2(n10569), .ZN(n8464) );
  INV_X1 U11146 ( .A(n8466), .ZN(n8467) );
  NAND2_X1 U11147 ( .A1(n8467), .A2(SI_2_), .ZN(n8468) );
  INV_X1 U11148 ( .A(n8685), .ZN(n8471) );
  NAND2_X1 U11149 ( .A1(n8472), .A2(SI_3_), .ZN(n8473) );
  INV_X1 U11150 ( .A(n8713), .ZN(n8474) );
  NAND2_X1 U11151 ( .A1(n8475), .A2(SI_4_), .ZN(n8476) );
  XNOR2_X1 U11152 ( .A(n8478), .B(SI_5_), .ZN(n8725) );
  INV_X1 U11153 ( .A(n8725), .ZN(n8477) );
  NAND2_X1 U11154 ( .A1(n8478), .A2(SI_5_), .ZN(n8479) );
  XNOR2_X1 U11155 ( .A(n8482), .B(SI_6_), .ZN(n8751) );
  INV_X1 U11156 ( .A(n8751), .ZN(n8481) );
  NAND2_X1 U11157 ( .A1(n8482), .A2(SI_6_), .ZN(n8483) );
  XNOR2_X1 U11158 ( .A(n8485), .B(SI_7_), .ZN(n8770) );
  INV_X1 U11159 ( .A(n8770), .ZN(n8484) );
  XNOR2_X1 U11160 ( .A(n8487), .B(SI_8_), .ZN(n8787) );
  INV_X1 U11161 ( .A(n8787), .ZN(n8486) );
  NAND2_X1 U11162 ( .A1(n8487), .A2(SI_8_), .ZN(n8488) );
  MUX2_X1 U11163 ( .A(n10679), .B(n10681), .S(n10572), .Z(n8489) );
  XNOR2_X1 U11164 ( .A(n8489), .B(SI_9_), .ZN(n8808) );
  INV_X1 U11165 ( .A(n8489), .ZN(n8490) );
  NAND2_X1 U11166 ( .A1(n8490), .A2(SI_9_), .ZN(n8491) );
  XNOR2_X1 U11167 ( .A(n8494), .B(SI_10_), .ZN(n8830) );
  INV_X1 U11168 ( .A(n8830), .ZN(n8493) );
  NAND2_X1 U11169 ( .A1(n8494), .A2(SI_10_), .ZN(n8851) );
  NAND2_X1 U11170 ( .A1(n8495), .A2(n10608), .ZN(n8866) );
  INV_X1 U11171 ( .A(n8866), .ZN(n8498) );
  INV_X1 U11172 ( .A(n8496), .ZN(n8497) );
  AOI21_X1 U11173 ( .B1(n8869), .B2(n8498), .A(n8497), .ZN(n8499) );
  MUX2_X1 U11174 ( .A(n10791), .B(n10788), .S(n10572), .Z(n8500) );
  NAND2_X1 U11175 ( .A1(n8500), .A2(n10800), .ZN(n8503) );
  INV_X1 U11176 ( .A(n8500), .ZN(n8501) );
  NAND2_X1 U11177 ( .A1(n8501), .A2(SI_13_), .ZN(n8502) );
  NOR2_X1 U11178 ( .A1(n8936), .A2(SI_14_), .ZN(n8508) );
  NAND2_X1 U11179 ( .A1(n8504), .A2(n10786), .ZN(n8509) );
  INV_X1 U11180 ( .A(n8504), .ZN(n8505) );
  NAND2_X1 U11181 ( .A1(n8505), .A2(SI_15_), .ZN(n8506) );
  NAND2_X1 U11182 ( .A1(n8936), .A2(SI_14_), .ZN(n8507) );
  NAND2_X1 U11183 ( .A1(n8510), .A2(n8509), .ZN(n8961) );
  MUX2_X1 U11184 ( .A(n10994), .B(n15692), .S(n10572), .Z(n8511) );
  NAND2_X1 U11185 ( .A1(n8511), .A2(n10835), .ZN(n8514) );
  INV_X1 U11186 ( .A(n8511), .ZN(n8512) );
  NAND2_X1 U11187 ( .A1(n8512), .A2(SI_16_), .ZN(n8513) );
  INV_X1 U11188 ( .A(n8516), .ZN(n8517) );
  NAND2_X1 U11189 ( .A1(n8517), .A2(SI_17_), .ZN(n8518) );
  NAND2_X1 U11190 ( .A1(n8523), .A2(SI_19_), .ZN(n9026) );
  MUX2_X1 U11191 ( .A(n11443), .B(n11442), .S(n10572), .Z(n9004) );
  INV_X1 U11192 ( .A(n9004), .ZN(n9021) );
  NAND2_X1 U11193 ( .A1(n9021), .A2(SI_18_), .ZN(n8521) );
  NAND3_X1 U11194 ( .A1(n9026), .A2(n11013), .A3(n9004), .ZN(n8525) );
  INV_X1 U11195 ( .A(n8523), .ZN(n8524) );
  NAND2_X1 U11196 ( .A1(n8524), .A2(n12934), .ZN(n9025) );
  MUX2_X1 U11197 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n10572), .Z(n9141) );
  INV_X1 U11198 ( .A(n9141), .ZN(n8527) );
  NAND2_X1 U11199 ( .A1(n8527), .A2(n11767), .ZN(n8528) );
  OAI21_X1 U11200 ( .B1(n9136), .B2(SI_20_), .A(n8528), .ZN(n8531) );
  AOI22_X1 U11201 ( .A1(n8529), .A2(n8528), .B1(n9141), .B2(SI_21_), .ZN(n8530) );
  INV_X1 U11202 ( .A(n9108), .ZN(n8532) );
  NAND2_X1 U11203 ( .A1(n8532), .A2(n11785), .ZN(n8533) );
  AND2_X1 U11204 ( .A1(n9124), .A2(SI_22_), .ZN(n8534) );
  AOI22_X1 U11205 ( .A1(n8534), .A2(n8533), .B1(n9108), .B2(SI_23_), .ZN(n8535) );
  MUX2_X1 U11206 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n10572), .Z(n9090) );
  NAND2_X1 U11207 ( .A1(n8536), .A2(SI_24_), .ZN(n8537) );
  NAND2_X1 U11208 ( .A1(n8538), .A2(n12451), .ZN(n8541) );
  INV_X1 U11209 ( .A(n8538), .ZN(n8539) );
  NAND2_X1 U11210 ( .A1(n8539), .A2(SI_25_), .ZN(n8540) );
  NAND2_X1 U11211 ( .A1(n8541), .A2(n8540), .ZN(n9075) );
  MUX2_X1 U11212 ( .A(n14451), .B(n12893), .S(n10572), .Z(n9179) );
  NAND2_X1 U11213 ( .A1(n8542), .A2(SI_27_), .ZN(n8543) );
  NAND2_X1 U11214 ( .A1(n8546), .A2(n13699), .ZN(n8550) );
  INV_X1 U11215 ( .A(n8546), .ZN(n8547) );
  NAND2_X1 U11216 ( .A1(n8547), .A2(SI_28_), .ZN(n8548) );
  NAND2_X1 U11217 ( .A1(n8550), .A2(n8548), .ZN(n9224) );
  INV_X1 U11218 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12938) );
  MUX2_X1 U11219 ( .A(n12938), .B(n12895), .S(n10572), .Z(n8551) );
  XNOR2_X1 U11220 ( .A(n8551), .B(SI_29_), .ZN(n9212) );
  NAND2_X1 U11221 ( .A1(n9213), .A2(n9212), .ZN(n8553) );
  NAND2_X1 U11222 ( .A1(n8551), .A2(n15690), .ZN(n8552) );
  NAND2_X1 U11223 ( .A1(n8554), .A2(SI_30_), .ZN(n9206) );
  INV_X1 U11224 ( .A(n8554), .ZN(n8555) );
  INV_X1 U11225 ( .A(SI_30_), .ZN(n13693) );
  NAND2_X1 U11226 ( .A1(n8555), .A2(n13693), .ZN(n8556) );
  NAND2_X1 U11227 ( .A1(n9206), .A2(n8556), .ZN(n8557) );
  NAND2_X1 U11228 ( .A1(n8558), .A2(n8557), .ZN(n8559) );
  NOR2_X1 U11229 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n8560) );
  NAND2_X1 U11230 ( .A1(n8586), .A2(n8560), .ZN(n8561) );
  INV_X2 U11231 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9323) );
  NAND4_X1 U11232 ( .A1(n8604), .A2(n8591), .A3(n8600), .A4(n9323), .ZN(n9308)
         );
  NOR2_X1 U11233 ( .A1(n8561), .A2(n9308), .ZN(n8575) );
  NOR2_X2 U11234 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8563) );
  NOR2_X2 U11235 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8562) );
  INV_X1 U11236 ( .A(n8584), .ZN(n8566) );
  INV_X1 U11237 ( .A(n8587), .ZN(n8567) );
  NOR2_X2 U11238 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n8585) );
  NOR2_X2 U11239 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8583) );
  NAND2_X1 U11240 ( .A1(n8585), .A2(n8583), .ZN(n8571) );
  NAND4_X1 U11241 ( .A1(n8575), .A2(n8574), .A3(n8573), .A4(n8572), .ZN(n8579)
         );
  INV_X1 U11242 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8576) );
  AND2_X2 U11243 ( .A1(n6408), .A2(n10572), .ZN(n8687) );
  NAND2_X1 U11244 ( .A1(n9125), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8581) );
  INV_X1 U11245 ( .A(n8601), .ZN(n8593) );
  NAND2_X1 U11246 ( .A1(n9313), .A2(n9311), .ZN(n9005) );
  NAND2_X1 U11247 ( .A1(n8603), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U11248 ( .A1(n14286), .A2(n9131), .ZN(n8621) );
  INV_X1 U11249 ( .A(n8624), .ZN(n12741) );
  OR2_X2 U11250 ( .A1(n8609), .A2(n14440), .ZN(n8610) );
  INV_X1 U11251 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14389) );
  INV_X1 U11252 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n14036) );
  OR2_X1 U11253 ( .A1(n8924), .A2(n14036), .ZN(n8611) );
  OAI211_X1 U11254 ( .C1(n8950), .C2(n14389), .A(n8612), .B(n8611), .ZN(n13928) );
  NAND2_X1 U11255 ( .A1(n9194), .A2(n13928), .ZN(n9266) );
  INV_X1 U11256 ( .A(n11896), .ZN(n9332) );
  NAND2_X1 U11257 ( .A1(n9332), .A2(n14031), .ZN(n10434) );
  INV_X1 U11258 ( .A(n10434), .ZN(n8613) );
  NAND2_X1 U11259 ( .A1(n8613), .A2(n11662), .ZN(n9300) );
  NAND2_X1 U11260 ( .A1(n11587), .A2(n11662), .ZN(n9497) );
  NAND4_X1 U11261 ( .A1(n9266), .A2(n9300), .A3(n8614), .A4(n9497), .ZN(n8619)
         );
  INV_X1 U11262 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14289) );
  OR2_X1 U11263 ( .A1(n8948), .A2(n14289), .ZN(n8618) );
  INV_X1 U11264 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n14044) );
  OR2_X1 U11265 ( .A1(n8924), .A2(n14044), .ZN(n8617) );
  INV_X1 U11266 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14392) );
  OR2_X1 U11267 ( .A1(n8950), .A2(n14392), .ZN(n8616) );
  AND3_X1 U11268 ( .A1(n8618), .A2(n8617), .A3(n8616), .ZN(n12918) );
  INV_X1 U11269 ( .A(n12918), .ZN(n13929) );
  NAND2_X1 U11270 ( .A1(n8619), .A2(n13929), .ZN(n8620) );
  NAND2_X1 U11271 ( .A1(n8621), .A2(n8620), .ZN(n9256) );
  INV_X1 U11272 ( .A(n9256), .ZN(n9265) );
  INV_X2 U11273 ( .A(n6410), .ZN(n8693) );
  CLKBUF_X3 U11274 ( .A(n8693), .Z(n9194) );
  NOR2_X1 U11275 ( .A1(n12918), .A2(n9194), .ZN(n8622) );
  AOI21_X1 U11276 ( .B1(n14286), .B2(n9194), .A(n8622), .ZN(n9257) );
  INV_X1 U11277 ( .A(n9257), .ZN(n9264) );
  NAND2_X1 U11278 ( .A1(n8706), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U11279 ( .A1(n8676), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8629) );
  INV_X1 U11280 ( .A(n8675), .ZN(n8627) );
  NAND2_X1 U11281 ( .A1(n8627), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U11282 ( .A1(n11896), .A2(n14031), .ZN(n8630) );
  NAND2_X1 U11283 ( .A1(n8630), .A2(n9337), .ZN(n8637) );
  INV_X1 U11284 ( .A(n15321), .ZN(n8634) );
  OAI21_X1 U11285 ( .B1(n10572), .B2(n8632), .A(n8631), .ZN(n8633) );
  NAND3_X1 U11286 ( .A1(n8965), .A2(n13954), .A3(n8636), .ZN(n8641) );
  NAND4_X1 U11287 ( .A1(n8638), .A2(n6517), .A3(n11407), .A4(n8637), .ZN(n8639) );
  AND2_X1 U11288 ( .A1(n8639), .A2(n6487), .ZN(n8640) );
  NAND2_X1 U11289 ( .A1(n8687), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8647) );
  XNOR2_X1 U11290 ( .A(n8642), .B(SI_1_), .ZN(n8644) );
  NAND2_X1 U11291 ( .A1(n9214), .A2(n9574), .ZN(n8646) );
  INV_X4 U11292 ( .A(n8690), .ZN(n10854) );
  INV_X1 U11293 ( .A(n8662), .ZN(n8659) );
  INV_X1 U11294 ( .A(n15322), .ZN(n10873) );
  NAND2_X1 U11295 ( .A1(n8676), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8651) );
  INV_X1 U11296 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n14281) );
  INV_X1 U11297 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U11298 ( .A1(n8693), .A2(n7158), .ZN(n8652) );
  INV_X1 U11299 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10863) );
  OR2_X1 U11300 ( .A1(n8673), .A2(n10863), .ZN(n8656) );
  INV_X1 U11301 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11614) );
  INV_X1 U11302 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8653) );
  OR2_X1 U11303 ( .A1(n8675), .A2(n8653), .ZN(n8654) );
  NAND2_X1 U11304 ( .A1(n6412), .A2(n13952), .ZN(n8668) );
  NAND2_X1 U11305 ( .A1(n8687), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8665) );
  NAND2_X1 U11306 ( .A1(n8659), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8660) );
  MUX2_X1 U11307 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8660), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n8663) );
  INV_X1 U11308 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U11309 ( .A1(n8662), .A2(n8661), .ZN(n8683) );
  INV_X1 U11310 ( .A(n15341), .ZN(n10875) );
  NAND2_X1 U11311 ( .A1(n10854), .A2(n10875), .ZN(n8664) );
  NAND2_X1 U11312 ( .A1(n8965), .A2(n11619), .ZN(n8667) );
  NAND2_X1 U11313 ( .A1(n8965), .A2(n13952), .ZN(n8669) );
  OAI22_X1 U11314 ( .A1(n8672), .A2(n8671), .B1(n8695), .B2(n8696), .ZN(n8699)
         );
  AOI22_X1 U11315 ( .A1(n6412), .A2(n7158), .B1(n8965), .B2(n14277), .ZN(n8670) );
  AOI21_X1 U11316 ( .B1(n8672), .B2(n8671), .A(n8670), .ZN(n8698) );
  INV_X1 U11317 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10865) );
  INV_X1 U11318 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U11319 ( .A1(n8676), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U11320 ( .A1(n6411), .A2(n13951), .ZN(n8692) );
  NAND2_X1 U11321 ( .A1(n8683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8682) );
  MUX2_X1 U11322 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8682), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8684) );
  NAND2_X1 U11323 ( .A1(n10564), .A2(n9214), .ZN(n8689) );
  NAND2_X1 U11324 ( .A1(n8687), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8688) );
  OAI211_X1 U11325 ( .C1(n8690), .C2(n10877), .A(n8689), .B(n8688), .ZN(n10391) );
  NAND2_X1 U11326 ( .A1(n8965), .A2(n10391), .ZN(n8691) );
  AND2_X1 U11327 ( .A1(n8692), .A2(n8691), .ZN(n8701) );
  NAND2_X1 U11328 ( .A1(n8693), .A2(n13951), .ZN(n8694) );
  OAI21_X1 U11329 ( .B1(n8965), .B2(n11414), .A(n8694), .ZN(n8700) );
  INV_X1 U11330 ( .A(n8700), .ZN(n8703) );
  INV_X1 U11331 ( .A(n8701), .ZN(n8702) );
  NAND2_X1 U11332 ( .A1(n8703), .A2(n8702), .ZN(n8704) );
  NAND2_X1 U11333 ( .A1(n8705), .A2(n8704), .ZN(n8722) );
  BUF_X2 U11334 ( .A(n8706), .Z(n9235) );
  NAND2_X1 U11335 ( .A1(n9235), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8712) );
  INV_X1 U11336 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8707) );
  OR2_X1 U11337 ( .A1(n8950), .A2(n8707), .ZN(n8711) );
  NAND2_X1 U11338 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8733) );
  OAI21_X1 U11339 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8733), .ZN(n11655) );
  OR2_X1 U11340 ( .A1(n9234), .A2(n11655), .ZN(n8710) );
  INV_X1 U11341 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U11342 ( .A1(n6412), .A2(n13950), .ZN(n8719) );
  XNOR2_X1 U11343 ( .A(n8713), .B(n8714), .ZN(n10565) );
  NAND2_X1 U11344 ( .A1(n10565), .A2(n9214), .ZN(n8717) );
  NAND2_X1 U11345 ( .A1(n8726), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8715) );
  AOI22_X1 U11346 ( .A1(n8687), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10854), 
        .B2(n10896), .ZN(n8716) );
  NAND2_X1 U11347 ( .A1(n8693), .A2(n15478), .ZN(n8718) );
  NAND2_X1 U11348 ( .A1(n8719), .A2(n8718), .ZN(n8723) );
  NAND2_X1 U11349 ( .A1(n8693), .A2(n13950), .ZN(n8720) );
  OAI21_X1 U11350 ( .B1(n11656), .B2(n8965), .A(n8720), .ZN(n8721) );
  INV_X1 U11351 ( .A(n8723), .ZN(n8724) );
  NAND2_X1 U11352 ( .A1(n10590), .A2(n9228), .ZN(n8730) );
  OAI21_X1 U11353 ( .B1(n8726), .B2(P2_IR_REG_4__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8727) );
  MUX2_X1 U11354 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8727), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8728) );
  INV_X1 U11355 ( .A(n9311), .ZN(n8871) );
  AND2_X1 U11356 ( .A1(n8728), .A2(n8871), .ZN(n13964) );
  AOI22_X1 U11357 ( .A1(n9125), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10854), 
        .B2(n13964), .ZN(n8729) );
  NAND2_X1 U11358 ( .A1(n8730), .A2(n8729), .ZN(n13821) );
  NAND2_X1 U11359 ( .A1(n13821), .A2(n9131), .ZN(n8741) );
  NAND2_X1 U11360 ( .A1(n6407), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8739) );
  INV_X1 U11361 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10885) );
  OR2_X1 U11362 ( .A1(n8924), .A2(n10885), .ZN(n8738) );
  INV_X1 U11363 ( .A(n8733), .ZN(n8731) );
  NAND2_X1 U11364 ( .A1(n8731), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8758) );
  INV_X1 U11365 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11366 ( .A1(n8733), .A2(n8732), .ZN(n8734) );
  NAND2_X1 U11367 ( .A1(n8758), .A2(n8734), .ZN(n13819) );
  OR2_X1 U11368 ( .A1(n9234), .A2(n13819), .ZN(n8737) );
  INV_X1 U11369 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8735) );
  OR2_X1 U11370 ( .A1(n8948), .A2(n8735), .ZN(n8736) );
  NAND2_X1 U11371 ( .A1(n9194), .A2(n13949), .ZN(n8740) );
  NAND2_X1 U11372 ( .A1(n8741), .A2(n8740), .ZN(n8746) );
  INV_X1 U11373 ( .A(n13949), .ZN(n11645) );
  NAND2_X1 U11374 ( .A1(n13821), .A2(n9244), .ZN(n8742) );
  OAI21_X1 U11375 ( .B1(n11645), .B2(n9194), .A(n8742), .ZN(n8743) );
  NAND2_X1 U11376 ( .A1(n8744), .A2(n8743), .ZN(n8750) );
  INV_X1 U11377 ( .A(n8745), .ZN(n8748) );
  INV_X1 U11378 ( .A(n8746), .ZN(n8747) );
  NAND2_X1 U11379 ( .A1(n8748), .A2(n8747), .ZN(n8749) );
  XNOR2_X1 U11380 ( .A(n8752), .B(n8751), .ZN(n10570) );
  NAND2_X1 U11381 ( .A1(n10570), .A2(n9228), .ZN(n8755) );
  NAND2_X1 U11382 ( .A1(n8871), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8753) );
  XNOR2_X1 U11383 ( .A(n8753), .B(P2_IR_REG_6__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U11384 ( .A1(n9125), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10854), 
        .B2(n11039), .ZN(n8754) );
  NAND2_X1 U11385 ( .A1(n8755), .A2(n8754), .ZN(n11856) );
  NAND2_X1 U11386 ( .A1(n11856), .A2(n9194), .ZN(n8766) );
  NAND2_X1 U11387 ( .A1(n6407), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8764) );
  INV_X1 U11388 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10888) );
  OR2_X1 U11389 ( .A1(n8924), .A2(n10888), .ZN(n8763) );
  INV_X1 U11390 ( .A(n8758), .ZN(n8756) );
  NAND2_X1 U11391 ( .A1(n8756), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8777) );
  INV_X1 U11392 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U11393 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  NAND2_X1 U11394 ( .A1(n8777), .A2(n8759), .ZN(n11854) );
  OR2_X1 U11395 ( .A1(n9234), .A2(n11854), .ZN(n8762) );
  INV_X1 U11396 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8760) );
  OR2_X1 U11397 ( .A1(n8948), .A2(n8760), .ZN(n8761) );
  NAND2_X1 U11398 ( .A1(n9131), .A2(n13948), .ZN(n8765) );
  NAND2_X1 U11399 ( .A1(n8766), .A2(n8765), .ZN(n8768) );
  AOI22_X1 U11400 ( .A1(n11856), .A2(n9131), .B1(n13948), .B2(n9194), .ZN(
        n8767) );
  XNOR2_X1 U11401 ( .A(n8771), .B(n8770), .ZN(n10594) );
  NAND2_X1 U11402 ( .A1(n10594), .A2(n9228), .ZN(n8774) );
  NAND2_X1 U11403 ( .A1(n8789), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8772) );
  XNOR2_X1 U11404 ( .A(n8772), .B(P2_IR_REG_7__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U11405 ( .A1(n9125), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10854), 
        .B2(n11042), .ZN(n8773) );
  NAND2_X2 U11406 ( .A1(n8774), .A2(n8773), .ZN(n11844) );
  NAND2_X1 U11407 ( .A1(n11844), .A2(n9131), .ZN(n8784) );
  NAND2_X1 U11408 ( .A1(n6407), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8782) );
  INV_X1 U11409 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11775) );
  OR2_X1 U11410 ( .A1(n8924), .A2(n11775), .ZN(n8781) );
  INV_X1 U11411 ( .A(n8777), .ZN(n8775) );
  INV_X1 U11412 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11413 ( .A1(n8777), .A2(n8776), .ZN(n8778) );
  NAND2_X1 U11414 ( .A1(n8816), .A2(n8778), .ZN(n11797) );
  OR2_X1 U11415 ( .A1(n9234), .A2(n11797), .ZN(n8780) );
  INV_X1 U11416 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11030) );
  OR2_X1 U11417 ( .A1(n8948), .A2(n11030), .ZN(n8779) );
  NAND2_X1 U11418 ( .A1(n13947), .A2(n9244), .ZN(n8783) );
  NAND2_X1 U11419 ( .A1(n8784), .A2(n8783), .ZN(n8786) );
  AOI22_X1 U11420 ( .A1(n11844), .A2(n9194), .B1(n9131), .B2(n13947), .ZN(
        n8785) );
  XNOR2_X1 U11421 ( .A(n8788), .B(n8787), .ZN(n10653) );
  NAND2_X1 U11422 ( .A1(n10653), .A2(n9228), .ZN(n8798) );
  INV_X1 U11423 ( .A(n8789), .ZN(n8791) );
  NAND2_X1 U11424 ( .A1(n8791), .A2(n8790), .ZN(n8793) );
  NAND2_X1 U11425 ( .A1(n8793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8792) );
  MUX2_X1 U11426 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8792), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8796) );
  INV_X1 U11427 ( .A(n8793), .ZN(n8795) );
  INV_X1 U11428 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11429 ( .A1(n8795), .A2(n8794), .ZN(n8832) );
  AOI22_X1 U11430 ( .A1(n9125), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10854), 
        .B2(n13975), .ZN(n8797) );
  NAND2_X1 U11431 ( .A1(n12159), .A2(n9194), .ZN(n8804) );
  NAND2_X1 U11432 ( .A1(n6407), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8802) );
  INV_X1 U11433 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n12375) );
  OR2_X1 U11434 ( .A1(n8924), .A2(n12375), .ZN(n8801) );
  INV_X1 U11435 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8815) );
  XNOR2_X1 U11436 ( .A(n8816), .B(n8815), .ZN(n13769) );
  OR2_X1 U11437 ( .A1(n9234), .A2(n13769), .ZN(n8800) );
  INV_X1 U11438 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n12156) );
  OR2_X1 U11439 ( .A1(n8948), .A2(n12156), .ZN(n8799) );
  OR2_X1 U11440 ( .A1(n12216), .A2(n9244), .ZN(n8803) );
  NAND2_X1 U11441 ( .A1(n8804), .A2(n8803), .ZN(n8806) );
  INV_X1 U11442 ( .A(n12216), .ZN(n13946) );
  AOI22_X1 U11443 ( .A1(n12159), .A2(n9131), .B1(n13946), .B2(n9194), .ZN(
        n8805) );
  INV_X1 U11444 ( .A(n8808), .ZN(n8809) );
  XNOR2_X1 U11445 ( .A(n8810), .B(n8809), .ZN(n10677) );
  NAND2_X1 U11446 ( .A1(n10677), .A2(n9228), .ZN(n8813) );
  NAND2_X1 U11447 ( .A1(n8832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8811) );
  XNOR2_X1 U11448 ( .A(n8811), .B(P2_IR_REG_9__SCAN_IN), .ZN(n15383) );
  AOI22_X1 U11449 ( .A1(n9125), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10854), 
        .B2(n15383), .ZN(n8812) );
  NAND2_X1 U11450 ( .A1(n13851), .A2(n9131), .ZN(n8825) );
  NAND2_X1 U11451 ( .A1(n6407), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8823) );
  INV_X1 U11452 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n12221) );
  OR2_X1 U11453 ( .A1(n8924), .A2(n12221), .ZN(n8822) );
  INV_X1 U11454 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8814) );
  OAI21_X1 U11455 ( .B1(n8816), .B2(n8815), .A(n8814), .ZN(n8819) );
  INV_X1 U11456 ( .A(n8816), .ZN(n8818) );
  INV_X1 U11457 ( .A(n8836), .ZN(n8838) );
  NAND2_X1 U11458 ( .A1(n8819), .A2(n8838), .ZN(n13849) );
  OR2_X1 U11459 ( .A1(n9234), .A2(n13849), .ZN(n8821) );
  INV_X1 U11460 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n12280) );
  OR2_X1 U11461 ( .A1(n8948), .A2(n12280), .ZN(n8820) );
  NAND2_X1 U11462 ( .A1(n13944), .A2(n8965), .ZN(n8824) );
  NAND2_X1 U11463 ( .A1(n8825), .A2(n8824), .ZN(n8828) );
  NAND2_X1 U11464 ( .A1(n13851), .A2(n9194), .ZN(n8826) );
  OAI21_X1 U11465 ( .B1(n12547), .B2(n9194), .A(n8826), .ZN(n8827) );
  INV_X1 U11466 ( .A(n8828), .ZN(n8829) );
  NAND2_X1 U11467 ( .A1(n10686), .A2(n9228), .ZN(n8835) );
  NAND2_X1 U11468 ( .A1(n8853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8833) );
  XNOR2_X1 U11469 ( .A(n8833), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15395) );
  AOI22_X1 U11470 ( .A1(n9125), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n15395), 
        .B2(n10854), .ZN(n8834) );
  NAND2_X1 U11471 ( .A1(n13753), .A2(n9194), .ZN(n8846) );
  NAND2_X1 U11472 ( .A1(n6407), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8844) );
  INV_X1 U11473 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n12551) );
  OR2_X1 U11474 ( .A1(n8924), .A2(n12551), .ZN(n8843) );
  INV_X1 U11475 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U11476 ( .A1(n8838), .A2(n8837), .ZN(n8839) );
  NAND2_X1 U11477 ( .A1(n8883), .A2(n8839), .ZN(n13751) );
  OR2_X1 U11478 ( .A1(n9234), .A2(n13751), .ZN(n8842) );
  INV_X1 U11479 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8840) );
  OR2_X1 U11480 ( .A1(n8948), .A2(n8840), .ZN(n8841) );
  OR2_X1 U11481 ( .A1(n12422), .A2(n9244), .ZN(n8845) );
  NAND2_X1 U11482 ( .A1(n8846), .A2(n8845), .ZN(n8849) );
  AOI21_X1 U11483 ( .B1(n8850), .B2(n8849), .A(n8847), .ZN(n8848) );
  NAND2_X1 U11484 ( .A1(n8866), .A2(n8852), .ZN(n8867) );
  XNOR2_X1 U11485 ( .A(n8868), .B(n8867), .ZN(n10730) );
  NAND2_X1 U11486 ( .A1(n10730), .A2(n9228), .ZN(n8856) );
  OAI21_X1 U11487 ( .B1(n8853), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8854) );
  XNOR2_X1 U11488 ( .A(n8854), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U11489 ( .A1(n11050), .A2(n10854), .B1(n9125), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U11490 ( .A1(n14382), .A2(n9131), .ZN(n8863) );
  NAND2_X1 U11491 ( .A1(n9235), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8861) );
  INV_X1 U11492 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8857) );
  OR2_X1 U11493 ( .A1(n8950), .A2(n8857), .ZN(n8860) );
  INV_X1 U11494 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8881) );
  XNOR2_X1 U11495 ( .A(n8883), .B(n8881), .ZN(n13890) );
  OR2_X1 U11496 ( .A1(n9234), .A2(n13890), .ZN(n8859) );
  INV_X1 U11497 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11035) );
  OR2_X1 U11498 ( .A1(n8948), .A2(n11035), .ZN(n8858) );
  NAND4_X1 U11499 ( .A1(n8861), .A2(n8860), .A3(n8859), .A4(n8858), .ZN(n13942) );
  NAND2_X1 U11500 ( .A1(n9194), .A2(n13942), .ZN(n8862) );
  INV_X1 U11501 ( .A(n13942), .ZN(n10408) );
  NAND2_X1 U11502 ( .A1(n14382), .A2(n8965), .ZN(n8864) );
  OAI21_X1 U11503 ( .B1(n10408), .B2(n9194), .A(n8864), .ZN(n8865) );
  XNOR2_X1 U11504 ( .A(n8870), .B(n8869), .ZN(n10792) );
  NAND2_X1 U11505 ( .A1(n10792), .A2(n9228), .ZN(n8879) );
  OR2_X1 U11506 ( .A1(n8872), .A2(n8871), .ZN(n8874) );
  NAND2_X1 U11507 ( .A1(n8874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8873) );
  MUX2_X1 U11508 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8873), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8877) );
  INV_X1 U11509 ( .A(n8874), .ZN(n8876) );
  NAND2_X1 U11510 ( .A1(n8876), .A2(n8875), .ZN(n8917) );
  NAND2_X1 U11511 ( .A1(n8877), .A2(n8917), .ZN(n12238) );
  INV_X1 U11512 ( .A(n12238), .ZN(n12247) );
  AOI22_X1 U11513 ( .A1(n9125), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10854), 
        .B2(n12247), .ZN(n8878) );
  NAND2_X1 U11514 ( .A1(n13793), .A2(n8965), .ZN(n8890) );
  NAND2_X1 U11515 ( .A1(n6407), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8888) );
  INV_X1 U11516 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12443) );
  OR2_X1 U11517 ( .A1(n8924), .A2(n12443), .ZN(n8887) );
  INV_X1 U11518 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8880) );
  OAI21_X1 U11519 ( .B1(n8883), .B2(n8881), .A(n8880), .ZN(n8884) );
  NAND2_X1 U11520 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n8882) );
  NAND2_X1 U11521 ( .A1(n8884), .A2(n8903), .ZN(n13790) );
  OR2_X1 U11522 ( .A1(n9234), .A2(n13790), .ZN(n8886) );
  INV_X1 U11523 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n12575) );
  OR2_X1 U11524 ( .A1(n8948), .A2(n12575), .ZN(n8885) );
  OR2_X1 U11525 ( .A1(n12583), .A2(n9244), .ZN(n8889) );
  NAND2_X1 U11526 ( .A1(n8890), .A2(n8889), .ZN(n8892) );
  AOI22_X1 U11527 ( .A1(n13793), .A2(n9131), .B1(n13941), .B2(n9194), .ZN(
        n8891) );
  AOI21_X1 U11528 ( .B1(n8893), .B2(n8892), .A(n8891), .ZN(n8895) );
  NOR2_X1 U11529 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  XNOR2_X1 U11530 ( .A(n8897), .B(n8896), .ZN(n10787) );
  NAND2_X1 U11531 ( .A1(n10787), .A2(n9228), .ZN(n8900) );
  NAND2_X1 U11532 ( .A1(n8917), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8898) );
  XNOR2_X1 U11533 ( .A(n8898), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15424) );
  AOI22_X1 U11534 ( .A1(n9125), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10854), 
        .B2(n15424), .ZN(n8899) );
  NAND2_X1 U11535 ( .A1(n12589), .A2(n9131), .ZN(n8910) );
  NAND2_X1 U11536 ( .A1(n6407), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8908) );
  INV_X1 U11537 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12590) );
  OR2_X1 U11538 ( .A1(n8924), .A2(n12590), .ZN(n8907) );
  INV_X1 U11539 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U11540 ( .A1(n8903), .A2(n8902), .ZN(n8904) );
  NAND2_X1 U11541 ( .A1(n8946), .A2(n8904), .ZN(n13865) );
  OR2_X1 U11542 ( .A1(n9234), .A2(n13865), .ZN(n8906) );
  INV_X1 U11543 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n12654) );
  OR2_X1 U11544 ( .A1(n8948), .A2(n12654), .ZN(n8905) );
  NAND2_X1 U11545 ( .A1(n13940), .A2(n9194), .ZN(n8909) );
  NAND2_X1 U11546 ( .A1(n8910), .A2(n8909), .ZN(n8913) );
  NAND2_X1 U11547 ( .A1(n12589), .A2(n9194), .ZN(n8911) );
  OAI21_X1 U11548 ( .B1(n13730), .B2(n9194), .A(n8911), .ZN(n8912) );
  INV_X1 U11549 ( .A(n8913), .ZN(n8914) );
  NAND2_X1 U11550 ( .A1(n8915), .A2(n10797), .ZN(n8935) );
  XNOR2_X1 U11551 ( .A(n8937), .B(n8936), .ZN(n10996) );
  NAND2_X1 U11552 ( .A1(n10996), .A2(n9228), .ZN(n8922) );
  OAI21_X1 U11553 ( .B1(n8917), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8918) );
  MUX2_X1 U11554 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8918), .S(
        P2_IR_REG_14__SCAN_IN), .Z(n8920) );
  AND2_X1 U11555 ( .A1(n8920), .A2(n8919), .ZN(n15437) );
  AOI22_X1 U11556 ( .A1(n9125), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n10854), 
        .B2(n15437), .ZN(n8921) );
  NAND2_X2 U11557 ( .A1(n8922), .A2(n8921), .ZN(n14377) );
  NAND2_X1 U11558 ( .A1(n14377), .A2(n8965), .ZN(n8931) );
  NAND2_X1 U11559 ( .A1(n6407), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8929) );
  INV_X1 U11560 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8923) );
  OR2_X1 U11561 ( .A1(n8924), .A2(n8923), .ZN(n8928) );
  XNOR2_X1 U11562 ( .A(n8946), .B(n8945), .ZN(n13727) );
  OR2_X1 U11563 ( .A1(n9234), .A2(n13727), .ZN(n8927) );
  INV_X1 U11564 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8925) );
  OR2_X1 U11565 ( .A1(n8948), .A2(n8925), .ZN(n8926) );
  OR2_X1 U11566 ( .A1(n12584), .A2(n9244), .ZN(n8930) );
  NAND2_X1 U11567 ( .A1(n8931), .A2(n8930), .ZN(n8934) );
  NAND2_X1 U11568 ( .A1(n14377), .A2(n9131), .ZN(n8932) );
  OAI21_X1 U11569 ( .B1(n12584), .B2(n6411), .A(n8932), .ZN(n8933) );
  NAND2_X1 U11570 ( .A1(n11060), .A2(n9228), .ZN(n8943) );
  NAND2_X1 U11571 ( .A1(n8919), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8940) );
  MUX2_X1 U11572 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8940), .S(
        P2_IR_REG_15__SCAN_IN), .Z(n8941) );
  OR2_X1 U11573 ( .A1(n8919), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8983) );
  AOI22_X1 U11574 ( .A1(n9125), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n10854), 
        .B2(n13993), .ZN(n8942) );
  NAND2_X2 U11575 ( .A1(n8943), .A2(n8942), .ZN(n14433) );
  NAND2_X1 U11576 ( .A1(n14433), .A2(n9131), .ZN(n8956) );
  OAI21_X1 U11577 ( .B1(n8946), .B2(n8945), .A(n12252), .ZN(n8947) );
  AND2_X1 U11578 ( .A1(n8947), .A2(n8969), .ZN(n14257) );
  NAND2_X1 U11579 ( .A1(n9149), .A2(n14257), .ZN(n8954) );
  NAND2_X1 U11580 ( .A1(n9235), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8953) );
  INV_X1 U11581 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n12248) );
  OR2_X1 U11582 ( .A1(n8948), .A2(n12248), .ZN(n8952) );
  INV_X1 U11583 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8949) );
  OR2_X1 U11584 ( .A1(n8950), .A2(n8949), .ZN(n8951) );
  NAND4_X1 U11585 ( .A1(n8954), .A2(n8953), .A3(n8952), .A4(n8951), .ZN(n13938) );
  NAND2_X1 U11586 ( .A1(n9194), .A2(n13938), .ZN(n8955) );
  NAND2_X1 U11587 ( .A1(n8956), .A2(n8955), .ZN(n8958) );
  AOI22_X1 U11588 ( .A1(n14433), .A2(n9194), .B1(n9131), .B2(n13938), .ZN(
        n8957) );
  XNOR2_X1 U11589 ( .A(n8961), .B(n8960), .ZN(n10992) );
  NAND2_X1 U11590 ( .A1(n10992), .A2(n9228), .ZN(n8964) );
  NAND2_X1 U11591 ( .A1(n8983), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8962) );
  XNOR2_X1 U11592 ( .A(n8962), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14011) );
  AOI22_X1 U11593 ( .A1(n9125), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10854), 
        .B2(n14011), .ZN(n8963) );
  NAND2_X1 U11594 ( .A1(n14245), .A2(n8965), .ZN(n8975) );
  NAND2_X1 U11595 ( .A1(n9235), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8967) );
  NAND2_X1 U11596 ( .A1(n6407), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8966) );
  AND2_X1 U11597 ( .A1(n8967), .A2(n8966), .ZN(n8973) );
  INV_X1 U11598 ( .A(n8969), .ZN(n8968) );
  INV_X1 U11599 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n15656) );
  NAND2_X1 U11600 ( .A1(n8969), .A2(n15656), .ZN(n8970) );
  NAND2_X1 U11601 ( .A1(n8990), .A2(n8970), .ZN(n14240) );
  OR2_X1 U11602 ( .A1(n14240), .A2(n9234), .ZN(n8972) );
  NAND2_X1 U11603 ( .A1(n13937), .A2(n9131), .ZN(n8974) );
  NAND2_X1 U11604 ( .A1(n8975), .A2(n8974), .ZN(n8978) );
  AOI22_X1 U11605 ( .A1(n14245), .A2(n9131), .B1(n13937), .B2(n9194), .ZN(
        n8976) );
  AOI21_X1 U11606 ( .B1(n8979), .B2(n8978), .A(n8976), .ZN(n8977) );
  INV_X1 U11607 ( .A(n8977), .ZN(n8980) );
  XNOR2_X1 U11608 ( .A(n8981), .B(n8982), .ZN(n11089) );
  NAND2_X1 U11609 ( .A1(n11089), .A2(n9228), .ZN(n8987) );
  OAI21_X1 U11610 ( .B1(n8983), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8984) );
  MUX2_X1 U11611 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8984), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8985) );
  AND2_X1 U11612 ( .A1(n8985), .A2(n9005), .ZN(n15449) );
  AOI22_X1 U11613 ( .A1(n10854), .A2(n15449), .B1(n9125), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U11614 ( .A1(n14222), .A2(n9131), .ZN(n8996) );
  INV_X1 U11615 ( .A(n8990), .ZN(n8988) );
  INV_X1 U11616 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U11617 ( .A1(n8990), .A2(n8989), .ZN(n8991) );
  NAND2_X1 U11618 ( .A1(n9009), .A2(n8991), .ZN(n13825) );
  OR2_X1 U11619 ( .A1(n13825), .A2(n9234), .ZN(n8994) );
  AOI22_X1 U11620 ( .A1(n6407), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n9235), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8993) );
  INV_X1 U11621 ( .A(n14198), .ZN(n13936) );
  NAND2_X1 U11622 ( .A1(n13936), .A2(n9194), .ZN(n8995) );
  NAND2_X1 U11623 ( .A1(n8996), .A2(n8995), .ZN(n8998) );
  NAND2_X1 U11624 ( .A1(n8999), .A2(n8998), .ZN(n9002) );
  NAND2_X1 U11625 ( .A1(n14222), .A2(n9194), .ZN(n8997) );
  OAI21_X1 U11626 ( .B1(n14198), .B2(n9194), .A(n8997), .ZN(n9001) );
  INV_X1 U11627 ( .A(n9017), .ZN(n9020) );
  NAND2_X1 U11628 ( .A1(n9005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9006) );
  XNOR2_X1 U11629 ( .A(n9006), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14017) );
  AOI22_X1 U11630 ( .A1(n9125), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n10854), 
        .B2(n14017), .ZN(n9007) );
  NAND2_X1 U11631 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  AND2_X1 U11632 ( .A1(n9046), .A2(n9010), .ZN(n14208) );
  NAND2_X1 U11633 ( .A1(n14208), .A2(n9149), .ZN(n9013) );
  AOI22_X1 U11634 ( .A1(n6407), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n9235), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n9012) );
  NOR2_X1 U11635 ( .A1(n10421), .A2(n9244), .ZN(n9014) );
  AOI21_X1 U11636 ( .B1(n14209), .B2(n9194), .A(n9014), .ZN(n9016) );
  INV_X1 U11637 ( .A(n9016), .ZN(n9019) );
  OAI22_X1 U11638 ( .A1(n14352), .A2(n9244), .B1(n10421), .B2(n6412), .ZN(
        n9015) );
  NAND2_X1 U11639 ( .A1(n9022), .A2(n9021), .ZN(n9024) );
  OR2_X1 U11640 ( .A1(n9003), .A2(n11013), .ZN(n9023) );
  NAND2_X1 U11641 ( .A1(n9026), .A2(n9025), .ZN(n9027) );
  NAND2_X1 U11642 ( .A1(n11585), .A2(n9228), .ZN(n9030) );
  AOI22_X1 U11643 ( .A1(n9125), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n14031), 
        .B2(n10854), .ZN(n9029) );
  NAND2_X2 U11644 ( .A1(n9030), .A2(n9029), .ZN(n14179) );
  INV_X1 U11645 ( .A(n14179), .ZN(n14421) );
  XNOR2_X1 U11646 ( .A(n9046), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n14180) );
  NAND2_X1 U11647 ( .A1(n14180), .A2(n9149), .ZN(n9035) );
  INV_X1 U11648 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14347) );
  NAND2_X1 U11649 ( .A1(n9235), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U11650 ( .A1(n6407), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9031) );
  OAI211_X1 U11651 ( .C1(n8948), .C2(n14347), .A(n9032), .B(n9031), .ZN(n9033)
         );
  INV_X1 U11652 ( .A(n9033), .ZN(n9034) );
  OAI22_X1 U11653 ( .A1(n14421), .A2(n9244), .B1(n14200), .B2(n6412), .ZN(
        n9037) );
  AOI22_X1 U11654 ( .A1(n14179), .A2(n9194), .B1(n9131), .B2(n13934), .ZN(
        n9036) );
  XNOR2_X1 U11655 ( .A(n9137), .B(n9040), .ZN(n11661) );
  NAND2_X1 U11656 ( .A1(n11661), .A2(n9228), .ZN(n9042) );
  NAND2_X1 U11657 ( .A1(n9125), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9041) );
  NAND2_X2 U11658 ( .A1(n9042), .A2(n9041), .ZN(n14336) );
  AND2_X1 U11659 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n9043) );
  INV_X1 U11660 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n13760) );
  INV_X1 U11661 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9045) );
  OAI21_X1 U11662 ( .B1(n9046), .B2(n13760), .A(n9045), .ZN(n9047) );
  NAND2_X1 U11663 ( .A1(n9146), .A2(n9047), .ZN(n14164) );
  OR2_X1 U11664 ( .A1(n14164), .A2(n9234), .ZN(n9052) );
  INV_X1 U11665 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n14342) );
  NAND2_X1 U11666 ( .A1(n6407), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U11667 ( .A1(n9235), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9048) );
  OAI211_X1 U11668 ( .C1(n14342), .C2(n8948), .A(n9049), .B(n9048), .ZN(n9050)
         );
  INV_X1 U11669 ( .A(n9050), .ZN(n9051) );
  AOI22_X1 U11670 ( .A1(n14336), .A2(n9244), .B1(n9131), .B2(n13933), .ZN(
        n9053) );
  AOI22_X1 U11671 ( .A1(n14336), .A2(n9131), .B1(n13933), .B2(n9194), .ZN(
        n9055) );
  INV_X1 U11672 ( .A(n9053), .ZN(n9054) );
  XNOR2_X1 U11673 ( .A(n9056), .B(SI_26_), .ZN(n9057) );
  NAND2_X1 U11674 ( .A1(n12596), .A2(n9214), .ZN(n9060) );
  NAND2_X1 U11675 ( .A1(n9125), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9059) );
  INV_X1 U11676 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13778) );
  INV_X1 U11677 ( .A(n9148), .ZN(n9062) );
  AND2_X1 U11678 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n9061) );
  INV_X1 U11679 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13838) );
  NAND2_X1 U11680 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n9063) );
  INV_X1 U11681 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9065) );
  INV_X1 U11682 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9064) );
  OAI21_X1 U11683 ( .B1(n9094), .B2(n9065), .A(n9064), .ZN(n9066) );
  NAND2_X1 U11684 ( .A1(n14068), .A2(n9149), .ZN(n9072) );
  INV_X1 U11685 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U11686 ( .A1(n6407), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9068) );
  NAND2_X1 U11687 ( .A1(n9235), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9067) );
  OAI211_X1 U11688 ( .C1(n9069), .C2(n8948), .A(n9068), .B(n9067), .ZN(n9070)
         );
  INV_X1 U11689 ( .A(n9070), .ZN(n9071) );
  OR2_X1 U11690 ( .A1(n14070), .A2(n9131), .ZN(n9074) );
  NAND2_X1 U11691 ( .A1(n14083), .A2(n9131), .ZN(n9073) );
  NAND2_X1 U11692 ( .A1(n9074), .A2(n9073), .ZN(n9172) );
  XNOR2_X1 U11693 ( .A(n9076), .B(n9075), .ZN(n12381) );
  NAND2_X1 U11694 ( .A1(n12381), .A2(n9228), .ZN(n9078) );
  NAND2_X1 U11695 ( .A1(n9125), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9077) );
  XNOR2_X1 U11696 ( .A(n9094), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14088) );
  NAND2_X1 U11697 ( .A1(n14088), .A2(n9149), .ZN(n9084) );
  INV_X1 U11698 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U11699 ( .A1(n6407), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U11700 ( .A1(n9235), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9079) );
  OAI211_X1 U11701 ( .C1(n9081), .C2(n8948), .A(n9080), .B(n9079), .ZN(n9082)
         );
  INV_X1 U11702 ( .A(n9082), .ZN(n9083) );
  NOR2_X1 U11703 ( .A1(n13913), .A2(n9131), .ZN(n9085) );
  AOI21_X1 U11704 ( .B1(n14089), .B2(n9131), .A(n9085), .ZN(n9169) );
  NAND2_X1 U11705 ( .A1(n14089), .A2(n9194), .ZN(n9087) );
  OR2_X1 U11706 ( .A1(n13913), .A2(n9244), .ZN(n9086) );
  NAND2_X1 U11707 ( .A1(n9087), .A2(n9086), .ZN(n9168) );
  NAND2_X1 U11708 ( .A1(n9169), .A2(n9168), .ZN(n9088) );
  NAND2_X1 U11709 ( .A1(n9177), .A2(n9088), .ZN(n9199) );
  XNOR2_X1 U11710 ( .A(n9089), .B(n9090), .ZN(n12138) );
  NAND2_X1 U11711 ( .A1(n12138), .A2(n9228), .ZN(n9092) );
  NAND2_X1 U11712 ( .A1(n9125), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U11713 ( .A1(n9114), .A2(n13838), .ZN(n9093) );
  NAND2_X1 U11714 ( .A1(n9094), .A2(n9093), .ZN(n14104) );
  OR2_X1 U11715 ( .A1(n14104), .A2(n9234), .ZN(n9100) );
  INV_X1 U11716 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U11717 ( .A1(n9235), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9096) );
  NAND2_X1 U11718 ( .A1(n6407), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9095) );
  OAI211_X1 U11719 ( .C1(n8948), .C2(n9097), .A(n9096), .B(n9095), .ZN(n9098)
         );
  INV_X1 U11720 ( .A(n9098), .ZN(n9099) );
  NOR2_X1 U11721 ( .A1(n14114), .A2(n9131), .ZN(n9101) );
  AOI21_X1 U11722 ( .B1(n14312), .B2(n9131), .A(n9101), .ZN(n9198) );
  NAND2_X1 U11723 ( .A1(n14312), .A2(n9194), .ZN(n9103) );
  NAND2_X1 U11724 ( .A1(n14081), .A2(n9131), .ZN(n9102) );
  NAND2_X1 U11725 ( .A1(n9103), .A2(n9102), .ZN(n9197) );
  AND2_X1 U11726 ( .A1(n9198), .A2(n9197), .ZN(n9104) );
  OR2_X1 U11727 ( .A1(n9199), .A2(n9104), .ZN(n9167) );
  NAND2_X1 U11728 ( .A1(n6660), .A2(n9124), .ZN(n9107) );
  NAND2_X1 U11729 ( .A1(n9105), .A2(SI_22_), .ZN(n9106) );
  NAND2_X1 U11730 ( .A1(n9107), .A2(n9106), .ZN(n9110) );
  XNOR2_X1 U11731 ( .A(n9108), .B(SI_23_), .ZN(n9109) );
  XNOR2_X2 U11732 ( .A(n9110), .B(n9109), .ZN(n11931) );
  NAND2_X1 U11733 ( .A1(n11931), .A2(n9228), .ZN(n9112) );
  NAND2_X1 U11734 ( .A1(n9125), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9111) );
  NAND2_X2 U11735 ( .A1(n9112), .A2(n9111), .ZN(n14122) );
  INV_X1 U11736 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13878) );
  INV_X1 U11737 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9113) );
  OAI21_X1 U11738 ( .B1(n9148), .B2(n13878), .A(n9113), .ZN(n9115) );
  NAND2_X1 U11739 ( .A1(n9115), .A2(n9114), .ZN(n13742) );
  OR2_X1 U11740 ( .A1(n13742), .A2(n9234), .ZN(n9120) );
  INV_X1 U11741 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14325) );
  NAND2_X1 U11742 ( .A1(n6407), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U11743 ( .A1(n9235), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9116) );
  OAI211_X1 U11744 ( .C1(n14325), .C2(n8948), .A(n9117), .B(n9116), .ZN(n9118)
         );
  INV_X1 U11745 ( .A(n9118), .ZN(n9119) );
  NOR2_X1 U11746 ( .A1(n13877), .A2(n9131), .ZN(n9121) );
  AOI21_X1 U11747 ( .B1(n14122), .B2(n9131), .A(n9121), .ZN(n9166) );
  NAND2_X1 U11748 ( .A1(n14122), .A2(n9244), .ZN(n9123) );
  NAND2_X1 U11749 ( .A1(n14098), .A2(n9131), .ZN(n9122) );
  NAND2_X1 U11750 ( .A1(n9123), .A2(n9122), .ZN(n9165) );
  XNOR2_X1 U11751 ( .A(n9897), .B(n9124), .ZN(n11895) );
  NAND2_X1 U11752 ( .A1(n11895), .A2(n9228), .ZN(n9127) );
  NAND2_X1 U11753 ( .A1(n9125), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9126) );
  XNOR2_X1 U11754 ( .A(n9148), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n14139) );
  INV_X1 U11755 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14330) );
  NAND2_X1 U11756 ( .A1(n6407), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U11757 ( .A1(n9235), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9128) );
  OAI211_X1 U11758 ( .C1(n14330), .C2(n8948), .A(n9129), .B(n9128), .ZN(n9130)
         );
  AOI21_X1 U11759 ( .B1(n14139), .B2(n9149), .A(n9130), .ZN(n14113) );
  NOR2_X1 U11760 ( .A1(n14113), .A2(n9131), .ZN(n9132) );
  AOI21_X1 U11761 ( .B1(n14138), .B2(n9131), .A(n9132), .ZN(n9163) );
  NAND2_X1 U11762 ( .A1(n14138), .A2(n9244), .ZN(n9134) );
  OR2_X1 U11763 ( .A1(n14113), .A2(n9244), .ZN(n9133) );
  NAND2_X1 U11764 ( .A1(n9134), .A2(n9133), .ZN(n9162) );
  AND2_X1 U11765 ( .A1(n9163), .A2(n9162), .ZN(n9135) );
  NAND2_X1 U11766 ( .A1(n9137), .A2(n9136), .ZN(n9140) );
  INV_X1 U11767 ( .A(n9039), .ZN(n9138) );
  NAND2_X1 U11768 ( .A1(n9138), .A2(SI_20_), .ZN(n9139) );
  XNOR2_X1 U11769 ( .A(n9141), .B(SI_21_), .ZN(n9142) );
  NAND2_X1 U11770 ( .A1(n11689), .A2(n9228), .ZN(n9145) );
  NAND2_X1 U11771 ( .A1(n9125), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U11772 ( .A1(n14151), .A2(n9131), .ZN(n9156) );
  NAND2_X1 U11773 ( .A1(n9146), .A2(n13778), .ZN(n9147) );
  AND2_X1 U11774 ( .A1(n9148), .A2(n9147), .ZN(n14152) );
  NAND2_X1 U11775 ( .A1(n14152), .A2(n9149), .ZN(n9154) );
  INV_X1 U11776 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n15668) );
  NAND2_X1 U11777 ( .A1(n9235), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U11778 ( .A1(n6407), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9150) );
  OAI211_X1 U11779 ( .C1(n15668), .C2(n8948), .A(n9151), .B(n9150), .ZN(n9152)
         );
  INV_X1 U11780 ( .A(n9152), .ZN(n9153) );
  NAND2_X1 U11781 ( .A1(n9154), .A2(n9153), .ZN(n13932) );
  NAND2_X1 U11782 ( .A1(n13932), .A2(n9194), .ZN(n9155) );
  AND2_X1 U11783 ( .A1(n13932), .A2(n9131), .ZN(n9157) );
  AOI21_X1 U11784 ( .B1(n14151), .B2(n9194), .A(n9157), .ZN(n9161) );
  NAND2_X1 U11785 ( .A1(n7862), .A2(n9158), .ZN(n9159) );
  OR3_X1 U11786 ( .A1(n9164), .A2(n9163), .A3(n9162), .ZN(n9205) );
  OR3_X1 U11787 ( .A1(n9167), .A2(n9166), .A3(n9165), .ZN(n9203) );
  INV_X1 U11788 ( .A(n9168), .ZN(n9171) );
  INV_X1 U11789 ( .A(n9169), .ZN(n9170) );
  AND2_X1 U11790 ( .A1(n9171), .A2(n9170), .ZN(n9176) );
  INV_X1 U11791 ( .A(n9172), .ZN(n9175) );
  INV_X1 U11792 ( .A(n9173), .ZN(n9174) );
  AOI22_X1 U11793 ( .A1(n9177), .A2(n9176), .B1(n9175), .B2(n9174), .ZN(n9202)
         );
  XNOR2_X1 U11794 ( .A(n9179), .B(SI_27_), .ZN(n9180) );
  XNOR2_X1 U11795 ( .A(n9178), .B(n9180), .ZN(n12892) );
  NAND2_X1 U11796 ( .A1(n12892), .A2(n9214), .ZN(n9182) );
  NAND2_X1 U11797 ( .A1(n9125), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9181) );
  INV_X1 U11798 ( .A(n9184), .ZN(n9183) );
  NAND2_X1 U11799 ( .A1(n9183), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9232) );
  INV_X1 U11800 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13713) );
  NAND2_X1 U11801 ( .A1(n9184), .A2(n13713), .ZN(n9185) );
  NAND2_X1 U11802 ( .A1(n9232), .A2(n9185), .ZN(n14057) );
  OR2_X1 U11803 ( .A1(n14057), .A2(n9234), .ZN(n9191) );
  INV_X1 U11804 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9188) );
  NAND2_X1 U11805 ( .A1(n6407), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9187) );
  NAND2_X1 U11806 ( .A1(n9235), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9186) );
  OAI211_X1 U11807 ( .C1(n9188), .C2(n8948), .A(n9187), .B(n9186), .ZN(n9189)
         );
  INV_X1 U11808 ( .A(n9189), .ZN(n9190) );
  AND2_X1 U11809 ( .A1(n14065), .A2(n9131), .ZN(n9192) );
  AOI21_X1 U11810 ( .B1(n14298), .B2(n9244), .A(n9192), .ZN(n9247) );
  NAND2_X1 U11811 ( .A1(n14298), .A2(n9131), .ZN(n9196) );
  NAND2_X1 U11812 ( .A1(n14065), .A2(n9194), .ZN(n9195) );
  NAND2_X1 U11813 ( .A1(n9196), .A2(n9195), .ZN(n9246) );
  NAND2_X1 U11814 ( .A1(n9247), .A2(n9246), .ZN(n9201) );
  OR3_X1 U11815 ( .A1(n9199), .A2(n9198), .A3(n9197), .ZN(n9200) );
  AND4_X1 U11816 ( .A1(n9203), .A2(n9202), .A3(n9201), .A4(n9200), .ZN(n9204)
         );
  MUX2_X1 U11817 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n10572), .Z(n9208) );
  XNOR2_X1 U11818 ( .A(n9208), .B(SI_31_), .ZN(n9209) );
  NAND2_X1 U11819 ( .A1(n14438), .A2(n9214), .ZN(n9211) );
  NAND2_X1 U11820 ( .A1(n9125), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9210) );
  NAND2_X1 U11821 ( .A1(n12894), .A2(n9214), .ZN(n9216) );
  NAND2_X1 U11822 ( .A1(n9125), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9215) );
  INV_X1 U11823 ( .A(n14292), .ZN(n12922) );
  INV_X1 U11824 ( .A(n9232), .ZN(n9217) );
  NAND2_X1 U11825 ( .A1(n9217), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12927) );
  OR2_X1 U11826 ( .A1(n12927), .A2(n9234), .ZN(n9222) );
  INV_X1 U11827 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n15716) );
  NAND2_X1 U11828 ( .A1(n6407), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U11829 ( .A1(n9235), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9218) );
  OAI211_X1 U11830 ( .C1(n15716), .C2(n8948), .A(n9219), .B(n9218), .ZN(n9220)
         );
  INV_X1 U11831 ( .A(n9220), .ZN(n9221) );
  NAND2_X1 U11832 ( .A1(n9222), .A2(n9221), .ZN(n13930) );
  INV_X1 U11833 ( .A(n13930), .ZN(n9223) );
  OAI22_X1 U11834 ( .A1(n12922), .A2(n9244), .B1(n9223), .B2(n6411), .ZN(n9255) );
  AOI22_X1 U11835 ( .A1(n14292), .A2(n9194), .B1(n9131), .B2(n13930), .ZN(
        n9254) );
  NOR2_X1 U11836 ( .A1(n9255), .A2(n9254), .ZN(n9253) );
  NAND2_X1 U11837 ( .A1(n9225), .A2(n9224), .ZN(n9226) );
  NAND2_X1 U11838 ( .A1(n9227), .A2(n9226), .ZN(n14443) );
  NAND2_X1 U11839 ( .A1(n14443), .A2(n9228), .ZN(n9230) );
  NAND2_X1 U11840 ( .A1(n9125), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U11841 ( .A1(n12678), .A2(n8965), .ZN(n9243) );
  INV_X1 U11842 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9231) );
  NAND2_X1 U11843 ( .A1(n9232), .A2(n9231), .ZN(n9233) );
  NAND2_X1 U11844 ( .A1(n12927), .A2(n9233), .ZN(n9496) );
  OR2_X1 U11845 ( .A1(n9496), .A2(n9234), .ZN(n9241) );
  INV_X1 U11846 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U11847 ( .A1(n6407), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9237) );
  NAND2_X1 U11848 ( .A1(n9235), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9236) );
  OAI211_X1 U11849 ( .C1(n9238), .C2(n8948), .A(n9237), .B(n9236), .ZN(n9239)
         );
  INV_X1 U11850 ( .A(n9239), .ZN(n9240) );
  NAND2_X1 U11851 ( .A1(n14050), .A2(n9131), .ZN(n9242) );
  NAND2_X1 U11852 ( .A1(n9243), .A2(n9242), .ZN(n9251) );
  INV_X1 U11853 ( .A(n9251), .ZN(n9249) );
  AND2_X1 U11854 ( .A1(n14050), .A2(n9244), .ZN(n9245) );
  AOI21_X1 U11855 ( .B1(n12678), .B2(n9131), .A(n9245), .ZN(n9252) );
  INV_X1 U11856 ( .A(n9252), .ZN(n9248) );
  OAI22_X1 U11857 ( .A1(n9249), .A2(n9248), .B1(n9247), .B2(n9246), .ZN(n9250)
         );
  NOR3_X1 U11858 ( .A1(n9294), .A2(n9253), .A3(n9250), .ZN(n9263) );
  AOI22_X1 U11859 ( .A1(n14387), .A2(n9194), .B1(n9131), .B2(n13928), .ZN(
        n9260) );
  INV_X1 U11860 ( .A(n9267), .ZN(n9259) );
  AOI22_X1 U11861 ( .A1(n9257), .A2(n9256), .B1(n9255), .B2(n9254), .ZN(n9258)
         );
  AOI21_X1 U11862 ( .B1(n9260), .B2(n9259), .A(n9258), .ZN(n9261) );
  INV_X1 U11863 ( .A(n9266), .ZN(n9268) );
  AOI211_X1 U11864 ( .C1(n6411), .C2(n14387), .A(n9268), .B(n9267), .ZN(n9270)
         );
  XNOR2_X1 U11865 ( .A(n14292), .B(n13930), .ZN(n12914) );
  INV_X1 U11866 ( .A(n12914), .ZN(n9293) );
  XNOR2_X1 U11867 ( .A(n14286), .B(n12918), .ZN(n9292) );
  NAND2_X1 U11868 ( .A1(n12678), .A2(n14050), .ZN(n12911) );
  OR2_X1 U11869 ( .A1(n12678), .A2(n14050), .ZN(n9271) );
  NAND2_X1 U11870 ( .A1(n12911), .A2(n9271), .ZN(n10435) );
  XNOR2_X1 U11871 ( .A(n14070), .B(n14083), .ZN(n14071) );
  OR2_X1 U11872 ( .A1(n14138), .A2(n14113), .ZN(n10426) );
  NAND2_X1 U11873 ( .A1(n14138), .A2(n14113), .ZN(n9272) );
  NAND2_X1 U11874 ( .A1(n10426), .A2(n9272), .ZN(n14127) );
  XNOR2_X1 U11875 ( .A(n14209), .B(n10421), .ZN(n14186) );
  XNOR2_X1 U11876 ( .A(n14222), .B(n14198), .ZN(n14220) );
  XNOR2_X1 U11877 ( .A(n14245), .B(n13937), .ZN(n14232) );
  INV_X1 U11878 ( .A(n14232), .ZN(n14233) );
  INV_X1 U11879 ( .A(n13938), .ZN(n13811) );
  XNOR2_X1 U11880 ( .A(n14433), .B(n13811), .ZN(n14258) );
  XNOR2_X1 U11881 ( .A(n14377), .B(n13939), .ZN(n12643) );
  NOR2_X1 U11882 ( .A1(n12589), .A2(n13730), .ZN(n10412) );
  NAND2_X1 U11883 ( .A1(n12589), .A2(n13730), .ZN(n10411) );
  INV_X1 U11884 ( .A(n10411), .ZN(n9273) );
  XNOR2_X1 U11885 ( .A(n11844), .B(n12152), .ZN(n11771) );
  INV_X1 U11886 ( .A(n11771), .ZN(n9279) );
  AND2_X1 U11887 ( .A1(n13954), .A2(n11407), .ZN(n11341) );
  OR2_X1 U11888 ( .A1(n11341), .A2(n10985), .ZN(n15469) );
  NAND2_X1 U11889 ( .A1(n13953), .A2(n12747), .ZN(n9275) );
  NAND2_X1 U11890 ( .A1(n10986), .A2(n11410), .ZN(n9276) );
  NOR2_X1 U11891 ( .A1(n15469), .A2(n9276), .ZN(n9277) );
  XNOR2_X1 U11892 ( .A(n13952), .B(n11619), .ZN(n11622) );
  NAND3_X1 U11893 ( .A1(n9279), .A2(n9278), .A3(n11859), .ZN(n9280) );
  XNOR2_X1 U11894 ( .A(n12159), .B(n12216), .ZN(n12151) );
  XNOR2_X1 U11895 ( .A(n13851), .B(n12547), .ZN(n12215) );
  NOR2_X1 U11896 ( .A1(n12582), .A2(n9281), .ZN(n9283) );
  XNOR2_X1 U11897 ( .A(n13793), .B(n12583), .ZN(n12436) );
  INV_X1 U11898 ( .A(n12436), .ZN(n9282) );
  XNOR2_X1 U11899 ( .A(n14382), .B(n13942), .ZN(n12430) );
  NAND4_X1 U11900 ( .A1(n12643), .A2(n9283), .A3(n9282), .A4(n12430), .ZN(
        n9284) );
  XNOR2_X1 U11901 ( .A(n14179), .B(n13934), .ZN(n14173) );
  NAND2_X1 U11902 ( .A1(n14159), .A2(n14173), .ZN(n9285) );
  XNOR2_X1 U11903 ( .A(n14312), .B(n14114), .ZN(n10429) );
  XNOR2_X1 U11904 ( .A(n14089), .B(n13913), .ZN(n14078) );
  OR2_X1 U11905 ( .A1(n14122), .A2(n14098), .ZN(n10380) );
  INV_X1 U11906 ( .A(n10380), .ZN(n9287) );
  AND2_X1 U11907 ( .A1(n14122), .A2(n14098), .ZN(n10381) );
  NAND2_X1 U11908 ( .A1(n14117), .A2(n14148), .ZN(n9288) );
  NOR2_X1 U11909 ( .A1(n14071), .A2(n9290), .ZN(n9291) );
  XNOR2_X1 U11910 ( .A(n14298), .B(n14065), .ZN(n14048) );
  XNOR2_X1 U11911 ( .A(n9295), .B(n14031), .ZN(n9298) );
  NAND2_X1 U11912 ( .A1(n9324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9297) );
  OR2_X1 U11913 ( .A1(n10855), .A2(P2_U3088), .ZN(n9331) );
  NOR3_X1 U11914 ( .A1(n9298), .A2(n8614), .A3(n9331), .ZN(n9299) );
  INV_X1 U11915 ( .A(n9300), .ZN(n9303) );
  NOR3_X1 U11916 ( .A1(n11690), .A2(n11587), .A3(n11662), .ZN(n9302) );
  INV_X1 U11917 ( .A(n9331), .ZN(n11932) );
  NAND2_X1 U11918 ( .A1(n9305), .A2(n7858), .ZN(n9334) );
  NAND2_X1 U11919 ( .A1(n11896), .A2(n7191), .ZN(n9306) );
  OAI211_X1 U11920 ( .C1(n14031), .C2(n11690), .A(n9306), .B(n9497), .ZN(n9307) );
  OR2_X1 U11921 ( .A1(n8587), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9309) );
  NOR2_X1 U11922 ( .A1(n9309), .A2(n9308), .ZN(n9310) );
  AND2_X1 U11923 ( .A1(n9311), .A2(n9310), .ZN(n9312) );
  NOR2_X1 U11924 ( .A1(n9317), .A2(n14440), .ZN(n9314) );
  MUX2_X1 U11925 ( .A(n14440), .B(n9314), .S(P2_IR_REG_25__SCAN_IN), .Z(n9315)
         );
  NAND2_X1 U11926 ( .A1(n9319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9320) );
  MUX2_X1 U11927 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9320), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9322) );
  NAND2_X1 U11928 ( .A1(n9322), .A2(n9321), .ZN(n12598) );
  NAND2_X1 U11929 ( .A1(n10855), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9327) );
  INV_X1 U11930 ( .A(n14449), .ZN(n12916) );
  INV_X1 U11931 ( .A(n10859), .ZN(n9329) );
  NAND4_X1 U11932 ( .A1(n15466), .A2(n12916), .A3(n14097), .A4(n9494), .ZN(
        n9330) );
  OAI211_X1 U11933 ( .C1(n9332), .C2(n9331), .A(n9330), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9333) );
  INV_X1 U11934 ( .A(n9337), .ZN(n9338) );
  XNOR2_X1 U11935 ( .A(n14122), .B(n9451), .ZN(n9439) );
  XNOR2_X1 U11936 ( .A(n14138), .B(n9451), .ZN(n9437) );
  NOR2_X4 U11937 ( .A1(n11408), .A2(n11410), .ZN(n14262) );
  NAND2_X1 U11938 ( .A1(n9349), .A2(n7158), .ZN(n9341) );
  XNOR2_X1 U11939 ( .A(n9340), .B(n9341), .ZN(n11472) );
  NAND2_X1 U11940 ( .A1(n11471), .A2(n11472), .ZN(n11470) );
  INV_X1 U11941 ( .A(n9340), .ZN(n9342) );
  NAND2_X1 U11942 ( .A1(n9342), .A2(n9341), .ZN(n9343) );
  XNOR2_X1 U11943 ( .A(n9344), .B(n15472), .ZN(n9346) );
  NAND2_X1 U11944 ( .A1(n9349), .A2(n13952), .ZN(n9345) );
  NAND2_X1 U11945 ( .A1(n9346), .A2(n9345), .ZN(n9348) );
  XNOR2_X1 U11946 ( .A(n9451), .B(n11414), .ZN(n9350) );
  NAND2_X1 U11947 ( .A1(n9349), .A2(n13951), .ZN(n9351) );
  INV_X1 U11948 ( .A(n9350), .ZN(n9353) );
  INV_X1 U11949 ( .A(n9351), .ZN(n9352) );
  NAND2_X1 U11950 ( .A1(n9353), .A2(n9352), .ZN(n9354) );
  XNOR2_X1 U11951 ( .A(n9451), .B(n11656), .ZN(n9355) );
  NAND2_X1 U11952 ( .A1(n14241), .A2(n13950), .ZN(n9356) );
  NAND2_X1 U11953 ( .A1(n9355), .A2(n9356), .ZN(n9360) );
  INV_X1 U11954 ( .A(n9355), .ZN(n9358) );
  INV_X1 U11955 ( .A(n9356), .ZN(n9357) );
  NAND2_X1 U11956 ( .A1(n9358), .A2(n9357), .ZN(n9359) );
  AND2_X1 U11957 ( .A1(n9360), .A2(n9359), .ZN(n11546) );
  NAND2_X1 U11958 ( .A1(n11545), .A2(n9360), .ZN(n13816) );
  XNOR2_X1 U11959 ( .A(n9454), .B(n13821), .ZN(n9361) );
  NAND2_X1 U11960 ( .A1(n14241), .A2(n13949), .ZN(n9362) );
  NAND2_X1 U11961 ( .A1(n9361), .A2(n9362), .ZN(n9366) );
  INV_X1 U11962 ( .A(n9361), .ZN(n9364) );
  INV_X1 U11963 ( .A(n9362), .ZN(n9363) );
  NAND2_X1 U11964 ( .A1(n9364), .A2(n9363), .ZN(n9365) );
  AND2_X1 U11965 ( .A1(n9366), .A2(n9365), .ZN(n13817) );
  NAND2_X1 U11966 ( .A1(n13816), .A2(n13817), .ZN(n13815) );
  NAND2_X1 U11967 ( .A1(n13815), .A2(n9366), .ZN(n11518) );
  XNOR2_X1 U11968 ( .A(n11856), .B(n9454), .ZN(n9367) );
  NAND2_X1 U11969 ( .A1(n9349), .A2(n13948), .ZN(n9368) );
  XNOR2_X1 U11970 ( .A(n9367), .B(n9368), .ZN(n11517) );
  INV_X1 U11971 ( .A(n9367), .ZN(n9370) );
  INV_X1 U11972 ( .A(n9368), .ZN(n9369) );
  NAND2_X1 U11973 ( .A1(n9370), .A2(n9369), .ZN(n9371) );
  XNOR2_X1 U11974 ( .A(n11844), .B(n9451), .ZN(n9374) );
  NAND2_X1 U11975 ( .A1(n13947), .A2(n14241), .ZN(n9372) );
  XNOR2_X1 U11976 ( .A(n9374), .B(n9372), .ZN(n11796) );
  INV_X1 U11977 ( .A(n9372), .ZN(n9373) );
  XNOR2_X1 U11978 ( .A(n12159), .B(n9454), .ZN(n9375) );
  NAND2_X1 U11979 ( .A1(n13946), .A2(n9349), .ZN(n9376) );
  NAND2_X1 U11980 ( .A1(n9375), .A2(n9376), .ZN(n9380) );
  INV_X1 U11981 ( .A(n9375), .ZN(n9378) );
  INV_X1 U11982 ( .A(n9376), .ZN(n9377) );
  NAND2_X1 U11983 ( .A1(n9378), .A2(n9377), .ZN(n9379) );
  NAND2_X1 U11984 ( .A1(n9380), .A2(n9379), .ZN(n13767) );
  XNOR2_X1 U11985 ( .A(n13851), .B(n9454), .ZN(n9381) );
  NAND2_X1 U11986 ( .A1(n13944), .A2(n9349), .ZN(n9382) );
  NAND2_X1 U11987 ( .A1(n9381), .A2(n9382), .ZN(n9386) );
  INV_X1 U11988 ( .A(n9381), .ZN(n9384) );
  INV_X1 U11989 ( .A(n9382), .ZN(n9383) );
  NAND2_X1 U11990 ( .A1(n9384), .A2(n9383), .ZN(n9385) );
  AND2_X1 U11991 ( .A1(n9386), .A2(n9385), .ZN(n13845) );
  XNOR2_X1 U11992 ( .A(n13753), .B(n9454), .ZN(n9388) );
  NAND2_X1 U11993 ( .A1(n13943), .A2(n9349), .ZN(n9387) );
  XNOR2_X1 U11994 ( .A(n9388), .B(n9387), .ZN(n13747) );
  XNOR2_X1 U11995 ( .A(n14382), .B(n9454), .ZN(n9389) );
  NAND2_X1 U11996 ( .A1(n14241), .A2(n13942), .ZN(n9390) );
  NAND2_X1 U11997 ( .A1(n9389), .A2(n9390), .ZN(n9394) );
  INV_X1 U11998 ( .A(n9389), .ZN(n9392) );
  INV_X1 U11999 ( .A(n9390), .ZN(n9391) );
  NAND2_X1 U12000 ( .A1(n9392), .A2(n9391), .ZN(n9393) );
  NAND2_X1 U12001 ( .A1(n9394), .A2(n9393), .ZN(n13885) );
  XNOR2_X1 U12002 ( .A(n13793), .B(n9454), .ZN(n9395) );
  NAND2_X1 U12003 ( .A1(n13941), .A2(n9349), .ZN(n9396) );
  NAND2_X1 U12004 ( .A1(n9395), .A2(n9396), .ZN(n13784) );
  INV_X1 U12005 ( .A(n9395), .ZN(n9398) );
  INV_X1 U12006 ( .A(n9396), .ZN(n9397) );
  NAND2_X1 U12007 ( .A1(n9398), .A2(n9397), .ZN(n13785) );
  XNOR2_X1 U12008 ( .A(n14377), .B(n9454), .ZN(n9400) );
  NAND2_X1 U12009 ( .A1(n13939), .A2(n9349), .ZN(n13723) );
  XNOR2_X1 U12010 ( .A(n12589), .B(n9454), .ZN(n9401) );
  NAND2_X1 U12011 ( .A1(n13940), .A2(n14241), .ZN(n9402) );
  AND2_X1 U12012 ( .A1(n9401), .A2(n9402), .ZN(n13720) );
  AOI21_X1 U12013 ( .B1(n9400), .B2(n13723), .A(n13720), .ZN(n9399) );
  NAND2_X1 U12014 ( .A1(n13719), .A2(n9399), .ZN(n9408) );
  INV_X1 U12015 ( .A(n9400), .ZN(n13724) );
  INV_X1 U12016 ( .A(n9401), .ZN(n9404) );
  INV_X1 U12017 ( .A(n9402), .ZN(n9403) );
  NAND2_X1 U12018 ( .A1(n9404), .A2(n9403), .ZN(n13722) );
  NAND2_X1 U12019 ( .A1(n13722), .A2(n13723), .ZN(n9406) );
  NOR2_X1 U12020 ( .A1(n13722), .A2(n13723), .ZN(n9405) );
  AOI21_X1 U12021 ( .B1(n13724), .B2(n9406), .A(n9405), .ZN(n9407) );
  XNOR2_X1 U12022 ( .A(n14433), .B(n9454), .ZN(n9411) );
  NAND2_X1 U12023 ( .A1(n14241), .A2(n13938), .ZN(n13923) );
  NAND2_X1 U12024 ( .A1(n9411), .A2(n13923), .ZN(n9409) );
  XNOR2_X1 U12025 ( .A(n14245), .B(n9454), .ZN(n13806) );
  NAND2_X1 U12026 ( .A1(n13937), .A2(n14241), .ZN(n13807) );
  NAND2_X1 U12027 ( .A1(n13806), .A2(n13807), .ZN(n13827) );
  AND2_X1 U12028 ( .A1(n9409), .A2(n13827), .ZN(n9410) );
  NAND2_X1 U12029 ( .A1(n13805), .A2(n9410), .ZN(n9416) );
  XNOR2_X1 U12030 ( .A(n14222), .B(n9451), .ZN(n9417) );
  INV_X1 U12031 ( .A(n9349), .ZN(n9447) );
  NOR2_X1 U12032 ( .A1(n14198), .A2(n9447), .ZN(n9418) );
  XNOR2_X1 U12033 ( .A(n9417), .B(n9418), .ZN(n13828) );
  INV_X1 U12034 ( .A(n9411), .ZN(n13804) );
  INV_X1 U12035 ( .A(n13923), .ZN(n9412) );
  NAND3_X1 U12036 ( .A1(n13827), .A2(n13804), .A3(n9412), .ZN(n9413) );
  OAI21_X1 U12037 ( .B1(n13806), .B2(n13807), .A(n9413), .ZN(n9414) );
  NOR2_X1 U12038 ( .A1(n13828), .A2(n9414), .ZN(n9415) );
  INV_X1 U12039 ( .A(n9417), .ZN(n9420) );
  INV_X1 U12040 ( .A(n9418), .ZN(n9419) );
  NAND2_X1 U12041 ( .A1(n9420), .A2(n9419), .ZN(n9421) );
  XNOR2_X1 U12042 ( .A(n14209), .B(n9451), .ZN(n9424) );
  NOR2_X1 U12043 ( .A1(n10421), .A2(n9447), .ZN(n9423) );
  XNOR2_X1 U12044 ( .A(n9424), .B(n9423), .ZN(n13895) );
  INV_X1 U12045 ( .A(n13895), .ZN(n9422) );
  XNOR2_X1 U12046 ( .A(n14179), .B(n9454), .ZN(n9425) );
  OR2_X1 U12047 ( .A1(n14200), .A2(n9447), .ZN(n9426) );
  NAND2_X1 U12048 ( .A1(n9425), .A2(n9426), .ZN(n13757) );
  INV_X1 U12049 ( .A(n9425), .ZN(n9428) );
  INV_X1 U12050 ( .A(n9426), .ZN(n9427) );
  NAND2_X1 U12051 ( .A1(n9428), .A2(n9427), .ZN(n13756) );
  XNOR2_X1 U12052 ( .A(n14336), .B(n9454), .ZN(n9429) );
  NAND2_X1 U12053 ( .A1(n13933), .A2(n9349), .ZN(n9430) );
  NAND2_X1 U12054 ( .A1(n9429), .A2(n9430), .ZN(n13854) );
  INV_X1 U12055 ( .A(n9429), .ZN(n9432) );
  INV_X1 U12056 ( .A(n9430), .ZN(n9431) );
  NAND2_X1 U12057 ( .A1(n9432), .A2(n9431), .ZN(n13855) );
  XNOR2_X1 U12058 ( .A(n14151), .B(n9451), .ZN(n9435) );
  NAND2_X1 U12059 ( .A1(n13932), .A2(n14241), .ZN(n9433) );
  XNOR2_X1 U12060 ( .A(n9435), .B(n9433), .ZN(n13776) );
  INV_X1 U12061 ( .A(n9433), .ZN(n9434) );
  NAND2_X1 U12062 ( .A1(n9435), .A2(n9434), .ZN(n9436) );
  OR2_X1 U12063 ( .A1(n14113), .A2(n9447), .ZN(n13734) );
  INV_X1 U12064 ( .A(n13734), .ZN(n13874) );
  NOR2_X1 U12065 ( .A1(n13877), .A2(n9447), .ZN(n9440) );
  INV_X1 U12066 ( .A(n9439), .ZN(n13737) );
  INV_X1 U12067 ( .A(n9440), .ZN(n13741) );
  XNOR2_X1 U12068 ( .A(n14312), .B(n9454), .ZN(n9444) );
  NAND2_X1 U12069 ( .A1(n14081), .A2(n14241), .ZN(n9443) );
  NOR2_X1 U12070 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  AOI21_X1 U12071 ( .B1(n9444), .B2(n9443), .A(n9445), .ZN(n13836) );
  INV_X1 U12072 ( .A(n9445), .ZN(n9446) );
  XNOR2_X1 U12073 ( .A(n14089), .B(n9454), .ZN(n9449) );
  OR2_X1 U12074 ( .A1(n13913), .A2(n9447), .ZN(n9448) );
  NOR2_X1 U12075 ( .A1(n9449), .A2(n9448), .ZN(n9450) );
  AOI21_X1 U12076 ( .B1(n9449), .B2(n9448), .A(n9450), .ZN(n13797) );
  XNOR2_X1 U12077 ( .A(n14070), .B(n9451), .ZN(n9460) );
  NAND2_X1 U12078 ( .A1(n14083), .A2(n14241), .ZN(n9461) );
  XNOR2_X1 U12079 ( .A(n9460), .B(n9461), .ZN(n13908) );
  XNOR2_X1 U12080 ( .A(n14298), .B(n9451), .ZN(n9459) );
  INV_X1 U12081 ( .A(n9459), .ZN(n9453) );
  AND2_X1 U12082 ( .A1(n14065), .A2(n9349), .ZN(n9458) );
  INV_X1 U12083 ( .A(n9458), .ZN(n9452) );
  NOR2_X1 U12084 ( .A1(n9453), .A2(n9452), .ZN(n13709) );
  NAND2_X1 U12085 ( .A1(n14050), .A2(n9349), .ZN(n9455) );
  XNOR2_X1 U12086 ( .A(n9455), .B(n9454), .ZN(n9456) );
  XNOR2_X1 U12087 ( .A(n12678), .B(n9456), .ZN(n9465) );
  NOR2_X1 U12088 ( .A1(n9459), .A2(n9458), .ZN(n13710) );
  INV_X1 U12089 ( .A(n9460), .ZN(n9463) );
  INV_X1 U12090 ( .A(n9461), .ZN(n9462) );
  NOR2_X1 U12091 ( .A1(n9463), .A2(n9462), .ZN(n13708) );
  NOR2_X1 U12092 ( .A1(n13710), .A2(n13708), .ZN(n9464) );
  NAND2_X1 U12093 ( .A1(n9465), .A2(n9464), .ZN(n9469) );
  OR3_X1 U12094 ( .A1(n13710), .A2(n13708), .A3(n9465), .ZN(n9467) );
  XNOR2_X1 U12095 ( .A(n13709), .B(n9465), .ZN(n9466) );
  OAI21_X1 U12096 ( .B1(n13906), .B2(n9469), .A(n9468), .ZN(n9488) );
  NAND2_X1 U12097 ( .A1(n12141), .A2(n12598), .ZN(n9474) );
  INV_X1 U12098 ( .A(n12598), .ZN(n9472) );
  XNOR2_X1 U12099 ( .A(n12141), .B(P2_B_REG_SCAN_IN), .ZN(n9470) );
  NAND2_X1 U12100 ( .A1(n12382), .A2(n9470), .ZN(n9471) );
  INV_X1 U12101 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15461) );
  NAND2_X1 U12102 ( .A1(n15458), .A2(n15461), .ZN(n9473) );
  INV_X1 U12103 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15464) );
  NAND2_X1 U12104 ( .A1(n15458), .A2(n15464), .ZN(n9476) );
  NAND2_X1 U12105 ( .A1(n12382), .A2(n12598), .ZN(n9475) );
  NAND2_X1 U12106 ( .A1(n9476), .A2(n9475), .ZN(n15465) );
  INV_X1 U12107 ( .A(n15465), .ZN(n9486) );
  NOR4_X1 U12108 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n9480) );
  NOR4_X1 U12109 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9479) );
  NOR4_X1 U12110 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n9478) );
  NOR4_X1 U12111 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n9477) );
  NAND4_X1 U12112 ( .A1(n9480), .A2(n9479), .A3(n9478), .A4(n9477), .ZN(n9485)
         );
  NOR2_X1 U12113 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .ZN(
        n15606) );
  NOR4_X1 U12114 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n9483) );
  NOR4_X1 U12115 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n9482) );
  NOR4_X1 U12116 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9481) );
  NAND4_X1 U12117 ( .A1(n15606), .A2(n9483), .A3(n9482), .A4(n9481), .ZN(n9484) );
  NAND2_X1 U12118 ( .A1(n9486), .A2(n10442), .ZN(n11402) );
  NOR2_X1 U12119 ( .A1(n15479), .A2(n10856), .ZN(n9487) );
  OAI21_X1 U12120 ( .B1(n9489), .B2(n9488), .A(n13872), .ZN(n9505) );
  NOR2_X1 U12121 ( .A1(n11408), .A2(n11662), .ZN(n11613) );
  NAND2_X1 U12122 ( .A1(n9495), .A2(n11613), .ZN(n9491) );
  NAND2_X1 U12123 ( .A1(n13930), .A2(n14082), .ZN(n9493) );
  NAND2_X1 U12124 ( .A1(n14065), .A2(n14097), .ZN(n9492) );
  AND2_X1 U12125 ( .A1(n9493), .A2(n9492), .ZN(n10438) );
  INV_X1 U12126 ( .A(n9496), .ZN(n12677) );
  NAND2_X1 U12127 ( .A1(n10856), .A2(n9497), .ZN(n11404) );
  NAND2_X1 U12128 ( .A1(n11404), .A2(n10855), .ZN(n9498) );
  INV_X1 U12129 ( .A(n10978), .ZN(n9501) );
  NAND2_X1 U12130 ( .A1(n9499), .A2(n10443), .ZN(n9500) );
  NAND2_X1 U12131 ( .A1(n9501), .A2(n9500), .ZN(n11339) );
  AOI22_X1 U12132 ( .A1(n12677), .A2(n13917), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9502) );
  OAI21_X1 U12133 ( .B1(n10438), .B2(n13919), .A(n9502), .ZN(n9503) );
  AOI21_X1 U12134 ( .B1(n12678), .B2(n13926), .A(n9503), .ZN(n9504) );
  NAND2_X1 U12135 ( .A1(n9505), .A2(n9504), .ZN(P2_U3192) );
  NOR2_X2 U12136 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9507) );
  NOR2_X2 U12137 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9506) );
  AND4_X2 U12138 ( .A1(n9508), .A2(n9507), .A3(n9506), .A4(n9675), .ZN(n9511)
         );
  AND2_X2 U12139 ( .A1(n9510), .A2(n9509), .ZN(n9622) );
  NOR2_X1 U12140 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n9516) );
  NOR2_X1 U12141 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9515) );
  NOR2_X1 U12142 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9518) );
  NOR2_X1 U12143 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n9517) );
  OR2_X1 U12144 ( .A1(n9551), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9758) );
  INV_X1 U12145 ( .A(n9758), .ZN(n9528) );
  NAND2_X1 U12146 ( .A1(n9528), .A2(n9527), .ZN(n9776) );
  INV_X1 U12147 ( .A(n9776), .ZN(n9530) );
  INV_X1 U12148 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U12149 ( .A1(n9530), .A2(n9529), .ZN(n9762) );
  INV_X1 U12150 ( .A(n9789), .ZN(n9532) );
  INV_X1 U12151 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9531) );
  NAND2_X1 U12152 ( .A1(n9532), .A2(n9531), .ZN(n9817) );
  OAI21_X1 U12153 ( .B1(n9807), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9533) );
  XNOR2_X1 U12154 ( .A(n9533), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14682) );
  AOI22_X1 U12155 ( .A1(n14682), .A2(n9848), .B1(n9849), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n9534) );
  INV_X1 U12156 ( .A(n9640), .ZN(n9536) );
  XNOR2_X1 U12157 ( .A(n9853), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14875) );
  XNOR2_X2 U12158 ( .A(n9539), .B(n15135), .ZN(n9542) );
  NAND2_X1 U12159 ( .A1(n14875), .A2(n9966), .ZN(n9548) );
  INV_X1 U12160 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14876) );
  NAND2_X2 U12161 ( .A1(n15144), .A2(n9543), .ZN(n10029) );
  NAND2_X1 U12162 ( .A1(n9985), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9545) );
  AND2_X4 U12163 ( .A1(n12896), .A2(n9542), .ZN(n10027) );
  NAND2_X1 U12164 ( .A1(n10027), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9544) );
  OAI211_X1 U12165 ( .C1(n14876), .C2(n6403), .A(n9545), .B(n9544), .ZN(n9546)
         );
  INV_X1 U12166 ( .A(n9546), .ZN(n9547) );
  INV_X1 U12167 ( .A(n12722), .ZN(n9844) );
  NAND2_X1 U12168 ( .A1(n9552), .A2(n9560), .ZN(n9553) );
  NAND2_X1 U12169 ( .A1(n9556), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U12170 ( .A1(n9559), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9561) );
  NAND2_X1 U12171 ( .A1(n9562), .A2(n12939), .ZN(n10019) );
  INV_X1 U12172 ( .A(n9562), .ZN(n9565) );
  NAND2_X1 U12173 ( .A1(n9565), .A2(n10923), .ZN(n9566) );
  MUX2_X1 U12174 ( .A(n14889), .B(n7159), .S(n10045), .Z(n9845) );
  NAND2_X1 U12175 ( .A1(n10572), .A2(SI_0_), .ZN(n9568) );
  NAND2_X1 U12176 ( .A1(n9568), .A2(n9567), .ZN(n9570) );
  AND2_X1 U12177 ( .A1(n9570), .A2(n9569), .ZN(n15152) );
  MUX2_X1 U12178 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15152), .S(n10660), .Z(n10935) );
  INV_X1 U12179 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11902) );
  INV_X1 U12180 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9571) );
  INV_X1 U12181 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15247) );
  NAND2_X1 U12182 ( .A1(n11909), .A2(n14626), .ZN(n10082) );
  NAND2_X1 U12183 ( .A1(n10082), .A2(n10749), .ZN(n9572) );
  NAND2_X1 U12184 ( .A1(n9572), .A2(n10942), .ZN(n9573) );
  NAND2_X1 U12185 ( .A1(n9573), .A2(n9837), .ZN(n9584) );
  NAND2_X1 U12186 ( .A1(n10942), .A2(n10045), .ZN(n9583) );
  INV_X1 U12187 ( .A(n9574), .ZN(n10589) );
  INV_X1 U12188 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n15249) );
  INV_X1 U12189 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9575) );
  OR2_X1 U12190 ( .A1(n10660), .A2(n10700), .ZN(n9576) );
  NAND2_X1 U12191 ( .A1(n10027), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9582) );
  INV_X1 U12192 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9577) );
  OR2_X1 U12193 ( .A1(n10026), .A2(n9577), .ZN(n9581) );
  INV_X1 U12194 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10701) );
  OR2_X1 U12195 ( .A1(n6402), .A2(n10701), .ZN(n9580) );
  INV_X1 U12196 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U12197 ( .A1(n12007), .A2(n11152), .ZN(n10943) );
  NAND4_X1 U12198 ( .A1(n9584), .A2(n9583), .A3(n10943), .A4(n10944), .ZN(
        n9606) );
  NAND2_X1 U12199 ( .A1(n10027), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9586) );
  INV_X1 U12200 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10704) );
  INV_X1 U12201 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10694) );
  OR2_X1 U12202 ( .A1(n10029), .A2(n10694), .ZN(n9585) );
  INV_X1 U12203 ( .A(n9597), .ZN(n9588) );
  INV_X1 U12204 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U12205 ( .A1(n9598), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9589) );
  MUX2_X1 U12206 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9589), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9590) );
  INV_X1 U12207 ( .A(n9622), .ZN(n9619) );
  NAND2_X1 U12208 ( .A1(n10027), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9596) );
  INV_X1 U12209 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11751) );
  OR2_X1 U12210 ( .A1(n10026), .A2(n11751), .ZN(n9595) );
  INV_X1 U12211 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11745) );
  OR2_X1 U12212 ( .A1(n6401), .A2(n11745), .ZN(n9594) );
  INV_X1 U12213 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10693) );
  OR2_X1 U12214 ( .A1(n10029), .A2(n10693), .ZN(n9593) );
  AND4_X2 U12215 ( .A1(n9596), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n14623)
         );
  OR2_X1 U12216 ( .A1(n10015), .A2(n10667), .ZN(n9601) );
  OR2_X1 U12217 ( .A1(n9592), .A2(n10668), .ZN(n9600) );
  OR2_X1 U12218 ( .A1(n10660), .A2(n10766), .ZN(n9599) );
  AND3_X4 U12219 ( .A1(n9601), .A2(n9600), .A3(n9599), .ZN(n11225) );
  NAND2_X1 U12220 ( .A1(n14623), .A2(n11225), .ZN(n11590) );
  NAND2_X2 U12221 ( .A1(n11590), .A2(n9602), .ZN(n10946) );
  NAND2_X1 U12222 ( .A1(n11152), .A2(n10045), .ZN(n9603) );
  NAND2_X1 U12223 ( .A1(n11152), .A2(n11218), .ZN(n10084) );
  NAND2_X1 U12224 ( .A1(n9604), .A2(n10084), .ZN(n9605) );
  NAND4_X1 U12225 ( .A1(n9606), .A2(n11941), .A3(n10946), .A4(n9605), .ZN(
        n9618) );
  OR2_X1 U12226 ( .A1(n9837), .A2(n14623), .ZN(n9610) );
  NAND2_X1 U12227 ( .A1(n9837), .A2(n14623), .ZN(n9609) );
  NAND2_X1 U12228 ( .A1(n9609), .A2(n11754), .ZN(n9607) );
  INV_X1 U12229 ( .A(n15234), .ZN(n11952) );
  AOI21_X1 U12230 ( .B1(n9608), .B2(n9607), .A(n11952), .ZN(n9614) );
  OAI21_X1 U12231 ( .B1(n9609), .B2(n14622), .A(n11754), .ZN(n9612) );
  NAND2_X1 U12232 ( .A1(n9610), .A2(n11225), .ZN(n9611) );
  AOI21_X1 U12233 ( .B1(n9612), .B2(n9611), .A(n15234), .ZN(n9613) );
  NAND3_X1 U12234 ( .A1(n10045), .A2(n11952), .A3(n14622), .ZN(n9616) );
  NAND3_X1 U12235 ( .A1(n9837), .A2(n11596), .A3(n15234), .ZN(n9615) );
  NAND2_X1 U12236 ( .A1(n10565), .A2(n9591), .ZN(n9625) );
  NAND2_X1 U12237 ( .A1(n9619), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9620) );
  MUX2_X1 U12238 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9620), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9623) );
  INV_X1 U12239 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U12240 ( .A1(n9622), .A2(n9621), .ZN(n9659) );
  NAND2_X1 U12241 ( .A1(n9623), .A2(n9659), .ZN(n10774) );
  INV_X1 U12242 ( .A(n10774), .ZN(n10706) );
  AOI22_X1 U12243 ( .A1(n9849), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9848), .B2(
        n10706), .ZN(n9624) );
  NAND2_X1 U12244 ( .A1(n9625), .A2(n9624), .ZN(n11607) );
  NAND2_X1 U12245 ( .A1(n10027), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9630) );
  OAI21_X1 U12246 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n9640), .ZN(n11960) );
  OR2_X1 U12247 ( .A1(n10026), .A2(n11960), .ZN(n9629) );
  INV_X1 U12248 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10705) );
  OR2_X1 U12249 ( .A1(n6402), .A2(n10705), .ZN(n9628) );
  INV_X1 U12250 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9626) );
  OR2_X1 U12251 ( .A1(n10029), .A2(n9626), .ZN(n9627) );
  NAND4_X1 U12252 ( .A1(n9630), .A2(n9629), .A3(n9628), .A4(n9627), .ZN(n14621) );
  MUX2_X1 U12253 ( .A(n6406), .B(n14621), .S(n10045), .Z(n9634) );
  NAND2_X1 U12254 ( .A1(n9633), .A2(n9634), .ZN(n9632) );
  MUX2_X1 U12255 ( .A(n14621), .B(n6406), .S(n10045), .Z(n9631) );
  NAND2_X1 U12256 ( .A1(n9632), .A2(n9631), .ZN(n9638) );
  INV_X1 U12257 ( .A(n9633), .ZN(n9636) );
  INV_X1 U12258 ( .A(n9634), .ZN(n9635) );
  NAND2_X1 U12259 ( .A1(n9636), .A2(n9635), .ZN(n9637) );
  NAND2_X1 U12260 ( .A1(n10027), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9645) );
  INV_X1 U12261 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10695) );
  OR2_X1 U12262 ( .A1(n10029), .A2(n10695), .ZN(n9644) );
  INV_X1 U12263 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U12264 ( .A1(n9640), .A2(n9639), .ZN(n9641) );
  NAND2_X1 U12265 ( .A1(n9653), .A2(n9641), .ZN(n12046) );
  OR2_X1 U12266 ( .A1(n10026), .A2(n12046), .ZN(n9643) );
  INV_X1 U12267 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n12041) );
  OR2_X1 U12268 ( .A1(n6402), .A2(n12041), .ZN(n9642) );
  NAND4_X1 U12269 ( .A1(n9645), .A2(n9644), .A3(n9643), .A4(n9642), .ZN(n14620) );
  NAND2_X1 U12270 ( .A1(n10590), .A2(n9591), .ZN(n9648) );
  NAND2_X1 U12271 ( .A1(n9659), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9646) );
  XNOR2_X1 U12272 ( .A(n9646), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U12273 ( .A1(n9849), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9848), .B2(
        n10707), .ZN(n9647) );
  NAND2_X1 U12274 ( .A1(n9648), .A2(n9647), .ZN(n12045) );
  MUX2_X1 U12275 ( .A(n14620), .B(n12045), .S(n10045), .Z(n9650) );
  MUX2_X1 U12276 ( .A(n14620), .B(n12045), .S(n9837), .Z(n9649) );
  NAND2_X1 U12277 ( .A1(n9985), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9658) );
  INV_X1 U12278 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9651) );
  OR2_X1 U12279 ( .A1(n9988), .A2(n9651), .ZN(n9657) );
  INV_X1 U12280 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9652) );
  NAND2_X1 U12281 ( .A1(n9653), .A2(n9652), .ZN(n9654) );
  NAND2_X1 U12282 ( .A1(n9667), .A2(n9654), .ZN(n12013) );
  OR2_X1 U12283 ( .A1(n10026), .A2(n12013), .ZN(n9656) );
  INV_X1 U12284 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n12011) );
  OR2_X1 U12285 ( .A1(n6402), .A2(n12011), .ZN(n9655) );
  NAND4_X1 U12286 ( .A1(n9658), .A2(n9657), .A3(n9656), .A4(n9655), .ZN(n14619) );
  NAND2_X1 U12287 ( .A1(n10570), .A2(n9591), .ZN(n9662) );
  NAND2_X1 U12288 ( .A1(n9674), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9660) );
  XNOR2_X1 U12289 ( .A(n9660), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U12290 ( .A1(n9849), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9848), .B2(
        n10738), .ZN(n9661) );
  NAND2_X1 U12291 ( .A1(n9662), .A2(n9661), .ZN(n12012) );
  BUF_X1 U12292 ( .A(n9837), .Z(n9975) );
  MUX2_X1 U12293 ( .A(n14619), .B(n12012), .S(n9975), .Z(n9664) );
  MUX2_X1 U12294 ( .A(n14619), .B(n12012), .S(n10045), .Z(n9663) );
  INV_X1 U12295 ( .A(n9664), .ZN(n9665) );
  NAND2_X1 U12296 ( .A1(n9985), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9673) );
  INV_X1 U12297 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9666) );
  OR2_X1 U12298 ( .A1(n9988), .A2(n9666), .ZN(n9672) );
  NAND2_X1 U12299 ( .A1(n9667), .A2(n10744), .ZN(n9668) );
  NAND2_X1 U12300 ( .A1(n9685), .A2(n9668), .ZN(n12114) );
  OR2_X1 U12301 ( .A1(n10026), .A2(n12114), .ZN(n9671) );
  INV_X1 U12302 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9669) );
  OR2_X1 U12303 ( .A1(n6402), .A2(n9669), .ZN(n9670) );
  NAND4_X1 U12304 ( .A1(n9673), .A2(n9672), .A3(n9671), .A4(n9670), .ZN(n14618) );
  NAND2_X1 U12305 ( .A1(n10594), .A2(n9591), .ZN(n9679) );
  INV_X1 U12306 ( .A(n9674), .ZN(n9676) );
  NAND2_X1 U12307 ( .A1(n9676), .A2(n9675), .ZN(n9691) );
  NAND2_X1 U12308 ( .A1(n9691), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9677) );
  XNOR2_X1 U12309 ( .A(n9677), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U12310 ( .A1(n9849), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9848), .B2(
        n10838), .ZN(n9678) );
  NAND2_X1 U12311 ( .A1(n9679), .A2(n9678), .ZN(n15301) );
  MUX2_X1 U12312 ( .A(n14618), .B(n15301), .S(n10045), .Z(n9682) );
  MUX2_X1 U12313 ( .A(n14618), .B(n15301), .S(n9975), .Z(n9680) );
  INV_X1 U12314 ( .A(n9682), .ZN(n9683) );
  NAND2_X1 U12315 ( .A1(n10027), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9690) );
  INV_X1 U12316 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10836) );
  OR2_X1 U12317 ( .A1(n10029), .A2(n10836), .ZN(n9689) );
  NAND2_X1 U12318 ( .A1(n9685), .A2(n9684), .ZN(n9686) );
  NAND2_X1 U12319 ( .A1(n9705), .A2(n9686), .ZN(n12102) );
  OR2_X1 U12320 ( .A1(n10026), .A2(n12102), .ZN(n9688) );
  INV_X1 U12321 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n12097) );
  OR2_X1 U12322 ( .A1(n6403), .A2(n12097), .ZN(n9687) );
  NAND4_X1 U12323 ( .A1(n9690), .A2(n9689), .A3(n9688), .A4(n9687), .ZN(n14617) );
  NAND2_X1 U12324 ( .A1(n10653), .A2(n9591), .ZN(n9696) );
  INV_X1 U12325 ( .A(n9691), .ZN(n9693) );
  INV_X1 U12326 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9692) );
  NAND2_X1 U12327 ( .A1(n9693), .A2(n9692), .ZN(n9711) );
  NAND2_X1 U12328 ( .A1(n9711), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9694) );
  XNOR2_X1 U12329 ( .A(n9694), .B(P1_IR_REG_8__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U12330 ( .A1(n9849), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9848), .B2(
        n11001), .ZN(n9695) );
  NAND2_X1 U12331 ( .A1(n9696), .A2(n9695), .ZN(n12101) );
  MUX2_X1 U12332 ( .A(n14617), .B(n12101), .S(n9837), .Z(n9700) );
  MUX2_X1 U12333 ( .A(n14617), .B(n12101), .S(n10045), .Z(n9697) );
  NAND2_X1 U12334 ( .A1(n9698), .A2(n9697), .ZN(n9703) );
  INV_X1 U12335 ( .A(n9699), .ZN(n9701) );
  NAND2_X1 U12336 ( .A1(n9701), .A2(n6780), .ZN(n9702) );
  NAND2_X1 U12337 ( .A1(n10027), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9710) );
  INV_X1 U12338 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11069) );
  OR2_X1 U12339 ( .A1(n10029), .A2(n11069), .ZN(n9709) );
  NAND2_X1 U12340 ( .A1(n9705), .A2(n9704), .ZN(n9706) );
  NAND2_X1 U12341 ( .A1(n9724), .A2(n9706), .ZN(n12057) );
  OR2_X1 U12342 ( .A1(n10026), .A2(n12057), .ZN(n9708) );
  INV_X1 U12343 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n12055) );
  OR2_X1 U12344 ( .A1(n6403), .A2(n12055), .ZN(n9707) );
  NAND4_X1 U12345 ( .A1(n9710), .A2(n9709), .A3(n9708), .A4(n9707), .ZN(n14616) );
  NAND2_X1 U12346 ( .A1(n10677), .A2(n9591), .ZN(n9718) );
  NAND2_X1 U12347 ( .A1(n9713), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9716) );
  INV_X1 U12348 ( .A(n9713), .ZN(n9715) );
  INV_X1 U12349 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9714) );
  NAND2_X1 U12350 ( .A1(n9715), .A2(n9714), .ZN(n9730) );
  AOI22_X1 U12351 ( .A1(n9849), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11002), 
        .B2(n9848), .ZN(n9717) );
  MUX2_X1 U12352 ( .A(n14616), .B(n12183), .S(n10045), .Z(n9721) );
  MUX2_X1 U12353 ( .A(n14616), .B(n12183), .S(n9975), .Z(n9719) );
  INV_X1 U12354 ( .A(n9721), .ZN(n9722) );
  NAND2_X1 U12355 ( .A1(n9985), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9729) );
  INV_X1 U12356 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15722) );
  OR2_X1 U12357 ( .A1(n9988), .A2(n15722), .ZN(n9728) );
  INV_X1 U12358 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U12359 ( .A1(n9724), .A2(n9723), .ZN(n9725) );
  NAND2_X1 U12360 ( .A1(n9740), .A2(n9725), .ZN(n12271) );
  OR2_X1 U12361 ( .A1(n10026), .A2(n12271), .ZN(n9727) );
  INV_X1 U12362 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12189) );
  OR2_X1 U12363 ( .A1(n6402), .A2(n12189), .ZN(n9726) );
  NAND4_X1 U12364 ( .A1(n9729), .A2(n9728), .A3(n9727), .A4(n9726), .ZN(n14615) );
  NAND2_X1 U12365 ( .A1(n10686), .A2(n9591), .ZN(n9733) );
  NAND2_X1 U12366 ( .A1(n9730), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9731) );
  XNOR2_X1 U12367 ( .A(n9731), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U12368 ( .A1(n11393), .A2(n9848), .B1(n9849), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9732) );
  MUX2_X1 U12369 ( .A(n14615), .B(n12295), .S(n9975), .Z(n9736) );
  MUX2_X1 U12370 ( .A(n14615), .B(n12295), .S(n10045), .Z(n9734) );
  NAND2_X1 U12371 ( .A1(n9735), .A2(n9734), .ZN(n9739) );
  INV_X1 U12372 ( .A(n9736), .ZN(n9737) );
  NAND2_X1 U12373 ( .A1(n9740), .A2(n11391), .ZN(n9741) );
  NAND2_X1 U12374 ( .A1(n9753), .A2(n9741), .ZN(n12536) );
  OR2_X1 U12375 ( .A1(n12536), .A2(n10026), .ZN(n9745) );
  NAND2_X1 U12376 ( .A1(n10027), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9744) );
  INV_X1 U12377 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n12292) );
  OR2_X1 U12378 ( .A1(n6403), .A2(n12292), .ZN(n9743) );
  INV_X1 U12379 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11677) );
  OR2_X1 U12380 ( .A1(n10029), .A2(n11677), .ZN(n9742) );
  NAND4_X1 U12381 ( .A1(n9745), .A2(n9744), .A3(n9743), .A4(n9742), .ZN(n14614) );
  NAND2_X1 U12382 ( .A1(n10730), .A2(n9591), .ZN(n9749) );
  NAND2_X1 U12383 ( .A1(n9551), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9746) );
  MUX2_X1 U12384 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9746), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n9747) );
  AOI22_X1 U12385 ( .A1(n9849), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9848), 
        .B2(n11680), .ZN(n9748) );
  MUX2_X1 U12386 ( .A(n14614), .B(n12532), .S(n10045), .Z(n9751) );
  MUX2_X1 U12387 ( .A(n14614), .B(n12532), .S(n9975), .Z(n9750) );
  INV_X1 U12388 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n15731) );
  NAND2_X1 U12389 ( .A1(n9753), .A2(n15731), .ZN(n9754) );
  NAND2_X1 U12390 ( .A1(n9771), .A2(n9754), .ZN(n14496) );
  INV_X1 U12391 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12461) );
  OAI22_X1 U12392 ( .A1(n14496), .A2(n10026), .B1(n6403), .B2(n12461), .ZN(
        n9757) );
  INV_X1 U12393 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11675) );
  NOR2_X1 U12394 ( .A1(n10029), .A2(n11675), .ZN(n9756) );
  INV_X1 U12395 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n15728) );
  NOR2_X1 U12396 ( .A1(n9988), .A2(n15728), .ZN(n9755) );
  NAND2_X1 U12397 ( .A1(n9758), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9759) );
  MUX2_X1 U12398 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9759), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n9760) );
  NAND2_X1 U12399 ( .A1(n9760), .A2(n9776), .ZN(n11684) );
  INV_X1 U12400 ( .A(n11684), .ZN(n11975) );
  AOI22_X1 U12401 ( .A1(n9849), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9848), 
        .B2(n11975), .ZN(n9761) );
  INV_X1 U12402 ( .A(n15097), .ZN(n14503) );
  MUX2_X1 U12403 ( .A(n12770), .B(n14503), .S(n10045), .Z(n9782) );
  MUX2_X1 U12404 ( .A(n14613), .B(n15097), .S(n9837), .Z(n9781) );
  NAND2_X1 U12405 ( .A1(n10996), .A2(n9591), .ZN(n9765) );
  NAND2_X1 U12406 ( .A1(n9762), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9763) );
  XNOR2_X1 U12407 ( .A(n9763), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12657) );
  AOI22_X1 U12408 ( .A1(n9849), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9848), 
        .B2(n12657), .ZN(n9764) );
  NAND2_X2 U12409 ( .A1(n9765), .A2(n9764), .ZN(n15085) );
  NAND2_X1 U12410 ( .A1(n9773), .A2(n9766), .ZN(n9767) );
  NAND2_X1 U12411 ( .A1(n9795), .A2(n9767), .ZN(n14947) );
  AOI22_X1 U12412 ( .A1(n10027), .A2(P1_REG0_REG_14__SCAN_IN), .B1(n9985), 
        .B2(P1_REG1_REG_14__SCAN_IN), .ZN(n9769) );
  INV_X1 U12413 ( .A(n6403), .ZN(n9984) );
  NAND2_X1 U12414 ( .A1(n9984), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9768) );
  OAI211_X1 U12415 ( .C1(n14947), .C2(n10026), .A(n9769), .B(n9768), .ZN(
        n14612) );
  INV_X1 U12416 ( .A(n14612), .ZN(n14555) );
  NAND2_X1 U12417 ( .A1(n15085), .A2(n14555), .ZN(n9800) );
  AND2_X2 U12418 ( .A1(n12687), .A2(n9800), .ZN(n14958) );
  NAND2_X1 U12419 ( .A1(n9771), .A2(n9770), .ZN(n9772) );
  NAND2_X1 U12420 ( .A1(n9773), .A2(n9772), .ZN(n14557) );
  AOI22_X1 U12421 ( .A1(n10027), .A2(P1_REG0_REG_13__SCAN_IN), .B1(n9985), 
        .B2(P1_REG1_REG_13__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U12422 ( .A1(n9984), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9774) );
  OAI211_X1 U12423 ( .C1(n14557), .C2(n10026), .A(n9775), .B(n9774), .ZN(
        n14963) );
  INV_X1 U12424 ( .A(n14963), .ZN(n12779) );
  NAND2_X1 U12425 ( .A1(n10787), .A2(n9591), .ZN(n9779) );
  NAND2_X1 U12426 ( .A1(n9776), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9777) );
  XNOR2_X1 U12427 ( .A(n9777), .B(P1_IR_REG_13__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U12428 ( .A1(n9849), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9848), 
        .B2(n12388), .ZN(n9778) );
  NAND2_X2 U12429 ( .A1(n9779), .A2(n9778), .ZN(n15092) );
  INV_X1 U12430 ( .A(n15092), .ZN(n14563) );
  MUX2_X1 U12431 ( .A(n12779), .B(n14563), .S(n10045), .Z(n9785) );
  MUX2_X1 U12432 ( .A(n14963), .B(n15092), .S(n9975), .Z(n9780) );
  AOI22_X1 U12433 ( .A1(n9782), .A2(n9781), .B1(n9785), .B2(n9780), .ZN(n9783)
         );
  NAND2_X1 U12434 ( .A1(n14963), .A2(n10045), .ZN(n9788) );
  INV_X1 U12435 ( .A(n9785), .ZN(n9787) );
  NAND2_X1 U12436 ( .A1(n15092), .A2(n9975), .ZN(n9786) );
  NAND2_X1 U12437 ( .A1(n11060), .A2(n9591), .ZN(n9793) );
  NAND2_X1 U12438 ( .A1(n9789), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9790) );
  MUX2_X1 U12439 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9790), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n9791) );
  NAND2_X1 U12440 ( .A1(n9791), .A2(n9817), .ZN(n12658) );
  AOI22_X1 U12441 ( .A1(n15264), .A2(n9848), .B1(n9849), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n9792) );
  NAND2_X2 U12442 ( .A1(n9793), .A2(n9792), .ZN(n15078) );
  INV_X1 U12443 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15260) );
  INV_X1 U12444 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U12445 ( .A1(n9795), .A2(n9794), .ZN(n9796) );
  NAND2_X1 U12446 ( .A1(n9821), .A2(n9796), .ZN(n14593) );
  OR2_X1 U12447 ( .A1(n14593), .A2(n10026), .ZN(n9798) );
  AOI22_X1 U12448 ( .A1(n10027), .A2(P1_REG0_REG_15__SCAN_IN), .B1(n9985), 
        .B2(P1_REG1_REG_15__SCAN_IN), .ZN(n9797) );
  OAI211_X1 U12449 ( .C1(n6402), .C2(n15260), .A(n9798), .B(n9797), .ZN(n14961) );
  INV_X1 U12450 ( .A(n14961), .ZN(n14917) );
  OR2_X2 U12451 ( .A1(n15078), .A2(n14917), .ZN(n12688) );
  NAND2_X1 U12452 ( .A1(n12688), .A2(n12687), .ZN(n9799) );
  NAND2_X1 U12453 ( .A1(n9799), .A2(n9975), .ZN(n9803) );
  NAND2_X1 U12454 ( .A1(n15078), .A2(n14917), .ZN(n10089) );
  NAND2_X1 U12455 ( .A1(n10089), .A2(n9800), .ZN(n9801) );
  NAND2_X1 U12456 ( .A1(n9801), .A2(n10045), .ZN(n9802) );
  NAND2_X1 U12457 ( .A1(n9803), .A2(n9802), .ZN(n9804) );
  NAND2_X1 U12458 ( .A1(n11089), .A2(n9591), .ZN(n9810) );
  NAND2_X1 U12459 ( .A1(n9807), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9808) );
  XNOR2_X1 U12460 ( .A(n9808), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14671) );
  AOI22_X1 U12461 ( .A1(n14671), .A2(n9848), .B1(n9849), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n9809) );
  NAND2_X1 U12462 ( .A1(n6555), .A2(n6848), .ZN(n9811) );
  NAND2_X1 U12463 ( .A1(n9853), .A2(n9811), .ZN(n14891) );
  INV_X1 U12464 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14892) );
  NAND2_X1 U12465 ( .A1(n9985), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U12466 ( .A1(n10027), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9812) );
  OAI211_X1 U12467 ( .C1(n14892), .C2(n6402), .A(n9813), .B(n9812), .ZN(n9814)
         );
  INV_X1 U12468 ( .A(n9814), .ZN(n9815) );
  NOR2_X1 U12469 ( .A1(n14898), .A2(n14610), .ZN(n12719) );
  NAND2_X1 U12470 ( .A1(n14898), .A2(n14610), .ZN(n12718) );
  INV_X1 U12471 ( .A(n12718), .ZN(n9829) );
  NAND2_X1 U12472 ( .A1(n10992), .A2(n9591), .ZN(n9820) );
  NAND2_X1 U12473 ( .A1(n9817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9818) );
  XNOR2_X1 U12474 ( .A(n9818), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14654) );
  AOI22_X1 U12475 ( .A1(n14654), .A2(n9848), .B1(n9849), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U12476 ( .A1(n9821), .A2(n12671), .ZN(n9822) );
  AND2_X1 U12477 ( .A1(n6555), .A2(n9822), .ZN(n14919) );
  NAND2_X1 U12478 ( .A1(n14919), .A2(n9966), .ZN(n9827) );
  INV_X1 U12479 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14908) );
  NAND2_X1 U12480 ( .A1(n10027), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9824) );
  NAND2_X1 U12481 ( .A1(n9985), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9823) );
  OAI211_X1 U12482 ( .C1(n14908), .C2(n6403), .A(n9824), .B(n9823), .ZN(n9825)
         );
  INV_X1 U12483 ( .A(n9825), .ZN(n9826) );
  AND2_X1 U12484 ( .A1(n14887), .A2(n10045), .ZN(n9828) );
  AOI21_X1 U12485 ( .B1(n15073), .B2(n9837), .A(n9828), .ZN(n9834) );
  MUX2_X1 U12486 ( .A(n14887), .B(n15073), .S(n10045), .Z(n9833) );
  OAI22_X1 U12487 ( .A1(n12719), .A2(n9829), .B1(n9834), .B2(n9833), .ZN(n9830) );
  INV_X1 U12488 ( .A(n9830), .ZN(n9832) );
  MUX2_X1 U12489 ( .A(n10089), .B(n12688), .S(n10045), .Z(n9831) );
  NOR2_X1 U12490 ( .A1(n14898), .A2(n14915), .ZN(n14868) );
  INV_X1 U12491 ( .A(n9833), .ZN(n9836) );
  NAND2_X1 U12492 ( .A1(n14898), .A2(n14915), .ZN(n12692) );
  INV_X1 U12493 ( .A(n12692), .ZN(n10081) );
  INV_X1 U12494 ( .A(n9834), .ZN(n9835) );
  OR4_X1 U12495 ( .A1(n14868), .A2(n9836), .A3(n10081), .A4(n9835), .ZN(n9841)
         );
  AND2_X1 U12496 ( .A1(n14610), .A2(n9837), .ZN(n9839) );
  OAI21_X1 U12497 ( .B1(n9837), .B2(n14610), .A(n14898), .ZN(n9838) );
  OAI21_X1 U12498 ( .B1(n9839), .B2(n14898), .A(n9838), .ZN(n9840) );
  NAND3_X1 U12499 ( .A1(n9842), .A2(n9841), .A3(n9840), .ZN(n9843) );
  OAI21_X1 U12500 ( .B1(n9844), .B2(n9845), .A(n9843), .ZN(n9847) );
  NAND2_X1 U12501 ( .A1(n15058), .A2(n14889), .ZN(n12720) );
  NAND2_X1 U12502 ( .A1(n9845), .A2(n12720), .ZN(n9846) );
  NAND2_X1 U12503 ( .A1(n9847), .A2(n9846), .ZN(n9860) );
  AOI22_X1 U12504 ( .A1(n9849), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9848), 
        .B2(n7274), .ZN(n9850) );
  INV_X1 U12505 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n14575) );
  INV_X1 U12506 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9852) );
  OAI21_X1 U12507 ( .B1(n9853), .B2(n14575), .A(n9852), .ZN(n9854) );
  NAND2_X1 U12508 ( .A1(n9854), .A2(n9864), .ZN(n14858) );
  OR2_X1 U12509 ( .A1(n14858), .A2(n10026), .ZN(n9859) );
  INV_X1 U12510 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14857) );
  NAND2_X1 U12511 ( .A1(n9985), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U12512 ( .A1(n10027), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9855) );
  OAI211_X1 U12513 ( .C1(n14857), .C2(n6403), .A(n9856), .B(n9855), .ZN(n9857)
         );
  INV_X1 U12514 ( .A(n9857), .ZN(n9858) );
  NAND2_X1 U12515 ( .A1(n9859), .A2(n9858), .ZN(n14609) );
  INV_X1 U12516 ( .A(n14609), .ZN(n14866) );
  OR2_X1 U12517 ( .A1(n14861), .A2(n14866), .ZN(n9861) );
  NAND2_X1 U12518 ( .A1(n9860), .A2(n14853), .ZN(n9863) );
  MUX2_X1 U12519 ( .A(n12694), .B(n9861), .S(n9975), .Z(n9862) );
  NAND2_X1 U12520 ( .A1(n9863), .A2(n9862), .ZN(n9874) );
  NAND2_X1 U12521 ( .A1(n9864), .A2(n14546), .ZN(n9865) );
  NAND2_X1 U12522 ( .A1(n9876), .A2(n9865), .ZN(n14842) );
  INV_X1 U12523 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15655) );
  NAND2_X1 U12524 ( .A1(n9985), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U12525 ( .A1(n9984), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9866) );
  OAI211_X1 U12526 ( .C1(n9988), .C2(n15655), .A(n9867), .B(n9866), .ZN(n9868)
         );
  INV_X1 U12527 ( .A(n9868), .ZN(n9869) );
  INV_X1 U12528 ( .A(n14825), .ZN(n14490) );
  NAND2_X1 U12529 ( .A1(n11661), .A2(n9591), .ZN(n9871) );
  OR2_X1 U12530 ( .A1(n9592), .A2(n12933), .ZN(n9870) );
  NAND2_X2 U12531 ( .A1(n9871), .A2(n9870), .ZN(n15043) );
  MUX2_X1 U12532 ( .A(n14490), .B(n14846), .S(n9837), .Z(n9873) );
  MUX2_X1 U12533 ( .A(n14825), .B(n15043), .S(n10045), .Z(n9872) );
  INV_X1 U12534 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U12535 ( .A1(n9876), .A2(n9875), .ZN(n9877) );
  AND2_X1 U12536 ( .A1(n9890), .A2(n9877), .ZN(n14831) );
  NAND2_X1 U12537 ( .A1(n14831), .A2(n9966), .ZN(n9883) );
  INV_X1 U12538 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U12539 ( .A1(n9985), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9879) );
  NAND2_X1 U12540 ( .A1(n10027), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9878) );
  OAI211_X1 U12541 ( .C1(n9880), .C2(n6402), .A(n9879), .B(n9878), .ZN(n9881)
         );
  INV_X1 U12542 ( .A(n9881), .ZN(n9882) );
  NAND2_X1 U12543 ( .A1(n11689), .A2(n9591), .ZN(n9885) );
  OR2_X1 U12544 ( .A1(n9592), .A2(n12941), .ZN(n9884) );
  NAND2_X2 U12545 ( .A1(n9885), .A2(n9884), .ZN(n15036) );
  MUX2_X1 U12546 ( .A(n14608), .B(n15036), .S(n9975), .Z(n9887) );
  INV_X1 U12547 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U12548 ( .A1(n9890), .A2(n9889), .ZN(n9891) );
  NAND2_X1 U12549 ( .A1(n9903), .A2(n9891), .ZN(n14813) );
  INV_X1 U12550 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14812) );
  NAND2_X1 U12551 ( .A1(n10027), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9893) );
  NAND2_X1 U12552 ( .A1(n9985), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9892) );
  OAI211_X1 U12553 ( .C1(n14812), .C2(n6402), .A(n9893), .B(n9892), .ZN(n9894)
         );
  INV_X1 U12554 ( .A(n9894), .ZN(n9895) );
  XNOR2_X1 U12555 ( .A(n9898), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15150) );
  MUX2_X1 U12556 ( .A(n14826), .B(n15030), .S(n9837), .Z(n9900) );
  MUX2_X1 U12557 ( .A(n14826), .B(n15030), .S(n10045), .Z(n9899) );
  INV_X1 U12558 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U12559 ( .A1(n9903), .A2(n9902), .ZN(n9904) );
  AND2_X1 U12560 ( .A1(n9921), .A2(n9904), .ZN(n14796) );
  NAND2_X1 U12561 ( .A1(n14796), .A2(n9966), .ZN(n9910) );
  INV_X1 U12562 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9907) );
  NAND2_X1 U12563 ( .A1(n9985), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9906) );
  NAND2_X1 U12564 ( .A1(n10027), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9905) );
  OAI211_X1 U12565 ( .C1(n9907), .C2(n6403), .A(n9906), .B(n9905), .ZN(n9908)
         );
  INV_X1 U12566 ( .A(n9908), .ZN(n9909) );
  NAND2_X1 U12567 ( .A1(n11931), .A2(n9591), .ZN(n9912) );
  OR2_X1 U12568 ( .A1(n9592), .A2(n15719), .ZN(n9911) );
  MUX2_X1 U12569 ( .A(n14607), .B(n15025), .S(n10045), .Z(n9916) );
  MUX2_X1 U12570 ( .A(n14607), .B(n15025), .S(n9837), .Z(n9913) );
  NAND2_X1 U12571 ( .A1(n9914), .A2(n9913), .ZN(n9919) );
  INV_X1 U12572 ( .A(n9915), .ZN(n9917) );
  INV_X1 U12573 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9920) );
  NAND2_X1 U12574 ( .A1(n9921), .A2(n9920), .ZN(n9922) );
  NAND2_X1 U12575 ( .A1(n9934), .A2(n9922), .ZN(n14538) );
  INV_X1 U12576 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U12577 ( .A1(n9985), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U12578 ( .A1(n10027), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9923) );
  OAI211_X1 U12579 ( .C1(n9925), .C2(n6403), .A(n9924), .B(n9923), .ZN(n9926)
         );
  INV_X1 U12580 ( .A(n9926), .ZN(n9927) );
  NAND2_X1 U12581 ( .A1(n12138), .A2(n9591), .ZN(n9930) );
  OR2_X1 U12582 ( .A1(n9592), .A2(n12140), .ZN(n9929) );
  MUX2_X1 U12583 ( .A(n14606), .B(n14781), .S(n9837), .Z(n9932) );
  MUX2_X1 U12584 ( .A(n14606), .B(n14781), .S(n10045), .Z(n9931) );
  INV_X1 U12585 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U12586 ( .A1(n9934), .A2(n9933), .ZN(n9935) );
  NAND2_X1 U12587 ( .A1(n14764), .A2(n9966), .ZN(n9941) );
  INV_X1 U12588 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U12589 ( .A1(n9985), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U12590 ( .A1(n10027), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9936) );
  OAI211_X1 U12591 ( .C1(n9938), .C2(n6402), .A(n9937), .B(n9936), .ZN(n9939)
         );
  INV_X1 U12592 ( .A(n9939), .ZN(n9940) );
  NAND2_X1 U12593 ( .A1(n12381), .A2(n9591), .ZN(n9943) );
  OR2_X1 U12594 ( .A1(n9592), .A2(n12386), .ZN(n9942) );
  MUX2_X1 U12595 ( .A(n14605), .B(n15012), .S(n10045), .Z(n9947) );
  NAND2_X1 U12596 ( .A1(n9946), .A2(n9947), .ZN(n9945) );
  MUX2_X1 U12597 ( .A(n14605), .B(n15012), .S(n9975), .Z(n9944) );
  NAND2_X1 U12598 ( .A1(n9945), .A2(n9944), .ZN(n9951) );
  INV_X1 U12599 ( .A(n9946), .ZN(n9949) );
  INV_X1 U12600 ( .A(n9947), .ZN(n9948) );
  INV_X1 U12601 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U12602 ( .A1(n9953), .A2(n9952), .ZN(n9954) );
  NAND2_X1 U12603 ( .A1(n14747), .A2(n9966), .ZN(n9960) );
  INV_X1 U12604 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U12605 ( .A1(n9985), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U12606 ( .A1(n10027), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9955) );
  OAI211_X1 U12607 ( .C1(n9957), .C2(n6402), .A(n9956), .B(n9955), .ZN(n9958)
         );
  INV_X1 U12608 ( .A(n9958), .ZN(n9959) );
  NAND2_X1 U12609 ( .A1(n12596), .A2(n9591), .ZN(n9962) );
  OR2_X1 U12610 ( .A1(n9592), .A2(n12738), .ZN(n9961) );
  MUX2_X1 U12611 ( .A(n14604), .B(n14750), .S(n9975), .Z(n9964) );
  MUX2_X1 U12612 ( .A(n14604), .B(n14750), .S(n10045), .Z(n9963) );
  NAND2_X1 U12613 ( .A1(n14736), .A2(n9966), .ZN(n9972) );
  INV_X1 U12614 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U12615 ( .A1(n10027), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U12616 ( .A1(n9985), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9967) );
  OAI211_X1 U12617 ( .C1(n6403), .C2(n9969), .A(n9968), .B(n9967), .ZN(n9970)
         );
  INV_X1 U12618 ( .A(n9970), .ZN(n9971) );
  NAND2_X1 U12619 ( .A1(n12892), .A2(n9591), .ZN(n9974) );
  OR2_X1 U12620 ( .A1(n9592), .A2(n12893), .ZN(n9973) );
  MUX2_X1 U12621 ( .A(n14603), .B(n14737), .S(n10045), .Z(n9977) );
  MUX2_X1 U12622 ( .A(n14603), .B(n14737), .S(n9975), .Z(n9976) );
  INV_X1 U12623 ( .A(n9982), .ZN(n9979) );
  AND2_X1 U12624 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9978) );
  NAND2_X1 U12625 ( .A1(n9979), .A2(n9978), .ZN(n14718) );
  INV_X1 U12626 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9981) );
  INV_X1 U12627 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9980) );
  OAI21_X1 U12628 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(n9983) );
  NAND2_X1 U12629 ( .A1(n14718), .A2(n9983), .ZN(n12703) );
  INV_X1 U12630 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n15624) );
  NAND2_X1 U12631 ( .A1(n9984), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U12632 ( .A1(n9985), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9986) );
  OAI211_X1 U12633 ( .C1(n9988), .C2(n15624), .A(n9987), .B(n9986), .ZN(n9989)
         );
  INV_X1 U12634 ( .A(n9989), .ZN(n9990) );
  NAND2_X1 U12635 ( .A1(n14443), .A2(n9591), .ZN(n9993) );
  OR2_X1 U12636 ( .A1(n9592), .A2(n15148), .ZN(n9992) );
  MUX2_X1 U12637 ( .A(n14708), .B(n14991), .S(n9837), .Z(n9997) );
  NAND2_X1 U12638 ( .A1(n9996), .A2(n9997), .ZN(n9995) );
  MUX2_X1 U12639 ( .A(n14708), .B(n14991), .S(n10045), .Z(n9994) );
  INV_X1 U12640 ( .A(n9996), .ZN(n9999) );
  INV_X1 U12641 ( .A(n9997), .ZN(n9998) );
  NAND2_X1 U12642 ( .A1(n14438), .A2(n9591), .ZN(n10001) );
  INV_X1 U12643 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15136) );
  OR2_X1 U12644 ( .A1(n9592), .A2(n15136), .ZN(n10000) );
  NAND2_X1 U12645 ( .A1(n10027), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n10005) );
  INV_X1 U12646 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10002) );
  OR2_X1 U12647 ( .A1(n10029), .A2(n10002), .ZN(n10004) );
  INV_X1 U12648 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14694) );
  OR2_X1 U12649 ( .A1(n6402), .A2(n14694), .ZN(n10003) );
  INV_X1 U12650 ( .A(n14697), .ZN(n14601) );
  XNOR2_X1 U12651 ( .A(n14699), .B(n14601), .ZN(n10078) );
  NAND2_X1 U12652 ( .A1(n10006), .A2(n10007), .ZN(n10008) );
  NAND2_X1 U12653 ( .A1(n10970), .A2(n10008), .ZN(n10009) );
  NAND2_X1 U12654 ( .A1(n10749), .A2(n7274), .ZN(n11742) );
  NAND2_X1 U12655 ( .A1(n10009), .A2(n11742), .ZN(n10067) );
  INV_X1 U12656 ( .A(n10067), .ZN(n10010) );
  NAND2_X1 U12657 ( .A1(n10078), .A2(n10010), .ZN(n10058) );
  NAND2_X1 U12658 ( .A1(n10011), .A2(n10923), .ZN(n10925) );
  INV_X1 U12659 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14702) );
  NAND2_X1 U12660 ( .A1(n10027), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n10014) );
  INV_X1 U12661 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10012) );
  OR2_X1 U12662 ( .A1(n10029), .A2(n10012), .ZN(n10013) );
  OAI211_X1 U12663 ( .C1(n6403), .C2(n14702), .A(n10014), .B(n10013), .ZN(
        n14713) );
  OAI21_X1 U12664 ( .B1(n14601), .B2(n10925), .A(n14713), .ZN(n10018) );
  INV_X1 U12665 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15145) );
  OR2_X1 U12666 ( .A1(n9592), .A2(n15145), .ZN(n10016) );
  MUX2_X1 U12667 ( .A(n10018), .B(n14974), .S(n10045), .Z(n10047) );
  INV_X1 U12668 ( .A(n10047), .ZN(n10025) );
  INV_X1 U12669 ( .A(n14974), .ZN(n14705) );
  NAND2_X1 U12670 ( .A1(n14705), .A2(n9975), .ZN(n10023) );
  NAND2_X1 U12671 ( .A1(n10045), .A2(n14601), .ZN(n10020) );
  NAND2_X1 U12672 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  NAND2_X1 U12673 ( .A1(n10021), .A2(n14713), .ZN(n10022) );
  NAND2_X1 U12674 ( .A1(n10023), .A2(n10022), .ZN(n10046) );
  INV_X1 U12675 ( .A(n10046), .ZN(n10024) );
  AND2_X1 U12676 ( .A1(n10025), .A2(n10024), .ZN(n10061) );
  OR2_X1 U12677 ( .A1(n14718), .A2(n10026), .ZN(n10035) );
  INV_X1 U12678 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n14717) );
  NAND2_X1 U12679 ( .A1(n10027), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n10031) );
  INV_X1 U12680 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10028) );
  OR2_X1 U12681 ( .A1(n10029), .A2(n10028), .ZN(n10030) );
  OAI211_X1 U12682 ( .C1(n14717), .C2(n6402), .A(n10031), .B(n10030), .ZN(
        n10033) );
  INV_X1 U12683 ( .A(n10033), .ZN(n10034) );
  NAND2_X1 U12684 ( .A1(n10035), .A2(n10034), .ZN(n14602) );
  NAND2_X1 U12685 ( .A1(n12894), .A2(n9591), .ZN(n10037) );
  OR2_X1 U12686 ( .A1(n9592), .A2(n12895), .ZN(n10036) );
  MUX2_X1 U12687 ( .A(n14602), .B(n14986), .S(n10045), .Z(n10048) );
  INV_X1 U12688 ( .A(n10048), .ZN(n10040) );
  INV_X1 U12689 ( .A(n14602), .ZN(n10079) );
  MUX2_X1 U12690 ( .A(n10079), .B(n10038), .S(n9975), .Z(n10049) );
  INV_X1 U12691 ( .A(n10049), .ZN(n10039) );
  NOR2_X1 U12692 ( .A1(n10040), .A2(n10039), .ZN(n10055) );
  NAND2_X1 U12693 ( .A1(n10099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10042) );
  XNOR2_X1 U12694 ( .A(n10042), .B(n10041), .ZN(n10114) );
  INV_X1 U12695 ( .A(n10114), .ZN(n10659) );
  NAND2_X1 U12696 ( .A1(n10659), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11210) );
  NAND2_X1 U12697 ( .A1(n14699), .A2(n10045), .ZN(n10065) );
  NAND2_X1 U12698 ( .A1(n12939), .A2(n10923), .ZN(n10096) );
  AND2_X1 U12699 ( .A1(n10067), .A2(n10096), .ZN(n10062) );
  AND2_X1 U12700 ( .A1(n10047), .A2(n10046), .ZN(n10056) );
  NOR2_X1 U12701 ( .A1(n10049), .A2(n10048), .ZN(n10076) );
  INV_X1 U12702 ( .A(n10076), .ZN(n10051) );
  NAND2_X1 U12703 ( .A1(n10051), .A2(n10050), .ZN(n10052) );
  NOR2_X1 U12704 ( .A1(n10060), .A2(n10052), .ZN(n10053) );
  INV_X1 U12705 ( .A(n10054), .ZN(n10077) );
  INV_X1 U12706 ( .A(n10055), .ZN(n10059) );
  INV_X1 U12707 ( .A(n10056), .ZN(n10057) );
  OAI22_X1 U12708 ( .A1(n10060), .A2(n10059), .B1(n10058), .B2(n10057), .ZN(
        n10075) );
  INV_X1 U12709 ( .A(n10061), .ZN(n10072) );
  INV_X1 U12710 ( .A(n10062), .ZN(n10063) );
  NOR3_X1 U12711 ( .A1(n6978), .A2(n14601), .A3(n10063), .ZN(n10066) );
  NOR3_X1 U12712 ( .A1(n10065), .A2(n14601), .A3(n10067), .ZN(n10064) );
  AOI21_X1 U12713 ( .B1(n10066), .B2(n10065), .A(n10064), .ZN(n10071) );
  XNOR2_X1 U12714 ( .A(n10068), .B(n10067), .ZN(n10069) );
  NAND4_X1 U12715 ( .A1(n10069), .A2(n6978), .A3(n14601), .A4(n10096), .ZN(
        n10070) );
  OAI211_X1 U12716 ( .C1(n10073), .C2(n10072), .A(n10071), .B(n10070), .ZN(
        n10074) );
  AOI211_X1 U12717 ( .C1(n10077), .C2(n10076), .A(n10075), .B(n10074), .ZN(
        n10119) );
  INV_X1 U12718 ( .A(n10078), .ZN(n10095) );
  XOR2_X1 U12719 ( .A(n14713), .B(n14705), .Z(n10094) );
  XNOR2_X1 U12720 ( .A(n14991), .B(n14732), .ZN(n12707) );
  INV_X1 U12721 ( .A(n14728), .ZN(n10093) );
  XNOR2_X1 U12722 ( .A(n14750), .B(n14765), .ZN(n14745) );
  XNOR2_X1 U12723 ( .A(n15012), .B(n14605), .ZN(n14760) );
  NAND2_X1 U12724 ( .A1(n12756), .A2(n14826), .ZN(n10080) );
  XNOR2_X1 U12725 ( .A(n12295), .B(n12289), .ZN(n12187) );
  INV_X1 U12726 ( .A(n14616), .ZN(n12182) );
  XNOR2_X1 U12727 ( .A(n12183), .B(n12182), .ZN(n11888) );
  INV_X1 U12728 ( .A(n14617), .ZN(n11886) );
  XNOR2_X1 U12729 ( .A(n12101), .B(n11886), .ZN(n12095) );
  XNOR2_X1 U12730 ( .A(n15301), .B(n14618), .ZN(n12119) );
  XNOR2_X1 U12731 ( .A(n12045), .B(n11600), .ZN(n12036) );
  AND2_X1 U12732 ( .A1(n10942), .A2(n10082), .ZN(n10927) );
  OR2_X1 U12733 ( .A1(n11152), .A2(n11218), .ZN(n10083) );
  NAND2_X1 U12734 ( .A1(n10084), .A2(n10083), .ZN(n11017) );
  NAND4_X1 U12735 ( .A1(n10927), .A2(n11941), .A3(n10946), .A4(n11017), .ZN(
        n10085) );
  NOR3_X1 U12736 ( .A1(n12036), .A2(n10085), .A3(n11957), .ZN(n10086) );
  XNOR2_X1 U12737 ( .A(n12012), .B(n14619), .ZN(n11878) );
  NAND3_X1 U12738 ( .A1(n12119), .A2(n10086), .A3(n11878), .ZN(n10087) );
  OR4_X1 U12739 ( .A1(n12187), .A2(n11888), .A3(n12095), .A4(n10087), .ZN(
        n10088) );
  XNOR2_X1 U12740 ( .A(n15092), .B(n14963), .ZN(n12507) );
  INV_X1 U12741 ( .A(n12507), .ZN(n12708) );
  XNOR2_X1 U12742 ( .A(n12532), .B(n14614), .ZN(n12286) );
  OR4_X1 U12743 ( .A1(n10088), .A2(n12457), .A3(n12708), .A4(n12298), .ZN(
        n10090) );
  INV_X1 U12744 ( .A(n14958), .ZN(n12711) );
  INV_X1 U12745 ( .A(n14887), .ZN(n12690) );
  XNOR2_X1 U12746 ( .A(n15073), .B(n12690), .ZN(n14913) );
  AND4_X1 U12747 ( .A1(n14853), .A2(n7863), .A3(n12689), .A4(n14870), .ZN(
        n10091) );
  XNOR2_X1 U12748 ( .A(n15036), .B(n14608), .ZN(n14824) );
  XNOR2_X1 U12749 ( .A(n15043), .B(n14490), .ZN(n14837) );
  INV_X1 U12750 ( .A(n14837), .ZN(n14839) );
  XNOR2_X1 U12751 ( .A(n14781), .B(n14798), .ZN(n12699) );
  INV_X1 U12752 ( .A(n10096), .ZN(n10097) );
  NAND3_X1 U12753 ( .A1(n10098), .A2(n10050), .A3(n10097), .ZN(n10118) );
  NAND2_X1 U12754 ( .A1(n10109), .A2(n10111), .ZN(n10105) );
  NAND2_X1 U12755 ( .A1(n10105), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10106) );
  MUX2_X1 U12756 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10106), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n10108) );
  INV_X1 U12757 ( .A(n10109), .ZN(n10110) );
  NAND2_X1 U12758 ( .A1(n10110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10112) );
  INV_X1 U12759 ( .A(n10115), .ZN(n10756) );
  AND2_X1 U12760 ( .A1(n10007), .A2(n14716), .ZN(n10952) );
  NAND4_X1 U12761 ( .A1(n11740), .A2(n10756), .A3(n14962), .A4(n11206), .ZN(
        n10116) );
  OAI211_X1 U12762 ( .C1(n15151), .C2(n11210), .A(n10116), .B(P1_B_REG_SCAN_IN), .ZN(n10117) );
  OAI211_X1 U12763 ( .C1(n10119), .C2(n11210), .A(n10118), .B(n10117), .ZN(
        n10120) );
  INV_X1 U12764 ( .A(n10123), .ZN(n10124) );
  AOI21_X1 U12765 ( .B1(n6491), .B2(n11095), .A(n10124), .ZN(n10251) );
  INV_X1 U12766 ( .A(n10126), .ZN(n10142) );
  AND2_X1 U12767 ( .A1(n10126), .A2(n10125), .ZN(n10137) );
  NAND2_X1 U12768 ( .A1(n15534), .A2(n12342), .ZN(n10301) );
  NAND3_X1 U12769 ( .A1(n10131), .A2(n10301), .A3(n10338), .ZN(n10129) );
  NAND2_X1 U12770 ( .A1(n10129), .A2(n10301), .ZN(n10127) );
  MUX2_X1 U12771 ( .A(n15527), .B(n10127), .S(n11704), .Z(n10128) );
  INV_X1 U12772 ( .A(n10128), .ZN(n10135) );
  INV_X1 U12773 ( .A(n10129), .ZN(n10130) );
  INV_X2 U12774 ( .A(n6456), .ZN(n10335) );
  OAI21_X1 U12775 ( .B1(n10135), .B2(n10134), .A(n10133), .ZN(n10136) );
  OAI21_X1 U12776 ( .B1(n11095), .B2(n10137), .A(n10136), .ZN(n10140) );
  OAI21_X1 U12777 ( .B1(n11724), .B2(n10458), .A(n10139), .ZN(n10138) );
  NOR2_X1 U12778 ( .A1(n10335), .A2(n12311), .ZN(n10144) );
  INV_X1 U12779 ( .A(n12311), .ZN(n15566) );
  NOR2_X1 U12780 ( .A1(n11095), .A2(n15566), .ZN(n10143) );
  MUX2_X1 U12781 ( .A(n10144), .B(n10143), .S(n12355), .Z(n10146) );
  INV_X1 U12782 ( .A(n12167), .ZN(n10145) );
  NAND2_X1 U12783 ( .A1(n10151), .A2(n10147), .ZN(n10150) );
  INV_X1 U12784 ( .A(n10465), .ZN(n12163) );
  NAND2_X1 U12785 ( .A1(n13126), .A2(n12163), .ZN(n10148) );
  NAND2_X1 U12786 ( .A1(n10152), .A2(n10148), .ZN(n10149) );
  MUX2_X1 U12787 ( .A(n10150), .B(n10149), .S(n10335), .Z(n10154) );
  MUX2_X1 U12788 ( .A(n10152), .B(n10151), .S(n10335), .Z(n10153) );
  MUX2_X1 U12789 ( .A(n10156), .B(n10155), .S(n10335), .Z(n10157) );
  INV_X1 U12790 ( .A(n10157), .ZN(n10158) );
  NOR2_X1 U12791 ( .A1(n10158), .A2(n11836), .ZN(n10164) );
  INV_X1 U12792 ( .A(n11804), .ZN(n10162) );
  MUX2_X1 U12793 ( .A(n10160), .B(n10159), .S(n10335), .Z(n10161) );
  INV_X1 U12794 ( .A(n10165), .ZN(n10167) );
  MUX2_X1 U12795 ( .A(n10167), .B(n10166), .S(n11095), .Z(n10168) );
  NOR2_X1 U12796 ( .A1(n12346), .A2(n13122), .ZN(n10171) );
  MUX2_X1 U12797 ( .A(n10171), .B(n10170), .S(n10335), .Z(n10173) );
  INV_X1 U12798 ( .A(n12491), .ZN(n10172) );
  NAND2_X1 U12799 ( .A1(n10180), .A2(n10176), .ZN(n10178) );
  OAI21_X1 U12800 ( .B1(n13073), .B2(n12495), .A(n10179), .ZN(n10177) );
  MUX2_X1 U12801 ( .A(n10178), .B(n10177), .S(n11095), .Z(n10182) );
  MUX2_X1 U12802 ( .A(n10180), .B(n10179), .S(n10335), .Z(n10181) );
  INV_X1 U12803 ( .A(n10185), .ZN(n10184) );
  OAI22_X1 U12804 ( .A1(n10191), .A2(n10190), .B1(n10189), .B2(n10532), .ZN(
        n10192) );
  AOI21_X1 U12805 ( .B1(n10196), .B2(n10195), .A(n10532), .ZN(n10198) );
  NAND2_X1 U12806 ( .A1(n13498), .A2(n11095), .ZN(n10197) );
  INV_X1 U12807 ( .A(n10200), .ZN(n10201) );
  AOI21_X1 U12808 ( .B1(n10214), .B2(n10201), .A(n10532), .ZN(n10202) );
  NAND2_X1 U12809 ( .A1(n10203), .A2(n10202), .ZN(n10213) );
  INV_X1 U12810 ( .A(n10210), .ZN(n10205) );
  NAND2_X1 U12811 ( .A1(n10206), .A2(n10532), .ZN(n10207) );
  INV_X1 U12812 ( .A(n10208), .ZN(n10209) );
  MUX2_X1 U12813 ( .A(n10210), .B(n10209), .S(n10335), .Z(n10211) );
  XNOR2_X1 U12814 ( .A(n13641), .B(n13454), .ZN(n10220) );
  NOR3_X1 U12815 ( .A1(n13450), .A2(n10215), .A3(n10532), .ZN(n10221) );
  NOR3_X1 U12816 ( .A1(n10216), .A2(n11095), .A3(n13470), .ZN(n10219) );
  NOR2_X1 U12817 ( .A1(n10217), .A2(n10532), .ZN(n10218) );
  NOR4_X1 U12818 ( .A1(n10221), .A2(n10220), .A3(n10219), .A4(n10218), .ZN(
        n10227) );
  NAND2_X1 U12819 ( .A1(n10222), .A2(n10532), .ZN(n10224) );
  INV_X1 U12820 ( .A(n13428), .ZN(n10223) );
  OAI211_X1 U12821 ( .C1(n10335), .C2(n10225), .A(n10224), .B(n10223), .ZN(
        n10226) );
  NAND3_X1 U12822 ( .A1(n13630), .A2(n13431), .A3(n11095), .ZN(n10229) );
  INV_X1 U12823 ( .A(n13383), .ZN(n10233) );
  NOR2_X1 U12824 ( .A1(n13369), .A2(n10233), .ZN(n10232) );
  MUX2_X1 U12825 ( .A(n10233), .B(n10232), .S(n10335), .Z(n10234) );
  AOI21_X1 U12826 ( .B1(n10235), .B2(n13401), .A(n10234), .ZN(n10240) );
  INV_X1 U12827 ( .A(n10236), .ZN(n10243) );
  MUX2_X1 U12828 ( .A(n10238), .B(n13372), .S(n10335), .Z(n10239) );
  NAND2_X1 U12829 ( .A1(n13118), .A2(n11095), .ZN(n10241) );
  NOR2_X1 U12830 ( .A1(n13615), .A2(n10241), .ZN(n10242) );
  NOR2_X1 U12831 ( .A1(n13350), .A2(n10242), .ZN(n10247) );
  NAND4_X1 U12832 ( .A1(n10250), .A2(n10247), .A3(n10243), .A4(n10532), .ZN(
        n10249) );
  INV_X1 U12833 ( .A(n10251), .ZN(n10246) );
  AOI22_X1 U12834 ( .A1(n10251), .A2(n10244), .B1(n10247), .B2(n11095), .ZN(
        n10245) );
  OAI21_X1 U12835 ( .B1(n10247), .B2(n10246), .A(n10245), .ZN(n10248) );
  INV_X1 U12836 ( .A(n13354), .ZN(n10258) );
  NAND2_X1 U12837 ( .A1(n10259), .A2(n10258), .ZN(n10289) );
  INV_X1 U12838 ( .A(n10252), .ZN(n10253) );
  INV_X1 U12839 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12743) );
  XNOR2_X1 U12840 ( .A(n12743), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n10260) );
  XNOR2_X1 U12841 ( .A(n10261), .B(n10260), .ZN(n13691) );
  NAND2_X1 U12842 ( .A1(n13691), .A2(n8357), .ZN(n10257) );
  OR2_X1 U12843 ( .A1(n10265), .A2(n13693), .ZN(n10256) );
  AND2_X2 U12844 ( .A1(n10257), .A2(n10256), .ZN(n13607) );
  AND2_X1 U12845 ( .A1(n13607), .A2(n12619), .ZN(n10320) );
  NOR2_X1 U12846 ( .A1(n10259), .A2(n10258), .ZN(n10280) );
  OAI22_X1 U12847 ( .A1(n10261), .A2(n10260), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n15145), .ZN(n10263) );
  XNOR2_X1 U12848 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .ZN(n10262) );
  XNOR2_X1 U12849 ( .A(n10263), .B(n10262), .ZN(n13685) );
  NAND2_X1 U12850 ( .A1(n13685), .A2(n8357), .ZN(n10267) );
  INV_X1 U12851 ( .A(SI_31_), .ZN(n10264) );
  OR2_X1 U12852 ( .A1(n10265), .A2(n10264), .ZN(n10266) );
  NAND2_X1 U12853 ( .A1(n10268), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U12854 ( .A1(n10269), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10272) );
  NAND2_X1 U12855 ( .A1(n10270), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10271) );
  AND3_X1 U12856 ( .A1(n10273), .A2(n10272), .A3(n10271), .ZN(n10274) );
  OR2_X1 U12857 ( .A1(n10286), .A2(n13335), .ZN(n10279) );
  INV_X1 U12858 ( .A(n13607), .ZN(n10277) );
  INV_X1 U12859 ( .A(n12619), .ZN(n10276) );
  NAND2_X1 U12860 ( .A1(n10277), .A2(n10276), .ZN(n10278) );
  NAND2_X1 U12861 ( .A1(n10279), .A2(n10278), .ZN(n10283) );
  AND2_X1 U12862 ( .A1(n10286), .A2(n13335), .ZN(n10321) );
  NOR2_X1 U12863 ( .A1(n10281), .A2(n10280), .ZN(n10297) );
  INV_X1 U12864 ( .A(n10297), .ZN(n10295) );
  INV_X1 U12865 ( .A(n13335), .ZN(n13117) );
  OAI211_X1 U12866 ( .C1(n13607), .C2(n13117), .A(n13313), .B(n10289), .ZN(
        n10282) );
  NOR2_X1 U12867 ( .A1(n10283), .A2(n10282), .ZN(n10294) );
  INV_X1 U12868 ( .A(n10283), .ZN(n10324) );
  OR2_X1 U12869 ( .A1(n10286), .A2(n13313), .ZN(n10285) );
  AND2_X1 U12870 ( .A1(n13117), .A2(n13321), .ZN(n10287) );
  NAND2_X1 U12871 ( .A1(n7174), .A2(n10287), .ZN(n10284) );
  NAND2_X1 U12872 ( .A1(n10285), .A2(n10284), .ZN(n10296) );
  INV_X1 U12873 ( .A(n10296), .ZN(n10292) );
  AOI211_X1 U12874 ( .C1(n13607), .C2(n10289), .A(n13313), .B(n10286), .ZN(
        n10291) );
  INV_X1 U12875 ( .A(n10287), .ZN(n10288) );
  AOI21_X1 U12876 ( .B1(n10295), .B2(n10294), .A(n10293), .ZN(n10300) );
  NAND2_X1 U12877 ( .A1(n10297), .A2(n10296), .ZN(n10299) );
  NOR2_X1 U12878 ( .A1(n10321), .A2(n10448), .ZN(n10298) );
  INV_X1 U12879 ( .A(n13401), .ZN(n10317) );
  INV_X1 U12880 ( .A(n10301), .ZN(n10302) );
  NAND3_X1 U12881 ( .A1(n11540), .A2(n11709), .A3(n11722), .ZN(n10305) );
  INV_X1 U12882 ( .A(n15530), .ZN(n10303) );
  NAND2_X1 U12883 ( .A1(n10303), .A2(n10466), .ZN(n10304) );
  NOR2_X1 U12884 ( .A1(n10305), .A2(n10304), .ZN(n10307) );
  NAND4_X1 U12885 ( .A1(n10307), .A2(n12167), .A3(n12306), .A4(n10306), .ZN(
        n10308) );
  OR3_X1 U12886 ( .A1(n10308), .A2(n11836), .A3(n11804), .ZN(n10309) );
  NOR2_X1 U12887 ( .A1(n10309), .A2(n7637), .ZN(n10310) );
  NAND4_X1 U12888 ( .A1(n10311), .A2(n12468), .A3(n12491), .A4(n10310), .ZN(
        n10312) );
  NOR2_X1 U12889 ( .A1(n12564), .A2(n10312), .ZN(n10313) );
  NAND4_X1 U12890 ( .A1(n13482), .A2(n13535), .A3(n10313), .A4(n7624), .ZN(
        n10314) );
  NAND4_X1 U12891 ( .A1(n13416), .A2(n7857), .A3(n13446), .A4(n13438), .ZN(
        n10316) );
  INV_X1 U12892 ( .A(n10321), .ZN(n10322) );
  XNOR2_X1 U12893 ( .A(n10325), .B(n13321), .ZN(n10327) );
  INV_X1 U12894 ( .A(n10451), .ZN(n10326) );
  NAND2_X1 U12895 ( .A1(n10327), .A2(n10326), .ZN(n10328) );
  OR2_X1 U12896 ( .A1(n11094), .A2(P3_U3151), .ZN(n11783) );
  INV_X1 U12897 ( .A(n11783), .ZN(n10329) );
  NOR3_X1 U12898 ( .A1(n10538), .A2(n13214), .A3(n13701), .ZN(n10331) );
  OAI21_X1 U12899 ( .B1(n11783), .B2(n10338), .A(P3_B_REG_SCAN_IN), .ZN(n10330) );
  OR2_X1 U12900 ( .A1(n10331), .A2(n10330), .ZN(n10332) );
  NAND2_X1 U12901 ( .A1(n10333), .A2(n10332), .ZN(P3_U3296) );
  NAND2_X1 U12902 ( .A1(n10335), .A2(n10334), .ZN(n11695) );
  INV_X1 U12903 ( .A(n11697), .ZN(n13684) );
  NAND2_X1 U12904 ( .A1(n11695), .A2(n13684), .ZN(n11699) );
  OAI211_X1 U12905 ( .C1(n10338), .C2(n10337), .A(n10336), .B(n10448), .ZN(
        n10339) );
  NAND2_X1 U12906 ( .A1(n10339), .A2(n11697), .ZN(n10340) );
  NAND2_X1 U12907 ( .A1(n11699), .A2(n10340), .ZN(n10341) );
  NAND2_X1 U12908 ( .A1(n10341), .A2(n10532), .ZN(n10344) );
  INV_X1 U12909 ( .A(n11699), .ZN(n10342) );
  NAND2_X1 U12910 ( .A1(n10342), .A2(n10531), .ZN(n10343) );
  NAND2_X1 U12911 ( .A1(n10344), .A2(n10343), .ZN(n10349) );
  NAND3_X1 U12912 ( .A1(n10347), .A2(n10346), .A3(n10345), .ZN(n10348) );
  INV_X1 U12913 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10351) );
  NAND2_X1 U12914 ( .A1(n10259), .A2(n13590), .ZN(n10352) );
  NAND2_X1 U12915 ( .A1(n7853), .A2(n10352), .ZN(P3_U3488) );
  NAND2_X1 U12916 ( .A1(n13954), .A2(n11345), .ZN(n10983) );
  NAND2_X1 U12917 ( .A1(n10353), .A2(n10983), .ZN(n10982) );
  NAND3_X1 U12918 ( .A1(n10982), .A2(n11079), .A3(n11080), .ZN(n10356) );
  INV_X1 U12919 ( .A(n13951), .ZN(n11644) );
  NAND2_X1 U12920 ( .A1(n11644), .A2(n11414), .ZN(n10357) );
  INV_X1 U12921 ( .A(n13950), .ZN(n10393) );
  NAND2_X1 U12922 ( .A1(n10393), .A2(n11656), .ZN(n10358) );
  OR2_X1 U12923 ( .A1(n13821), .A2(n13949), .ZN(n10359) );
  OR2_X1 U12924 ( .A1(n11856), .A2(n13948), .ZN(n10360) );
  OR2_X1 U12925 ( .A1(n11844), .A2(n13947), .ZN(n10361) );
  INV_X1 U12926 ( .A(n12151), .ZN(n12146) );
  NAND2_X1 U12927 ( .A1(n12159), .A2(n13946), .ZN(n12212) );
  NAND2_X1 U12928 ( .A1(n13851), .A2(n13944), .ZN(n12540) );
  OR2_X1 U12929 ( .A1(n13851), .A2(n13944), .ZN(n10362) );
  NAND2_X1 U12930 ( .A1(n13753), .A2(n13943), .ZN(n10363) );
  AND2_X1 U12931 ( .A1(n14382), .A2(n13942), .ZN(n10365) );
  NAND2_X1 U12932 ( .A1(n13793), .A2(n13941), .ZN(n10366) );
  AND2_X1 U12933 ( .A1(n12589), .A2(n13940), .ZN(n10367) );
  NAND2_X1 U12934 ( .A1(n14377), .A2(n13939), .ZN(n10368) );
  INV_X1 U12935 ( .A(n14258), .ZN(n10370) );
  NAND2_X1 U12936 ( .A1(n14222), .A2(n13936), .ZN(n14191) );
  NAND2_X1 U12937 ( .A1(n14245), .A2(n13937), .ZN(n14190) );
  AND2_X1 U12938 ( .A1(n14191), .A2(n14190), .ZN(n10371) );
  NAND2_X1 U12939 ( .A1(n14189), .A2(n10371), .ZN(n10373) );
  INV_X1 U12940 ( .A(n10421), .ZN(n13935) );
  OR2_X1 U12941 ( .A1(n14209), .A2(n13935), .ZN(n10374) );
  NAND2_X1 U12942 ( .A1(n14179), .A2(n13934), .ZN(n10375) );
  OR2_X1 U12943 ( .A1(n14179), .A2(n13934), .ZN(n10376) );
  NAND2_X1 U12944 ( .A1(n14336), .A2(n13933), .ZN(n10378) );
  INV_X1 U12945 ( .A(n14113), .ZN(n13931) );
  NAND2_X1 U12946 ( .A1(n14138), .A2(n13931), .ZN(n10379) );
  NAND2_X1 U12947 ( .A1(n14312), .A2(n14081), .ZN(n10382) );
  NAND2_X1 U12948 ( .A1(n14089), .A2(n14096), .ZN(n10384) );
  INV_X1 U12949 ( .A(n14048), .ZN(n14054) );
  NAND2_X1 U12950 ( .A1(n14298), .A2(n14065), .ZN(n10385) );
  INV_X1 U12951 ( .A(n10435), .ZN(n10386) );
  AND2_X1 U12952 ( .A1(n14031), .A2(n11662), .ZN(n10388) );
  NAND2_X1 U12953 ( .A1(n11896), .A2(n10388), .ZN(n15484) );
  NAND2_X1 U12954 ( .A1(n10984), .A2(n10389), .ZN(n11621) );
  NAND2_X1 U12955 ( .A1(n11621), .A2(n11622), .ZN(n11620) );
  INV_X1 U12956 ( .A(n13952), .ZN(n11476) );
  NAND2_X1 U12957 ( .A1(n11476), .A2(n11619), .ZN(n10390) );
  NAND2_X1 U12958 ( .A1(n11644), .A2(n11667), .ZN(n10392) );
  NAND2_X1 U12959 ( .A1(n10393), .A2(n15478), .ZN(n10394) );
  NAND2_X1 U12960 ( .A1(n13821), .A2(n11645), .ZN(n10395) );
  INV_X1 U12961 ( .A(n13948), .ZN(n10396) );
  NAND2_X1 U12962 ( .A1(n11856), .A2(n10396), .ZN(n10397) );
  OR2_X1 U12963 ( .A1(n11844), .A2(n12152), .ZN(n10398) );
  NAND2_X1 U12964 ( .A1(n11844), .A2(n12152), .ZN(n10399) );
  OR2_X1 U12965 ( .A1(n12159), .A2(n12216), .ZN(n10400) );
  NAND2_X1 U12966 ( .A1(n12148), .A2(n10400), .ZN(n12214) );
  AOI22_X1 U12967 ( .A1(n13753), .A2(n12422), .B1(n12547), .B2(n13851), .ZN(
        n10401) );
  NAND2_X1 U12968 ( .A1(n12214), .A2(n10401), .ZN(n10407) );
  OR2_X1 U12969 ( .A1(n13851), .A2(n12547), .ZN(n12418) );
  NAND2_X1 U12970 ( .A1(n12418), .A2(n12422), .ZN(n10404) );
  NAND2_X1 U12971 ( .A1(n13943), .A2(n13944), .ZN(n10402) );
  NOR2_X1 U12972 ( .A1(n13851), .A2(n10402), .ZN(n10403) );
  AOI21_X1 U12973 ( .B1(n12555), .B2(n10404), .A(n10403), .ZN(n10405) );
  NAND2_X1 U12974 ( .A1(n14382), .A2(n10408), .ZN(n10409) );
  OR2_X1 U12975 ( .A1(n13793), .A2(n12583), .ZN(n10410) );
  OR2_X1 U12976 ( .A1(n14377), .A2(n12584), .ZN(n10413) );
  NAND2_X1 U12977 ( .A1(n12635), .A2(n10413), .ZN(n10415) );
  NAND2_X1 U12978 ( .A1(n14377), .A2(n12584), .ZN(n10414) );
  OR2_X1 U12979 ( .A1(n14433), .A2(n13811), .ZN(n10416) );
  OR2_X1 U12980 ( .A1(n14245), .A2(n10417), .ZN(n10418) );
  NOR2_X1 U12981 ( .A1(n14222), .A2(n14198), .ZN(n10420) );
  NAND2_X1 U12982 ( .A1(n14222), .A2(n14198), .ZN(n10419) );
  INV_X1 U12983 ( .A(n13933), .ZN(n10423) );
  NAND2_X1 U12984 ( .A1(n14336), .A2(n10423), .ZN(n10424) );
  INV_X1 U12985 ( .A(n13932), .ZN(n13876) );
  NAND2_X1 U12986 ( .A1(n14122), .A2(n13877), .ZN(n10427) );
  OR2_X1 U12987 ( .A1(n14122), .A2(n13877), .ZN(n10428) );
  NAND2_X1 U12988 ( .A1(n14312), .A2(n14114), .ZN(n14077) );
  NAND2_X1 U12989 ( .A1(n14089), .A2(n13913), .ZN(n14063) );
  AOI22_X1 U12990 ( .A1(n14070), .A2(n14083), .B1(n14404), .B2(n14096), .ZN(
        n10430) );
  INV_X1 U12991 ( .A(n14083), .ZN(n13800) );
  INV_X1 U12992 ( .A(n14065), .ZN(n10431) );
  AND2_X1 U12993 ( .A1(n14298), .A2(n10431), .ZN(n10432) );
  NAND2_X1 U12994 ( .A1(n8614), .A2(n11410), .ZN(n10433) );
  OAI21_X1 U12995 ( .B1(n10436), .B2(n10435), .A(n14252), .ZN(n10437) );
  NAND2_X1 U12997 ( .A1(n11616), .A2(n15472), .ZN(n11615) );
  INV_X1 U12998 ( .A(n13821), .ZN(n11632) );
  INV_X1 U12999 ( .A(n11856), .ZN(n15488) );
  INV_X1 U13000 ( .A(n14377), .ZN(n12642) );
  NAND2_X1 U13001 ( .A1(n14150), .A2(n14411), .ZN(n14135) );
  OR2_X2 U13002 ( .A1(n14135), .A2(n14122), .ZN(n14119) );
  AOI21_X1 U13003 ( .B1(n14052), .B2(n12678), .A(n14363), .ZN(n10441) );
  NAND2_X1 U13004 ( .A1(n10441), .A2(n12923), .ZN(n12681) );
  OAI21_X1 U13005 ( .B1(n12684), .B2(n14386), .A(n6499), .ZN(n14395) );
  NAND2_X1 U13006 ( .A1(n10443), .A2(n15465), .ZN(n10976) );
  NAND2_X1 U13007 ( .A1(n15500), .A2(n9238), .ZN(n10446) );
  INV_X1 U13008 ( .A(n12678), .ZN(n14398) );
  NAND2_X1 U13009 ( .A1(n10447), .A2(n7854), .ZN(P2_U3527) );
  NAND2_X1 U13010 ( .A1(n11704), .A2(n11555), .ZN(n10449) );
  XNOR2_X1 U13011 ( .A(n13552), .B(n10509), .ZN(n12903) );
  NOR2_X1 U13012 ( .A1(n12903), .A2(n13379), .ZN(n12898) );
  AOI21_X1 U13013 ( .B1(n12903), .B2(n13379), .A(n12898), .ZN(n10514) );
  XNOR2_X1 U13014 ( .A(n13635), .B(n6400), .ZN(n12953) );
  XNOR2_X1 U13015 ( .A(n12346), .B(n6399), .ZN(n10476) );
  XNOR2_X1 U13016 ( .A(n10459), .B(n10452), .ZN(n10461) );
  INV_X1 U13017 ( .A(n10453), .ZN(n10457) );
  NOR2_X1 U13018 ( .A1(n10459), .A2(n15526), .ZN(n10456) );
  XNOR2_X1 U13019 ( .A(n10459), .B(n10458), .ZN(n10460) );
  XNOR2_X1 U13020 ( .A(n10460), .B(n15536), .ZN(n11560) );
  NAND2_X1 U13021 ( .A1(n11559), .A2(n11560), .ZN(n11558) );
  XNOR2_X1 U13022 ( .A(n10461), .B(n13128), .ZN(n12352) );
  NAND2_X1 U13023 ( .A1(n10460), .A2(n11724), .ZN(n12353) );
  XNOR2_X1 U13024 ( .A(n6399), .B(n12311), .ZN(n10462) );
  NAND2_X1 U13025 ( .A1(n10462), .A2(n12355), .ZN(n10463) );
  OAI21_X1 U13026 ( .B1(n10462), .B2(n12355), .A(n10463), .ZN(n12123) );
  INV_X1 U13027 ( .A(n10463), .ZN(n10464) );
  XNOR2_X1 U13028 ( .A(n6399), .B(n10465), .ZN(n10467) );
  XNOR2_X1 U13029 ( .A(n10467), .B(n12328), .ZN(n11759) );
  XNOR2_X1 U13030 ( .A(n6399), .B(n12338), .ZN(n10470) );
  XNOR2_X1 U13031 ( .A(n10470), .B(n12205), .ZN(n12478) );
  XNOR2_X1 U13032 ( .A(n10466), .B(n10509), .ZN(n12204) );
  XNOR2_X1 U13033 ( .A(n6399), .B(n11717), .ZN(n12202) );
  NAND2_X1 U13034 ( .A1(n10467), .A2(n12328), .ZN(n12200) );
  OAI21_X1 U13035 ( .B1(n12202), .B2(n13125), .A(n12200), .ZN(n10468) );
  NOR4_X1 U13036 ( .A1(n11758), .A2(n12478), .A3(n12204), .A4(n10468), .ZN(
        n10475) );
  INV_X1 U13037 ( .A(n12478), .ZN(n10469) );
  AND2_X1 U13038 ( .A1(n12202), .A2(n13125), .ZN(n12203) );
  AOI21_X1 U13039 ( .B1(n10469), .B2(n12203), .A(n12204), .ZN(n10473) );
  INV_X1 U13040 ( .A(n12204), .ZN(n12476) );
  AOI21_X1 U13041 ( .B1(n10469), .B2(n13124), .A(n12476), .ZN(n10472) );
  INV_X1 U13042 ( .A(n10470), .ZN(n10471) );
  OAI22_X1 U13043 ( .A1(n10473), .A2(n10472), .B1(n13034), .B2(n10471), .ZN(
        n10474) );
  XNOR2_X1 U13044 ( .A(n6400), .B(n13038), .ZN(n10477) );
  XNOR2_X1 U13045 ( .A(n10477), .B(n13123), .ZN(n13030) );
  XNOR2_X1 U13046 ( .A(n10476), .B(n13033), .ZN(n10550) );
  INV_X1 U13047 ( .A(n13123), .ZN(n12233) );
  NAND2_X1 U13048 ( .A1(n10477), .A2(n12233), .ZN(n10551) );
  XNOR2_X1 U13049 ( .A(n13601), .B(n10509), .ZN(n12977) );
  XNOR2_X1 U13050 ( .A(n12988), .B(n6400), .ZN(n12982) );
  AOI22_X1 U13051 ( .A1(n12982), .A2(n13076), .B1(n13073), .B2(n12977), .ZN(
        n10478) );
  INV_X1 U13052 ( .A(n12982), .ZN(n10480) );
  XNOR2_X1 U13053 ( .A(n13058), .B(n6399), .ZN(n10481) );
  NAND2_X1 U13054 ( .A1(n10481), .A2(n12948), .ZN(n13051) );
  NAND2_X1 U13055 ( .A1(n13053), .A2(n13051), .ZN(n10483) );
  INV_X1 U13056 ( .A(n10481), .ZN(n10482) );
  NAND2_X1 U13057 ( .A1(n10482), .A2(n13537), .ZN(n13052) );
  NAND2_X1 U13058 ( .A1(n10483), .A2(n13052), .ZN(n12945) );
  XNOR2_X1 U13059 ( .A(n13680), .B(n6400), .ZN(n10484) );
  XNOR2_X1 U13060 ( .A(n10484), .B(n13121), .ZN(n12946) );
  XNOR2_X1 U13061 ( .A(n13669), .B(n10459), .ZN(n10485) );
  XNOR2_X1 U13062 ( .A(n10485), .B(n13538), .ZN(n13106) );
  XNOR2_X1 U13063 ( .A(n13585), .B(n10509), .ZN(n13003) );
  INV_X1 U13064 ( .A(n13003), .ZN(n10486) );
  XNOR2_X1 U13065 ( .A(n13660), .B(n6400), .ZN(n10487) );
  XNOR2_X1 U13066 ( .A(n10487), .B(n13487), .ZN(n13011) );
  INV_X1 U13067 ( .A(n10487), .ZN(n10488) );
  NAND2_X1 U13068 ( .A1(n10488), .A2(n13487), .ZN(n10489) );
  XNOR2_X1 U13069 ( .A(n13580), .B(n6400), .ZN(n13081) );
  NAND2_X1 U13070 ( .A1(n13081), .A2(n13501), .ZN(n10490) );
  NAND2_X1 U13071 ( .A1(n13083), .A2(n10490), .ZN(n10493) );
  INV_X1 U13072 ( .A(n13081), .ZN(n10491) );
  NAND2_X1 U13073 ( .A1(n10491), .A2(n13469), .ZN(n10492) );
  NAND2_X1 U13074 ( .A1(n10493), .A2(n10492), .ZN(n12964) );
  XNOR2_X1 U13075 ( .A(n13462), .B(n6399), .ZN(n10494) );
  XNOR2_X1 U13076 ( .A(n10494), .B(n13085), .ZN(n12963) );
  NAND2_X1 U13077 ( .A1(n10494), .A2(n13488), .ZN(n10495) );
  XNOR2_X1 U13078 ( .A(n13646), .B(n6399), .ZN(n10496) );
  XNOR2_X1 U13079 ( .A(n10496), .B(n13470), .ZN(n13043) );
  INV_X1 U13080 ( .A(n10496), .ZN(n10497) );
  NAND2_X1 U13081 ( .A1(n10497), .A2(n13470), .ZN(n10498) );
  XNOR2_X1 U13082 ( .A(n13641), .B(n6400), .ZN(n10499) );
  NAND2_X1 U13083 ( .A1(n10499), .A2(n13454), .ZN(n10500) );
  OAI21_X1 U13084 ( .B1(n10499), .B2(n13454), .A(n10500), .ZN(n12971) );
  OAI21_X1 U13085 ( .B1(n13418), .B2(n12953), .A(n12954), .ZN(n10504) );
  XNOR2_X1 U13086 ( .A(n13630), .B(n6399), .ZN(n12956) );
  AOI22_X1 U13087 ( .A1(n12956), .A2(n13431), .B1(n13418), .B2(n12953), .ZN(
        n10503) );
  XNOR2_X1 U13088 ( .A(n13565), .B(n10509), .ZN(n10501) );
  NOR2_X1 U13089 ( .A1(n10501), .A2(n13119), .ZN(n12995) );
  AOI21_X1 U13090 ( .B1(n10501), .B2(n13119), .A(n12995), .ZN(n13019) );
  OAI21_X1 U13091 ( .B1(n13431), .B2(n12956), .A(n13019), .ZN(n10502) );
  XNOR2_X1 U13092 ( .A(n12992), .B(n6399), .ZN(n10505) );
  NAND2_X1 U13093 ( .A1(n10505), .A2(n13404), .ZN(n10508) );
  INV_X1 U13094 ( .A(n10505), .ZN(n10506) );
  NAND2_X1 U13095 ( .A1(n10506), .A2(n13378), .ZN(n10507) );
  AND2_X1 U13096 ( .A1(n10508), .A2(n10507), .ZN(n12994) );
  NAND2_X1 U13097 ( .A1(n12993), .A2(n10508), .ZN(n13093) );
  XNOR2_X1 U13098 ( .A(n13615), .B(n10509), .ZN(n10510) );
  NOR2_X1 U13099 ( .A1(n10510), .A2(n13118), .ZN(n10511) );
  AOI21_X1 U13100 ( .B1(n10510), .B2(n13118), .A(n10511), .ZN(n13094) );
  NAND2_X1 U13101 ( .A1(n13093), .A2(n13094), .ZN(n13092) );
  INV_X1 U13102 ( .A(n10511), .ZN(n10512) );
  NAND2_X1 U13103 ( .A1(n13092), .A2(n10512), .ZN(n10513) );
  NAND2_X1 U13104 ( .A1(n10513), .A2(n10514), .ZN(n12909) );
  OAI21_X1 U13105 ( .B1(n10514), .B2(n10513), .A(n12909), .ZN(n10518) );
  NAND3_X1 U13106 ( .A1(n10529), .A2(n10527), .A3(n15567), .ZN(n10515) );
  OAI21_X1 U13107 ( .B1(n10524), .B2(n10525), .A(n10515), .ZN(n10517) );
  INV_X1 U13108 ( .A(n11098), .ZN(n10516) );
  NAND2_X1 U13109 ( .A1(n10518), .A2(n13095), .ZN(n10544) );
  INV_X1 U13110 ( .A(n13552), .ZN(n13366) );
  NOR2_X1 U13111 ( .A1(n10527), .A2(n15507), .ZN(n10519) );
  INV_X1 U13112 ( .A(n10522), .ZN(n10520) );
  NAND2_X1 U13113 ( .A1(n10537), .A2(n10520), .ZN(n10521) );
  NAND2_X1 U13114 ( .A1(n10537), .A2(n10522), .ZN(n10523) );
  INV_X1 U13115 ( .A(n10524), .ZN(n10526) );
  NAND2_X1 U13116 ( .A1(n10526), .A2(n10525), .ZN(n10534) );
  INV_X1 U13117 ( .A(n10527), .ZN(n10528) );
  NAND2_X1 U13118 ( .A1(n10529), .A2(n10528), .ZN(n10533) );
  INV_X1 U13119 ( .A(n10530), .ZN(n10547) );
  NAND4_X1 U13120 ( .A1(n10534), .A2(n10533), .A3(n10547), .A4(n11696), .ZN(
        n10535) );
  NAND2_X1 U13121 ( .A1(n10535), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13122 ( .A1(n13364), .A2(n13111), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10539) );
  OAI21_X1 U13123 ( .B1(n13387), .B2(n13098), .A(n10539), .ZN(n10540) );
  AOI21_X1 U13124 ( .B1(n12633), .B2(n13100), .A(n10540), .ZN(n10541) );
  INV_X1 U13125 ( .A(n10542), .ZN(n10543) );
  NAND2_X1 U13126 ( .A1(n10544), .A2(n10543), .ZN(P3_U3154) );
  AND2_X1 U13127 ( .A1(n10545), .A2(n10855), .ZN(n10858) );
  INV_X1 U13128 ( .A(n10587), .ZN(n10546) );
  INV_X1 U13129 ( .A(n10548), .ZN(n10553) );
  AOI21_X1 U13130 ( .B1(n10549), .B2(n10551), .A(n10550), .ZN(n10552) );
  NOR3_X1 U13131 ( .A1(n10553), .A2(n10552), .A3(n13115), .ZN(n10558) );
  NOR2_X1 U13132 ( .A1(n13103), .A2(n12346), .ZN(n10557) );
  AND2_X1 U13133 ( .A1(n13045), .A2(n12344), .ZN(n10556) );
  NAND2_X1 U13134 ( .A1(n13107), .A2(n13123), .ZN(n10554) );
  NAND2_X1 U13135 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n12072)
         );
  OAI211_X1 U13136 ( .C1(n13073), .C2(n13109), .A(n10554), .B(n12072), .ZN(
        n10555) );
  OR4_X1 U13137 ( .A1(n10558), .A2(n10557), .A3(n10556), .A4(n10555), .ZN(
        P3_U3157) );
  INV_X1 U13138 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10560) );
  NAND2_X1 U13139 ( .A1(n10559), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10630) );
  AOI21_X1 U13140 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n10560), .A(n7182), .ZN(
        n10561) );
  INV_X1 U13141 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15636) );
  NOR2_X1 U13142 ( .A1(n10561), .A2(n15636), .ZN(n15756) );
  AOI21_X1 U13143 ( .B1(n10561), .B2(n15636), .A(n15756), .ZN(SUB_1596_U53) );
  NAND2_X1 U13144 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_STATE_REG_SCAN_IN), .ZN(
        n10562) );
  OAI21_X1 U13145 ( .B1(n10563), .B2(P3_STATE_REG_SCAN_IN), .A(n10562), .ZN(
        P3_U3295) );
  AND2_X1 U13146 ( .A1(n10572), .A2(P2_U3088), .ZN(n14445) );
  INV_X2 U13147 ( .A(n14445), .ZN(n12742) );
  OAI222_X1 U13148 ( .A1(n12742), .A2(n7178), .B1(n14447), .B2(n6871), .C1(
        P2_U3088), .C2(n10877), .ZN(P2_U3324) );
  INV_X1 U13149 ( .A(n10565), .ZN(n10669) );
  INV_X1 U13150 ( .A(n10896), .ZN(n10884) );
  OAI222_X1 U13151 ( .A1(n12742), .A2(n10566), .B1(n14447), .B2(n10669), .C1(
        P2_U3088), .C2(n10884), .ZN(P2_U3323) );
  AND2_X1 U13152 ( .A1(n10567), .A2(P1_U3086), .ZN(n11934) );
  INV_X2 U13153 ( .A(n11934), .ZN(n15149) );
  OAI222_X1 U13154 ( .A1(n15149), .A2(n10568), .B1(n15141), .B2(n6871), .C1(
        P1_U3086), .C2(n14639), .ZN(P1_U3352) );
  OAI222_X1 U13155 ( .A1(n10700), .A2(P1_U3086), .B1(n15141), .B2(n10589), 
        .C1(n10569), .C2(n15149), .ZN(P1_U3354) );
  INV_X1 U13156 ( .A(n10570), .ZN(n10671) );
  INV_X1 U13157 ( .A(n11039), .ZN(n10904) );
  OAI222_X1 U13158 ( .A1(n12742), .A2(n10571), .B1(n14447), .B2(n10671), .C1(
        P2_U3088), .C2(n10904), .ZN(P2_U3321) );
  INV_X1 U13159 ( .A(n6622), .ZN(n13705) );
  OAI222_X1 U13160 ( .A1(n11421), .A2(P3_U3151), .B1(n13707), .B2(n10574), 
        .C1(n10573), .C2(n13705), .ZN(P3_U3289) );
  INV_X1 U13161 ( .A(n10575), .ZN(n10577) );
  INV_X1 U13162 ( .A(SI_8_), .ZN(n10576) );
  OAI222_X1 U13163 ( .A1(n11914), .A2(P3_U3151), .B1(n13707), .B2(n10577), 
        .C1(n10576), .C2(n13705), .ZN(P3_U3287) );
  OAI222_X1 U13164 ( .A1(n13140), .A2(P3_U3151), .B1(n13707), .B2(n10579), 
        .C1(n10578), .C2(n13705), .ZN(P3_U3285) );
  NAND2_X1 U13165 ( .A1(n12384), .A2(P1_B_REG_SCAN_IN), .ZN(n10581) );
  INV_X1 U13166 ( .A(n12139), .ZN(n10580) );
  MUX2_X1 U13167 ( .A(n10581), .B(P1_B_REG_SCAN_IN), .S(n10580), .Z(n10582) );
  INV_X1 U13168 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13169 ( .A1(n12740), .A2(n12384), .ZN(n10917) );
  INV_X1 U13170 ( .A(n10917), .ZN(n10584) );
  AOI22_X1 U13171 ( .A1(n15596), .A2(n10585), .B1(n10587), .B2(n10584), .ZN(
        P1_U3446) );
  INV_X1 U13172 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n15651) );
  NAND2_X1 U13173 ( .A1(n12740), .A2(n12139), .ZN(n10919) );
  INV_X1 U13174 ( .A(n10919), .ZN(n10586) );
  AOI22_X1 U13175 ( .A1(n15596), .A2(n15651), .B1(n10587), .B2(n10586), .ZN(
        P1_U3445) );
  OAI222_X1 U13176 ( .A1(P2_U3088), .A2(n15322), .B1(n14447), .B2(n10589), 
        .C1(n10588), .C2(n12742), .ZN(P2_U3326) );
  INV_X1 U13177 ( .A(n10590), .ZN(n10675) );
  INV_X1 U13178 ( .A(n13964), .ZN(n10591) );
  OAI222_X1 U13179 ( .A1(n12742), .A2(n10592), .B1(n14447), .B2(n10675), .C1(
        P2_U3088), .C2(n10591), .ZN(P2_U3322) );
  OAI222_X1 U13180 ( .A1(n12742), .A2(n10593), .B1(n14447), .B2(n10667), .C1(
        P2_U3088), .C2(n15341), .ZN(P2_U3325) );
  INV_X1 U13181 ( .A(n10594), .ZN(n10673) );
  INV_X1 U13182 ( .A(n11042), .ZN(n15368) );
  OAI222_X1 U13183 ( .A1(n12742), .A2(n10595), .B1(n14447), .B2(n10673), .C1(
        P2_U3088), .C2(n15368), .ZN(P2_U3320) );
  INV_X1 U13184 ( .A(n13707), .ZN(n11781) );
  AOI222_X1 U13185 ( .A1(n10597), .A2(n11781), .B1(n10596), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n6622), .ZN(n10598) );
  INV_X1 U13186 ( .A(n10598), .ZN(P3_U3291) );
  AOI222_X1 U13187 ( .A1(n10599), .A2(n11781), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11263), .C1(SI_5_), .C2(n6622), .ZN(n10600) );
  INV_X1 U13188 ( .A(n10600), .ZN(P3_U3290) );
  AOI222_X1 U13189 ( .A1(n10601), .A2(n11781), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n7497), .C1(SI_2_), .C2(n6622), .ZN(n10602) );
  INV_X1 U13190 ( .A(n10602), .ZN(P3_U3293) );
  AOI222_X1 U13191 ( .A1(n10603), .A2(n11781), .B1(SI_7_), .B2(n6622), .C1(
        n11427), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10604) );
  INV_X1 U13192 ( .A(n10604), .ZN(P3_U3288) );
  AOI222_X1 U13193 ( .A1(n10605), .A2(n11781), .B1(SI_3_), .B2(n6622), .C1(
        n11281), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10606) );
  INV_X1 U13194 ( .A(n10606), .ZN(P3_U3292) );
  OAI222_X1 U13195 ( .A1(P3_U3151), .A2(n13155), .B1(n13705), .B2(n10608), 
        .C1(n13707), .C2(n10607), .ZN(P3_U3284) );
  NAND2_X1 U13196 ( .A1(n13683), .A2(P3_D_REG_0__SCAN_IN), .ZN(n10609) );
  OAI21_X1 U13197 ( .B1(n13683), .B2(n10610), .A(n10609), .ZN(P3_U3376) );
  INV_X1 U13198 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10611) );
  NAND2_X1 U13199 ( .A1(n10611), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U13200 ( .A1(n10613), .A2(n10612), .ZN(n10631) );
  NAND2_X1 U13201 ( .A1(n10614), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10617) );
  INV_X1 U13202 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10615) );
  NAND2_X1 U13203 ( .A1(n10615), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U13204 ( .A1(n10626), .A2(n7368), .ZN(n10618) );
  NAND2_X1 U13205 ( .A1(n10618), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10619) );
  INV_X1 U13206 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10620) );
  INV_X1 U13207 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10623) );
  XNOR2_X1 U13208 ( .A(n10644), .B(n10623), .ZN(n15153) );
  NAND2_X1 U13209 ( .A1(n10624), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n10625) );
  NAND2_X1 U13210 ( .A1(n10626), .A2(n10625), .ZN(n15753) );
  OAI21_X1 U13211 ( .B1(n10629), .B2(n10628), .A(n10627), .ZN(n10637) );
  NAND2_X1 U13212 ( .A1(n10631), .A2(n10630), .ZN(n10632) );
  NAND2_X1 U13213 ( .A1(n10633), .A2(n10632), .ZN(n10634) );
  NAND2_X1 U13214 ( .A1(n10634), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10636) );
  XOR2_X1 U13215 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10634), .Z(n15755) );
  NAND2_X1 U13216 ( .A1(n15756), .A2(n15755), .ZN(n10635) );
  NAND2_X1 U13217 ( .A1(n10636), .A2(n10635), .ZN(n10638) );
  NAND2_X1 U13218 ( .A1(n10637), .A2(n10638), .ZN(n15230) );
  INV_X1 U13219 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15232) );
  NAND2_X1 U13220 ( .A1(n15230), .A2(n15232), .ZN(n10641) );
  INV_X1 U13221 ( .A(n10637), .ZN(n10640) );
  INV_X1 U13222 ( .A(n10638), .ZN(n10639) );
  NAND2_X1 U13223 ( .A1(n10640), .A2(n10639), .ZN(n15231) );
  AND2_X1 U13224 ( .A1(n10641), .A2(n15231), .ZN(n15752) );
  OAI21_X1 U13225 ( .B1(n15753), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n15752), .ZN(
        n10643) );
  NAND2_X1 U13226 ( .A1(n15753), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U13227 ( .A1(n10643), .A2(n10642), .ZN(n15154) );
  AND2_X1 U13228 ( .A1(n10644), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10645) );
  INV_X1 U13229 ( .A(n10647), .ZN(n10648) );
  NAND2_X1 U13230 ( .A1(n10651), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n10652) );
  NAND2_X1 U13231 ( .A1(n11128), .A2(n10652), .ZN(SUB_1596_U58) );
  INV_X1 U13232 ( .A(n10653), .ZN(n10656) );
  INV_X1 U13233 ( .A(n11001), .ZN(n10849) );
  OAI222_X1 U13234 ( .A1(n15149), .A2(n10654), .B1(n15141), .B2(n10656), .C1(
        P1_U3086), .C2(n10849), .ZN(P1_U3347) );
  INV_X1 U13235 ( .A(n13975), .ZN(n10655) );
  OAI222_X1 U13236 ( .A1(n12742), .A2(n10657), .B1(n14447), .B2(n10656), .C1(
        P2_U3088), .C2(n10655), .ZN(P2_U3319) );
  INV_X1 U13237 ( .A(n11740), .ZN(n10658) );
  NAND2_X1 U13238 ( .A1(n10658), .A2(n11210), .ZN(n10697) );
  OR2_X1 U13239 ( .A1(n10970), .A2(n10659), .ZN(n10661) );
  AND2_X1 U13240 ( .A1(n10661), .A2(n10660), .ZN(n10696) );
  INV_X1 U13241 ( .A(n10696), .ZN(n10662) );
  NOR2_X1 U13242 ( .A1(n15255), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U13243 ( .A1(n11922), .A2(P3_U3151), .B1(n13707), .B2(n10664), 
        .C1(n10663), .C2(n13705), .ZN(P3_U3286) );
  OAI222_X1 U13244 ( .A1(n7124), .A2(P3_U3151), .B1(n13707), .B2(n10666), .C1(
        n10665), .C2(n13705), .ZN(P3_U3294) );
  OAI222_X1 U13245 ( .A1(n15149), .A2(n10668), .B1(n15141), .B2(n10667), .C1(
        P1_U3086), .C2(n10766), .ZN(P1_U3353) );
  OAI222_X1 U13246 ( .A1(n15149), .A2(n10670), .B1(n15141), .B2(n10669), .C1(
        P1_U3086), .C2(n10774), .ZN(P1_U3351) );
  INV_X1 U13247 ( .A(n10738), .ZN(n10715) );
  OAI222_X1 U13248 ( .A1(n15149), .A2(n10672), .B1(n15141), .B2(n10671), .C1(
        P1_U3086), .C2(n10715), .ZN(P1_U3349) );
  INV_X1 U13249 ( .A(n10838), .ZN(n10841) );
  OAI222_X1 U13250 ( .A1(n15149), .A2(n10674), .B1(n15141), .B2(n10673), .C1(
        P1_U3086), .C2(n10841), .ZN(P1_U3348) );
  INV_X1 U13251 ( .A(n10707), .ZN(n10722) );
  OAI222_X1 U13252 ( .A1(n15149), .A2(n10676), .B1(n15141), .B2(n10675), .C1(
        P1_U3086), .C2(n10722), .ZN(P1_U3350) );
  INV_X1 U13253 ( .A(n10677), .ZN(n10680) );
  INV_X1 U13254 ( .A(n15383), .ZN(n10678) );
  OAI222_X1 U13255 ( .A1(n12742), .A2(n10679), .B1(n14447), .B2(n10680), .C1(
        P2_U3088), .C2(n10678), .ZN(P2_U3318) );
  OAI222_X1 U13256 ( .A1(n15149), .A2(n10681), .B1(n15141), .B2(n10680), .C1(
        P1_U3086), .C2(n11070), .ZN(P1_U3346) );
  INV_X1 U13257 ( .A(n10682), .ZN(n10683) );
  OAI222_X1 U13258 ( .A1(P3_U3151), .A2(n13180), .B1(n13705), .B2(n10684), 
        .C1(n13707), .C2(n10683), .ZN(P3_U3283) );
  NAND2_X1 U13259 ( .A1(n13130), .A2(P3_DATAO_REG_11__SCAN_IN), .ZN(n10685) );
  OAI21_X1 U13260 ( .B1(n13130), .B2(n13073), .A(n10685), .ZN(P3_U3502) );
  INV_X1 U13261 ( .A(n10686), .ZN(n10689) );
  INV_X1 U13262 ( .A(n15395), .ZN(n10687) );
  OAI222_X1 U13263 ( .A1(n12742), .A2(n10688), .B1(n14447), .B2(n10689), .C1(
        P2_U3088), .C2(n10687), .ZN(P2_U3317) );
  INV_X1 U13264 ( .A(n11393), .ZN(n11388) );
  OAI222_X1 U13265 ( .A1(n15149), .A2(n10690), .B1(n15141), .B2(n10689), .C1(
        P1_U3086), .C2(n11388), .ZN(P1_U3345) );
  INV_X1 U13266 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10691) );
  MUX2_X1 U13267 ( .A(n10691), .B(P1_REG1_REG_6__SCAN_IN), .S(n10738), .Z(
        n10699) );
  MUX2_X1 U13268 ( .A(n9578), .B(P1_REG1_REG_1__SCAN_IN), .S(n10700), .Z(
        n14629) );
  AND2_X1 U13269 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n14628) );
  NAND2_X1 U13270 ( .A1(n14629), .A2(n14628), .ZN(n14627) );
  INV_X1 U13271 ( .A(n10700), .ZN(n14634) );
  NAND2_X1 U13272 ( .A1(n14634), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10692) );
  NAND2_X1 U13273 ( .A1(n14627), .A2(n10692), .ZN(n10764) );
  MUX2_X1 U13274 ( .A(n10693), .B(P1_REG1_REG_2__SCAN_IN), .S(n10766), .Z(
        n10765) );
  NAND2_X1 U13275 ( .A1(n10764), .A2(n10765), .ZN(n10763) );
  OAI21_X1 U13276 ( .B1(n10766), .B2(n10693), .A(n10763), .ZN(n14643) );
  MUX2_X1 U13277 ( .A(n10694), .B(P1_REG1_REG_3__SCAN_IN), .S(n14639), .Z(
        n14644) );
  MUX2_X1 U13278 ( .A(n9626), .B(P1_REG1_REG_4__SCAN_IN), .S(n10774), .Z(
        n10778) );
  XNOR2_X1 U13279 ( .A(n10707), .B(n10695), .ZN(n10720) );
  NAND2_X1 U13280 ( .A1(n6465), .A2(n10720), .ZN(n10719) );
  OAI21_X1 U13281 ( .B1(n10707), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10719), .ZN(
        n10698) );
  NAND2_X1 U13282 ( .A1(n10697), .A2(n10696), .ZN(n15258) );
  NOR2_X1 U13283 ( .A1(n10698), .A2(n10699), .ZN(n10734) );
  AOI211_X1 U13284 ( .C1(n10699), .C2(n10698), .A(n14687), .B(n10734), .ZN(
        n10718) );
  MUX2_X1 U13285 ( .A(n10701), .B(P1_REG2_REG_1__SCAN_IN), .S(n10700), .Z(
        n14632) );
  AND2_X1 U13286 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10702) );
  NAND2_X1 U13287 ( .A1(n14632), .A2(n10702), .ZN(n14631) );
  NAND2_X1 U13288 ( .A1(n14634), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10703) );
  NAND2_X1 U13289 ( .A1(n14631), .A2(n10703), .ZN(n10761) );
  MUX2_X1 U13290 ( .A(n11745), .B(P1_REG2_REG_2__SCAN_IN), .S(n10766), .Z(
        n10762) );
  NAND2_X1 U13291 ( .A1(n10761), .A2(n10762), .ZN(n10760) );
  INV_X1 U13292 ( .A(n10760), .ZN(n14647) );
  NOR2_X1 U13293 ( .A1(n10766), .A2(n11745), .ZN(n14646) );
  MUX2_X1 U13294 ( .A(n10704), .B(P1_REG2_REG_3__SCAN_IN), .S(n14639), .Z(
        n14645) );
  MUX2_X1 U13295 ( .A(n10705), .B(P1_REG2_REG_4__SCAN_IN), .S(n10774), .Z(
        n10775) );
  MUX2_X1 U13296 ( .A(n12041), .B(P1_REG2_REG_5__SCAN_IN), .S(n10707), .Z(
        n10724) );
  NOR2_X1 U13297 ( .A1(n10722), .A2(n12041), .ZN(n10710) );
  MUX2_X1 U13298 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n12011), .S(n10738), .Z(
        n10709) );
  OAI21_X1 U13299 ( .B1(n10723), .B2(n10710), .A(n10709), .ZN(n10741) );
  INV_X1 U13300 ( .A(n10741), .ZN(n10712) );
  OR2_X1 U13301 ( .A1(n10115), .A2(n15146), .ZN(n10708) );
  NOR3_X1 U13302 ( .A1(n10723), .A2(n10710), .A3(n10709), .ZN(n10711) );
  NOR3_X1 U13303 ( .A1(n10712), .A2(n14677), .A3(n10711), .ZN(n10717) );
  INV_X1 U13304 ( .A(n15146), .ZN(n10928) );
  NAND2_X1 U13305 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11204) );
  INV_X1 U13306 ( .A(n11204), .ZN(n10713) );
  AOI21_X1 U13307 ( .B1(n15255), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10713), .ZN(
        n10714) );
  OAI21_X1 U13308 ( .B1(n14686), .B2(n10715), .A(n10714), .ZN(n10716) );
  OR3_X1 U13309 ( .A1(n10718), .A2(n10717), .A3(n10716), .ZN(P1_U3249) );
  OAI21_X1 U13310 ( .B1(n10720), .B2(n6465), .A(n10719), .ZN(n10728) );
  NAND2_X1 U13311 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11365) );
  NAND2_X1 U13312 ( .A1(n15255), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n10721) );
  OAI211_X1 U13313 ( .C1(n14686), .C2(n10722), .A(n11365), .B(n10721), .ZN(
        n10727) );
  AOI211_X1 U13314 ( .C1(n10725), .C2(n10724), .A(n10723), .B(n14677), .ZN(
        n10726) );
  AOI211_X1 U13315 ( .C1(n15266), .C2(n10728), .A(n10727), .B(n10726), .ZN(
        n10729) );
  INV_X1 U13316 ( .A(n10729), .ZN(P1_U3248) );
  INV_X1 U13317 ( .A(n10730), .ZN(n10732) );
  INV_X1 U13318 ( .A(n11680), .ZN(n11678) );
  OAI222_X1 U13319 ( .A1(n15149), .A2(n10731), .B1(n15141), .B2(n10732), .C1(
        P1_U3086), .C2(n11678), .ZN(P1_U3344) );
  INV_X1 U13320 ( .A(n11050), .ZN(n15406) );
  OAI222_X1 U13321 ( .A1(n12742), .A2(n10733), .B1(n14447), .B2(n10732), .C1(
        P2_U3088), .C2(n15406), .ZN(P2_U3316) );
  INV_X1 U13322 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10735) );
  MUX2_X1 U13323 ( .A(n10735), .B(P1_REG1_REG_7__SCAN_IN), .S(n10838), .Z(
        n10736) );
  AOI211_X1 U13324 ( .C1(n10737), .C2(n10736), .A(n14687), .B(n10837), .ZN(
        n10748) );
  NAND2_X1 U13325 ( .A1(n10738), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10740) );
  MUX2_X1 U13326 ( .A(n9669), .B(P1_REG2_REG_7__SCAN_IN), .S(n10838), .Z(
        n10739) );
  AOI21_X1 U13327 ( .B1(n10741), .B2(n10740), .A(n10739), .ZN(n10844) );
  INV_X1 U13328 ( .A(n10844), .ZN(n10743) );
  NAND3_X1 U13329 ( .A1(n10741), .A2(n10740), .A3(n10739), .ZN(n10742) );
  NAND3_X1 U13330 ( .A1(n10743), .A2(n15267), .A3(n10742), .ZN(n10746) );
  NOR2_X1 U13331 ( .A1(n10744), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11537) );
  AOI21_X1 U13332 ( .B1(n15255), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n11537), .ZN(
        n10745) );
  OAI211_X1 U13333 ( .C1(n14686), .C2(n10841), .A(n10746), .B(n10745), .ZN(
        n10747) );
  OR2_X1 U13334 ( .A1(n10748), .A2(n10747), .ZN(P1_U3250) );
  NAND2_X4 U13335 ( .A1(n11168), .A2(n14906), .ZN(n12855) );
  INV_X1 U13336 ( .A(n11207), .ZN(n10752) );
  NAND2_X1 U13337 ( .A1(n11176), .A2(n14626), .ZN(n10754) );
  NAND2_X1 U13338 ( .A1(n10752), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10753) );
  OAI211_X1 U13339 ( .C1(n12755), .C2(n11909), .A(n10754), .B(n10753), .ZN(
        n11153) );
  NAND2_X1 U13340 ( .A1(n10755), .A2(n11153), .ZN(n11156) );
  OAI21_X1 U13341 ( .B1(n10755), .B2(n11153), .A(n11156), .ZN(n10973) );
  NAND2_X1 U13342 ( .A1(n10973), .A2(n10115), .ZN(n10759) );
  NAND2_X1 U13343 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14630) );
  AOI21_X1 U13344 ( .B1(n10756), .B2(n14630), .A(n15146), .ZN(n10758) );
  OR2_X1 U13345 ( .A1(n10115), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10757) );
  AND2_X1 U13346 ( .A1(n10757), .A2(n10928), .ZN(n15248) );
  NOR2_X1 U13347 ( .A1(n15248), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n15252) );
  AOI211_X1 U13348 ( .C1(n10759), .C2(n10758), .A(n15252), .B(n14611), .ZN(
        n10783) );
  OAI211_X1 U13349 ( .C1(n10762), .C2(n10761), .A(n15267), .B(n10760), .ZN(
        n10771) );
  OAI211_X1 U13350 ( .C1(n10765), .C2(n10764), .A(n15266), .B(n10763), .ZN(
        n10770) );
  AOI22_X1 U13351 ( .A1(n15255), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10769) );
  INV_X1 U13352 ( .A(n14686), .ZN(n15263) );
  INV_X1 U13353 ( .A(n10766), .ZN(n10767) );
  NAND2_X1 U13354 ( .A1(n15263), .A2(n10767), .ZN(n10768) );
  NAND4_X1 U13355 ( .A1(n10771), .A2(n10770), .A3(n10769), .A4(n10768), .ZN(
        n10772) );
  OR2_X1 U13356 ( .A1(n10783), .A2(n10772), .ZN(P1_U3245) );
  NAND2_X1 U13357 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n11382) );
  NAND2_X1 U13358 ( .A1(n15255), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10773) );
  OAI211_X1 U13359 ( .C1(n14686), .C2(n10774), .A(n11382), .B(n10773), .ZN(
        n10782) );
  XNOR2_X1 U13360 ( .A(n10776), .B(n10775), .ZN(n10780) );
  OAI211_X1 U13361 ( .C1(n10778), .C2(n10777), .A(n15266), .B(n7288), .ZN(
        n10779) );
  OAI21_X1 U13362 ( .B1(n14677), .B2(n10780), .A(n10779), .ZN(n10781) );
  OR3_X1 U13363 ( .A1(n10783), .A2(n10782), .A3(n10781), .ZN(P1_U3247) );
  INV_X1 U13364 ( .A(n10784), .ZN(n10785) );
  OAI222_X1 U13365 ( .A1(P3_U3151), .A2(n7411), .B1(n13705), .B2(n10786), .C1(
        n13707), .C2(n10785), .ZN(P3_U3280) );
  INV_X1 U13366 ( .A(n10787), .ZN(n10790) );
  INV_X1 U13367 ( .A(n12388), .ZN(n12391) );
  OAI222_X1 U13368 ( .A1(n15149), .A2(n10788), .B1(n15141), .B2(n10790), .C1(
        n12391), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U13369 ( .A(n15424), .ZN(n10789) );
  OAI222_X1 U13370 ( .A1(n12742), .A2(n10791), .B1(n14447), .B2(n10790), .C1(
        n10789), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U13371 ( .A(n10792), .ZN(n10794) );
  OAI222_X1 U13372 ( .A1(n12742), .A2(n10793), .B1(n14447), .B2(n10794), .C1(
        n12238), .C2(P2_U3088), .ZN(P2_U3315) );
  OAI222_X1 U13373 ( .A1(n15149), .A2(n10795), .B1(n15141), .B2(n10794), .C1(
        n11684), .C2(P1_U3086), .ZN(P1_U3343) );
  OAI222_X1 U13374 ( .A1(P3_U3151), .A2(n13221), .B1(n13705), .B2(n10797), 
        .C1(n13707), .C2(n10796), .ZN(P3_U3281) );
  INV_X1 U13375 ( .A(n13213), .ZN(n13183) );
  INV_X1 U13376 ( .A(n10798), .ZN(n10799) );
  OAI222_X1 U13377 ( .A1(P3_U3151), .A2(n13183), .B1(n13705), .B2(n10800), 
        .C1(n13707), .C2(n10799), .ZN(P3_U3282) );
  NOR2_X1 U13378 ( .A1(n13683), .A2(n10801), .ZN(n10803) );
  CLKBUF_X1 U13379 ( .A(n10803), .Z(n10827) );
  INV_X1 U13380 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10802) );
  NOR2_X1 U13381 ( .A1(n10827), .A2(n10802), .ZN(P3_U3249) );
  INV_X1 U13382 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10804) );
  NOR2_X1 U13383 ( .A1(n10827), .A2(n10804), .ZN(P3_U3237) );
  INV_X1 U13384 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10805) );
  NOR2_X1 U13385 ( .A1(n10827), .A2(n10805), .ZN(P3_U3247) );
  INV_X1 U13386 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10806) );
  NOR2_X1 U13387 ( .A1(n10827), .A2(n10806), .ZN(P3_U3256) );
  INV_X1 U13388 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10807) );
  NOR2_X1 U13389 ( .A1(n10827), .A2(n10807), .ZN(P3_U3248) );
  INV_X1 U13390 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n15652) );
  NOR2_X1 U13391 ( .A1(n10803), .A2(n15652), .ZN(P3_U3242) );
  INV_X1 U13392 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10808) );
  NOR2_X1 U13393 ( .A1(n10803), .A2(n10808), .ZN(P3_U3243) );
  INV_X1 U13394 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10809) );
  NOR2_X1 U13395 ( .A1(n10803), .A2(n10809), .ZN(P3_U3238) );
  INV_X1 U13396 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10810) );
  NOR2_X1 U13397 ( .A1(n10827), .A2(n10810), .ZN(P3_U3253) );
  INV_X1 U13398 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10811) );
  NOR2_X1 U13399 ( .A1(n10803), .A2(n10811), .ZN(P3_U3262) );
  INV_X1 U13400 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10812) );
  NOR2_X1 U13401 ( .A1(n10803), .A2(n10812), .ZN(P3_U3244) );
  INV_X1 U13402 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10813) );
  NOR2_X1 U13403 ( .A1(n10803), .A2(n10813), .ZN(P3_U3245) );
  INV_X1 U13404 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10814) );
  NOR2_X1 U13405 ( .A1(n10827), .A2(n10814), .ZN(P3_U3246) );
  INV_X1 U13406 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10815) );
  NOR2_X1 U13407 ( .A1(n10827), .A2(n10815), .ZN(P3_U3255) );
  INV_X1 U13408 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10816) );
  NOR2_X1 U13409 ( .A1(n10803), .A2(n10816), .ZN(P3_U3240) );
  INV_X1 U13410 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10817) );
  NOR2_X1 U13411 ( .A1(n10803), .A2(n10817), .ZN(P3_U3239) );
  INV_X1 U13412 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10818) );
  NOR2_X1 U13413 ( .A1(n10827), .A2(n10818), .ZN(P3_U3261) );
  INV_X1 U13414 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10819) );
  NOR2_X1 U13415 ( .A1(n10827), .A2(n10819), .ZN(P3_U3251) );
  INV_X1 U13416 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10820) );
  NOR2_X1 U13417 ( .A1(n10827), .A2(n10820), .ZN(P3_U3252) );
  INV_X1 U13418 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10821) );
  NOR2_X1 U13419 ( .A1(n10803), .A2(n10821), .ZN(P3_U3236) );
  INV_X1 U13420 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10822) );
  NOR2_X1 U13421 ( .A1(n10803), .A2(n10822), .ZN(P3_U3235) );
  INV_X1 U13422 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10823) );
  NOR2_X1 U13423 ( .A1(n10827), .A2(n10823), .ZN(P3_U3263) );
  INV_X1 U13424 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10824) );
  NOR2_X1 U13425 ( .A1(n10827), .A2(n10824), .ZN(P3_U3259) );
  INV_X1 U13426 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10825) );
  NOR2_X1 U13427 ( .A1(n10827), .A2(n10825), .ZN(P3_U3257) );
  INV_X1 U13428 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10826) );
  NOR2_X1 U13429 ( .A1(n10827), .A2(n10826), .ZN(P3_U3250) );
  INV_X1 U13430 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n15669) );
  NOR2_X1 U13431 ( .A1(n10827), .A2(n15669), .ZN(P3_U3254) );
  INV_X1 U13432 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10828) );
  NOR2_X1 U13433 ( .A1(n10803), .A2(n10828), .ZN(P3_U3260) );
  INV_X1 U13434 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10829) );
  NOR2_X1 U13435 ( .A1(n10827), .A2(n10829), .ZN(P3_U3234) );
  INV_X1 U13436 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10830) );
  NOR2_X1 U13437 ( .A1(n10827), .A2(n10830), .ZN(P3_U3241) );
  INV_X1 U13438 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10831) );
  NOR2_X1 U13439 ( .A1(n10827), .A2(n10831), .ZN(P3_U3258) );
  INV_X1 U13440 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n15721) );
  NAND2_X1 U13441 ( .A1(P3_U3897), .A2(n12205), .ZN(n10832) );
  OAI21_X1 U13442 ( .B1(P3_U3897), .B2(n15721), .A(n10832), .ZN(P3_U3499) );
  INV_X1 U13443 ( .A(n13259), .ZN(n13274) );
  INV_X1 U13444 ( .A(n10833), .ZN(n10834) );
  OAI222_X1 U13445 ( .A1(P3_U3151), .A2(n13274), .B1(n13705), .B2(n10835), 
        .C1(n13707), .C2(n10834), .ZN(P3_U3279) );
  XNOR2_X1 U13446 ( .A(n11001), .B(n10836), .ZN(n10840) );
  OAI21_X1 U13447 ( .B1(n10840), .B2(n10839), .A(n10999), .ZN(n10852) );
  NOR2_X1 U13448 ( .A1(n10841), .A2(n9669), .ZN(n10843) );
  MUX2_X1 U13449 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n12097), .S(n11001), .Z(
        n10842) );
  OAI21_X1 U13450 ( .B1(n10844), .B2(n10843), .A(n10842), .ZN(n11005) );
  INV_X1 U13451 ( .A(n11005), .ZN(n10846) );
  NOR3_X1 U13452 ( .A1(n10844), .A2(n10843), .A3(n10842), .ZN(n10845) );
  NOR3_X1 U13453 ( .A1(n10846), .A2(n10845), .A3(n14677), .ZN(n10851) );
  AND2_X1 U13454 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10847) );
  AOI21_X1 U13455 ( .B1(n15255), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n10847), .ZN(
        n10848) );
  OAI21_X1 U13456 ( .B1(n14686), .B2(n10849), .A(n10848), .ZN(n10850) );
  AOI211_X1 U13457 ( .C1(n10852), .C2(n15266), .A(n10851), .B(n10850), .ZN(
        n10853) );
  INV_X1 U13458 ( .A(n10853), .ZN(P1_U3251) );
  AOI21_X1 U13459 ( .B1(n10856), .B2(n10855), .A(n10854), .ZN(n10857) );
  OR2_X1 U13460 ( .A1(n10858), .A2(n10857), .ZN(n10860) );
  NAND2_X1 U13461 ( .A1(n10860), .A2(n10859), .ZN(n15323) );
  NOR2_X2 U13462 ( .A1(n15323), .A2(P2_U3088), .ZN(n15450) );
  INV_X1 U13463 ( .A(n15450), .ZN(n15405) );
  NAND2_X1 U13464 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n11548) );
  INV_X1 U13465 ( .A(n11548), .ZN(n10872) );
  NOR2_X1 U13466 ( .A1(n10859), .A2(P2_U3088), .ZN(n14444) );
  NAND2_X1 U13467 ( .A1(n10860), .A2(n14444), .ZN(n10879) );
  INV_X1 U13468 ( .A(n10879), .ZN(n10861) );
  AND2_X1 U13469 ( .A1(n15321), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n15332) );
  NAND2_X1 U13470 ( .A1(n15331), .A2(n15332), .ZN(n15330) );
  NAND2_X1 U13471 ( .A1(n10873), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U13472 ( .A1(n15330), .A2(n10862), .ZN(n15344) );
  MUX2_X1 U13473 ( .A(n10863), .B(P2_REG2_REG_2__SCAN_IN), .S(n15341), .Z(
        n15345) );
  NAND2_X1 U13474 ( .A1(n15344), .A2(n15345), .ZN(n15343) );
  NAND2_X1 U13475 ( .A1(n10875), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10864) );
  NAND2_X1 U13476 ( .A1(n15343), .A2(n10864), .ZN(n15358) );
  MUX2_X1 U13477 ( .A(n10865), .B(P2_REG2_REG_3__SCAN_IN), .S(n10877), .Z(
        n15359) );
  OR2_X1 U13478 ( .A1(n10877), .A2(n10865), .ZN(n10869) );
  NAND2_X1 U13479 ( .A1(n15357), .A2(n10869), .ZN(n10867) );
  INV_X1 U13480 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11650) );
  MUX2_X1 U13481 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11650), .S(n10896), .Z(
        n10866) );
  MUX2_X1 U13482 ( .A(n11650), .B(P2_REG2_REG_4__SCAN_IN), .S(n10896), .Z(
        n10868) );
  NAND3_X1 U13483 ( .A1(n15357), .A2(n10869), .A3(n10868), .ZN(n10870) );
  AND3_X1 U13484 ( .A1(n15451), .A2(n13957), .A3(n10870), .ZN(n10871) );
  AOI211_X1 U13485 ( .C1(n15336), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n10872), .B(
        n10871), .ZN(n10883) );
  MUX2_X1 U13486 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n8708), .S(n10896), .Z(
        n10881) );
  INV_X1 U13487 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n12745) );
  AND2_X1 U13488 ( .A1(n15321), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n15326) );
  NAND2_X1 U13489 ( .A1(n10873), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10874) );
  INV_X1 U13490 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n15497) );
  NAND2_X1 U13491 ( .A1(n15338), .A2(n15339), .ZN(n15337) );
  NAND2_X1 U13492 ( .A1(n10875), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10876) );
  INV_X1 U13493 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n15637) );
  MUX2_X1 U13494 ( .A(n15637), .B(P2_REG1_REG_3__SCAN_IN), .S(n10877), .Z(
        n15351) );
  INV_X1 U13495 ( .A(n10877), .ZN(n15352) );
  NAND2_X1 U13496 ( .A1(n15352), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10878) );
  NAND2_X1 U13497 ( .A1(n15349), .A2(n10878), .ZN(n10880) );
  NOR2_X2 U13498 ( .A1(n10879), .A2(n12916), .ZN(n15402) );
  NAND2_X1 U13499 ( .A1(n10880), .A2(n10881), .ZN(n10898) );
  OAI211_X1 U13500 ( .C1(n10881), .C2(n10880), .A(n15402), .B(n10898), .ZN(
        n10882) );
  OAI211_X1 U13501 ( .C1(n15405), .C2(n10884), .A(n10883), .B(n10882), .ZN(
        P2_U3218) );
  NAND2_X1 U13502 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n11519) );
  INV_X1 U13503 ( .A(n11519), .ZN(n10895) );
  NAND2_X1 U13504 ( .A1(n10896), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n13956) );
  NAND2_X1 U13505 ( .A1(n13957), .A2(n13956), .ZN(n10887) );
  MUX2_X1 U13506 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10885), .S(n13964), .Z(
        n10886) );
  NAND2_X1 U13507 ( .A1(n13964), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10892) );
  NAND2_X1 U13508 ( .A1(n13959), .A2(n10892), .ZN(n10890) );
  MUX2_X1 U13509 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10888), .S(n11039), .Z(
        n10889) );
  NAND2_X1 U13510 ( .A1(n10890), .A2(n10889), .ZN(n11041) );
  MUX2_X1 U13511 ( .A(n10888), .B(P2_REG2_REG_6__SCAN_IN), .S(n11039), .Z(
        n10891) );
  NAND3_X1 U13512 ( .A1(n13959), .A2(n10892), .A3(n10891), .ZN(n10893) );
  AND3_X1 U13513 ( .A1(n15451), .A2(n11041), .A3(n10893), .ZN(n10894) );
  AOI211_X1 U13514 ( .C1(n15336), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n10895), .B(
        n10894), .ZN(n10903) );
  MUX2_X1 U13515 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n8760), .S(n11039), .Z(
        n10901) );
  NAND2_X1 U13516 ( .A1(n10896), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10897) );
  NAND2_X1 U13517 ( .A1(n10898), .A2(n10897), .ZN(n13962) );
  MUX2_X1 U13518 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n8735), .S(n13964), .Z(
        n13963) );
  NAND2_X1 U13519 ( .A1(n13962), .A2(n13963), .ZN(n13961) );
  NAND2_X1 U13520 ( .A1(n13964), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U13521 ( .A1(n10900), .A2(n10901), .ZN(n11029) );
  OAI211_X1 U13522 ( .C1(n10901), .C2(n10900), .A(n15402), .B(n11029), .ZN(
        n10902) );
  OAI211_X1 U13523 ( .C1(n15405), .C2(n10904), .A(n10903), .B(n10902), .ZN(
        P2_U3220) );
  NOR2_X1 U13524 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n15605) );
  NOR4_X1 U13525 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10907) );
  NOR4_X1 U13526 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n10906) );
  NOR4_X1 U13527 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n10905) );
  AND4_X1 U13528 ( .A1(n15605), .A2(n10907), .A3(n10906), .A4(n10905), .ZN(
        n10913) );
  NOR4_X1 U13529 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n10911) );
  NOR4_X1 U13530 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n10910) );
  NOR4_X1 U13531 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n10909) );
  NOR4_X1 U13532 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n10908) );
  AND4_X1 U13533 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .ZN(
        n10912) );
  NAND2_X1 U13534 ( .A1(n10913), .A2(n10912), .ZN(n10964) );
  INV_X1 U13535 ( .A(n10964), .ZN(n10914) );
  NAND2_X1 U13536 ( .A1(n11740), .A2(n10914), .ZN(n10916) );
  INV_X1 U13537 ( .A(n11206), .ZN(n10915) );
  OR2_X1 U13538 ( .A1(n14893), .A2(n14716), .ZN(n10967) );
  INV_X1 U13539 ( .A(n11748), .ZN(n11739) );
  NAND2_X1 U13540 ( .A1(n15151), .A2(n14716), .ZN(n10921) );
  NOR2_X1 U13541 ( .A1(n10921), .A2(n10920), .ZN(n10922) );
  NOR2_X1 U13542 ( .A1(n10923), .A2(n14716), .ZN(n10924) );
  OR2_X1 U13543 ( .A1(n10006), .A2(n14716), .ZN(n10926) );
  INV_X1 U13544 ( .A(n10927), .ZN(n11906) );
  OAI21_X1 U13545 ( .B1(n15297), .B2(n15308), .A(n11906), .ZN(n10931) );
  NOR2_X1 U13546 ( .A1(n11152), .A2(n14916), .ZN(n11900) );
  INV_X1 U13547 ( .A(n11746), .ZN(n10954) );
  AND2_X1 U13548 ( .A1(n10954), .A2(n10935), .ZN(n10929) );
  NOR2_X1 U13549 ( .A1(n11900), .A2(n10929), .ZN(n10930) );
  AND2_X1 U13550 ( .A1(n10931), .A2(n10930), .ZN(n15275) );
  NAND2_X1 U13551 ( .A1(n15314), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10932) );
  OAI21_X1 U13552 ( .B1(n15314), .B2(n15275), .A(n10932), .ZN(P1_U3528) );
  INV_X1 U13553 ( .A(n13295), .ZN(n13299) );
  INV_X1 U13554 ( .A(n10933), .ZN(n10934) );
  OAI222_X1 U13555 ( .A1(P3_U3151), .A2(n13299), .B1(n13705), .B2(n15626), 
        .C1(n13707), .C2(n10934), .ZN(P3_U3278) );
  NAND2_X1 U13556 ( .A1(n14626), .A2(n10935), .ZN(n11014) );
  NAND2_X1 U13557 ( .A1(n11014), .A2(n11152), .ZN(n10936) );
  NAND2_X1 U13558 ( .A1(n10937), .A2(n10936), .ZN(n10940) );
  INV_X1 U13559 ( .A(n10940), .ZN(n10938) );
  NAND2_X1 U13560 ( .A1(n10938), .A2(n10946), .ZN(n10941) );
  INV_X1 U13561 ( .A(n10946), .ZN(n10939) );
  INV_X1 U13562 ( .A(n15282), .ZN(n15061) );
  NAND2_X1 U13563 ( .A1(n10943), .A2(n10942), .ZN(n10945) );
  AND2_X2 U13564 ( .A1(n10945), .A2(n10944), .ZN(n10947) );
  OAI21_X1 U13565 ( .B1(n10947), .B2(n10946), .A(n11595), .ZN(n10951) );
  OAI22_X1 U13566 ( .A1(n11596), .A2(n14916), .B1(n11152), .B2(n14918), .ZN(
        n10950) );
  INV_X1 U13567 ( .A(n14873), .ZN(n10948) );
  NOR2_X1 U13568 ( .A1(n11757), .A2(n10948), .ZN(n10949) );
  AOI211_X1 U13569 ( .C1(n15308), .C2(n10951), .A(n10950), .B(n10949), .ZN(
        n11744) );
  INV_X1 U13570 ( .A(n10952), .ZN(n10953) );
  INV_X1 U13571 ( .A(n11016), .ZN(n10955) );
  OAI211_X1 U13572 ( .C1(n10955), .C2(n11225), .A(n14949), .B(n11949), .ZN(
        n11752) );
  INV_X1 U13573 ( .A(n11752), .ZN(n10956) );
  AOI21_X1 U13574 ( .B1(n15302), .B2(n11754), .A(n10956), .ZN(n10957) );
  OAI211_X1 U13575 ( .C1(n11757), .C2(n15061), .A(n11744), .B(n10957), .ZN(
        n10960) );
  NAND2_X1 U13576 ( .A1(n10960), .A2(n15316), .ZN(n10958) );
  OAI21_X1 U13577 ( .B1(n15316), .B2(n10693), .A(n10958), .ZN(P1_U3530) );
  INV_X1 U13578 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U13579 ( .A1(n10960), .A2(n15310), .ZN(n10961) );
  OAI21_X1 U13580 ( .B1(n15310), .B2(n10962), .A(n10961), .ZN(P1_U3465) );
  NOR2_X1 U13581 ( .A1(n11748), .A2(n11736), .ZN(n10968) );
  INV_X1 U13582 ( .A(n10963), .ZN(n10965) );
  NAND2_X1 U13583 ( .A1(n10965), .A2(n10964), .ZN(n10966) );
  NAND2_X1 U13584 ( .A1(n10968), .A2(n10966), .ZN(n10969) );
  NAND2_X1 U13585 ( .A1(n10969), .A2(n10967), .ZN(n11208) );
  NAND2_X1 U13586 ( .A1(n10968), .A2(n11738), .ZN(n14595) );
  INV_X1 U13587 ( .A(n14556), .ZN(n14576) );
  INV_X1 U13588 ( .A(n11152), .ZN(n14625) );
  INV_X1 U13589 ( .A(n10969), .ZN(n10972) );
  AND3_X1 U13590 ( .A1(n11740), .A2(n10970), .A3(n15065), .ZN(n10971) );
  AOI22_X1 U13591 ( .A1(n14576), .A2(n14625), .B1(n14589), .B2(n10973), .ZN(
        n10975) );
  NAND2_X1 U13592 ( .A1(n15236), .A2(n11206), .ZN(n11228) );
  NAND2_X1 U13593 ( .A1(n11228), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10974) );
  OAI211_X1 U13594 ( .C1(n14600), .C2(n11909), .A(n10975), .B(n10974), .ZN(
        P1_U3232) );
  INV_X1 U13595 ( .A(n15462), .ZN(n10977) );
  INV_X1 U13596 ( .A(n15484), .ZN(n15476) );
  OAI21_X1 U13597 ( .B1(n10353), .B2(n10983), .A(n10982), .ZN(n14274) );
  AOI211_X1 U13598 ( .C1(n11345), .C2(n14277), .A(n11616), .B(n14363), .ZN(
        n14272) );
  OAI21_X1 U13599 ( .B1(n10986), .B2(n10985), .A(n10984), .ZN(n10987) );
  NAND2_X1 U13600 ( .A1(n10987), .A2(n14252), .ZN(n10990) );
  AOI22_X1 U13601 ( .A1(n14097), .A2(n13954), .B1(n14082), .B2(n13952), .ZN(
        n10989) );
  INV_X1 U13602 ( .A(n11864), .ZN(n14202) );
  NAND2_X1 U13603 ( .A1(n14274), .A2(n14202), .ZN(n10988) );
  NAND3_X1 U13604 ( .A1(n10990), .A2(n10989), .A3(n10988), .ZN(n14279) );
  AOI211_X1 U13605 ( .C1(n15476), .C2(n14274), .A(n14272), .B(n14279), .ZN(
        n12744) );
  MUX2_X1 U13606 ( .A(n8648), .B(n12744), .S(n15494), .Z(n10991) );
  OAI21_X1 U13607 ( .B1(n12747), .B2(n14428), .A(n10991), .ZN(P2_U3433) );
  INV_X1 U13608 ( .A(n10992), .ZN(n10995) );
  INV_X1 U13609 ( .A(n14011), .ZN(n10993) );
  OAI222_X1 U13610 ( .A1(n12742), .A2(n10994), .B1(n14447), .B2(n10995), .C1(
        n10993), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13611 ( .A(n14654), .ZN(n14657) );
  OAI222_X1 U13612 ( .A1(n15149), .A2(n15692), .B1(n15141), .B2(n10995), .C1(
        n14657), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13613 ( .A(n10996), .ZN(n10997) );
  INV_X1 U13614 ( .A(n15437), .ZN(n12242) );
  OAI222_X1 U13615 ( .A1(n12742), .A2(n15714), .B1(n14447), .B2(n10997), .C1(
        n12242), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13616 ( .A(n12657), .ZN(n12664) );
  OAI222_X1 U13617 ( .A1(n15149), .A2(n10998), .B1(n15141), .B2(n10997), .C1(
        n12664), .C2(P1_U3086), .ZN(P1_U3341) );
  XNOR2_X1 U13618 ( .A(n11002), .B(n11069), .ZN(n11071) );
  OAI21_X1 U13619 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n11001), .A(n10999), .ZN(
        n11072) );
  XOR2_X1 U13620 ( .A(n11071), .B(n11072), .Z(n11010) );
  AND2_X1 U13621 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n11992) );
  NOR2_X1 U13622 ( .A1(n14686), .A2(n11070), .ZN(n11000) );
  AOI211_X1 U13623 ( .C1(n15255), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n11992), .B(
        n11000), .ZN(n11009) );
  NAND2_X1 U13624 ( .A1(n11001), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11004) );
  MUX2_X1 U13625 ( .A(n12055), .B(P1_REG2_REG_9__SCAN_IN), .S(n11002), .Z(
        n11003) );
  AOI21_X1 U13626 ( .B1(n11005), .B2(n11004), .A(n11003), .ZN(n11064) );
  INV_X1 U13627 ( .A(n11064), .ZN(n11007) );
  NAND3_X1 U13628 ( .A1(n11005), .A2(n11004), .A3(n11003), .ZN(n11006) );
  NAND3_X1 U13629 ( .A1(n11007), .A2(n15267), .A3(n11006), .ZN(n11008) );
  OAI211_X1 U13630 ( .C1(n11010), .C2(n14687), .A(n11009), .B(n11008), .ZN(
        P1_U3252) );
  INV_X1 U13631 ( .A(n13324), .ZN(n13317) );
  INV_X1 U13632 ( .A(n11011), .ZN(n11012) );
  OAI222_X1 U13633 ( .A1(P3_U3151), .A2(n13317), .B1(n13705), .B2(n11013), 
        .C1(n13707), .C2(n11012), .ZN(P3_U3277) );
  XNOR2_X1 U13634 ( .A(n11017), .B(n11014), .ZN(n12009) );
  OR2_X1 U13635 ( .A1(n11909), .A2(n11218), .ZN(n11015) );
  NAND2_X1 U13636 ( .A1(n11016), .A2(n11015), .ZN(n11022) );
  NOR2_X1 U13637 ( .A1(n11022), .A2(n14906), .ZN(n11999) );
  NAND2_X1 U13638 ( .A1(n11017), .A2(n14626), .ZN(n11018) );
  AOI21_X1 U13639 ( .B1(n11018), .B2(n15308), .A(n14962), .ZN(n12004) );
  INV_X1 U13640 ( .A(n12004), .ZN(n11020) );
  NOR2_X1 U13641 ( .A1(n14623), .A2(n14916), .ZN(n11019) );
  AOI21_X1 U13642 ( .B1(n11020), .B2(n14626), .A(n11019), .ZN(n12002) );
  INV_X1 U13643 ( .A(n12002), .ZN(n11021) );
  AOI211_X1 U13644 ( .C1(n15302), .C2(n12007), .A(n11999), .B(n11021), .ZN(
        n11024) );
  XNOR2_X1 U13645 ( .A(n11022), .B(n11152), .ZN(n12003) );
  OR3_X1 U13646 ( .A1(n12003), .A2(n12004), .A3(n15007), .ZN(n11023) );
  OAI211_X1 U13647 ( .C1(n15304), .C2(n12009), .A(n11024), .B(n11023), .ZN(
        n11026) );
  NAND2_X1 U13648 ( .A1(n11026), .A2(n15316), .ZN(n11025) );
  OAI21_X1 U13649 ( .B1(n15316), .B2(n9578), .A(n11025), .ZN(P1_U3529) );
  INV_X1 U13650 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15700) );
  NAND2_X1 U13651 ( .A1(n11026), .A2(n15310), .ZN(n11027) );
  OAI21_X1 U13652 ( .B1(n15310), .B2(n15700), .A(n11027), .ZN(P1_U3462) );
  XNOR2_X1 U13653 ( .A(n12238), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n11037) );
  NAND2_X1 U13654 ( .A1(n11039), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U13655 ( .A1(n11029), .A2(n11028), .ZN(n15364) );
  XNOR2_X1 U13656 ( .A(n11042), .B(n11030), .ZN(n15365) );
  NAND2_X1 U13657 ( .A1(n15364), .A2(n15365), .ZN(n15363) );
  NAND2_X1 U13658 ( .A1(n11042), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11031) );
  NAND2_X1 U13659 ( .A1(n15363), .A2(n11031), .ZN(n13973) );
  XNOR2_X1 U13660 ( .A(n13975), .B(n12156), .ZN(n13974) );
  XNOR2_X1 U13661 ( .A(n15383), .B(n12280), .ZN(n15380) );
  NAND2_X1 U13662 ( .A1(n13975), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n15377) );
  AND2_X1 U13663 ( .A1(n15380), .A2(n15377), .ZN(n11032) );
  NAND2_X1 U13664 ( .A1(n15378), .A2(n11032), .ZN(n15379) );
  OR2_X1 U13665 ( .A1(n15383), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11033) );
  XNOR2_X1 U13666 ( .A(n15395), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n15392) );
  NAND2_X1 U13667 ( .A1(n15395), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11034) );
  XNOR2_X1 U13668 ( .A(n11050), .B(n11035), .ZN(n15403) );
  NAND2_X1 U13669 ( .A1(n11036), .A2(n11037), .ZN(n12246) );
  OAI21_X1 U13670 ( .B1(n11037), .B2(n11036), .A(n12246), .ZN(n11058) );
  INV_X1 U13671 ( .A(n15336), .ZN(n15457) );
  INV_X1 U13672 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n12607) );
  NAND2_X1 U13673 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n13789)
         );
  NAND2_X1 U13674 ( .A1(n15450), .A2(n12247), .ZN(n11038) );
  OAI211_X1 U13675 ( .C1(n15457), .C2(n12607), .A(n13789), .B(n11038), .ZN(
        n11057) );
  NAND2_X1 U13676 ( .A1(n11039), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n11040) );
  NAND2_X1 U13677 ( .A1(n11041), .A2(n11040), .ZN(n15371) );
  MUX2_X1 U13678 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11775), .S(n11042), .Z(
        n15372) );
  NAND2_X1 U13679 ( .A1(n11042), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13977) );
  NAND2_X1 U13680 ( .A1(n15370), .A2(n13977), .ZN(n11044) );
  MUX2_X1 U13681 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n12375), .S(n13975), .Z(
        n11043) );
  NAND2_X1 U13682 ( .A1(n11044), .A2(n11043), .ZN(n13979) );
  NAND2_X1 U13683 ( .A1(n13975), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11045) );
  MUX2_X1 U13684 ( .A(n12221), .B(P2_REG2_REG_9__SCAN_IN), .S(n15383), .Z(
        n11046) );
  OR2_X1 U13685 ( .A1(n15383), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n11047) );
  MUX2_X1 U13686 ( .A(n12551), .B(P2_REG2_REG_10__SCAN_IN), .S(n15395), .Z(
        n15397) );
  NAND2_X1 U13687 ( .A1(n15395), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11048) );
  NAND2_X1 U13688 ( .A1(n15398), .A2(n11048), .ZN(n15410) );
  INV_X1 U13689 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11049) );
  MUX2_X1 U13690 ( .A(n11049), .B(P2_REG2_REG_11__SCAN_IN), .S(n11050), .Z(
        n15409) );
  OR2_X1 U13691 ( .A1(n11050), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11053) );
  NAND2_X1 U13692 ( .A1(n15413), .A2(n11053), .ZN(n11051) );
  MUX2_X1 U13693 ( .A(n12443), .B(P2_REG2_REG_12__SCAN_IN), .S(n12238), .Z(
        n11052) );
  NAND2_X1 U13694 ( .A1(n11051), .A2(n11052), .ZN(n12240) );
  INV_X1 U13695 ( .A(n11052), .ZN(n11054) );
  NAND3_X1 U13696 ( .A1(n15413), .A2(n11054), .A3(n11053), .ZN(n11055) );
  AOI21_X1 U13697 ( .B1(n12240), .B2(n11055), .A(n15411), .ZN(n11056) );
  AOI211_X1 U13698 ( .C1(n11058), .C2(n15402), .A(n11057), .B(n11056), .ZN(
        n11059) );
  INV_X1 U13699 ( .A(n11059), .ZN(P2_U3226) );
  INV_X1 U13700 ( .A(n11060), .ZN(n11077) );
  OAI222_X1 U13701 ( .A1(n15149), .A2(n11061), .B1(n15141), .B2(n11077), .C1(
        n12658), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U13702 ( .A(n15255), .ZN(n15271) );
  INV_X1 U13703 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U13704 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12269)
         );
  OAI21_X1 U13705 ( .B1(n15271), .B2(n11578), .A(n12269), .ZN(n11068) );
  NOR2_X1 U13706 ( .A1(n11070), .A2(n12055), .ZN(n11063) );
  MUX2_X1 U13707 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n12189), .S(n11393), .Z(
        n11062) );
  INV_X1 U13708 ( .A(n11396), .ZN(n11066) );
  NOR3_X1 U13709 ( .A1(n11064), .A2(n11063), .A3(n11062), .ZN(n11065) );
  NOR3_X1 U13710 ( .A1(n11066), .A2(n11065), .A3(n14677), .ZN(n11067) );
  AOI211_X1 U13711 ( .C1(n15263), .C2(n11393), .A(n11068), .B(n11067), .ZN(
        n11076) );
  XOR2_X1 U13712 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n11393), .Z(n11073) );
  NAND2_X1 U13713 ( .A1(n11074), .A2(n11073), .ZN(n11386) );
  OAI211_X1 U13714 ( .C1(n11074), .C2(n11073), .A(n11386), .B(n15266), .ZN(
        n11075) );
  NAND2_X1 U13715 ( .A1(n11076), .A2(n11075), .ZN(P1_U3253) );
  OAI222_X1 U13716 ( .A1(n12742), .A2(n11078), .B1(n14447), .B2(n11077), .C1(
        n7246), .C2(P2_U3088), .ZN(P2_U3312) );
  NAND2_X1 U13717 ( .A1(n10982), .A2(n11079), .ZN(n11612) );
  INV_X1 U13718 ( .A(n11622), .ZN(n11611) );
  NAND2_X1 U13719 ( .A1(n11612), .A2(n11611), .ZN(n11610) );
  NAND3_X1 U13720 ( .A1(n11610), .A2(n7117), .A3(n11080), .ZN(n11082) );
  NAND2_X1 U13721 ( .A1(n11082), .A2(n11081), .ZN(n11673) );
  NAND2_X1 U13722 ( .A1(n11615), .A2(n11667), .ZN(n11083) );
  NAND3_X1 U13723 ( .A1(n11651), .A2(n14262), .A3(n11083), .ZN(n11669) );
  INV_X1 U13724 ( .A(n11669), .ZN(n11086) );
  XNOR2_X1 U13725 ( .A(n11084), .B(n7753), .ZN(n11085) );
  AOI22_X1 U13726 ( .A1(n14097), .A2(n13952), .B1(n14082), .B2(n13950), .ZN(
        n11350) );
  OAI21_X1 U13727 ( .B1(n11085), .B2(n14217), .A(n11350), .ZN(n11670) );
  AOI211_X1 U13728 ( .C1(n14366), .C2(n11673), .A(n11086), .B(n11670), .ZN(
        n11417) );
  OAI22_X1 U13729 ( .A1(n14428), .A2(n11414), .B1(n15494), .B2(n8674), .ZN(
        n11087) );
  INV_X1 U13730 ( .A(n11087), .ZN(n11088) );
  OAI21_X1 U13731 ( .B1(n11417), .B2(n15492), .A(n11088), .ZN(P2_U3439) );
  INV_X1 U13732 ( .A(n11089), .ZN(n11092) );
  INV_X1 U13733 ( .A(n14671), .ZN(n14669) );
  OAI222_X1 U13734 ( .A1(n15149), .A2(n11090), .B1(n15141), .B2(n11092), .C1(
        n14669), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13735 ( .A(n15449), .ZN(n11091) );
  OAI222_X1 U13736 ( .A1(n12742), .A2(n11093), .B1(n14447), .B2(n11092), .C1(
        n11091), .C2(P2_U3088), .ZN(P2_U3310) );
  NAND2_X1 U13737 ( .A1(n11095), .A2(n11094), .ZN(n11097) );
  NAND2_X1 U13738 ( .A1(n11097), .A2(n6404), .ZN(n11110) );
  INV_X1 U13739 ( .A(n11110), .ZN(n11099) );
  NAND2_X1 U13740 ( .A1(n11098), .A2(n11783), .ZN(n11111) );
  NAND2_X1 U13741 ( .A1(n11099), .A2(n11111), .ZN(n11112) );
  INV_X1 U13742 ( .A(n13701), .ZN(n11100) );
  MUX2_X1 U13743 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n13703), .Z(n11235) );
  INV_X1 U13744 ( .A(n7124), .ZN(n11102) );
  MUX2_X1 U13745 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n13703), .Z(n11256) );
  XNOR2_X1 U13746 ( .A(n11255), .B(n11256), .ZN(n11257) );
  XNOR2_X1 U13747 ( .A(n11258), .B(n11257), .ZN(n11125) );
  NOR2_X2 U13748 ( .A1(n11112), .A2(n11103), .ZN(n13311) );
  INV_X1 U13749 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n12086) );
  NOR2_X1 U13750 ( .A1(n12086), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U13751 ( .A1(n11104), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11106) );
  INV_X1 U13752 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15547) );
  INV_X1 U13753 ( .A(n11106), .ZN(n11107) );
  NOR2_X1 U13754 ( .A1(n11290), .A2(n11107), .ZN(n11108) );
  AOI21_X1 U13755 ( .B1(n11109), .B2(n11108), .A(n11247), .ZN(n11123) );
  AOI22_X1 U13756 ( .A1(n15503), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11122) );
  INV_X1 U13757 ( .A(n11112), .ZN(n11113) );
  INV_X1 U13758 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n11114) );
  NAND2_X1 U13759 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n11115), .ZN(n11232) );
  INV_X1 U13760 ( .A(n11232), .ZN(n11116) );
  OAI21_X1 U13761 ( .B1(n7124), .B2(n11116), .A(n7860), .ZN(n11284) );
  INV_X1 U13762 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11117) );
  OAI21_X1 U13763 ( .B1(n11119), .B2(n11118), .A(n11241), .ZN(n11120) );
  NAND2_X1 U13764 ( .A1(n13322), .A2(n11120), .ZN(n11121) );
  OAI211_X1 U13765 ( .C1(n13164), .C2(n11123), .A(n11122), .B(n11121), .ZN(
        n11124) );
  AOI21_X1 U13766 ( .B1(n13329), .B2(n11125), .A(n11124), .ZN(n11126) );
  OAI21_X1 U13767 ( .B1(n11255), .B2(n13314), .A(n11126), .ZN(P3_U3184) );
  NAND2_X1 U13768 ( .A1(n11129), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n11130) );
  NAND2_X1 U13769 ( .A1(n11131), .A2(n11130), .ZN(n11140) );
  XNOR2_X1 U13770 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n11132) );
  XNOR2_X1 U13771 ( .A(n11140), .B(n11132), .ZN(n15156) );
  INV_X1 U13772 ( .A(n11133), .ZN(n11134) );
  NAND2_X1 U13773 ( .A1(n11134), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n11135) );
  INV_X1 U13774 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n11137) );
  INV_X1 U13775 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n11138) );
  NAND2_X1 U13776 ( .A1(n11138), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n11139) );
  NAND2_X1 U13777 ( .A1(n11140), .A2(n11139), .ZN(n11143) );
  INV_X1 U13778 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n11141) );
  NAND2_X1 U13779 ( .A1(n11141), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n11142) );
  INV_X1 U13780 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n11144) );
  XNOR2_X1 U13781 ( .A(n11149), .B(n11144), .ZN(n11151) );
  INV_X1 U13782 ( .A(n11151), .ZN(n11145) );
  XNOR2_X1 U13783 ( .A(n11145), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15158) );
  NAND2_X1 U13784 ( .A1(n15157), .A2(n15158), .ZN(n11148) );
  NAND2_X1 U13785 ( .A1(n11146), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n11147) );
  NOR2_X1 U13786 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n11149), .ZN(n11150) );
  XNOR2_X1 U13787 ( .A(n11453), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n11450) );
  XNOR2_X1 U13788 ( .A(n11451), .B(n11450), .ZN(n11446) );
  INV_X1 U13789 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n13970) );
  XNOR2_X1 U13790 ( .A(n11445), .B(n13970), .ZN(SUB_1596_U55) );
  OAI22_X1 U13791 ( .A1(n12855), .A2(n11152), .B1(n11218), .B2(n12857), .ZN(
        n11157) );
  INV_X1 U13792 ( .A(n11153), .ZN(n11154) );
  NAND2_X1 U13793 ( .A1(n11154), .A2(n12866), .ZN(n11155) );
  NAND2_X1 U13794 ( .A1(n11156), .A2(n11155), .ZN(n11217) );
  NAND2_X1 U13795 ( .A1(n11216), .A2(n11217), .ZN(n11161) );
  INV_X1 U13796 ( .A(n11157), .ZN(n11158) );
  NAND2_X1 U13797 ( .A1(n11159), .A2(n11158), .ZN(n11160) );
  NAND2_X1 U13798 ( .A1(n11161), .A2(n11160), .ZN(n11224) );
  OAI22_X1 U13799 ( .A1(n14623), .A2(n12857), .B1(n12755), .B2(n11225), .ZN(
        n11162) );
  XNOR2_X1 U13800 ( .A(n11162), .B(n12875), .ZN(n11165) );
  OAI22_X1 U13801 ( .A1(n12855), .A2(n14623), .B1(n11225), .B2(n12857), .ZN(
        n11163) );
  XNOR2_X1 U13802 ( .A(n11165), .B(n11163), .ZN(n11223) );
  NAND2_X1 U13803 ( .A1(n11224), .A2(n11223), .ZN(n11167) );
  INV_X1 U13804 ( .A(n11163), .ZN(n11164) );
  NAND2_X1 U13805 ( .A1(n11165), .A2(n11164), .ZN(n11166) );
  NAND2_X1 U13806 ( .A1(n11167), .A2(n11166), .ZN(n15239) );
  NAND2_X1 U13807 ( .A1(n12871), .A2(n15234), .ZN(n11170) );
  NAND2_X1 U13808 ( .A1(n11176), .A2(n14622), .ZN(n11169) );
  NAND2_X1 U13809 ( .A1(n11170), .A2(n11169), .ZN(n11171) );
  OAI22_X1 U13810 ( .A1(n12855), .A2(n11596), .B1(n11952), .B2(n12857), .ZN(
        n11173) );
  NAND2_X1 U13811 ( .A1(n11354), .A2(n11174), .ZN(n15238) );
  NAND2_X1 U13812 ( .A1(n12877), .A2(n14621), .ZN(n11178) );
  CLKBUF_X3 U13813 ( .A(n11176), .Z(n12872) );
  NAND2_X1 U13814 ( .A1(n12872), .A2(n6406), .ZN(n11177) );
  AND2_X1 U13815 ( .A1(n11178), .A2(n11177), .ZN(n11355) );
  NAND2_X1 U13816 ( .A1(n12871), .A2(n6406), .ZN(n11180) );
  NAND2_X1 U13817 ( .A1(n11176), .A2(n14621), .ZN(n11179) );
  NAND2_X1 U13818 ( .A1(n11180), .A2(n11179), .ZN(n11181) );
  NAND2_X1 U13819 ( .A1(n12045), .A2(n12871), .ZN(n11185) );
  NAND2_X1 U13820 ( .A1(n12872), .A2(n14620), .ZN(n11184) );
  NAND2_X1 U13821 ( .A1(n11185), .A2(n11184), .ZN(n11186) );
  XNOR2_X1 U13822 ( .A(n11186), .B(n12875), .ZN(n11359) );
  NAND2_X1 U13823 ( .A1(n12877), .A2(n14620), .ZN(n11188) );
  NAND2_X1 U13824 ( .A1(n12045), .A2(n12872), .ZN(n11187) );
  AND2_X1 U13825 ( .A1(n11188), .A2(n11187), .ZN(n11358) );
  AOI22_X1 U13826 ( .A1(n11359), .A2(n11358), .B1(n11355), .B2(n11377), .ZN(
        n11189) );
  INV_X1 U13827 ( .A(n11359), .ZN(n11191) );
  INV_X1 U13828 ( .A(n11358), .ZN(n11190) );
  NAND2_X1 U13829 ( .A1(n11191), .A2(n11190), .ZN(n11192) );
  NAND2_X1 U13830 ( .A1(n12012), .A2(n12871), .ZN(n11195) );
  NAND2_X1 U13831 ( .A1(n12872), .A2(n14619), .ZN(n11194) );
  NAND2_X1 U13832 ( .A1(n11195), .A2(n11194), .ZN(n11196) );
  XNOR2_X1 U13833 ( .A(n11196), .B(n12866), .ZN(n11202) );
  INV_X1 U13834 ( .A(n11202), .ZN(n11200) );
  NAND2_X1 U13835 ( .A1(n12012), .A2(n12872), .ZN(n11198) );
  NAND2_X1 U13836 ( .A1(n12877), .A2(n14619), .ZN(n11197) );
  NAND2_X1 U13837 ( .A1(n11198), .A2(n11197), .ZN(n11201) );
  INV_X1 U13838 ( .A(n11201), .ZN(n11199) );
  AND2_X1 U13839 ( .A1(n11202), .A2(n11201), .ZN(n11526) );
  NOR2_X1 U13840 ( .A1(n7859), .A2(n11526), .ZN(n11203) );
  XNOR2_X1 U13841 ( .A(n11525), .B(n11203), .ZN(n11215) );
  INV_X1 U13842 ( .A(n14618), .ZN(n11882) );
  NOR2_X1 U13843 ( .A1(n14595), .A2(n14918), .ZN(n14560) );
  NAND2_X1 U13844 ( .A1(n14560), .A2(n14620), .ZN(n11205) );
  OAI211_X1 U13845 ( .C1(n11882), .C2(n14556), .A(n11205), .B(n11204), .ZN(
        n11213) );
  NAND3_X1 U13846 ( .A1(n11208), .A2(n11207), .A3(n11206), .ZN(n11209) );
  NAND2_X1 U13847 ( .A1(n11209), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11211) );
  NOR2_X1 U13848 ( .A1(n15246), .A2(n12013), .ZN(n11212) );
  AOI211_X1 U13849 ( .C1(n14586), .C2(n12012), .A(n11213), .B(n11212), .ZN(
        n11214) );
  OAI21_X1 U13850 ( .B1(n11215), .B2(n15237), .A(n11214), .ZN(P1_U3239) );
  XOR2_X1 U13851 ( .A(n11217), .B(n11216), .Z(n11222) );
  INV_X1 U13852 ( .A(n14560), .ZN(n14579) );
  OAI22_X1 U13853 ( .A1(n14579), .A2(n6900), .B1(n14623), .B2(n14556), .ZN(
        n11220) );
  NOR2_X1 U13854 ( .A1(n14600), .A2(n11218), .ZN(n11219) );
  AOI211_X1 U13855 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n11228), .A(n11220), .B(
        n11219), .ZN(n11221) );
  OAI21_X1 U13856 ( .B1(n15237), .B2(n11222), .A(n11221), .ZN(P1_U3222) );
  XOR2_X1 U13857 ( .A(n11224), .B(n11223), .Z(n11230) );
  OAI22_X1 U13858 ( .A1(n14579), .A2(n11152), .B1(n11596), .B2(n14556), .ZN(
        n11227) );
  NOR2_X1 U13859 ( .A1(n14600), .A2(n11225), .ZN(n11226) );
  AOI211_X1 U13860 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n11228), .A(n11227), .B(
        n11226), .ZN(n11229) );
  OAI21_X1 U13861 ( .B1(n15237), .B2(n11230), .A(n11229), .ZN(P1_U3237) );
  NAND3_X1 U13862 ( .A1(n13164), .A2(n13283), .A3(n13303), .ZN(n11234) );
  AOI22_X1 U13863 ( .A1(n15503), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11231) );
  OAI21_X1 U13864 ( .B1(n13283), .B2(n11232), .A(n11231), .ZN(n11233) );
  AOI21_X1 U13865 ( .B1(n11286), .B2(n11234), .A(n11233), .ZN(n11238) );
  AOI22_X1 U13866 ( .A1(n13311), .A2(P3_REG2_REG_0__SCAN_IN), .B1(n13329), 
        .B2(n11235), .ZN(n11236) );
  MUX2_X1 U13867 ( .A(n11236), .B(n13314), .S(P3_IR_REG_0__SCAN_IN), .Z(n11237) );
  NAND2_X1 U13868 ( .A1(n11238), .A2(n11237), .ZN(P3_U3182) );
  OR2_X1 U13869 ( .A1(n7497), .A2(n11114), .ZN(n11240) );
  NAND2_X1 U13870 ( .A1(n11242), .A2(n7495), .ZN(n11243) );
  NAND2_X1 U13871 ( .A1(n11244), .A2(n11243), .ZN(n11325) );
  INV_X1 U13872 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11245) );
  MUX2_X1 U13873 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n11245), .S(n11327), .Z(
        n11326) );
  NAND2_X1 U13874 ( .A1(n11327), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n11246) );
  XNOR2_X1 U13875 ( .A(n11299), .B(n11263), .ZN(n11298) );
  XOR2_X1 U13876 ( .A(n11298), .B(P3_REG1_REG_5__SCAN_IN), .Z(n11271) );
  INV_X1 U13877 ( .A(n11248), .ZN(n11328) );
  XNOR2_X1 U13878 ( .A(n11327), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n11329) );
  OAI21_X1 U13879 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11250), .A(n11315), .ZN(
        n11251) );
  NAND2_X1 U13880 ( .A1(n11251), .A2(n13311), .ZN(n11252) );
  NAND2_X1 U13881 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11760) );
  OAI211_X1 U13882 ( .C1(n11253), .C2(n13291), .A(n11252), .B(n11760), .ZN(
        n11254) );
  AOI21_X1 U13883 ( .B1(n11263), .B2(n13293), .A(n11254), .ZN(n11270) );
  OAI22_X1 U13884 ( .A1(n11258), .A2(n11257), .B1(n11256), .B2(n11255), .ZN(
        n11272) );
  MUX2_X1 U13885 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13703), .Z(n11259) );
  XNOR2_X1 U13886 ( .A(n11259), .B(n11281), .ZN(n11273) );
  INV_X1 U13887 ( .A(n11259), .ZN(n11260) );
  AOI22_X1 U13888 ( .A1(n11272), .A2(n11273), .B1(n11281), .B2(n11260), .ZN(
        n11323) );
  MUX2_X1 U13889 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13703), .Z(n11261) );
  XNOR2_X1 U13890 ( .A(n11261), .B(n11327), .ZN(n11324) );
  MUX2_X1 U13891 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13703), .Z(n11262) );
  NAND2_X1 U13892 ( .A1(n11262), .A2(n7505), .ZN(n11266) );
  INV_X1 U13893 ( .A(n11262), .ZN(n11264) );
  NAND2_X1 U13894 ( .A1(n11264), .A2(n11263), .ZN(n11310) );
  NOR2_X1 U13895 ( .A1(n11311), .A2(n7394), .ZN(n11268) );
  AOI21_X1 U13896 ( .B1(n11310), .B2(n11266), .A(n6706), .ZN(n11267) );
  OAI21_X1 U13897 ( .B1(n11268), .B2(n11267), .A(n13329), .ZN(n11269) );
  OAI211_X1 U13898 ( .C1(n11271), .C2(n13283), .A(n11270), .B(n11269), .ZN(
        P3_U3187) );
  XOR2_X1 U13899 ( .A(n11273), .B(n11272), .Z(n11283) );
  XOR2_X1 U13900 ( .A(n11274), .B(P3_REG1_REG_3__SCAN_IN), .Z(n11279) );
  AOI22_X1 U13901 ( .A1(n15503), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n11278) );
  OAI21_X1 U13902 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n11275), .A(n11330), .ZN(
        n11276) );
  NAND2_X1 U13903 ( .A1(n13311), .A2(n11276), .ZN(n11277) );
  OAI211_X1 U13904 ( .C1(n13283), .C2(n11279), .A(n11278), .B(n11277), .ZN(
        n11280) );
  AOI21_X1 U13905 ( .B1(n11281), .B2(n13293), .A(n11280), .ZN(n11282) );
  OAI21_X1 U13906 ( .B1(n11283), .B2(n13303), .A(n11282), .ZN(P3_U3185) );
  OAI21_X1 U13907 ( .B1(n7123), .B2(P3_REG1_REG_1__SCAN_IN), .A(n11285), .ZN(
        n11295) );
  XOR2_X1 U13908 ( .A(n11287), .B(n11286), .Z(n11289) );
  AOI22_X1 U13909 ( .A1(n15503), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11288) );
  OAI21_X1 U13910 ( .B1(n13303), .B2(n11289), .A(n11288), .ZN(n11294) );
  AOI21_X1 U13911 ( .B1(n15547), .B2(n11291), .A(n11290), .ZN(n11292) );
  NOR2_X1 U13912 ( .A1(n13164), .A2(n11292), .ZN(n11293) );
  AOI211_X1 U13913 ( .C1(n13322), .C2(n11295), .A(n11294), .B(n11293), .ZN(
        n11296) );
  OAI21_X1 U13914 ( .B1(n7124), .B2(n13314), .A(n11296), .ZN(P3_U3183) );
  INV_X1 U13915 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11304) );
  MUX2_X1 U13916 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n11304), .S(n11421), .Z(
        n11303) );
  NAND2_X1 U13917 ( .A1(n11298), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n11301) );
  NAND2_X1 U13918 ( .A1(n11299), .A2(n7505), .ZN(n11300) );
  OAI21_X1 U13919 ( .B1(n11303), .B2(n11302), .A(n11419), .ZN(n11321) );
  INV_X1 U13920 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11715) );
  MUX2_X1 U13921 ( .A(n11715), .B(n11304), .S(n13703), .Z(n11306) );
  INV_X1 U13922 ( .A(n11421), .ZN(n11305) );
  NAND2_X1 U13923 ( .A1(n11306), .A2(n11305), .ZN(n11425) );
  INV_X1 U13924 ( .A(n11306), .ZN(n11307) );
  NAND2_X1 U13925 ( .A1(n11307), .A2(n11421), .ZN(n11308) );
  NAND2_X1 U13926 ( .A1(n11425), .A2(n11308), .ZN(n11309) );
  INV_X1 U13927 ( .A(n11432), .ZN(n11313) );
  NAND3_X1 U13928 ( .A1(n11311), .A2(n11310), .A3(n11309), .ZN(n11312) );
  AOI21_X1 U13929 ( .B1(n11313), .B2(n11312), .A(n13303), .ZN(n11320) );
  XNOR2_X1 U13930 ( .A(n11421), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n11314) );
  AND3_X1 U13931 ( .A1(n11315), .A2(n11314), .A3(n6457), .ZN(n11316) );
  OAI21_X1 U13932 ( .B1(n11420), .B2(n11316), .A(n13311), .ZN(n11318) );
  AND2_X1 U13933 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n12330) );
  AOI21_X1 U13934 ( .B1(n15503), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n12330), .ZN(
        n11317) );
  OAI211_X1 U13935 ( .C1(n13314), .C2(n11421), .A(n11318), .B(n11317), .ZN(
        n11319) );
  AOI211_X1 U13936 ( .C1(n13322), .C2(n11321), .A(n11320), .B(n11319), .ZN(
        n11322) );
  INV_X1 U13937 ( .A(n11322), .ZN(P3_U3188) );
  XOR2_X1 U13938 ( .A(n11324), .B(n11323), .Z(n11338) );
  NOR2_X1 U13939 ( .A1(n13314), .A2(n11327), .ZN(n11335) );
  AND3_X1 U13940 ( .A1(n11330), .A2(n11329), .A3(n11328), .ZN(n11331) );
  OAI21_X1 U13941 ( .B1(n11332), .B2(n11331), .A(n13311), .ZN(n11333) );
  NAND2_X1 U13942 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n12125) );
  OAI211_X1 U13943 ( .C1(n7149), .C2(n13291), .A(n11333), .B(n12125), .ZN(
        n11334) );
  AOI211_X1 U13944 ( .C1(n13322), .C2(n11336), .A(n11335), .B(n11334), .ZN(
        n11337) );
  OAI21_X1 U13945 ( .B1(n11338), .B2(n13303), .A(n11337), .ZN(P3_U3186) );
  INV_X1 U13946 ( .A(n7158), .ZN(n11623) );
  NOR2_X1 U13947 ( .A1(n11339), .A2(P2_U3088), .ZN(n11474) );
  INV_X1 U13948 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11343) );
  AOI21_X1 U13949 ( .B1(n11341), .B2(n14241), .A(n11340), .ZN(n11342) );
  OAI22_X1 U13950 ( .A1(n11474), .A2(n11343), .B1(n13921), .B2(n11342), .ZN(
        n11344) );
  AOI21_X1 U13951 ( .B1(n11345), .B2(n13926), .A(n11344), .ZN(n11346) );
  OAI21_X1 U13952 ( .B1(n11623), .B2(n13900), .A(n11346), .ZN(P2_U3204) );
  XNOR2_X1 U13953 ( .A(n11348), .B(n11347), .ZN(n11353) );
  INV_X1 U13954 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15353) );
  AOI22_X1 U13955 ( .A1(n13917), .A2(n15353), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11349) );
  OAI21_X1 U13956 ( .B1(n11350), .B2(n13919), .A(n11349), .ZN(n11351) );
  AOI21_X1 U13957 ( .B1(n11667), .B2(n13926), .A(n11351), .ZN(n11352) );
  OAI21_X1 U13958 ( .B1(n11353), .B2(n13921), .A(n11352), .ZN(P2_U3190) );
  NAND2_X1 U13959 ( .A1(n15242), .A2(n11354), .ZN(n11357) );
  INV_X1 U13960 ( .A(n11355), .ZN(n11356) );
  NAND2_X1 U13961 ( .A1(n11357), .A2(n11356), .ZN(n11374) );
  NOR2_X1 U13962 ( .A1(n11357), .A2(n11356), .ZN(n11376) );
  AOI21_X1 U13963 ( .B1(n11377), .B2(n11374), .A(n11376), .ZN(n11361) );
  XNOR2_X1 U13964 ( .A(n11359), .B(n11358), .ZN(n11360) );
  XNOR2_X1 U13965 ( .A(n11361), .B(n11360), .ZN(n11362) );
  NAND2_X1 U13966 ( .A1(n11362), .A2(n14589), .ZN(n11368) );
  AND2_X1 U13967 ( .A1(n12045), .A2(n15302), .ZN(n15292) );
  NAND2_X1 U13968 ( .A1(n14960), .A2(n14619), .ZN(n11364) );
  NAND2_X1 U13969 ( .A1(n14962), .A2(n14621), .ZN(n11363) );
  AND2_X1 U13970 ( .A1(n11364), .A2(n11363), .ZN(n12039) );
  OAI21_X1 U13971 ( .B1(n14595), .B2(n12039), .A(n11365), .ZN(n11366) );
  AOI21_X1 U13972 ( .B1(n15236), .B2(n15292), .A(n11366), .ZN(n11367) );
  OAI211_X1 U13973 ( .C1(n15246), .C2(n12046), .A(n11368), .B(n11367), .ZN(
        P1_U3227) );
  INV_X1 U13974 ( .A(n11369), .ZN(n11370) );
  NOR3_X1 U13975 ( .A1(n11540), .A2(n13586), .A3(n11370), .ZN(n11371) );
  AOI21_X1 U13976 ( .B1(n15537), .B2(n13129), .A(n11371), .ZN(n12339) );
  INV_X1 U13977 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11372) );
  MUX2_X1 U13978 ( .A(n12339), .B(n11372), .S(n15583), .Z(n11373) );
  OAI21_X1 U13979 ( .B1(n12342), .B2(n13681), .A(n11373), .ZN(P3_U3390) );
  INV_X1 U13980 ( .A(n11374), .ZN(n11375) );
  NOR2_X1 U13981 ( .A1(n11376), .A2(n11375), .ZN(n11378) );
  XNOR2_X1 U13982 ( .A(n11378), .B(n11377), .ZN(n11379) );
  NAND2_X1 U13983 ( .A1(n11379), .A2(n14589), .ZN(n11385) );
  AND2_X1 U13984 ( .A1(n6406), .A2(n15302), .ZN(n15284) );
  NAND2_X1 U13985 ( .A1(n14960), .A2(n14620), .ZN(n11381) );
  NAND2_X1 U13986 ( .A1(n14962), .A2(n14622), .ZN(n11380) );
  AND2_X1 U13987 ( .A1(n11381), .A2(n11380), .ZN(n15287) );
  OAI21_X1 U13988 ( .B1(n14595), .B2(n15287), .A(n11382), .ZN(n11383) );
  AOI21_X1 U13989 ( .B1(n15236), .B2(n15284), .A(n11383), .ZN(n11384) );
  OAI211_X1 U13990 ( .C1(n15246), .C2(n11960), .A(n11385), .B(n11384), .ZN(
        P1_U3230) );
  XNOR2_X1 U13991 ( .A(n11680), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n11390) );
  INV_X1 U13992 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11387) );
  AOI21_X1 U13993 ( .B1(n11390), .B2(n11389), .A(n11676), .ZN(n11401) );
  NOR2_X1 U13994 ( .A1(n11391), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12533) );
  NOR2_X1 U13995 ( .A1(n14686), .A2(n11678), .ZN(n11392) );
  AOI211_X1 U13996 ( .C1(n15255), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n12533), 
        .B(n11392), .ZN(n11400) );
  NAND2_X1 U13997 ( .A1(n11393), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11395) );
  MUX2_X1 U13998 ( .A(n12292), .B(P1_REG2_REG_11__SCAN_IN), .S(n11680), .Z(
        n11394) );
  INV_X1 U13999 ( .A(n11679), .ZN(n11398) );
  NAND3_X1 U14000 ( .A1(n11396), .A2(n11395), .A3(n11394), .ZN(n11397) );
  NAND3_X1 U14001 ( .A1(n11398), .A2(n15267), .A3(n11397), .ZN(n11399) );
  OAI211_X1 U14002 ( .C1(n11401), .C2(n14687), .A(n11400), .B(n11399), .ZN(
        P1_U3254) );
  INV_X1 U14003 ( .A(n11402), .ZN(n11403) );
  AND3_X1 U14004 ( .A1(n15462), .A2(n11404), .A3(n11403), .ZN(n11405) );
  NAND2_X1 U14005 ( .A1(n15466), .A2(n11405), .ZN(n11406) );
  INV_X1 U14006 ( .A(n14242), .ZN(n14280) );
  NOR2_X1 U14007 ( .A1(n11408), .A2(n11407), .ZN(n15468) );
  OAI21_X1 U14008 ( .B1(n14202), .B2(n14252), .A(n15469), .ZN(n11409) );
  OAI21_X1 U14009 ( .B1(n11623), .B2(n14199), .A(n11409), .ZN(n15467) );
  AOI21_X1 U14010 ( .B1(n11410), .B2(n15468), .A(n15467), .ZN(n11413) );
  NAND2_X1 U14011 ( .A1(n14242), .A2(n11664), .ZN(n11660) );
  INV_X1 U14012 ( .A(n11660), .ZN(n14275) );
  AOI22_X1 U14013 ( .A1(n14275), .A2(n15469), .B1(n14273), .B2(n15468), .ZN(
        n11412) );
  AOI22_X1 U14014 ( .A1(n14280), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n14276), 
        .B2(P2_REG3_REG_0__SCAN_IN), .ZN(n11411) );
  OAI211_X1 U14015 ( .C1(n14280), .C2(n11413), .A(n11412), .B(n11411), .ZN(
        P2_U3265) );
  OAI22_X1 U14016 ( .A1(n14362), .A2(n11414), .B1(n15502), .B2(n15637), .ZN(
        n11415) );
  INV_X1 U14017 ( .A(n11415), .ZN(n11416) );
  OAI21_X1 U14018 ( .B1(n11417), .B2(n15500), .A(n11416), .ZN(P2_U3502) );
  NAND2_X1 U14019 ( .A1(n11421), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11418) );
  INV_X1 U14020 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n12415) );
  XNOR2_X1 U14021 ( .A(n11481), .B(n12415), .ZN(n11439) );
  INV_X1 U14022 ( .A(n11492), .ZN(n11423) );
  OAI21_X1 U14023 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n11424), .A(n11423), .ZN(
        n11437) );
  INV_X1 U14024 ( .A(n11425), .ZN(n11431) );
  INV_X1 U14025 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n12365) );
  MUX2_X1 U14026 ( .A(n12365), .B(n12415), .S(n13703), .Z(n11426) );
  NAND2_X1 U14027 ( .A1(n11426), .A2(n11427), .ZN(n11485) );
  INV_X1 U14028 ( .A(n11426), .ZN(n11428) );
  NAND2_X1 U14029 ( .A1(n11428), .A2(n6897), .ZN(n11429) );
  AND2_X1 U14030 ( .A1(n11485), .A2(n11429), .ZN(n11430) );
  OR3_X1 U14031 ( .A1(n11432), .A2(n11431), .A3(n11430), .ZN(n11433) );
  AOI21_X1 U14032 ( .B1(n11486), .B2(n11433), .A(n13303), .ZN(n11436) );
  NAND2_X1 U14033 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n12206) );
  NAND2_X1 U14034 ( .A1(n15503), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n11434) );
  OAI211_X1 U14035 ( .C1(n13314), .C2(n6897), .A(n12206), .B(n11434), .ZN(
        n11435) );
  AOI211_X1 U14036 ( .C1(n11437), .C2(n13311), .A(n11436), .B(n11435), .ZN(
        n11438) );
  OAI21_X1 U14037 ( .B1(n11439), .B2(n13283), .A(n11438), .ZN(P3_U3189) );
  INV_X1 U14038 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n15689) );
  NAND2_X1 U14039 ( .A1(n13065), .A2(P3_U3897), .ZN(n11440) );
  OAI21_X1 U14040 ( .B1(P3_U3897), .B2(n15689), .A(n11440), .ZN(P3_U3512) );
  INV_X1 U14041 ( .A(n11441), .ZN(n11444) );
  INV_X1 U14042 ( .A(n14682), .ZN(n14672) );
  OAI222_X1 U14043 ( .A1(n15149), .A2(n11442), .B1(n15141), .B2(n11444), .C1(
        n14672), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U14044 ( .A(n14017), .ZN(n14012) );
  OAI222_X1 U14045 ( .A1(P2_U3088), .A2(n14012), .B1(n14447), .B2(n11444), 
        .C1(n11443), .C2(n12742), .ZN(P2_U3309) );
  INV_X1 U14046 ( .A(n11446), .ZN(n11447) );
  OR2_X1 U14047 ( .A1(n11448), .A2(n11447), .ZN(n11449) );
  XOR2_X1 U14048 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), .Z(
        n11454) );
  XNOR2_X1 U14049 ( .A(n11580), .B(n11454), .ZN(n11455) );
  NAND2_X1 U14050 ( .A1(n11575), .A2(n11574), .ZN(n11457) );
  XNOR2_X1 U14051 ( .A(n11457), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  INV_X1 U14052 ( .A(SI_22_), .ZN(n11458) );
  AOI22_X1 U14053 ( .A1(n11459), .A2(P3_STATE_REG_SCAN_IN), .B1(n11458), .B2(
        n6622), .ZN(n11460) );
  OAI21_X1 U14054 ( .B1(n11461), .B2(n13707), .A(n11460), .ZN(n11462) );
  INV_X1 U14055 ( .A(n11462), .ZN(P3_U3273) );
  OAI21_X1 U14056 ( .B1(n11465), .B2(n11464), .A(n11463), .ZN(n11468) );
  OAI22_X1 U14057 ( .A1(n13905), .A2(n15472), .B1(n11474), .B2(n11614), .ZN(
        n11467) );
  OAI22_X1 U14058 ( .A1(n13900), .A2(n11644), .B1(n11623), .B2(n13912), .ZN(
        n11466) );
  AOI211_X1 U14059 ( .C1(n13872), .C2(n11468), .A(n11467), .B(n11466), .ZN(
        n11469) );
  INV_X1 U14060 ( .A(n11469), .ZN(P2_U3209) );
  OAI21_X1 U14061 ( .B1(n11472), .B2(n11471), .A(n11470), .ZN(n11479) );
  INV_X1 U14062 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11473) );
  OAI22_X1 U14063 ( .A1(n13905), .A2(n12747), .B1(n11474), .B2(n11473), .ZN(
        n11478) );
  INV_X1 U14064 ( .A(n13954), .ZN(n11475) );
  OAI22_X1 U14065 ( .A1(n13900), .A2(n11476), .B1(n11475), .B2(n13912), .ZN(
        n11477) );
  AOI211_X1 U14066 ( .C1(n13872), .C2(n11479), .A(n11478), .B(n11477), .ZN(
        n11480) );
  INV_X1 U14067 ( .A(n11480), .ZN(P2_U3194) );
  INV_X1 U14068 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n12336) );
  XNOR2_X1 U14069 ( .A(n11914), .B(n12336), .ZN(n11910) );
  NAND2_X1 U14070 ( .A1(n11482), .A2(n6897), .ZN(n11483) );
  NAND2_X1 U14071 ( .A1(n11484), .A2(n11483), .ZN(n11911) );
  XOR2_X1 U14072 ( .A(n11911), .B(n11910), .Z(n11498) );
  MUX2_X1 U14073 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13703), .Z(n11915) );
  XNOR2_X1 U14074 ( .A(n11915), .B(n11921), .ZN(n11487) );
  OAI21_X1 U14075 ( .B1(n11488), .B2(n11487), .A(n11913), .ZN(n11496) );
  NAND2_X1 U14076 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n12481) );
  NAND2_X1 U14077 ( .A1(n15503), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n11489) );
  OAI211_X1 U14078 ( .C1(n13314), .C2(n11914), .A(n12481), .B(n11489), .ZN(
        n11495) );
  INV_X1 U14079 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12133) );
  XNOR2_X1 U14080 ( .A(n11914), .B(n12133), .ZN(n11490) );
  OR3_X1 U14081 ( .A1(n11492), .A2(n11491), .A3(n11490), .ZN(n11493) );
  AOI21_X1 U14082 ( .B1(n11920), .B2(n11493), .A(n13164), .ZN(n11494) );
  AOI211_X1 U14083 ( .C1(n13329), .C2(n11496), .A(n11495), .B(n11494), .ZN(
        n11497) );
  OAI21_X1 U14084 ( .B1(n11498), .B2(n13283), .A(n11497), .ZN(P3_U3190) );
  OR2_X1 U14085 ( .A1(n11500), .A2(n11499), .ZN(n11502) );
  INV_X1 U14086 ( .A(n11637), .ZN(n11510) );
  OAI21_X1 U14087 ( .B1(n11654), .B2(n11632), .A(n14262), .ZN(n11503) );
  NOR2_X1 U14088 ( .A1(n11503), .A2(n11853), .ZN(n11634) );
  OAI21_X1 U14089 ( .B1(n11506), .B2(n11505), .A(n11504), .ZN(n11507) );
  NAND2_X1 U14090 ( .A1(n11507), .A2(n14252), .ZN(n11509) );
  AOI22_X1 U14091 ( .A1(n14097), .A2(n13950), .B1(n14082), .B2(n13948), .ZN(
        n11508) );
  OAI211_X1 U14092 ( .C1(n11637), .C2(n11864), .A(n11509), .B(n11508), .ZN(
        n11630) );
  AOI211_X1 U14093 ( .C1(n15476), .C2(n11510), .A(n11634), .B(n11630), .ZN(
        n11516) );
  INV_X1 U14094 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11511) );
  OAI22_X1 U14095 ( .A1(n14428), .A2(n11632), .B1(n15494), .B2(n11511), .ZN(
        n11512) );
  INV_X1 U14096 ( .A(n11512), .ZN(n11513) );
  OAI21_X1 U14097 ( .B1(n11516), .B2(n15492), .A(n11513), .ZN(P2_U3445) );
  OAI22_X1 U14098 ( .A1(n14362), .A2(n11632), .B1(n15502), .B2(n8735), .ZN(
        n11514) );
  INV_X1 U14099 ( .A(n11514), .ZN(n11515) );
  OAI21_X1 U14100 ( .B1(n11516), .B2(n15500), .A(n11515), .ZN(P2_U3504) );
  XNOR2_X1 U14101 ( .A(n11518), .B(n11517), .ZN(n11524) );
  OAI21_X1 U14102 ( .B1(n13891), .B2(n11854), .A(n11519), .ZN(n11520) );
  AOI21_X1 U14103 ( .B1(n13909), .B2(n13947), .A(n11520), .ZN(n11521) );
  OAI21_X1 U14104 ( .B1(n11645), .B2(n13912), .A(n11521), .ZN(n11522) );
  AOI21_X1 U14105 ( .B1(n11856), .B2(n13926), .A(n11522), .ZN(n11523) );
  OAI21_X1 U14106 ( .B1(n11524), .B2(n13921), .A(n11523), .ZN(P2_U3211) );
  INV_X1 U14107 ( .A(n15301), .ZN(n12115) );
  NAND2_X1 U14108 ( .A1(n15301), .A2(n12871), .ZN(n11529) );
  NAND2_X1 U14109 ( .A1(n12872), .A2(n14618), .ZN(n11528) );
  NAND2_X1 U14110 ( .A1(n11529), .A2(n11528), .ZN(n11530) );
  XNOR2_X1 U14111 ( .A(n11530), .B(n12866), .ZN(n11823) );
  NOR2_X1 U14112 ( .A1(n12855), .A2(n11882), .ZN(n11531) );
  AOI21_X1 U14113 ( .B1(n15301), .B2(n11176), .A(n11531), .ZN(n11821) );
  XNOR2_X1 U14114 ( .A(n11823), .B(n11821), .ZN(n11532) );
  OAI211_X1 U14115 ( .C1(n11533), .C2(n11532), .A(n11825), .B(n14589), .ZN(
        n11539) );
  INV_X1 U14116 ( .A(n14595), .ZN(n15241) );
  NAND2_X1 U14117 ( .A1(n14960), .A2(n14617), .ZN(n11535) );
  NAND2_X1 U14118 ( .A1(n14962), .A2(n14619), .ZN(n11534) );
  NAND2_X1 U14119 ( .A1(n11535), .A2(n11534), .ZN(n15300) );
  NOR2_X1 U14120 ( .A1(n15246), .A2(n12114), .ZN(n11536) );
  AOI211_X1 U14121 ( .C1(n15241), .C2(n15300), .A(n11537), .B(n11536), .ZN(
        n11538) );
  OAI211_X1 U14122 ( .C1(n12115), .C2(n14600), .A(n11539), .B(n11538), .ZN(
        P1_U3213) );
  NOR2_X1 U14123 ( .A1(n13045), .A2(P3_U3151), .ZN(n11573) );
  INV_X1 U14124 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11544) );
  INV_X1 U14125 ( .A(n11540), .ZN(n11542) );
  OAI22_X1 U14126 ( .A1(n15515), .A2(n13109), .B1(n13103), .B2(n12342), .ZN(
        n11541) );
  AOI21_X1 U14127 ( .B1(n13095), .B2(n11542), .A(n11541), .ZN(n11543) );
  OAI21_X1 U14128 ( .B1(n11573), .B2(n11544), .A(n11543), .ZN(P3_U3172) );
  OAI21_X1 U14129 ( .B1(n11547), .B2(n11546), .A(n11545), .ZN(n11552) );
  NAND2_X1 U14130 ( .A1(n13926), .A2(n15478), .ZN(n11549) );
  OAI211_X1 U14131 ( .C1(n13891), .C2(n11655), .A(n11549), .B(n11548), .ZN(
        n11551) );
  OAI22_X1 U14132 ( .A1(n13900), .A2(n11645), .B1(n11644), .B2(n13912), .ZN(
        n11550) );
  AOI211_X1 U14133 ( .C1(n11552), .C2(n13872), .A(n11551), .B(n11550), .ZN(
        n11553) );
  INV_X1 U14134 ( .A(n11553), .ZN(P2_U3202) );
  INV_X1 U14135 ( .A(n11554), .ZN(n11557) );
  OAI222_X1 U14136 ( .A1(n13707), .A2(n11557), .B1(n13705), .B2(n11556), .C1(
        P3_U3151), .C2(n11555), .ZN(P3_U3275) );
  INV_X1 U14137 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15508) );
  OAI21_X1 U14138 ( .B1(n11560), .B2(n11559), .A(n11558), .ZN(n11561) );
  NAND2_X1 U14139 ( .A1(n11561), .A2(n13095), .ZN(n11564) );
  OAI22_X1 U14140 ( .A1(n15514), .A2(n13109), .B1(n13103), .B2(n15505), .ZN(
        n11562) );
  AOI21_X1 U14141 ( .B1(n13107), .B2(n13129), .A(n11562), .ZN(n11563) );
  OAI211_X1 U14142 ( .C1(n11573), .C2(n15508), .A(n11564), .B(n11563), .ZN(
        P3_U3177) );
  INV_X1 U14143 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11572) );
  NAND3_X1 U14144 ( .A1(n15527), .A2(n15530), .A3(n6399), .ZN(n11565) );
  OAI211_X1 U14145 ( .C1(n11567), .C2(n15531), .A(n11566), .B(n11565), .ZN(
        n11568) );
  NAND2_X1 U14146 ( .A1(n11568), .A2(n13095), .ZN(n11571) );
  OAI22_X1 U14147 ( .A1(n11724), .A2(n13109), .B1(n13103), .B2(n15526), .ZN(
        n11569) );
  AOI21_X1 U14148 ( .B1(n13107), .B2(n15534), .A(n11569), .ZN(n11570) );
  OAI211_X1 U14149 ( .C1(n11573), .C2(n11572), .A(n11571), .B(n11570), .ZN(
        P3_U3162) );
  NAND2_X1 U14150 ( .A1(n11574), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11576) );
  INV_X1 U14151 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11577) );
  NAND2_X1 U14152 ( .A1(n11577), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U14153 ( .A1(n11578), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11579) );
  NAND2_X1 U14154 ( .A1(n12026), .A2(n11579), .ZN(n12025) );
  NAND2_X1 U14155 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(n11580), .ZN(n11582) );
  NOR2_X1 U14156 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(n11580), .ZN(n11581) );
  INV_X1 U14157 ( .A(n12024), .ZN(n11583) );
  XNOR2_X1 U14158 ( .A(n12025), .B(n11583), .ZN(n12021) );
  XNOR2_X1 U14159 ( .A(n12021), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(n11584) );
  XNOR2_X1 U14160 ( .A(n12022), .B(n11584), .ZN(SUB_1596_U70) );
  INV_X1 U14161 ( .A(n11585), .ZN(n11588) );
  OAI222_X1 U14162 ( .A1(n15149), .A2(n11586), .B1(n15141), .B2(n11588), .C1(
        P1_U3086), .C2(n14716), .ZN(P1_U3336) );
  INV_X1 U14163 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11589) );
  OAI222_X1 U14164 ( .A1(n12742), .A2(n11589), .B1(n14447), .B2(n11588), .C1(
        n11587), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U14165 ( .A(n11941), .ZN(n11938) );
  OR2_X1 U14166 ( .A1(n14622), .A2(n15234), .ZN(n11591) );
  NAND2_X1 U14167 ( .A1(n12035), .A2(n12036), .ZN(n12034) );
  OR2_X1 U14168 ( .A1(n12045), .A2(n14620), .ZN(n11592) );
  NAND2_X1 U14169 ( .A1(n12034), .A2(n11592), .ZN(n11593) );
  OAI21_X1 U14170 ( .B1(n11593), .B2(n11602), .A(n11870), .ZN(n11606) );
  INV_X1 U14171 ( .A(n11606), .ZN(n12020) );
  OAI22_X1 U14172 ( .A1(n11882), .A2(n14916), .B1(n11600), .B2(n14918), .ZN(
        n11605) );
  NAND2_X1 U14173 ( .A1(n11754), .A2(n14623), .ZN(n11594) );
  NAND2_X1 U14174 ( .A1(n11596), .A2(n15234), .ZN(n11597) );
  NAND2_X1 U14175 ( .A1(n6862), .A2(n6406), .ZN(n11598) );
  OR2_X1 U14176 ( .A1(n12045), .A2(n11600), .ZN(n11599) );
  NAND2_X1 U14177 ( .A1(n12045), .A2(n11600), .ZN(n11601) );
  XNOR2_X1 U14178 ( .A(n11879), .B(n11602), .ZN(n11603) );
  NOR2_X1 U14179 ( .A1(n11603), .A2(n15007), .ZN(n11604) );
  AOI211_X1 U14180 ( .C1(n14873), .C2(n11606), .A(n11605), .B(n11604), .ZN(
        n12010) );
  INV_X1 U14181 ( .A(n6406), .ZN(n11963) );
  AOI211_X1 U14182 ( .C1(n12012), .C2(n12042), .A(n14893), .B(n12111), .ZN(
        n12016) );
  AOI21_X1 U14183 ( .B1(n15302), .B2(n12012), .A(n12016), .ZN(n11608) );
  OAI211_X1 U14184 ( .C1(n12020), .C2(n15061), .A(n12010), .B(n11608), .ZN(
        n15112) );
  NAND2_X1 U14185 ( .A1(n15112), .A2(n15310), .ZN(n11609) );
  OAI21_X1 U14186 ( .B1(n15310), .B2(n9651), .A(n11609), .ZN(P1_U3477) );
  OAI21_X1 U14187 ( .B1(n11612), .B2(n11611), .A(n11610), .ZN(n15475) );
  INV_X1 U14188 ( .A(n15475), .ZN(n11629) );
  OAI22_X1 U14189 ( .A1(n14242), .A2(n10863), .B1(n11614), .B2(n14239), .ZN(
        n11618) );
  OAI211_X1 U14190 ( .C1(n11616), .C2(n15472), .A(n11615), .B(n14262), .ZN(
        n15471) );
  NOR2_X1 U14191 ( .A1(n14266), .A2(n15471), .ZN(n11617) );
  AOI211_X1 U14192 ( .C1(n14278), .C2(n11619), .A(n11618), .B(n11617), .ZN(
        n11628) );
  OAI21_X1 U14193 ( .B1(n11622), .B2(n11621), .A(n11620), .ZN(n11625) );
  OAI22_X1 U14194 ( .A1(n14199), .A2(n11644), .B1(n11623), .B2(n14197), .ZN(
        n11624) );
  AOI21_X1 U14195 ( .B1(n11625), .B2(n14252), .A(n11624), .ZN(n11626) );
  OAI21_X1 U14196 ( .B1(n11629), .B2(n11864), .A(n11626), .ZN(n15473) );
  NAND2_X1 U14197 ( .A1(n15473), .A2(n14242), .ZN(n11627) );
  OAI211_X1 U14198 ( .C1(n11629), .C2(n11660), .A(n11628), .B(n11627), .ZN(
        P2_U3263) );
  MUX2_X1 U14199 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11630), .S(n14242), .Z(
        n11631) );
  INV_X1 U14200 ( .A(n11631), .ZN(n11636) );
  OAI22_X1 U14201 ( .A1(n14226), .A2(n11632), .B1(n14239), .B2(n13819), .ZN(
        n11633) );
  AOI21_X1 U14202 ( .B1(n14273), .B2(n11634), .A(n11633), .ZN(n11635) );
  OAI211_X1 U14203 ( .C1(n11637), .C2(n11660), .A(n11636), .B(n11635), .ZN(
        P2_U3260) );
  OAI21_X1 U14204 ( .B1(n11640), .B2(n11639), .A(n11638), .ZN(n11646) );
  INV_X1 U14205 ( .A(n11646), .ZN(n15482) );
  OAI21_X1 U14206 ( .B1(n11643), .B2(n11642), .A(n11641), .ZN(n11649) );
  OAI22_X1 U14207 ( .A1(n14199), .A2(n11645), .B1(n11644), .B2(n14197), .ZN(
        n11648) );
  AND2_X1 U14208 ( .A1(n11646), .A2(n14202), .ZN(n11647) );
  AOI211_X1 U14209 ( .C1(n14252), .C2(n11649), .A(n11648), .B(n11647), .ZN(
        n15481) );
  MUX2_X1 U14210 ( .A(n11650), .B(n15481), .S(n14242), .Z(n11659) );
  NAND2_X1 U14211 ( .A1(n11651), .A2(n15478), .ZN(n11652) );
  NAND2_X1 U14212 ( .A1(n11652), .A2(n14262), .ZN(n11653) );
  NOR2_X1 U14213 ( .A1(n11654), .A2(n11653), .ZN(n15477) );
  OAI22_X1 U14214 ( .A1(n14226), .A2(n11656), .B1(n14239), .B2(n11655), .ZN(
        n11657) );
  AOI21_X1 U14215 ( .B1(n14273), .B2(n15477), .A(n11657), .ZN(n11658) );
  OAI211_X1 U14216 ( .C1(n15482), .C2(n11660), .A(n11659), .B(n11658), .ZN(
        P2_U3261) );
  INV_X1 U14217 ( .A(n11661), .ZN(n12932) );
  OAI222_X1 U14218 ( .A1(n12742), .A2(n11663), .B1(P2_U3088), .B2(n11662), 
        .C1(n14447), .C2(n12932), .ZN(P2_U3307) );
  INV_X1 U14219 ( .A(n11664), .ZN(n11665) );
  NAND2_X1 U14220 ( .A1(n11864), .A2(n11665), .ZN(n11666) );
  AOI22_X1 U14221 ( .A1(n14278), .A2(n11667), .B1(n15353), .B2(n14276), .ZN(
        n11668) );
  OAI21_X1 U14222 ( .B1(n14266), .B2(n11669), .A(n11668), .ZN(n11672) );
  MUX2_X1 U14223 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11670), .S(n14242), .Z(
        n11671) );
  AOI211_X1 U14224 ( .C1(n14268), .C2(n11673), .A(n11672), .B(n11671), .ZN(
        n11674) );
  INV_X1 U14225 ( .A(n11674), .ZN(P2_U3262) );
  XNOR2_X1 U14226 ( .A(n11684), .B(n11675), .ZN(n11970) );
  XOR2_X1 U14227 ( .A(n11970), .B(n11971), .Z(n11688) );
  MUX2_X1 U14228 ( .A(n12461), .B(P1_REG2_REG_12__SCAN_IN), .S(n11684), .Z(
        n11682) );
  OAI21_X1 U14229 ( .B1(n11682), .B2(n11681), .A(n11974), .ZN(n11686) );
  NAND2_X1 U14230 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14497)
         );
  NAND2_X1 U14231 ( .A1(n15255), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n11683) );
  OAI211_X1 U14232 ( .C1(n14686), .C2(n11684), .A(n14497), .B(n11683), .ZN(
        n11685) );
  AOI21_X1 U14233 ( .B1(n11686), .B2(n15267), .A(n11685), .ZN(n11687) );
  OAI21_X1 U14234 ( .B1(n11688), .B2(n14687), .A(n11687), .ZN(P1_U3255) );
  INV_X1 U14235 ( .A(n11689), .ZN(n12940) );
  OAI222_X1 U14236 ( .A1(n12742), .A2(n11691), .B1(n14447), .B2(n12940), .C1(
        n11690), .C2(P2_U3088), .ZN(P2_U3306) );
  OR2_X1 U14237 ( .A1(n11692), .A2(n11709), .ZN(n11693) );
  NAND2_X1 U14238 ( .A1(n11694), .A2(n11693), .ZN(n15580) );
  INV_X1 U14239 ( .A(n15580), .ZN(n11720) );
  NAND2_X1 U14240 ( .A1(n11696), .A2(n11695), .ZN(n11698) );
  NAND2_X1 U14241 ( .A1(n11698), .A2(n11697), .ZN(n11700) );
  AND2_X1 U14242 ( .A1(n11700), .A2(n11699), .ZN(n11701) );
  NAND2_X1 U14243 ( .A1(n11702), .A2(n11701), .ZN(n11716) );
  INV_X1 U14244 ( .A(n15507), .ZN(n15543) );
  NAND2_X1 U14245 ( .A1(n15507), .A2(n11704), .ZN(n12302) );
  INV_X1 U14246 ( .A(n12302), .ZN(n15523) );
  INV_X1 U14247 ( .A(n15545), .ZN(n12136) );
  INV_X1 U14248 ( .A(n15521), .ZN(n15528) );
  NAND2_X1 U14249 ( .A1(n15580), .A2(n15528), .ZN(n11714) );
  AOI22_X1 U14250 ( .A1(n15537), .A2(n13124), .B1(n15535), .B2(n13126), .ZN(
        n11713) );
  OR2_X1 U14251 ( .A1(n11705), .A2(n12167), .ZN(n12169) );
  INV_X1 U14252 ( .A(n11708), .ZN(n11706) );
  NAND2_X1 U14253 ( .A1(n12169), .A2(n11706), .ZN(n11707) );
  NAND2_X1 U14254 ( .A1(n11707), .A2(n11709), .ZN(n11711) );
  NOR2_X1 U14255 ( .A1(n11709), .A2(n11708), .ZN(n11710) );
  NAND2_X1 U14256 ( .A1(n12169), .A2(n11710), .ZN(n11787) );
  NAND3_X1 U14257 ( .A1(n11711), .A2(n15532), .A3(n11787), .ZN(n11712) );
  AND3_X1 U14258 ( .A1(n11714), .A2(n11713), .A3(n11712), .ZN(n15582) );
  MUX2_X1 U14259 ( .A(n11715), .B(n15582), .S(n15524), .Z(n11719) );
  OR2_X1 U14260 ( .A1(n11716), .A2(n15507), .ZN(n12166) );
  NOR2_X1 U14261 ( .A1(n15567), .A2(n11717), .ZN(n15578) );
  AOI22_X1 U14262 ( .A1(n12084), .A2(n15578), .B1(n15544), .B2(n12323), .ZN(
        n11718) );
  OAI211_X1 U14263 ( .C1(n11720), .C2(n12136), .A(n11719), .B(n11718), .ZN(
        P3_U3227) );
  OAI21_X1 U14264 ( .B1(n11723), .B2(n11722), .A(n11721), .ZN(n15562) );
  INV_X1 U14265 ( .A(n15562), .ZN(n11735) );
  INV_X1 U14266 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11732) );
  OAI22_X1 U14267 ( .A1(n15516), .A2(n11724), .B1(n12355), .B2(n15513), .ZN(
        n11731) );
  INV_X1 U14268 ( .A(n11725), .ZN(n11729) );
  AOI21_X1 U14269 ( .B1(n15510), .B2(n11727), .A(n11726), .ZN(n11728) );
  NOR3_X1 U14270 ( .A1(n11729), .A2(n11728), .A3(n13522), .ZN(n11730) );
  AOI211_X1 U14271 ( .C1(n15528), .C2(n15562), .A(n11731), .B(n11730), .ZN(
        n15559) );
  MUX2_X1 U14272 ( .A(n11732), .B(n15559), .S(n15524), .Z(n11734) );
  NOR2_X1 U14273 ( .A1(n15567), .A2(n12354), .ZN(n15561) );
  AOI22_X1 U14274 ( .A1(n12084), .A2(n15561), .B1(n15544), .B2(n12356), .ZN(
        n11733) );
  OAI211_X1 U14275 ( .C1(n11735), .C2(n12136), .A(n11734), .B(n11733), .ZN(
        P3_U3230) );
  INV_X1 U14276 ( .A(n11736), .ZN(n11737) );
  NAND2_X1 U14277 ( .A1(n11738), .A2(n11737), .ZN(n11750) );
  INV_X1 U14278 ( .A(n11742), .ZN(n11743) );
  AND2_X1 U14279 ( .A1(n14940), .A2(n11743), .ZN(n14879) );
  INV_X1 U14280 ( .A(n14879), .ZN(n12019) );
  MUX2_X1 U14281 ( .A(n11745), .B(n11744), .S(n14940), .Z(n11756) );
  NOR2_X1 U14282 ( .A1(n11746), .A2(n10007), .ZN(n11747) );
  NAND2_X1 U14283 ( .A1(n11748), .A2(n14716), .ZN(n11749) );
  OAI22_X1 U14284 ( .A1(n14953), .A2(n11752), .B1(n11751), .B2(n14946), .ZN(
        n11753) );
  AOI21_X1 U14285 ( .B1(n14956), .B2(n11754), .A(n11753), .ZN(n11755) );
  OAI211_X1 U14286 ( .C1(n11757), .C2(n12019), .A(n11756), .B(n11755), .ZN(
        P1_U3291) );
  AOI21_X1 U14287 ( .B1(n6602), .B2(n11759), .A(n11758), .ZN(n11764) );
  AOI22_X1 U14288 ( .A1(n13107), .A2(n13127), .B1(n13100), .B2(n13125), .ZN(
        n11761) );
  OAI211_X1 U14289 ( .C1(n13103), .C2(n12163), .A(n11761), .B(n11760), .ZN(
        n11762) );
  AOI21_X1 U14290 ( .B1(n12164), .B2(n13045), .A(n11762), .ZN(n11763) );
  OAI21_X1 U14291 ( .B1(n11764), .B2(n13115), .A(n11763), .ZN(P3_U3167) );
  INV_X1 U14292 ( .A(n11765), .ZN(n11768) );
  OAI222_X1 U14293 ( .A1(n13707), .A2(n11768), .B1(n13705), .B2(n11767), .C1(
        P3_U3151), .C2(n11766), .ZN(P3_U3274) );
  OAI21_X1 U14294 ( .B1(n6685), .B2(n11771), .A(n11769), .ZN(n11815) );
  INV_X1 U14295 ( .A(n11815), .ZN(n11780) );
  XNOR2_X1 U14296 ( .A(n11772), .B(n11771), .ZN(n11773) );
  AOI22_X1 U14297 ( .A1(n13946), .A2(n14082), .B1(n14097), .B2(n13948), .ZN(
        n11798) );
  OAI21_X1 U14298 ( .B1(n11773), .B2(n14217), .A(n11798), .ZN(n11813) );
  INV_X1 U14299 ( .A(n11813), .ZN(n11774) );
  MUX2_X1 U14300 ( .A(n11775), .B(n11774), .S(n14242), .Z(n11779) );
  AOI21_X1 U14301 ( .B1(n11852), .B2(n11844), .A(n14363), .ZN(n11776) );
  AND2_X1 U14302 ( .A1(n11776), .A2(n6614), .ZN(n11814) );
  OAI22_X1 U14303 ( .A1(n14226), .A2(n6837), .B1(n14239), .B2(n11797), .ZN(
        n11777) );
  AOI21_X1 U14304 ( .B1(n14273), .B2(n11814), .A(n11777), .ZN(n11778) );
  OAI211_X1 U14305 ( .C1(n11780), .C2(n14248), .A(n11779), .B(n11778), .ZN(
        P2_U3258) );
  NAND2_X1 U14306 ( .A1(n11782), .A2(n11781), .ZN(n11784) );
  OAI211_X1 U14307 ( .C1(n11785), .C2(n13705), .A(n11784), .B(n11783), .ZN(
        P3_U3272) );
  NAND2_X1 U14308 ( .A1(n11787), .A2(n11786), .ZN(n11788) );
  XNOR2_X1 U14309 ( .A(n11788), .B(n11791), .ZN(n11789) );
  OAI222_X1 U14310 ( .A1(n15513), .A2(n13034), .B1(n15516), .B2(n11790), .C1(
        n11789), .C2(n13522), .ZN(n12362) );
  AOI21_X1 U14311 ( .B1(n13586), .B2(n12366), .A(n12362), .ZN(n12414) );
  XNOR2_X1 U14312 ( .A(n11792), .B(n11791), .ZN(n12417) );
  OR2_X1 U14313 ( .A1(n12417), .A2(n13673), .ZN(n11794) );
  NAND2_X1 U14314 ( .A1(n15583), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n11793) );
  OAI211_X1 U14315 ( .C1(n12414), .C2(n15583), .A(n11794), .B(n11793), .ZN(
        P3_U3411) );
  XNOR2_X1 U14316 ( .A(n11795), .B(n11796), .ZN(n11802) );
  NAND2_X1 U14317 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15367) );
  OAI21_X1 U14318 ( .B1(n13891), .B2(n11797), .A(n15367), .ZN(n11800) );
  NOR2_X1 U14319 ( .A1(n13919), .A2(n11798), .ZN(n11799) );
  AOI211_X1 U14320 ( .C1(n11844), .C2(n13926), .A(n11800), .B(n11799), .ZN(
        n11801) );
  OAI21_X1 U14321 ( .B1(n11802), .B2(n13921), .A(n11801), .ZN(P2_U3185) );
  XNOR2_X1 U14322 ( .A(n11803), .B(n11804), .ZN(n12628) );
  AOI22_X1 U14323 ( .A1(n13670), .A2(n13038), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n15583), .ZN(n11812) );
  NOR2_X1 U14324 ( .A1(n11839), .A2(n7645), .ZN(n11838) );
  INV_X1 U14325 ( .A(n11838), .ZN(n11806) );
  AOI21_X1 U14326 ( .B1(n11806), .B2(n11805), .A(n11804), .ZN(n11810) );
  OR2_X1 U14327 ( .A1(n11838), .A2(n11807), .ZN(n12230) );
  NAND2_X1 U14328 ( .A1(n12230), .A2(n15532), .ZN(n11809) );
  AOI22_X1 U14329 ( .A1(n15537), .A2(n13122), .B1(n15535), .B2(n12205), .ZN(
        n11808) );
  OAI21_X1 U14330 ( .B1(n11810), .B2(n11809), .A(n11808), .ZN(n12625) );
  NAND2_X1 U14331 ( .A1(n12625), .A2(n15585), .ZN(n11811) );
  OAI211_X1 U14332 ( .C1(n12628), .C2(n13673), .A(n11812), .B(n11811), .ZN(
        P3_U3417) );
  AOI211_X1 U14333 ( .C1(n14366), .C2(n11815), .A(n11814), .B(n11813), .ZN(
        n11847) );
  INV_X1 U14334 ( .A(n14428), .ZN(n14434) );
  AOI22_X1 U14335 ( .A1(n14434), .A2(n11844), .B1(P2_REG0_REG_7__SCAN_IN), 
        .B2(n15492), .ZN(n11816) );
  OAI21_X1 U14336 ( .B1(n11847), .B2(n15492), .A(n11816), .ZN(P2_U3451) );
  NAND2_X1 U14337 ( .A1(n12101), .A2(n12871), .ZN(n11818) );
  NAND2_X1 U14338 ( .A1(n12872), .A2(n14617), .ZN(n11817) );
  NAND2_X1 U14339 ( .A1(n11818), .A2(n11817), .ZN(n11819) );
  XNOR2_X1 U14340 ( .A(n11819), .B(n12875), .ZN(n11983) );
  NOR2_X1 U14341 ( .A1(n12855), .A2(n11886), .ZN(n11820) );
  AOI21_X1 U14342 ( .B1(n12101), .B2(n11176), .A(n11820), .ZN(n11982) );
  XNOR2_X1 U14343 ( .A(n11983), .B(n11982), .ZN(n11829) );
  INV_X1 U14344 ( .A(n11821), .ZN(n11822) );
  NAND2_X1 U14345 ( .A1(n11823), .A2(n11822), .ZN(n11824) );
  INV_X1 U14346 ( .A(n11985), .ZN(n11827) );
  AOI21_X1 U14347 ( .B1(n11829), .B2(n11828), .A(n11827), .ZN(n11835) );
  INV_X1 U14348 ( .A(n12101), .ZN(n12103) );
  NOR2_X1 U14349 ( .A1(n12103), .A2(n15065), .ZN(n15108) );
  NAND2_X1 U14350 ( .A1(n14960), .A2(n14616), .ZN(n11831) );
  NAND2_X1 U14351 ( .A1(n14962), .A2(n14618), .ZN(n11830) );
  NAND2_X1 U14352 ( .A1(n11831), .A2(n11830), .ZN(n15106) );
  AOI22_X1 U14353 ( .A1(n15241), .A2(n15106), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11832) );
  OAI21_X1 U14354 ( .B1(n15246), .B2(n12102), .A(n11832), .ZN(n11833) );
  AOI21_X1 U14355 ( .B1(n15236), .B2(n15108), .A(n11833), .ZN(n11834) );
  OAI21_X1 U14356 ( .B1(n11835), .B2(n15237), .A(n11834), .ZN(P1_U3221) );
  INV_X1 U14357 ( .A(n13555), .ZN(n15579) );
  XNOR2_X1 U14358 ( .A(n11837), .B(n11836), .ZN(n12130) );
  AOI21_X1 U14359 ( .B1(n7645), .B2(n11839), .A(n11838), .ZN(n11842) );
  NAND2_X1 U14360 ( .A1(n12130), .A2(n15528), .ZN(n11841) );
  AOI22_X1 U14361 ( .A1(n15537), .A2(n13123), .B1(n15535), .B2(n13124), .ZN(
        n11840) );
  OAI211_X1 U14362 ( .C1(n13522), .C2(n11842), .A(n11841), .B(n11840), .ZN(
        n12131) );
  AOI21_X1 U14363 ( .B1(n15579), .B2(n12130), .A(n12131), .ZN(n12335) );
  AOI22_X1 U14364 ( .A1(n13670), .A2(n12480), .B1(n15583), .B2(
        P3_REG0_REG_8__SCAN_IN), .ZN(n11843) );
  OAI21_X1 U14365 ( .B1(n12335), .B2(n15583), .A(n11843), .ZN(P3_U3414) );
  NAND2_X1 U14366 ( .A1(n15500), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11846) );
  INV_X1 U14367 ( .A(n14362), .ZN(n14374) );
  NAND2_X1 U14368 ( .A1(n14374), .A2(n11844), .ZN(n11845) );
  OAI211_X1 U14369 ( .C1(n11847), .C2(n15500), .A(n11846), .B(n11845), .ZN(
        P2_U3506) );
  OR2_X1 U14370 ( .A1(n11849), .A2(n11848), .ZN(n11850) );
  INV_X1 U14371 ( .A(n15485), .ZN(n11867) );
  OAI211_X1 U14372 ( .C1(n11853), .C2(n15488), .A(n14262), .B(n11852), .ZN(
        n15486) );
  INV_X1 U14373 ( .A(n11854), .ZN(n11855) );
  AOI22_X1 U14374 ( .A1(n14278), .A2(n11856), .B1(n14276), .B2(n11855), .ZN(
        n11857) );
  OAI21_X1 U14375 ( .B1(n14266), .B2(n15486), .A(n11857), .ZN(n11866) );
  OAI21_X1 U14376 ( .B1(n11860), .B2(n11859), .A(n11858), .ZN(n11861) );
  NAND2_X1 U14377 ( .A1(n11861), .A2(n14252), .ZN(n11863) );
  AOI22_X1 U14378 ( .A1(n13947), .A2(n14082), .B1(n14097), .B2(n13949), .ZN(
        n11862) );
  OAI211_X1 U14379 ( .C1(n15485), .C2(n11864), .A(n11863), .B(n11862), .ZN(
        n15491) );
  MUX2_X1 U14380 ( .A(n15491), .B(P2_REG2_REG_6__SCAN_IN), .S(n14280), .Z(
        n11865) );
  AOI211_X1 U14381 ( .C1(n14275), .C2(n11867), .A(n11866), .B(n11865), .ZN(
        n11868) );
  INV_X1 U14382 ( .A(n11868), .ZN(P2_U3259) );
  OR2_X1 U14383 ( .A1(n12012), .A2(n14619), .ZN(n11869) );
  INV_X1 U14384 ( .A(n12119), .ZN(n12108) );
  NAND2_X1 U14385 ( .A1(n12109), .A2(n12108), .ZN(n12107) );
  OR2_X1 U14386 ( .A1(n15301), .A2(n14618), .ZN(n11871) );
  OR2_X1 U14387 ( .A1(n12101), .A2(n14617), .ZN(n11872) );
  OAI21_X1 U14388 ( .B1(n11873), .B2(n11888), .A(n12177), .ZN(n12051) );
  AOI21_X1 U14389 ( .B1(n12098), .B2(n12183), .A(n14893), .ZN(n11874) );
  NAND2_X1 U14390 ( .A1(n11874), .A2(n6795), .ZN(n12056) );
  NAND2_X1 U14391 ( .A1(n14960), .A2(n14615), .ZN(n11876) );
  NAND2_X1 U14392 ( .A1(n14962), .A2(n14617), .ZN(n11875) );
  NAND2_X1 U14393 ( .A1(n11876), .A2(n11875), .ZN(n12052) );
  INV_X1 U14394 ( .A(n12052), .ZN(n11877) );
  NAND2_X1 U14395 ( .A1(n12183), .A2(n15302), .ZN(n11997) );
  NAND3_X1 U14396 ( .A1(n12056), .A2(n11877), .A3(n11997), .ZN(n11891) );
  INV_X1 U14397 ( .A(n14619), .ZN(n11880) );
  NAND2_X1 U14398 ( .A1(n12012), .A2(n11880), .ZN(n11881) );
  NAND2_X1 U14399 ( .A1(n12118), .A2(n12119), .ZN(n11884) );
  NAND2_X1 U14400 ( .A1(n15301), .A2(n11882), .ZN(n11883) );
  OR2_X1 U14401 ( .A1(n12101), .A2(n11886), .ZN(n11887) );
  NAND2_X1 U14402 ( .A1(n11889), .A2(n11888), .ZN(n11890) );
  AOI21_X1 U14403 ( .B1(n12185), .B2(n11890), .A(n15007), .ZN(n12053) );
  AOI211_X1 U14404 ( .C1(n15297), .C2(n12051), .A(n11891), .B(n12053), .ZN(
        n11894) );
  NAND2_X1 U14405 ( .A1(n15309), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11892) );
  OAI21_X1 U14406 ( .B1(n11894), .B2(n15309), .A(n11892), .ZN(P1_U3486) );
  NAND2_X1 U14407 ( .A1(n15314), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11893) );
  OAI21_X1 U14408 ( .B1(n11894), .B2(n15314), .A(n11893), .ZN(P1_U3537) );
  INV_X1 U14409 ( .A(n11895), .ZN(n11897) );
  OAI222_X1 U14410 ( .A1(n12742), .A2(n11898), .B1(n14447), .B2(n11897), .C1(
        n11896), .C2(P2_U3088), .ZN(P2_U3305) );
  NOR3_X1 U14411 ( .A1(n11909), .A2(n14893), .A3(n7274), .ZN(n11899) );
  OAI21_X1 U14412 ( .B1(n11900), .B2(n11899), .A(n14940), .ZN(n11901) );
  OAI21_X1 U14413 ( .B1(n14946), .B2(n11902), .A(n11901), .ZN(n11903) );
  AOI21_X1 U14414 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14920), .A(n11903), .ZN(
        n11908) );
  NAND2_X1 U14415 ( .A1(n14940), .A2(n15308), .ZN(n14754) );
  INV_X1 U14416 ( .A(n11904), .ZN(n11905) );
  OAI21_X1 U14417 ( .B1(n14864), .B2(n14841), .A(n11906), .ZN(n11907) );
  OAI211_X1 U14418 ( .C1(n14937), .C2(n11909), .A(n11908), .B(n11907), .ZN(
        P1_U3293) );
  NAND2_X1 U14419 ( .A1(n11914), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11912) );
  INV_X1 U14420 ( .A(n11922), .ZN(n12067) );
  XOR2_X1 U14421 ( .A(n12066), .B(P3_REG1_REG_9__SCAN_IN), .Z(n11930) );
  MUX2_X1 U14422 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13703), .Z(n11916) );
  NOR2_X1 U14423 ( .A1(n11916), .A2(n11922), .ZN(n12068) );
  NAND2_X1 U14424 ( .A1(n11916), .A2(n11922), .ZN(n12069) );
  INV_X1 U14425 ( .A(n12069), .ZN(n11917) );
  NOR2_X1 U14426 ( .A1(n12068), .A2(n11917), .ZN(n11918) );
  XNOR2_X1 U14427 ( .A(n12070), .B(n11918), .ZN(n11928) );
  NAND2_X1 U14428 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n13032) );
  NAND2_X1 U14429 ( .A1(n15503), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11919) );
  OAI211_X1 U14430 ( .C1(n13314), .C2(n11922), .A(n13032), .B(n11919), .ZN(
        n11927) );
  NAND2_X1 U14431 ( .A1(n11923), .A2(n11922), .ZN(n12075) );
  NAND2_X1 U14432 ( .A1(n11924), .A2(n7509), .ZN(n11925) );
  AOI21_X1 U14433 ( .B1(n12077), .B2(n11925), .A(n13164), .ZN(n11926) );
  AOI211_X1 U14434 ( .C1(n11928), .C2(n13329), .A(n11927), .B(n11926), .ZN(
        n11929) );
  OAI21_X1 U14435 ( .B1(n11930), .B2(n13283), .A(n11929), .ZN(P3_U3191) );
  INV_X1 U14436 ( .A(n11931), .ZN(n11936) );
  AOI21_X1 U14437 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14445), .A(n11932), 
        .ZN(n11933) );
  OAI21_X1 U14438 ( .B1(n11936), .B2(n14447), .A(n11933), .ZN(P2_U3304) );
  AOI21_X1 U14439 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n11934), .A(n10050), 
        .ZN(n11935) );
  OAI21_X1 U14440 ( .B1(n11936), .B2(n15141), .A(n11935), .ZN(P1_U3332) );
  OAI21_X1 U14441 ( .B1(n11939), .B2(n11938), .A(n11937), .ZN(n15281) );
  OAI21_X1 U14442 ( .B1(n11942), .B2(n11941), .A(n11940), .ZN(n11943) );
  NAND2_X1 U14443 ( .A1(n11943), .A2(n15308), .ZN(n11948) );
  OR2_X1 U14444 ( .A1(n14623), .A2(n14918), .ZN(n11945) );
  NAND2_X1 U14445 ( .A1(n14960), .A2(n14621), .ZN(n11944) );
  NAND2_X1 U14446 ( .A1(n11945), .A2(n11944), .ZN(n15240) );
  INV_X1 U14447 ( .A(n15240), .ZN(n11947) );
  NAND2_X1 U14448 ( .A1(n15281), .A2(n14873), .ZN(n11946) );
  NAND3_X1 U14449 ( .A1(n11948), .A2(n11947), .A3(n11946), .ZN(n15280) );
  MUX2_X1 U14450 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n15280), .S(n14940), .Z(
        n11954) );
  AOI211_X1 U14451 ( .C1(n15234), .C2(n11949), .A(n14893), .B(n11959), .ZN(
        n15276) );
  INV_X1 U14452 ( .A(n14946), .ZN(n14934) );
  INV_X1 U14453 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U14454 ( .A1(n15276), .A2(n14924), .B1(n14934), .B2(n11950), .ZN(
        n11951) );
  OAI21_X1 U14455 ( .B1(n11952), .B2(n14937), .A(n11951), .ZN(n11953) );
  AOI211_X1 U14456 ( .C1(n14879), .C2(n15281), .A(n11954), .B(n11953), .ZN(
        n11955) );
  INV_X1 U14457 ( .A(n11955), .ZN(P1_U3290) );
  OAI21_X1 U14458 ( .B1(n11958), .B2(n11957), .A(n11956), .ZN(n15290) );
  OAI211_X1 U14459 ( .C1(n11959), .C2(n11963), .A(n12044), .B(n14949), .ZN(
        n15285) );
  OAI22_X1 U14460 ( .A1(n15285), .A2(n14953), .B1(n11960), .B2(n14946), .ZN(
        n11961) );
  AOI21_X1 U14461 ( .B1(n14920), .B2(P1_REG2_REG_4__SCAN_IN), .A(n11961), .ZN(
        n11962) );
  OAI21_X1 U14462 ( .B1(n11963), .B2(n14937), .A(n11962), .ZN(n11968) );
  OAI21_X1 U14463 ( .B1(n11965), .B2(n6860), .A(n11964), .ZN(n11966) );
  NAND2_X1 U14464 ( .A1(n11966), .A2(n15308), .ZN(n15288) );
  AOI21_X1 U14465 ( .B1(n15288), .B2(n15287), .A(n14920), .ZN(n11967) );
  AOI211_X1 U14466 ( .C1(n14841), .C2(n15290), .A(n11968), .B(n11967), .ZN(
        n11969) );
  INV_X1 U14467 ( .A(n11969), .ZN(P1_U3289) );
  XNOR2_X1 U14468 ( .A(n12388), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11973) );
  NOR2_X1 U14469 ( .A1(n11972), .A2(n11973), .ZN(n12387) );
  AOI211_X1 U14470 ( .C1(n11973), .C2(n11972), .A(n14687), .B(n12387), .ZN(
        n11981) );
  OAI21_X1 U14471 ( .B1(n11975), .B2(P1_REG2_REG_12__SCAN_IN), .A(n11974), 
        .ZN(n11977) );
  INV_X1 U14472 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n15702) );
  MUX2_X1 U14473 ( .A(n15702), .B(P1_REG2_REG_13__SCAN_IN), .S(n12388), .Z(
        n11976) );
  NOR2_X1 U14474 ( .A1(n11977), .A2(n11976), .ZN(n12397) );
  AOI211_X1 U14475 ( .C1(n11977), .C2(n11976), .A(n14677), .B(n12397), .ZN(
        n11980) );
  NAND2_X1 U14476 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14554)
         );
  NAND2_X1 U14477 ( .A1(n15255), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n11978) );
  OAI211_X1 U14478 ( .C1(n14686), .C2(n12391), .A(n14554), .B(n11978), .ZN(
        n11979) );
  OR3_X1 U14479 ( .A1(n11981), .A2(n11980), .A3(n11979), .ZN(P1_U3256) );
  INV_X1 U14480 ( .A(n15236), .ZN(n11998) );
  NAND2_X1 U14481 ( .A1(n11983), .A2(n11982), .ZN(n11984) );
  NAND2_X1 U14482 ( .A1(n12183), .A2(n12871), .ZN(n11987) );
  NAND2_X1 U14483 ( .A1(n12872), .A2(n14616), .ZN(n11986) );
  NAND2_X1 U14484 ( .A1(n11987), .A2(n11986), .ZN(n11988) );
  XNOR2_X1 U14485 ( .A(n11988), .B(n12866), .ZN(n12260) );
  NOR2_X1 U14486 ( .A1(n12855), .A2(n12182), .ZN(n11989) );
  AOI21_X1 U14487 ( .B1(n12183), .B2(n11176), .A(n11989), .ZN(n12258) );
  XNOR2_X1 U14488 ( .A(n12260), .B(n12258), .ZN(n11990) );
  OAI211_X1 U14489 ( .C1(n11991), .C2(n11990), .A(n12262), .B(n14589), .ZN(
        n11996) );
  AOI21_X1 U14490 ( .B1(n15241), .B2(n12052), .A(n11992), .ZN(n11993) );
  OAI21_X1 U14491 ( .B1(n15246), .B2(n12057), .A(n11993), .ZN(n11994) );
  INV_X1 U14492 ( .A(n11994), .ZN(n11995) );
  OAI211_X1 U14493 ( .C1(n11998), .C2(n11997), .A(n11996), .B(n11995), .ZN(
        P1_U3231) );
  AOI22_X1 U14494 ( .A1(n14924), .A2(n11999), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14934), .ZN(n12001) );
  OR2_X1 U14495 ( .A1(n14940), .A2(n10701), .ZN(n12000) );
  OAI211_X1 U14496 ( .C1(n14920), .C2(n12002), .A(n12001), .B(n12000), .ZN(
        n12006) );
  NOR3_X1 U14497 ( .A1(n14754), .A2(n12004), .A3(n12003), .ZN(n12005) );
  AOI211_X1 U14498 ( .C1(n14956), .C2(n12007), .A(n12006), .B(n12005), .ZN(
        n12008) );
  OAI21_X1 U14499 ( .B1(n14969), .B2(n12009), .A(n12008), .ZN(P1_U3292) );
  MUX2_X1 U14500 ( .A(n12011), .B(n12010), .S(n14940), .Z(n12018) );
  INV_X1 U14501 ( .A(n12012), .ZN(n12014) );
  OAI22_X1 U14502 ( .A1(n14937), .A2(n12014), .B1(n12013), .B2(n14946), .ZN(
        n12015) );
  AOI21_X1 U14503 ( .B1(n12016), .B2(n14924), .A(n12015), .ZN(n12017) );
  OAI211_X1 U14504 ( .C1(n12020), .C2(n12019), .A(n12018), .B(n12017), .ZN(
        P1_U3287) );
  NAND2_X1 U14505 ( .A1(n12022), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n12023) );
  INV_X1 U14506 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n12027) );
  NAND2_X1 U14507 ( .A1(n12027), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n12408) );
  INV_X1 U14508 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n12028) );
  NAND2_X1 U14509 ( .A1(n12028), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n12029) );
  AND2_X1 U14510 ( .A1(n12408), .A2(n12029), .ZN(n12406) );
  INV_X1 U14511 ( .A(n12406), .ZN(n12030) );
  XNOR2_X1 U14512 ( .A(n12407), .B(n12030), .ZN(n12031) );
  NAND2_X1 U14513 ( .A1(n12405), .A2(n12404), .ZN(n12033) );
  XNOR2_X1 U14514 ( .A(n12033), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U14515 ( .B1(n12035), .B2(n12036), .A(n12034), .ZN(n15296) );
  INV_X1 U14516 ( .A(n15296), .ZN(n12050) );
  XNOR2_X1 U14517 ( .A(n12037), .B(n12036), .ZN(n12038) );
  NOR2_X1 U14518 ( .A1(n12038), .A2(n15007), .ZN(n15294) );
  INV_X1 U14519 ( .A(n12039), .ZN(n15291) );
  NOR2_X1 U14520 ( .A1(n15294), .A2(n15291), .ZN(n12040) );
  MUX2_X1 U14521 ( .A(n12041), .B(n12040), .S(n14940), .Z(n12049) );
  INV_X1 U14522 ( .A(n12042), .ZN(n12043) );
  AOI211_X1 U14523 ( .C1(n12045), .C2(n12044), .A(n14906), .B(n12043), .ZN(
        n15293) );
  OAI22_X1 U14524 ( .A1(n14937), .A2(n6760), .B1(n14946), .B2(n12046), .ZN(
        n12047) );
  AOI21_X1 U14525 ( .B1(n15293), .B2(n14924), .A(n12047), .ZN(n12048) );
  OAI211_X1 U14526 ( .C1(n14969), .C2(n12050), .A(n12049), .B(n12048), .ZN(
        P1_U3288) );
  INV_X1 U14527 ( .A(n12051), .ZN(n12063) );
  NOR2_X1 U14528 ( .A1(n12053), .A2(n12052), .ZN(n12054) );
  MUX2_X1 U14529 ( .A(n12055), .B(n12054), .S(n14940), .Z(n12062) );
  INV_X1 U14530 ( .A(n12056), .ZN(n12060) );
  INV_X1 U14531 ( .A(n12183), .ZN(n12058) );
  OAI22_X1 U14532 ( .A1(n12058), .A2(n14937), .B1(n14946), .B2(n12057), .ZN(
        n12059) );
  AOI21_X1 U14533 ( .B1(n12060), .B2(n14924), .A(n12059), .ZN(n12061) );
  OAI211_X1 U14534 ( .C1(n14969), .C2(n12063), .A(n12062), .B(n12061), .ZN(
        P1_U3284) );
  INV_X1 U14535 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12064) );
  XNOR2_X1 U14536 ( .A(n13140), .B(n12064), .ZN(n13131) );
  XOR2_X1 U14537 ( .A(n13131), .B(n13132), .Z(n12083) );
  MUX2_X1 U14538 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13703), .Z(n13135) );
  XNOR2_X1 U14539 ( .A(n13135), .B(n13140), .ZN(n13136) );
  XNOR2_X1 U14540 ( .A(n13137), .B(n13136), .ZN(n12081) );
  NAND2_X1 U14541 ( .A1(n15503), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n12071) );
  OAI211_X1 U14542 ( .C1(n13314), .C2(n13140), .A(n12072), .B(n12071), .ZN(
        n12080) );
  INV_X1 U14543 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n13142) );
  XNOR2_X1 U14544 ( .A(n13140), .B(n13142), .ZN(n12074) );
  INV_X1 U14545 ( .A(n12074), .ZN(n12076) );
  NAND3_X1 U14546 ( .A1(n12077), .A2(n12076), .A3(n12075), .ZN(n12078) );
  AOI21_X1 U14547 ( .B1(n13141), .B2(n12078), .A(n13164), .ZN(n12079) );
  AOI211_X1 U14548 ( .C1(n13329), .C2(n12081), .A(n12080), .B(n12079), .ZN(
        n12082) );
  OAI21_X1 U14549 ( .B1(n12083), .B2(n13283), .A(n12082), .ZN(P3_U3192) );
  AOI22_X1 U14550 ( .A1(n13519), .A2(n12085), .B1(n15544), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n12088) );
  MUX2_X1 U14551 ( .A(n12086), .B(n12339), .S(n15524), .Z(n12087) );
  NAND2_X1 U14552 ( .A1(n12088), .A2(n12087), .ZN(P3_U3233) );
  OAI21_X1 U14553 ( .B1(n12090), .B2(n12095), .A(n12089), .ZN(n12091) );
  INV_X1 U14554 ( .A(n12091), .ZN(n15111) );
  INV_X1 U14555 ( .A(n12092), .ZN(n12093) );
  AOI211_X1 U14556 ( .C1(n12095), .C2(n12094), .A(n15007), .B(n12093), .ZN(
        n15109) );
  NOR2_X1 U14557 ( .A1(n15109), .A2(n15106), .ZN(n12096) );
  MUX2_X1 U14558 ( .A(n12097), .B(n12096), .S(n14940), .Z(n12106) );
  INV_X1 U14559 ( .A(n12112), .ZN(n12100) );
  INV_X1 U14560 ( .A(n12098), .ZN(n12099) );
  AOI211_X1 U14561 ( .C1(n12101), .C2(n12100), .A(n14906), .B(n12099), .ZN(
        n15107) );
  OAI22_X1 U14562 ( .A1(n14937), .A2(n12103), .B1(n12102), .B2(n14946), .ZN(
        n12104) );
  AOI21_X1 U14563 ( .B1(n15107), .B2(n14924), .A(n12104), .ZN(n12105) );
  OAI211_X1 U14564 ( .C1(n15111), .C2(n14969), .A(n12106), .B(n12105), .ZN(
        P1_U3285) );
  OAI21_X1 U14565 ( .B1(n12109), .B2(n12108), .A(n12107), .ZN(n12110) );
  INV_X1 U14566 ( .A(n12110), .ZN(n15305) );
  OAI21_X1 U14567 ( .B1(n12111), .B2(n12115), .A(n14949), .ZN(n12113) );
  NOR2_X1 U14568 ( .A1(n12113), .A2(n12112), .ZN(n15299) );
  MUX2_X1 U14569 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n15300), .S(n14940), .Z(
        n12117) );
  OAI22_X1 U14570 ( .A1(n14937), .A2(n12115), .B1(n14946), .B2(n12114), .ZN(
        n12116) );
  AOI211_X1 U14571 ( .C1(n15299), .C2(n14924), .A(n12117), .B(n12116), .ZN(
        n12121) );
  XNOR2_X1 U14572 ( .A(n12118), .B(n12119), .ZN(n15307) );
  NAND2_X1 U14573 ( .A1(n15307), .A2(n14864), .ZN(n12120) );
  OAI211_X1 U14574 ( .C1(n15305), .C2(n14969), .A(n12121), .B(n12120), .ZN(
        P1_U3286) );
  AOI21_X1 U14575 ( .B1(n12124), .B2(n12123), .A(n12122), .ZN(n12129) );
  AOI22_X1 U14576 ( .A1(n13107), .A2(n13128), .B1(n13100), .B2(n13126), .ZN(
        n12126) );
  OAI211_X1 U14577 ( .C1(n13103), .C2(n15566), .A(n12126), .B(n12125), .ZN(
        n12127) );
  AOI21_X1 U14578 ( .B1(n12310), .B2(n13111), .A(n12127), .ZN(n12128) );
  OAI21_X1 U14579 ( .B1(n12129), .B2(n13115), .A(n12128), .ZN(P3_U3170) );
  INV_X1 U14580 ( .A(n12130), .ZN(n12137) );
  INV_X1 U14581 ( .A(n12131), .ZN(n12132) );
  MUX2_X1 U14582 ( .A(n12133), .B(n12132), .S(n15524), .Z(n12135) );
  AOI22_X1 U14583 ( .A1(n13519), .A2(n12480), .B1(n15544), .B2(n12485), .ZN(
        n12134) );
  OAI211_X1 U14584 ( .C1(n12137), .C2(n12136), .A(n12135), .B(n12134), .ZN(
        P3_U3225) );
  INV_X1 U14585 ( .A(n12138), .ZN(n12142) );
  OAI222_X1 U14586 ( .A1(n15149), .A2(n12140), .B1(n15141), .B2(n12142), .C1(
        n12139), .C2(P1_U3086), .ZN(P1_U3331) );
  OAI222_X1 U14587 ( .A1(n12742), .A2(n12143), .B1(n14447), .B2(n12142), .C1(
        n12141), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U14588 ( .A(n12213), .ZN(n12144) );
  AOI21_X1 U14589 ( .B1(n12146), .B2(n12145), .A(n12144), .ZN(n12372) );
  INV_X1 U14590 ( .A(n12222), .ZN(n12147) );
  AOI211_X1 U14591 ( .C1(n12159), .C2(n6614), .A(n14363), .B(n12147), .ZN(
        n12377) );
  INV_X1 U14592 ( .A(n12148), .ZN(n12149) );
  AOI211_X1 U14593 ( .C1(n12151), .C2(n12150), .A(n14217), .B(n12149), .ZN(
        n12155) );
  NAND2_X1 U14594 ( .A1(n13944), .A2(n14082), .ZN(n12154) );
  OR2_X1 U14595 ( .A1(n12152), .A2(n14197), .ZN(n12153) );
  NAND2_X1 U14596 ( .A1(n12154), .A2(n12153), .ZN(n13772) );
  OR2_X1 U14597 ( .A1(n12155), .A2(n13772), .ZN(n12373) );
  AOI211_X1 U14598 ( .C1(n12372), .C2(n14366), .A(n12377), .B(n12373), .ZN(
        n12161) );
  OAI22_X1 U14599 ( .A1(n14362), .A2(n10439), .B1(n15502), .B2(n12156), .ZN(
        n12157) );
  INV_X1 U14600 ( .A(n12157), .ZN(n12158) );
  OAI21_X1 U14601 ( .B1(n12161), .B2(n15500), .A(n12158), .ZN(P2_U3507) );
  AOI22_X1 U14602 ( .A1(n14434), .A2(n12159), .B1(P2_REG0_REG_8__SCAN_IN), 
        .B2(n15492), .ZN(n12160) );
  OAI21_X1 U14603 ( .B1(n12161), .B2(n15492), .A(n12160), .ZN(P2_U3454) );
  XNOR2_X1 U14604 ( .A(n12162), .B(n12167), .ZN(n15573) );
  OR2_X1 U14605 ( .A1(n15567), .A2(n12163), .ZN(n15572) );
  INV_X1 U14606 ( .A(n12164), .ZN(n12165) );
  OAI22_X1 U14607 ( .A1(n12166), .A2(n15572), .B1(n12165), .B2(n15509), .ZN(
        n12175) );
  NAND2_X1 U14608 ( .A1(n15573), .A2(n15528), .ZN(n12173) );
  AOI22_X1 U14609 ( .A1(n15537), .A2(n13125), .B1(n15535), .B2(n13127), .ZN(
        n12172) );
  NAND2_X1 U14610 ( .A1(n11705), .A2(n12167), .ZN(n12168) );
  NAND2_X1 U14611 ( .A1(n12169), .A2(n12168), .ZN(n12170) );
  NAND2_X1 U14612 ( .A1(n12170), .A2(n15532), .ZN(n12171) );
  NAND3_X1 U14613 ( .A1(n12173), .A2(n12172), .A3(n12171), .ZN(n15576) );
  MUX2_X1 U14614 ( .A(n15576), .B(P3_REG2_REG_5__SCAN_IN), .S(n15549), .Z(
        n12174) );
  AOI211_X1 U14615 ( .C1(n15573), .C2(n15545), .A(n12175), .B(n12174), .ZN(
        n12176) );
  INV_X1 U14616 ( .A(n12176), .ZN(P3_U3228) );
  OAI21_X1 U14617 ( .B1(n12178), .B2(n12187), .A(n12297), .ZN(n12319) );
  AOI21_X1 U14618 ( .B1(n6795), .B2(n12295), .A(n14893), .ZN(n12181) );
  NAND2_X1 U14619 ( .A1(n14960), .A2(n14614), .ZN(n12270) );
  INV_X1 U14620 ( .A(n12270), .ZN(n12180) );
  AOI21_X1 U14621 ( .B1(n12181), .B2(n12291), .A(n12180), .ZN(n12315) );
  NAND2_X1 U14622 ( .A1(n12183), .A2(n12182), .ZN(n12184) );
  INV_X1 U14623 ( .A(n12187), .ZN(n12186) );
  NAND2_X1 U14624 ( .A1(n12188), .A2(n12187), .ZN(n12316) );
  NAND3_X1 U14625 ( .A1(n12285), .A2(n14864), .A3(n12316), .ZN(n12193) );
  NOR2_X1 U14626 ( .A1(n14940), .A2(n12189), .ZN(n12191) );
  NAND2_X1 U14627 ( .A1(n14962), .A2(n14616), .ZN(n12314) );
  OAI22_X1 U14628 ( .A1(n14920), .A2(n12314), .B1(n12271), .B2(n14946), .ZN(
        n12190) );
  AOI211_X1 U14629 ( .C1(n14956), .C2(n12295), .A(n12191), .B(n12190), .ZN(
        n12192) );
  OAI211_X1 U14630 ( .C1(n12315), .C2(n14953), .A(n12193), .B(n12192), .ZN(
        n12194) );
  AOI21_X1 U14631 ( .B1(n14841), .B2(n12319), .A(n12194), .ZN(n12195) );
  INV_X1 U14632 ( .A(n12195), .ZN(P1_U3283) );
  INV_X1 U14633 ( .A(n12196), .ZN(n12198) );
  OAI222_X1 U14634 ( .A1(n12199), .A2(P3_U3151), .B1(n13707), .B2(n12198), 
        .C1(n12197), .C2(n13705), .ZN(P3_U3271) );
  INV_X1 U14635 ( .A(n11758), .ZN(n12201) );
  NAND2_X1 U14636 ( .A1(n12201), .A2(n12200), .ZN(n12325) );
  XNOR2_X1 U14637 ( .A(n12202), .B(n13125), .ZN(n12326) );
  NOR2_X1 U14638 ( .A1(n12325), .A2(n12326), .ZN(n12324) );
  NOR2_X1 U14639 ( .A1(n12324), .A2(n12203), .ZN(n12477) );
  XNOR2_X1 U14640 ( .A(n12477), .B(n12204), .ZN(n12211) );
  AOI22_X1 U14641 ( .A1(n13107), .A2(n13125), .B1(n13100), .B2(n12205), .ZN(
        n12207) );
  OAI211_X1 U14642 ( .C1(n13103), .C2(n12208), .A(n12207), .B(n12206), .ZN(
        n12209) );
  AOI21_X1 U14643 ( .B1(n12363), .B2(n13111), .A(n12209), .ZN(n12210) );
  OAI21_X1 U14644 ( .B1(n12211), .B2(n13115), .A(n12210), .ZN(P3_U3153) );
  XNOR2_X1 U14645 ( .A(n12542), .B(n12215), .ZN(n12278) );
  INV_X1 U14646 ( .A(n12278), .ZN(n12226) );
  INV_X1 U14647 ( .A(n12215), .ZN(n12541) );
  NAND2_X1 U14648 ( .A1(n12214), .A2(n12541), .ZN(n12419) );
  OAI211_X1 U14649 ( .C1(n12214), .C2(n12541), .A(n12419), .B(n14252), .ZN(
        n12219) );
  NAND2_X1 U14650 ( .A1(n13943), .A2(n14082), .ZN(n12218) );
  OR2_X1 U14651 ( .A1(n12216), .A2(n14197), .ZN(n12217) );
  AND2_X1 U14652 ( .A1(n12218), .A2(n12217), .ZN(n13847) );
  NAND2_X1 U14653 ( .A1(n12219), .A2(n13847), .ZN(n12276) );
  INV_X1 U14654 ( .A(n12276), .ZN(n12220) );
  MUX2_X1 U14655 ( .A(n12221), .B(n12220), .S(n14242), .Z(n12225) );
  AOI211_X1 U14656 ( .C1(n13851), .C2(n12222), .A(n14363), .B(n12552), .ZN(
        n12277) );
  INV_X1 U14657 ( .A(n13851), .ZN(n12281) );
  OAI22_X1 U14658 ( .A1(n14226), .A2(n12281), .B1(n14239), .B2(n13849), .ZN(
        n12223) );
  AOI21_X1 U14659 ( .B1(n12277), .B2(n14273), .A(n12223), .ZN(n12224) );
  OAI211_X1 U14660 ( .C1(n14248), .C2(n12226), .A(n12225), .B(n12224), .ZN(
        P2_U3256) );
  XNOR2_X1 U14661 ( .A(n12228), .B(n7637), .ZN(n12343) );
  NOR2_X1 U14662 ( .A1(n12346), .A2(n15567), .ZN(n12234) );
  NAND2_X1 U14663 ( .A1(n12230), .A2(n12229), .ZN(n12231) );
  XNOR2_X1 U14664 ( .A(n12231), .B(n7637), .ZN(n12232) );
  OAI222_X1 U14665 ( .A1(n15513), .A2(n13073), .B1(n15516), .B2(n12233), .C1(
        n12232), .C2(n13522), .ZN(n12348) );
  AOI211_X1 U14666 ( .C1(n15569), .C2(n12343), .A(n12234), .B(n12348), .ZN(
        n12237) );
  NAND2_X1 U14667 ( .A1(n15593), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n12235) );
  OAI21_X1 U14668 ( .B1(n12237), .B2(n15593), .A(n12235), .ZN(P3_U3469) );
  NAND2_X1 U14669 ( .A1(n15583), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n12236) );
  OAI21_X1 U14670 ( .B1(n12237), .B2(n15583), .A(n12236), .ZN(P3_U3420) );
  NAND2_X1 U14671 ( .A1(n12238), .A2(n12443), .ZN(n12239) );
  MUX2_X1 U14672 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n12590), .S(n15424), .Z(
        n15426) );
  NAND2_X1 U14673 ( .A1(n15424), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12241) );
  NAND2_X1 U14674 ( .A1(n15425), .A2(n12241), .ZN(n12243) );
  NAND2_X1 U14675 ( .A1(n15438), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n12245) );
  NAND2_X1 U14676 ( .A1(n12243), .A2(n15437), .ZN(n12244) );
  NAND2_X1 U14677 ( .A1(n12245), .A2(n12244), .ZN(n13984) );
  XNOR2_X1 U14678 ( .A(n13984), .B(n7246), .ZN(n13983) );
  XNOR2_X1 U14679 ( .A(n13983), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n12257) );
  OAI21_X1 U14680 ( .B1(n12247), .B2(P2_REG1_REG_12__SCAN_IN), .A(n12246), 
        .ZN(n15420) );
  XNOR2_X1 U14681 ( .A(n15424), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n15421) );
  NOR2_X1 U14682 ( .A1(n15420), .A2(n15421), .ZN(n15419) );
  XNOR2_X1 U14683 ( .A(n15437), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15433) );
  INV_X1 U14684 ( .A(n12249), .ZN(n12251) );
  NOR2_X1 U14685 ( .A1(n12249), .A2(n12248), .ZN(n13991) );
  INV_X1 U14686 ( .A(n13991), .ZN(n12250) );
  OAI211_X1 U14687 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n12251), .A(n12250), 
        .B(n15402), .ZN(n12256) );
  NOR2_X1 U14688 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12252), .ZN(n12254) );
  INV_X1 U14689 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15182) );
  NOR2_X1 U14690 ( .A1(n15457), .A2(n15182), .ZN(n12253) );
  AOI211_X1 U14691 ( .C1(n15450), .C2(n13993), .A(n12254), .B(n12253), .ZN(
        n12255) );
  OAI211_X1 U14692 ( .C1(n12257), .C2(n15411), .A(n12256), .B(n12255), .ZN(
        P2_U3229) );
  INV_X1 U14693 ( .A(n12258), .ZN(n12259) );
  NAND2_X1 U14694 ( .A1(n12260), .A2(n12259), .ZN(n12261) );
  NAND2_X1 U14695 ( .A1(n12295), .A2(n12871), .ZN(n12264) );
  NAND2_X1 U14696 ( .A1(n12872), .A2(n14615), .ZN(n12263) );
  NAND2_X1 U14697 ( .A1(n12264), .A2(n12263), .ZN(n12265) );
  XNOR2_X1 U14698 ( .A(n12265), .B(n12866), .ZN(n12527) );
  NOR2_X1 U14699 ( .A1(n12855), .A2(n12289), .ZN(n12266) );
  AOI21_X1 U14700 ( .B1(n12295), .B2(n11176), .A(n12266), .ZN(n12525) );
  XNOR2_X1 U14701 ( .A(n12527), .B(n12525), .ZN(n12267) );
  OAI211_X1 U14702 ( .C1(n12268), .C2(n12267), .A(n12529), .B(n14589), .ZN(
        n12275) );
  OAI21_X1 U14703 ( .B1(n14595), .B2(n12270), .A(n12269), .ZN(n12273) );
  NOR2_X1 U14704 ( .A1(n15246), .A2(n12271), .ZN(n12272) );
  AOI211_X1 U14705 ( .C1(n14560), .C2(n14616), .A(n12273), .B(n12272), .ZN(
        n12274) );
  OAI211_X1 U14706 ( .C1(n12179), .C2(n14600), .A(n12275), .B(n12274), .ZN(
        P1_U3217) );
  AOI211_X1 U14707 ( .C1(n14366), .C2(n12278), .A(n12277), .B(n12276), .ZN(
        n12284) );
  AOI22_X1 U14708 ( .A1(n14434), .A2(n13851), .B1(P2_REG0_REG_9__SCAN_IN), 
        .B2(n15492), .ZN(n12279) );
  OAI21_X1 U14709 ( .B1(n12284), .B2(n15492), .A(n12279), .ZN(P2_U3457) );
  OAI22_X1 U14710 ( .A1(n14362), .A2(n12281), .B1(n15502), .B2(n12280), .ZN(
        n12282) );
  INV_X1 U14711 ( .A(n12282), .ZN(n12283) );
  OAI21_X1 U14712 ( .B1(n12284), .B2(n15500), .A(n12283), .ZN(P2_U3508) );
  OR2_X1 U14713 ( .A1(n12295), .A2(n12289), .ZN(n12287) );
  NAND3_X1 U14714 ( .A1(n12285), .A2(n12298), .A3(n12287), .ZN(n12288) );
  AND3_X1 U14715 ( .A1(n12505), .A2(n15308), .A3(n12288), .ZN(n12290) );
  OAI22_X1 U14716 ( .A1(n12770), .A2(n14916), .B1(n12289), .B2(n14918), .ZN(
        n12534) );
  NOR2_X1 U14717 ( .A1(n12290), .A2(n12534), .ZN(n15104) );
  AOI211_X1 U14718 ( .C1(n12532), .C2(n12291), .A(n14893), .B(n12514), .ZN(
        n15102) );
  NOR2_X1 U14719 ( .A1(n6793), .A2(n14937), .ZN(n12294) );
  OAI22_X1 U14720 ( .A1(n14940), .A2(n12292), .B1(n12536), .B2(n14946), .ZN(
        n12293) );
  AOI211_X1 U14721 ( .C1(n15102), .C2(n14924), .A(n12294), .B(n12293), .ZN(
        n12301) );
  OR2_X1 U14722 ( .A1(n12295), .A2(n14615), .ZN(n12296) );
  OAI21_X1 U14723 ( .B1(n12299), .B2(n12298), .A(n6644), .ZN(n15100) );
  NAND2_X1 U14724 ( .A1(n15100), .A2(n14841), .ZN(n12300) );
  OAI211_X1 U14725 ( .C1(n15104), .C2(n14920), .A(n12301), .B(n12300), .ZN(
        P1_U3282) );
  NAND2_X1 U14726 ( .A1(n15521), .A2(n12302), .ZN(n12303) );
  XNOR2_X1 U14727 ( .A(n12305), .B(n12304), .ZN(n15564) );
  INV_X1 U14728 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n12309) );
  XNOR2_X1 U14729 ( .A(n12307), .B(n12306), .ZN(n12308) );
  AOI222_X1 U14730 ( .A1(n15532), .A2(n12308), .B1(n13126), .B2(n15537), .C1(
        n13128), .C2(n15535), .ZN(n15565) );
  MUX2_X1 U14731 ( .A(n12309), .B(n15565), .S(n15524), .Z(n12313) );
  AOI22_X1 U14732 ( .A1(n13519), .A2(n12311), .B1(n15544), .B2(n12310), .ZN(
        n12312) );
  OAI211_X1 U14733 ( .C1(n13529), .C2(n15564), .A(n12313), .B(n12312), .ZN(
        P3_U3229) );
  OAI211_X1 U14734 ( .C1(n12179), .C2(n15065), .A(n12315), .B(n12314), .ZN(
        n12318) );
  AND3_X1 U14735 ( .A1(n12285), .A2(n15308), .A3(n12316), .ZN(n12317) );
  AOI211_X1 U14736 ( .C1(n15297), .C2(n12319), .A(n12318), .B(n12317), .ZN(
        n12322) );
  NAND2_X1 U14737 ( .A1(n15314), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n12320) );
  OAI21_X1 U14738 ( .B1(n12322), .B2(n15314), .A(n12320), .ZN(P1_U3538) );
  NAND2_X1 U14739 ( .A1(n15309), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n12321) );
  OAI21_X1 U14740 ( .B1(n12322), .B2(n15309), .A(n12321), .ZN(P1_U3489) );
  INV_X1 U14741 ( .A(n12323), .ZN(n12334) );
  AOI211_X1 U14742 ( .C1(n12326), .C2(n12325), .A(n13115), .B(n12324), .ZN(
        n12327) );
  INV_X1 U14743 ( .A(n12327), .ZN(n12333) );
  OAI22_X1 U14744 ( .A1(n12328), .A2(n13098), .B1(n13109), .B2(n12483), .ZN(
        n12329) );
  AOI211_X1 U14745 ( .C1(n13112), .C2(n12331), .A(n12330), .B(n12329), .ZN(
        n12332) );
  OAI211_X1 U14746 ( .C1(n12334), .C2(n13088), .A(n12333), .B(n12332), .ZN(
        P3_U3179) );
  MUX2_X1 U14747 ( .A(n12336), .B(n12335), .S(n15595), .Z(n12337) );
  OAI21_X1 U14748 ( .B1(n12338), .B2(n13597), .A(n12337), .ZN(P3_U3467) );
  INV_X1 U14749 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n12340) );
  MUX2_X1 U14750 ( .A(n12340), .B(n12339), .S(n15595), .Z(n12341) );
  OAI21_X1 U14751 ( .B1(n12342), .B2(n13597), .A(n12341), .ZN(P3_U3459) );
  INV_X1 U14752 ( .A(n12343), .ZN(n12350) );
  AOI22_X1 U14753 ( .A1(n15549), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15544), 
        .B2(n12344), .ZN(n12345) );
  OAI21_X1 U14754 ( .B1(n13534), .B2(n12346), .A(n12345), .ZN(n12347) );
  AOI21_X1 U14755 ( .B1(n12348), .B2(n15524), .A(n12347), .ZN(n12349) );
  OAI21_X1 U14756 ( .B1(n12350), .B2(n13529), .A(n12349), .ZN(P3_U3223) );
  NAND2_X1 U14757 ( .A1(n12351), .A2(n13095), .ZN(n12361) );
  AOI21_X1 U14758 ( .B1(n11558), .B2(n12353), .A(n12352), .ZN(n12360) );
  OAI22_X1 U14759 ( .A1(n12355), .A2(n13109), .B1(n13103), .B2(n12354), .ZN(
        n12358) );
  MUX2_X1 U14760 ( .A(P3_U3151), .B(n13111), .S(n12356), .Z(n12357) );
  AOI211_X1 U14761 ( .C1(n13107), .C2(n15536), .A(n12358), .B(n12357), .ZN(
        n12359) );
  OAI21_X1 U14762 ( .B1(n12361), .B2(n12360), .A(n12359), .ZN(P3_U3158) );
  AOI21_X1 U14763 ( .B1(n15544), .B2(n12363), .A(n12362), .ZN(n12364) );
  MUX2_X1 U14764 ( .A(n12365), .B(n12364), .S(n15524), .Z(n12368) );
  NAND2_X1 U14765 ( .A1(n13519), .A2(n12366), .ZN(n12367) );
  OAI211_X1 U14766 ( .C1(n12417), .C2(n13529), .A(n12368), .B(n12367), .ZN(
        P3_U3226) );
  INV_X1 U14767 ( .A(n12625), .ZN(n12369) );
  MUX2_X1 U14768 ( .A(n7509), .B(n12369), .S(n15524), .Z(n12371) );
  AOI22_X1 U14769 ( .A1(n13519), .A2(n13038), .B1(n15544), .B2(n13037), .ZN(
        n12370) );
  OAI211_X1 U14770 ( .C1(n12628), .C2(n13529), .A(n12371), .B(n12370), .ZN(
        P3_U3224) );
  INV_X1 U14771 ( .A(n12372), .ZN(n12380) );
  INV_X1 U14772 ( .A(n12373), .ZN(n12374) );
  MUX2_X1 U14773 ( .A(n12375), .B(n12374), .S(n14242), .Z(n12379) );
  OAI22_X1 U14774 ( .A1(n14226), .A2(n10439), .B1(n14239), .B2(n13769), .ZN(
        n12376) );
  AOI21_X1 U14775 ( .B1(n12377), .B2(n14273), .A(n12376), .ZN(n12378) );
  OAI211_X1 U14776 ( .C1(n14248), .C2(n12380), .A(n12379), .B(n12378), .ZN(
        P2_U3257) );
  INV_X1 U14777 ( .A(n12381), .ZN(n12385) );
  OAI222_X1 U14778 ( .A1(n12742), .A2(n12383), .B1(n14447), .B2(n12385), .C1(
        n12382), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U14779 ( .A1(n15149), .A2(n12386), .B1(n15141), .B2(n12385), .C1(
        n12384), .C2(P1_U3086), .ZN(P1_U3330) );
  XOR2_X1 U14780 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n12657), .Z(n12390) );
  OAI21_X1 U14781 ( .B1(n12390), .B2(n12389), .A(n12656), .ZN(n12402) );
  NOR2_X1 U14782 ( .A1(n12391), .A2(n15702), .ZN(n12395) );
  INV_X1 U14783 ( .A(n12395), .ZN(n12393) );
  INV_X1 U14784 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n12665) );
  MUX2_X1 U14785 ( .A(n12665), .B(P1_REG2_REG_14__SCAN_IN), .S(n12657), .Z(
        n12392) );
  NAND2_X1 U14786 ( .A1(n12393), .A2(n12392), .ZN(n12396) );
  MUX2_X1 U14787 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n12665), .S(n12657), .Z(
        n12394) );
  OAI21_X1 U14788 ( .B1(n12397), .B2(n12395), .A(n12394), .ZN(n12663) );
  OAI211_X1 U14789 ( .C1(n12397), .C2(n12396), .A(n12663), .B(n15267), .ZN(
        n12400) );
  NAND2_X1 U14790 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14465)
         );
  INV_X1 U14791 ( .A(n14465), .ZN(n12398) );
  AOI21_X1 U14792 ( .B1(n15255), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n12398), 
        .ZN(n12399) );
  OAI211_X1 U14793 ( .C1(n14686), .C2(n12664), .A(n12400), .B(n12399), .ZN(
        n12401) );
  AOI21_X1 U14794 ( .B1(n12402), .B2(n15266), .A(n12401), .ZN(n12403) );
  INV_X1 U14795 ( .A(n12403), .ZN(P1_U3257) );
  INV_X1 U14796 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15607) );
  NAND2_X1 U14797 ( .A1(n12407), .A2(n12406), .ZN(n12409) );
  NAND2_X1 U14798 ( .A1(n12409), .A2(n12408), .ZN(n12612) );
  INV_X1 U14799 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n13160) );
  XNOR2_X1 U14800 ( .A(n13160), .B(P1_ADDR_REG_12__SCAN_IN), .ZN(n12611) );
  INV_X1 U14801 ( .A(n12611), .ZN(n12410) );
  XNOR2_X1 U14802 ( .A(n12612), .B(n12410), .ZN(n12411) );
  NAND2_X1 U14803 ( .A1(n12412), .A2(n12411), .ZN(n12609) );
  NAND2_X1 U14804 ( .A1(n12608), .A2(n12609), .ZN(n12413) );
  XNOR2_X1 U14805 ( .A(n12413), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  MUX2_X1 U14806 ( .A(n12415), .B(n12414), .S(n15595), .Z(n12416) );
  OAI21_X1 U14807 ( .B1(n13592), .B2(n12417), .A(n12416), .ZN(P3_U3466) );
  AND2_X1 U14808 ( .A1(n12419), .A2(n12418), .ZN(n12545) );
  NOR2_X1 U14809 ( .A1(n12545), .A2(n12546), .ZN(n12544) );
  AOI21_X1 U14810 ( .B1(n12555), .B2(n13943), .A(n12544), .ZN(n12421) );
  OAI21_X1 U14811 ( .B1(n12421), .B2(n12430), .A(n12420), .ZN(n12425) );
  NAND2_X1 U14812 ( .A1(n13941), .A2(n14082), .ZN(n12424) );
  OR2_X1 U14813 ( .A1(n12422), .A2(n14197), .ZN(n12423) );
  NAND2_X1 U14814 ( .A1(n12424), .A2(n12423), .ZN(n13887) );
  AOI21_X1 U14815 ( .B1(n12425), .B2(n14252), .A(n13887), .ZN(n14384) );
  INV_X1 U14816 ( .A(n12440), .ZN(n12426) );
  AOI211_X1 U14817 ( .C1(n14382), .C2(n12554), .A(n14363), .B(n12426), .ZN(
        n14381) );
  INV_X1 U14818 ( .A(n13890), .ZN(n12427) );
  AOI22_X1 U14819 ( .A1(n14264), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n14276), 
        .B2(n12427), .ZN(n12428) );
  OAI21_X1 U14820 ( .B1(n7443), .B2(n14226), .A(n12428), .ZN(n12432) );
  XOR2_X1 U14821 ( .A(n12429), .B(n12430), .Z(n14385) );
  NOR2_X1 U14822 ( .A1(n14385), .A2(n14248), .ZN(n12431) );
  AOI211_X1 U14823 ( .C1(n14381), .C2(n14273), .A(n12432), .B(n12431), .ZN(
        n12433) );
  OAI21_X1 U14824 ( .B1(n14384), .B2(n14264), .A(n12433), .ZN(P2_U3254) );
  XNOR2_X1 U14825 ( .A(n12434), .B(n12436), .ZN(n12571) );
  INV_X1 U14826 ( .A(n12571), .ZN(n12448) );
  NAND2_X1 U14827 ( .A1(n12437), .A2(n12436), .ZN(n12438) );
  NAND3_X1 U14828 ( .A1(n12435), .A2(n14252), .A3(n12438), .ZN(n12439) );
  AOI22_X1 U14829 ( .A1(n13940), .A2(n14082), .B1(n14097), .B2(n13942), .ZN(
        n13788) );
  NAND2_X1 U14830 ( .A1(n12439), .A2(n13788), .ZN(n12574) );
  NAND2_X1 U14831 ( .A1(n12574), .A2(n14242), .ZN(n12447) );
  NAND2_X1 U14832 ( .A1(n12440), .A2(n13793), .ZN(n12441) );
  NAND2_X1 U14833 ( .A1(n12441), .A2(n14262), .ZN(n12442) );
  NOR2_X1 U14834 ( .A1(n12587), .A2(n12442), .ZN(n12572) );
  OAI22_X1 U14835 ( .A1(n14242), .A2(n12443), .B1(n13790), .B2(n14239), .ZN(
        n12445) );
  NOR2_X1 U14836 ( .A1(n7444), .A2(n14226), .ZN(n12444) );
  AOI211_X1 U14837 ( .C1(n12572), .C2(n14273), .A(n12445), .B(n12444), .ZN(
        n12446) );
  OAI211_X1 U14838 ( .C1(n12448), .C2(n14248), .A(n12447), .B(n12446), .ZN(
        P2_U3253) );
  INV_X1 U14839 ( .A(n12449), .ZN(n12450) );
  OAI222_X1 U14840 ( .A1(P3_U3151), .A2(n12452), .B1(n13705), .B2(n12451), 
        .C1(n13707), .C2(n12450), .ZN(P3_U3270) );
  OR2_X1 U14841 ( .A1(n12532), .A2(n14614), .ZN(n12453) );
  OAI21_X1 U14842 ( .B1(n12455), .B2(n12457), .A(n12502), .ZN(n12456) );
  INV_X1 U14843 ( .A(n12456), .ZN(n15099) );
  INV_X1 U14844 ( .A(n14614), .ZN(n12523) );
  OR2_X1 U14845 ( .A1(n12532), .A2(n12523), .ZN(n12503) );
  AOI21_X1 U14846 ( .B1(n12505), .B2(n12503), .A(n12457), .ZN(n12510) );
  NAND3_X1 U14847 ( .A1(n12505), .A2(n12457), .A3(n12503), .ZN(n12458) );
  NAND2_X1 U14848 ( .A1(n12458), .A2(n15308), .ZN(n12459) );
  AOI22_X1 U14849 ( .A1(n14963), .A2(n14960), .B1(n14962), .B2(n14614), .ZN(
        n14498) );
  OAI21_X1 U14850 ( .B1(n12510), .B2(n12459), .A(n14498), .ZN(n15095) );
  XNOR2_X1 U14851 ( .A(n12514), .B(n15097), .ZN(n12460) );
  AND2_X1 U14852 ( .A1(n12460), .A2(n14949), .ZN(n15096) );
  NAND2_X1 U14853 ( .A1(n15096), .A2(n14924), .ZN(n12464) );
  OAI22_X1 U14854 ( .A1(n14940), .A2(n12461), .B1(n14496), .B2(n14946), .ZN(
        n12462) );
  AOI21_X1 U14855 ( .B1(n15097), .B2(n14956), .A(n12462), .ZN(n12463) );
  NAND2_X1 U14856 ( .A1(n12464), .A2(n12463), .ZN(n12465) );
  AOI21_X1 U14857 ( .B1(n15095), .B2(n14940), .A(n12465), .ZN(n12466) );
  OAI21_X1 U14858 ( .B1(n15099), .B2(n14969), .A(n12466), .ZN(P1_U3281) );
  XOR2_X1 U14859 ( .A(n12467), .B(n12468), .Z(n12632) );
  AOI22_X1 U14860 ( .A1(n13519), .A2(n12988), .B1(n15544), .B2(n12987), .ZN(
        n12475) );
  INV_X1 U14861 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12473) );
  AOI21_X1 U14862 ( .B1(n12469), .B2(n12468), .A(n13522), .ZN(n12472) );
  OAI22_X1 U14863 ( .A1(n15516), .A2(n13073), .B1(n12948), .B2(n15513), .ZN(
        n12470) );
  AOI21_X1 U14864 ( .B1(n12472), .B2(n12471), .A(n12470), .ZN(n12629) );
  MUX2_X1 U14865 ( .A(n12473), .B(n12629), .S(n15524), .Z(n12474) );
  OAI211_X1 U14866 ( .C1(n12632), .C2(n13529), .A(n12475), .B(n12474), .ZN(
        P3_U3221) );
  MUX2_X1 U14867 ( .A(n12483), .B(n12477), .S(n12476), .Z(n12479) );
  XNOR2_X1 U14868 ( .A(n12479), .B(n12478), .ZN(n12487) );
  AOI22_X1 U14869 ( .A1(n13100), .A2(n13123), .B1(n13112), .B2(n12480), .ZN(
        n12482) );
  OAI211_X1 U14870 ( .C1(n12483), .C2(n13098), .A(n12482), .B(n12481), .ZN(
        n12484) );
  AOI21_X1 U14871 ( .B1(n12485), .B2(n13045), .A(n12484), .ZN(n12486) );
  OAI21_X1 U14872 ( .B1(n12487), .B2(n13115), .A(n12486), .ZN(P3_U3161) );
  XNOR2_X1 U14873 ( .A(n12488), .B(n12491), .ZN(n12489) );
  AOI222_X1 U14874 ( .A1(n15532), .A2(n12489), .B1(n10479), .B2(n15537), .C1(
        n13122), .C2(n15535), .ZN(n13599) );
  OAI21_X1 U14875 ( .B1(n12492), .B2(n12491), .A(n12490), .ZN(n13598) );
  INV_X1 U14876 ( .A(n13529), .ZN(n13543) );
  NAND2_X1 U14877 ( .A1(n13598), .A2(n13543), .ZN(n12497) );
  INV_X1 U14878 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n13145) );
  INV_X1 U14879 ( .A(n13078), .ZN(n12493) );
  OAI22_X1 U14880 ( .A1(n15524), .A2(n13145), .B1(n12493), .B2(n15509), .ZN(
        n12494) );
  AOI21_X1 U14881 ( .B1(n13519), .B2(n12495), .A(n12494), .ZN(n12496) );
  OAI211_X1 U14882 ( .C1(n15549), .C2(n13599), .A(n12497), .B(n12496), .ZN(
        P3_U3222) );
  INV_X1 U14883 ( .A(n12629), .ZN(n12498) );
  MUX2_X1 U14884 ( .A(P3_REG0_REG_12__SCAN_IN), .B(n12498), .S(n15585), .Z(
        n12499) );
  AOI21_X1 U14885 ( .B1(n13670), .B2(n12988), .A(n12499), .ZN(n12500) );
  OAI21_X1 U14886 ( .B1(n12632), .B2(n13673), .A(n12500), .ZN(P3_U3426) );
  OR2_X1 U14887 ( .A1(n15097), .A2(n14613), .ZN(n12501) );
  XNOR2_X1 U14888 ( .A(n12709), .B(n12507), .ZN(n15094) );
  OR2_X1 U14889 ( .A1(n15097), .A2(n12770), .ZN(n12504) );
  NAND2_X1 U14890 ( .A1(n12708), .A2(n12504), .ZN(n12509) );
  NAND2_X1 U14891 ( .A1(n15097), .A2(n12770), .ZN(n12506) );
  AND2_X1 U14892 ( .A1(n12507), .A2(n12506), .ZN(n12508) );
  OAI211_X1 U14893 ( .C1(n12510), .C2(n12509), .A(n15308), .B(n12686), .ZN(
        n12512) );
  AOI22_X1 U14894 ( .A1(n14612), .A2(n14960), .B1(n14962), .B2(n14613), .ZN(
        n12511) );
  NAND2_X1 U14895 ( .A1(n12512), .A2(n12511), .ZN(n15090) );
  NOR2_X1 U14896 ( .A1(n14946), .A2(n14557), .ZN(n12513) );
  OAI21_X1 U14897 ( .B1(n15090), .B2(n12513), .A(n14940), .ZN(n12519) );
  NAND2_X1 U14898 ( .A1(n12514), .A2(n14503), .ZN(n12515) );
  AOI21_X1 U14899 ( .B1(n12515), .B2(n15092), .A(n14893), .ZN(n12516) );
  AND2_X1 U14900 ( .A1(n12516), .A2(n14948), .ZN(n15091) );
  OAI22_X1 U14901 ( .A1(n14563), .A2(n14937), .B1(n14940), .B2(n15702), .ZN(
        n12517) );
  AOI21_X1 U14902 ( .B1(n15091), .B2(n14924), .A(n12517), .ZN(n12518) );
  OAI211_X1 U14903 ( .C1(n15094), .C2(n14969), .A(n12519), .B(n12518), .ZN(
        P1_U3280) );
  NAND2_X1 U14904 ( .A1(n12532), .A2(n12871), .ZN(n12521) );
  NAND2_X1 U14905 ( .A1(n12872), .A2(n14614), .ZN(n12520) );
  NAND2_X1 U14906 ( .A1(n12521), .A2(n12520), .ZN(n12522) );
  XNOR2_X1 U14907 ( .A(n12522), .B(n12875), .ZN(n12765) );
  NOR2_X1 U14908 ( .A1(n12855), .A2(n12523), .ZN(n12524) );
  AOI21_X1 U14909 ( .B1(n12532), .B2(n11176), .A(n12524), .ZN(n12764) );
  XNOR2_X1 U14910 ( .A(n12765), .B(n12764), .ZN(n12531) );
  INV_X1 U14911 ( .A(n12525), .ZN(n12526) );
  NAND2_X1 U14912 ( .A1(n12527), .A2(n12526), .ZN(n12528) );
  AOI21_X1 U14913 ( .B1(n12531), .B2(n12530), .A(n12766), .ZN(n12539) );
  AND2_X1 U14914 ( .A1(n12532), .A2(n15302), .ZN(n15101) );
  AOI21_X1 U14915 ( .B1(n15241), .B2(n12534), .A(n12533), .ZN(n12535) );
  OAI21_X1 U14916 ( .B1(n15246), .B2(n12536), .A(n12535), .ZN(n12537) );
  AOI21_X1 U14917 ( .B1(n15101), .B2(n15236), .A(n12537), .ZN(n12538) );
  OAI21_X1 U14918 ( .B1(n12539), .B2(n15237), .A(n12538), .ZN(P1_U3236) );
  OAI21_X1 U14919 ( .B1(n12542), .B2(n12541), .A(n12540), .ZN(n12543) );
  XNOR2_X1 U14920 ( .A(n12543), .B(n12546), .ZN(n12599) );
  AOI211_X1 U14921 ( .C1(n12546), .C2(n12545), .A(n14217), .B(n12544), .ZN(
        n12550) );
  OR2_X1 U14922 ( .A1(n12547), .A2(n14197), .ZN(n12549) );
  NAND2_X1 U14923 ( .A1(n14082), .A2(n13942), .ZN(n12548) );
  NAND2_X1 U14924 ( .A1(n12549), .A2(n12548), .ZN(n13749) );
  NOR2_X1 U14925 ( .A1(n12550), .A2(n13749), .ZN(n12600) );
  MUX2_X1 U14926 ( .A(n12551), .B(n12600), .S(n14242), .Z(n12558) );
  OR2_X1 U14927 ( .A1(n12552), .A2(n12555), .ZN(n12553) );
  AND3_X1 U14928 ( .A1(n12554), .A2(n14262), .A3(n12553), .ZN(n12602) );
  OAI22_X1 U14929 ( .A1(n12555), .A2(n14226), .B1(n14239), .B2(n13751), .ZN(
        n12556) );
  AOI21_X1 U14930 ( .B1(n12602), .B2(n14273), .A(n12556), .ZN(n12557) );
  OAI211_X1 U14931 ( .C1(n12599), .C2(n14248), .A(n12558), .B(n12557), .ZN(
        P2_U3255) );
  INV_X1 U14932 ( .A(n12559), .ZN(n12561) );
  OAI222_X1 U14933 ( .A1(n12562), .A2(P3_U3151), .B1(n13707), .B2(n12561), 
        .C1(n12560), .C2(n13705), .ZN(P3_U3269) );
  XOR2_X1 U14934 ( .A(n12563), .B(n12564), .Z(n12624) );
  AOI22_X1 U14935 ( .A1(n13519), .A2(n13058), .B1(n15544), .B2(n13057), .ZN(
        n12570) );
  INV_X1 U14936 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12568) );
  XNOR2_X1 U14937 ( .A(n12565), .B(n12564), .ZN(n12566) );
  OAI222_X1 U14938 ( .A1(n15513), .A2(n13524), .B1(n15516), .B2(n13076), .C1(
        n12566), .C2(n13522), .ZN(n12621) );
  INV_X1 U14939 ( .A(n12621), .ZN(n12567) );
  MUX2_X1 U14940 ( .A(n12568), .B(n12567), .S(n15524), .Z(n12569) );
  OAI211_X1 U14941 ( .C1(n12624), .C2(n13529), .A(n12570), .B(n12569), .ZN(
        P3_U3220) );
  AND2_X1 U14942 ( .A1(n12571), .A2(n14366), .ZN(n12573) );
  NOR3_X1 U14943 ( .A1(n12574), .A2(n12573), .A3(n12572), .ZN(n12578) );
  MUX2_X1 U14944 ( .A(n12578), .B(n12575), .S(n15500), .Z(n12576) );
  OAI21_X1 U14945 ( .B1(n7444), .B2(n14362), .A(n12576), .ZN(P2_U3511) );
  INV_X1 U14946 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n12577) );
  MUX2_X1 U14947 ( .A(n12578), .B(n12577), .S(n15492), .Z(n12579) );
  OAI21_X1 U14948 ( .B1(n7444), .B2(n14428), .A(n12579), .ZN(P2_U3466) );
  XOR2_X1 U14949 ( .A(n12580), .B(n12582), .Z(n12650) );
  INV_X1 U14950 ( .A(n12650), .ZN(n12595) );
  XOR2_X1 U14951 ( .A(n12581), .B(n12582), .Z(n12586) );
  OAI22_X1 U14952 ( .A1(n14199), .A2(n12584), .B1(n12583), .B2(n14197), .ZN(
        n13867) );
  INV_X1 U14953 ( .A(n13867), .ZN(n12585) );
  OAI21_X1 U14954 ( .B1(n12586), .B2(n14217), .A(n12585), .ZN(n12648) );
  NAND2_X1 U14955 ( .A1(n12648), .A2(n14242), .ZN(n12594) );
  INV_X1 U14956 ( .A(n12587), .ZN(n12588) );
  AOI211_X1 U14957 ( .C1(n12589), .C2(n12588), .A(n14363), .B(n12637), .ZN(
        n12649) );
  NOR2_X1 U14958 ( .A1(n13870), .A2(n14226), .ZN(n12592) );
  OAI22_X1 U14959 ( .A1(n14242), .A2(n12590), .B1(n13865), .B2(n14239), .ZN(
        n12591) );
  AOI211_X1 U14960 ( .C1(n12649), .C2(n14273), .A(n12592), .B(n12591), .ZN(
        n12593) );
  OAI211_X1 U14961 ( .C1(n12595), .C2(n14248), .A(n12594), .B(n12593), .ZN(
        P2_U3252) );
  INV_X1 U14962 ( .A(n12596), .ZN(n12739) );
  OAI222_X1 U14963 ( .A1(n12598), .A2(P2_U3088), .B1(n14447), .B2(n12739), 
        .C1(n12597), .C2(n12742), .ZN(P2_U3301) );
  INV_X1 U14964 ( .A(n12599), .ZN(n12603) );
  INV_X1 U14965 ( .A(n12600), .ZN(n12601) );
  AOI211_X1 U14966 ( .C1(n14366), .C2(n12603), .A(n12602), .B(n12601), .ZN(
        n12606) );
  AOI22_X1 U14967 ( .A1(n14434), .A2(n13753), .B1(P2_REG0_REG_10__SCAN_IN), 
        .B2(n15492), .ZN(n12604) );
  OAI21_X1 U14968 ( .B1(n12606), .B2(n15492), .A(n12604), .ZN(P2_U3460) );
  AOI22_X1 U14969 ( .A1(n14374), .A2(n13753), .B1(P2_REG1_REG_10__SCAN_IN), 
        .B2(n15500), .ZN(n12605) );
  OAI21_X1 U14970 ( .B1(n12606), .B2(n15500), .A(n12605), .ZN(P2_U3509) );
  XOR2_X1 U14971 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .Z(n12613) );
  XNOR2_X1 U14972 ( .A(n15163), .B(n12613), .ZN(n12614) );
  NAND2_X1 U14973 ( .A1(n15160), .A2(n15159), .ZN(n12616) );
  XNOR2_X1 U14974 ( .A(n12616), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  MUX2_X1 U14975 ( .A(P3_REG0_REG_13__SCAN_IN), .B(n12621), .S(n15585), .Z(
        n12617) );
  AOI21_X1 U14976 ( .B1(n13670), .B2(n13058), .A(n12617), .ZN(n12618) );
  OAI21_X1 U14977 ( .B1(n12624), .B2(n13673), .A(n12618), .ZN(P3_U3429) );
  INV_X1 U14978 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n15703) );
  NAND2_X1 U14979 ( .A1(n12619), .A2(P3_U3897), .ZN(n12620) );
  OAI21_X1 U14980 ( .B1(P3_U3897), .B2(n15703), .A(n12620), .ZN(P3_U3521) );
  MUX2_X1 U14981 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n12621), .S(n15595), .Z(
        n12622) );
  AOI21_X1 U14982 ( .B1(n13590), .B2(n13058), .A(n12622), .ZN(n12623) );
  OAI21_X1 U14983 ( .B1(n12624), .B2(n13592), .A(n12623), .ZN(P3_U3472) );
  MUX2_X1 U14984 ( .A(P3_REG1_REG_9__SCAN_IN), .B(n12625), .S(n15595), .Z(
        n12626) );
  AOI21_X1 U14985 ( .B1(n13590), .B2(n13038), .A(n12626), .ZN(n12627) );
  OAI21_X1 U14986 ( .B1(n13592), .B2(n12628), .A(n12627), .ZN(P3_U3468) );
  INV_X1 U14987 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n13153) );
  MUX2_X1 U14988 ( .A(n13153), .B(n12629), .S(n15595), .Z(n12631) );
  NAND2_X1 U14989 ( .A1(n13590), .A2(n12988), .ZN(n12630) );
  OAI211_X1 U14990 ( .C1(n12632), .C2(n13592), .A(n12631), .B(n12630), .ZN(
        P3_U3471) );
  INV_X1 U14991 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n15705) );
  NAND2_X1 U14992 ( .A1(n12633), .A2(P3_U3897), .ZN(n12634) );
  OAI21_X1 U14993 ( .B1(P3_U3897), .B2(n15705), .A(n12634), .ZN(P3_U3519) );
  XNOR2_X1 U14994 ( .A(n12635), .B(n12643), .ZN(n12636) );
  AOI222_X1 U14995 ( .A1(n14252), .A2(n12636), .B1(n13938), .B2(n14082), .C1(
        n13940), .C2(n14097), .ZN(n14379) );
  INV_X1 U14996 ( .A(n12637), .ZN(n12639) );
  INV_X1 U14997 ( .A(n14260), .ZN(n12638) );
  AOI211_X1 U14998 ( .C1(n14377), .C2(n12639), .A(n14363), .B(n12638), .ZN(
        n14376) );
  INV_X1 U14999 ( .A(n13727), .ZN(n12640) );
  AOI22_X1 U15000 ( .A1(n14264), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n14276), 
        .B2(n12640), .ZN(n12641) );
  OAI21_X1 U15001 ( .B1(n12642), .B2(n14226), .A(n12641), .ZN(n12646) );
  XNOR2_X1 U15002 ( .A(n12644), .B(n12643), .ZN(n14380) );
  NOR2_X1 U15003 ( .A1(n14380), .A2(n14248), .ZN(n12645) );
  AOI211_X1 U15004 ( .C1(n14376), .C2(n14273), .A(n12646), .B(n12645), .ZN(
        n12647) );
  OAI21_X1 U15005 ( .B1(n14379), .B2(n14280), .A(n12647), .ZN(P2_U3251) );
  INV_X1 U15006 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n12651) );
  AOI211_X1 U15007 ( .C1(n12650), .C2(n14366), .A(n12649), .B(n12648), .ZN(
        n12653) );
  MUX2_X1 U15008 ( .A(n12651), .B(n12653), .S(n15494), .Z(n12652) );
  OAI21_X1 U15009 ( .B1(n13870), .B2(n14428), .A(n12652), .ZN(P2_U3469) );
  MUX2_X1 U15010 ( .A(n12654), .B(n12653), .S(n15502), .Z(n12655) );
  OAI21_X1 U15011 ( .B1(n13870), .B2(n14362), .A(n12655), .ZN(P2_U3512) );
  XNOR2_X1 U15012 ( .A(n14654), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12662) );
  XNOR2_X1 U15013 ( .A(n12659), .B(n12658), .ZN(n15262) );
  NOR2_X1 U15014 ( .A1(n12661), .A2(n12662), .ZN(n14653) );
  AOI211_X1 U15015 ( .C1(n12662), .C2(n12661), .A(n14687), .B(n14653), .ZN(
        n12675) );
  OAI21_X1 U15016 ( .B1(n12665), .B2(n12664), .A(n12663), .ZN(n12666) );
  NOR2_X1 U15017 ( .A1(n12666), .A2(n15264), .ZN(n12667) );
  AOI21_X1 U15018 ( .B1(n15264), .B2(n12666), .A(n12667), .ZN(n15261) );
  NAND2_X1 U15019 ( .A1(n15261), .A2(n15260), .ZN(n15259) );
  INV_X1 U15020 ( .A(n12667), .ZN(n12668) );
  NAND2_X1 U15021 ( .A1(n15259), .A2(n12668), .ZN(n12670) );
  MUX2_X1 U15022 ( .A(n14908), .B(P1_REG2_REG_16__SCAN_IN), .S(n14654), .Z(
        n12669) );
  NOR2_X1 U15023 ( .A1(n12670), .A2(n12669), .ZN(n14660) );
  AOI211_X1 U15024 ( .C1(n12670), .C2(n12669), .A(n14677), .B(n14660), .ZN(
        n12674) );
  NOR2_X1 U15025 ( .A1(n12671), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14517) );
  AOI21_X1 U15026 ( .B1(n15255), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14517), 
        .ZN(n12672) );
  OAI21_X1 U15027 ( .B1(n14686), .B2(n14657), .A(n12672), .ZN(n12673) );
  OR3_X1 U15028 ( .A1(n12675), .A2(n12674), .A3(n12673), .ZN(P1_U3259) );
  AOI22_X1 U15029 ( .A1(n12677), .A2(n14276), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14264), .ZN(n12680) );
  NAND2_X1 U15030 ( .A1(n12678), .A2(n14278), .ZN(n12679) );
  OAI211_X1 U15031 ( .C1(n12681), .C2(n14266), .A(n12680), .B(n12679), .ZN(
        n12682) );
  AOI21_X1 U15032 ( .B1(n7139), .B2(n14242), .A(n12682), .ZN(n12683) );
  OAI21_X1 U15033 ( .B1(n14248), .B2(n12684), .A(n12683), .ZN(P2_U3237) );
  OR2_X1 U15034 ( .A1(n15092), .A2(n12779), .ZN(n12685) );
  NAND2_X1 U15035 ( .A1(n15073), .A2(n12690), .ZN(n12691) );
  INV_X1 U15036 ( .A(n15058), .ZN(n14877) );
  AOI22_X1 U15037 ( .A1(n14870), .A2(n14868), .B1(n14877), .B2(n14889), .ZN(
        n12693) );
  INV_X1 U15038 ( .A(n14608), .ZN(n14567) );
  OR2_X1 U15039 ( .A1(n15036), .A2(n14567), .ZN(n12695) );
  NAND2_X1 U15040 ( .A1(n14794), .A2(n14793), .ZN(n12698) );
  INV_X1 U15041 ( .A(n14607), .ZN(n14568) );
  NAND2_X1 U15042 ( .A1(n15025), .A2(n14568), .ZN(n12697) );
  INV_X1 U15043 ( .A(n14605), .ZN(n12856) );
  NAND2_X1 U15044 ( .A1(n15012), .A2(n12856), .ZN(n12700) );
  NAND2_X1 U15045 ( .A1(n14750), .A2(n14765), .ZN(n12702) );
  NOR2_X1 U15046 ( .A1(n14750), .A2(n14765), .ZN(n12701) );
  NAND2_X1 U15047 ( .A1(n14726), .A2(n14728), .ZN(n14725) );
  INV_X1 U15048 ( .A(n14737), .ZN(n15000) );
  INV_X1 U15049 ( .A(n15078), .ZN(n14938) );
  INV_X1 U15050 ( .A(n15073), .ZN(n14909) );
  INV_X1 U15051 ( .A(n14781), .ZN(n14784) );
  INV_X1 U15052 ( .A(n15012), .ZN(n14768) );
  INV_X1 U15053 ( .A(n14750), .ZN(n15003) );
  AOI211_X1 U15054 ( .C1(n14991), .C2(n6413), .A(n14906), .B(n14692), .ZN(
        n14994) );
  AOI22_X1 U15055 ( .A1(n14603), .A2(n14962), .B1(n14602), .B2(n14960), .ZN(
        n14992) );
  NAND2_X1 U15056 ( .A1(n14991), .A2(n14956), .ZN(n12705) );
  INV_X1 U15057 ( .A(n12703), .ZN(n12882) );
  AOI22_X1 U15058 ( .A1(n12882), .A2(n14934), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n14920), .ZN(n12704) );
  OAI211_X1 U15059 ( .C1(n14992), .C2(n14920), .A(n12705), .B(n12704), .ZN(
        n12706) );
  AOI21_X1 U15060 ( .B1(n14994), .B2(n14924), .A(n12706), .ZN(n12737) );
  INV_X1 U15061 ( .A(n12707), .ZN(n12735) );
  NAND2_X1 U15062 ( .A1(n15085), .A2(n14612), .ZN(n12710) );
  INV_X1 U15063 ( .A(n12710), .ZN(n14926) );
  NOR2_X1 U15064 ( .A1(n12711), .A2(n14926), .ZN(n12713) );
  NOR2_X1 U15065 ( .A1(n15078), .A2(n14961), .ZN(n12712) );
  AOI21_X1 U15066 ( .B1(n14927), .B2(n12713), .A(n12712), .ZN(n12714) );
  NAND2_X1 U15067 ( .A1(n15073), .A2(n14887), .ZN(n12716) );
  OR2_X1 U15068 ( .A1(n15073), .A2(n14887), .ZN(n12717) );
  INV_X1 U15069 ( .A(n12720), .ZN(n12721) );
  INV_X1 U15070 ( .A(n14853), .ZN(n12723) );
  OR2_X1 U15071 ( .A1(n6628), .A2(n14609), .ZN(n12724) );
  NAND2_X1 U15072 ( .A1(n15043), .A2(n14825), .ZN(n14804) );
  NAND2_X1 U15073 ( .A1(n14804), .A2(n14567), .ZN(n12727) );
  INV_X1 U15074 ( .A(n14804), .ZN(n12726) );
  AOI22_X1 U15075 ( .A1(n15036), .A2(n12727), .B1(n12726), .B2(n14608), .ZN(
        n12728) );
  AND2_X2 U15076 ( .A1(n12728), .A2(n14806), .ZN(n14789) );
  NOR2_X1 U15077 ( .A1(n15036), .A2(n14608), .ZN(n14805) );
  NAND2_X1 U15078 ( .A1(n12756), .A2(n14797), .ZN(n14790) );
  OAI21_X1 U15079 ( .B1(n15025), .B2(n14607), .A(n14790), .ZN(n12729) );
  AOI21_X1 U15080 ( .B1(n14789), .B2(n14805), .A(n12729), .ZN(n12730) );
  OR2_X1 U15081 ( .A1(n14781), .A2(n14606), .ZN(n12731) );
  NAND2_X1 U15082 ( .A1(n15012), .A2(n14605), .ZN(n12732) );
  NAND2_X1 U15083 ( .A1(n14750), .A2(n14604), .ZN(n12733) );
  AOI21_X1 U15084 ( .B1(n12735), .B2(n12734), .A(n14710), .ZN(n14995) );
  NAND2_X1 U15085 ( .A1(n14995), .A2(n14841), .ZN(n12736) );
  OAI211_X1 U15086 ( .C1(n14997), .C2(n14754), .A(n12737), .B(n12736), .ZN(
        P1_U3265) );
  OAI222_X1 U15087 ( .A1(n12740), .A2(P1_U3086), .B1(n15141), .B2(n12739), 
        .C1(n12738), .C2(n15149), .ZN(P1_U3329) );
  OAI222_X1 U15088 ( .A1(n14447), .A2(n15143), .B1(P2_U3088), .B2(n12741), 
        .C1(n12743), .C2(n12742), .ZN(P2_U3297) );
  MUX2_X1 U15089 ( .A(n12745), .B(n12744), .S(n15502), .Z(n12746) );
  OAI21_X1 U15090 ( .B1(n12747), .B2(n14362), .A(n12746), .ZN(P2_U3500) );
  NAND2_X1 U15091 ( .A1(n14991), .A2(n12872), .ZN(n12749) );
  NAND2_X1 U15092 ( .A1(n14708), .A2(n12877), .ZN(n12748) );
  NAND2_X1 U15093 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  XNOR2_X1 U15094 ( .A(n12750), .B(n12875), .ZN(n12753) );
  NOR2_X1 U15095 ( .A1(n14732), .A2(n12857), .ZN(n12751) );
  AOI21_X1 U15096 ( .B1(n14991), .B2(n12871), .A(n12751), .ZN(n12752) );
  XNOR2_X1 U15097 ( .A(n12753), .B(n12752), .ZN(n12885) );
  INV_X1 U15098 ( .A(n12885), .ZN(n12754) );
  NAND2_X1 U15099 ( .A1(n12754), .A2(n14589), .ZN(n12891) );
  OAI22_X1 U15100 ( .A1(n12756), .A2(n12857), .B1(n14797), .B2(n12855), .ZN(
        n12837) );
  INV_X1 U15101 ( .A(n12837), .ZN(n12840) );
  OAI22_X1 U15102 ( .A1(n12756), .A2(n12755), .B1(n14797), .B2(n12857), .ZN(
        n12757) );
  XNOR2_X1 U15103 ( .A(n12757), .B(n12866), .ZN(n12838) );
  INV_X1 U15104 ( .A(n12838), .ZN(n12839) );
  AOI22_X1 U15105 ( .A1(n15036), .A2(n12872), .B1(n12877), .B2(n14608), .ZN(
        n12836) );
  NAND2_X1 U15106 ( .A1(n15036), .A2(n12871), .ZN(n12759) );
  NAND2_X1 U15107 ( .A1(n14608), .A2(n12872), .ZN(n12758) );
  NAND2_X1 U15108 ( .A1(n12759), .A2(n12758), .ZN(n12760) );
  XNOR2_X1 U15109 ( .A(n12760), .B(n12866), .ZN(n12834) );
  INV_X1 U15110 ( .A(n12834), .ZN(n12835) );
  AOI22_X1 U15111 ( .A1(n15043), .A2(n12872), .B1(n12877), .B2(n14825), .ZN(
        n12833) );
  NAND2_X1 U15112 ( .A1(n15043), .A2(n12871), .ZN(n12762) );
  NAND2_X1 U15113 ( .A1(n14825), .A2(n12872), .ZN(n12761) );
  NAND2_X1 U15114 ( .A1(n12762), .A2(n12761), .ZN(n12763) );
  XNOR2_X1 U15115 ( .A(n12763), .B(n12866), .ZN(n12831) );
  INV_X1 U15116 ( .A(n12831), .ZN(n12832) );
  NAND2_X1 U15117 ( .A1(n15097), .A2(n12871), .ZN(n12768) );
  NAND2_X1 U15118 ( .A1(n12872), .A2(n14613), .ZN(n12767) );
  NAND2_X1 U15119 ( .A1(n12768), .A2(n12767), .ZN(n12769) );
  XNOR2_X1 U15120 ( .A(n12769), .B(n12866), .ZN(n12774) );
  NOR2_X1 U15121 ( .A1(n12855), .A2(n12770), .ZN(n12771) );
  AOI21_X1 U15122 ( .B1(n15097), .B2(n11176), .A(n12771), .ZN(n12772) );
  XNOR2_X1 U15123 ( .A(n12774), .B(n12772), .ZN(n14495) );
  INV_X1 U15124 ( .A(n12772), .ZN(n12773) );
  NAND2_X1 U15125 ( .A1(n12774), .A2(n12773), .ZN(n12775) );
  NAND2_X1 U15126 ( .A1(n14494), .A2(n12775), .ZN(n14553) );
  NAND2_X1 U15127 ( .A1(n15092), .A2(n12871), .ZN(n12777) );
  NAND2_X1 U15128 ( .A1(n14963), .A2(n12872), .ZN(n12776) );
  NAND2_X1 U15129 ( .A1(n12777), .A2(n12776), .ZN(n12778) );
  XNOR2_X1 U15130 ( .A(n12778), .B(n12866), .ZN(n12783) );
  NOR2_X1 U15131 ( .A1(n12779), .A2(n12855), .ZN(n12780) );
  AOI21_X1 U15132 ( .B1(n15092), .B2(n11176), .A(n12780), .ZN(n12781) );
  XNOR2_X1 U15133 ( .A(n12783), .B(n12781), .ZN(n14552) );
  NAND2_X1 U15134 ( .A1(n14553), .A2(n14552), .ZN(n14551) );
  INV_X1 U15135 ( .A(n12781), .ZN(n12782) );
  NAND2_X1 U15136 ( .A1(n12783), .A2(n12782), .ZN(n12784) );
  NAND2_X1 U15137 ( .A1(n14551), .A2(n12784), .ZN(n14463) );
  NAND2_X1 U15138 ( .A1(n15085), .A2(n12871), .ZN(n12786) );
  NAND2_X1 U15139 ( .A1(n14612), .A2(n12872), .ZN(n12785) );
  NAND2_X1 U15140 ( .A1(n12786), .A2(n12785), .ZN(n12787) );
  XNOR2_X1 U15141 ( .A(n12787), .B(n12875), .ZN(n12790) );
  AND2_X1 U15142 ( .A1(n14612), .A2(n12877), .ZN(n12788) );
  AOI21_X1 U15143 ( .B1(n15085), .B2(n11176), .A(n12788), .ZN(n12789) );
  XNOR2_X1 U15144 ( .A(n12790), .B(n12789), .ZN(n14464) );
  NAND2_X1 U15145 ( .A1(n12790), .A2(n12789), .ZN(n12791) );
  NAND2_X1 U15146 ( .A1(n15078), .A2(n12871), .ZN(n12793) );
  NAND2_X1 U15147 ( .A1(n14961), .A2(n12872), .ZN(n12792) );
  NAND2_X1 U15148 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  XNOR2_X1 U15149 ( .A(n12794), .B(n12875), .ZN(n14514) );
  NAND2_X1 U15150 ( .A1(n15078), .A2(n12872), .ZN(n12796) );
  NAND2_X1 U15151 ( .A1(n14961), .A2(n12877), .ZN(n12795) );
  AND2_X1 U15152 ( .A1(n12796), .A2(n12795), .ZN(n14512) );
  NAND2_X1 U15153 ( .A1(n15073), .A2(n12871), .ZN(n12798) );
  NAND2_X1 U15154 ( .A1(n14887), .A2(n12872), .ZN(n12797) );
  NAND2_X1 U15155 ( .A1(n12798), .A2(n12797), .ZN(n12799) );
  XNOR2_X1 U15156 ( .A(n12799), .B(n12866), .ZN(n14511) );
  NAND2_X1 U15157 ( .A1(n15073), .A2(n12872), .ZN(n12801) );
  NAND2_X1 U15158 ( .A1(n14887), .A2(n12877), .ZN(n12800) );
  NAND2_X1 U15159 ( .A1(n12801), .A2(n12800), .ZN(n14510) );
  NAND2_X1 U15160 ( .A1(n14511), .A2(n14510), .ZN(n12804) );
  OAI21_X1 U15161 ( .B1(n14514), .B2(n14512), .A(n12804), .ZN(n12802) );
  INV_X1 U15162 ( .A(n12802), .ZN(n12803) );
  NAND3_X1 U15163 ( .A1(n12804), .A2(n14514), .A3(n14512), .ZN(n12807) );
  INV_X1 U15164 ( .A(n14511), .ZN(n12806) );
  INV_X1 U15165 ( .A(n14510), .ZN(n12805) );
  NAND2_X1 U15166 ( .A1(n12806), .A2(n12805), .ZN(n14523) );
  NAND2_X1 U15167 ( .A1(n14898), .A2(n12871), .ZN(n12809) );
  NAND2_X1 U15168 ( .A1(n14610), .A2(n12872), .ZN(n12808) );
  NAND2_X1 U15169 ( .A1(n12809), .A2(n12808), .ZN(n12810) );
  XNOR2_X1 U15170 ( .A(n12810), .B(n12866), .ZN(n12815) );
  AND2_X1 U15171 ( .A1(n14610), .A2(n12877), .ZN(n12811) );
  AOI21_X1 U15172 ( .B1(n14898), .B2(n11176), .A(n12811), .ZN(n12813) );
  XNOR2_X1 U15173 ( .A(n12815), .B(n12813), .ZN(n14524) );
  NAND2_X1 U15174 ( .A1(n12812), .A2(n14524), .ZN(n14527) );
  INV_X1 U15175 ( .A(n12813), .ZN(n12814) );
  OR2_X1 U15176 ( .A1(n12815), .A2(n12814), .ZN(n12816) );
  INV_X1 U15177 ( .A(n14889), .ZN(n14530) );
  OAI22_X1 U15178 ( .A1(n14877), .A2(n12857), .B1(n14530), .B2(n12855), .ZN(
        n12820) );
  NAND2_X1 U15179 ( .A1(n15058), .A2(n12871), .ZN(n12818) );
  NAND2_X1 U15180 ( .A1(n14889), .A2(n12872), .ZN(n12817) );
  NAND2_X1 U15181 ( .A1(n12818), .A2(n12817), .ZN(n12819) );
  XNOR2_X1 U15182 ( .A(n12819), .B(n12866), .ZN(n12821) );
  INV_X1 U15183 ( .A(n12820), .ZN(n12823) );
  INV_X1 U15184 ( .A(n12821), .ZN(n12822) );
  NAND2_X1 U15185 ( .A1(n14861), .A2(n12871), .ZN(n12825) );
  NAND2_X1 U15186 ( .A1(n14609), .A2(n12872), .ZN(n12824) );
  AND2_X1 U15187 ( .A1(n14609), .A2(n12877), .ZN(n12827) );
  AOI21_X1 U15188 ( .B1(n14861), .B2(n11176), .A(n12827), .ZN(n12829) );
  INV_X1 U15189 ( .A(n12828), .ZN(n12830) );
  XNOR2_X1 U15190 ( .A(n12831), .B(n12833), .ZN(n14544) );
  XOR2_X1 U15191 ( .A(n12836), .B(n12834), .Z(n14487) );
  XNOR2_X1 U15192 ( .A(n12838), .B(n12837), .ZN(n14565) );
  AOI22_X1 U15193 ( .A1(n15025), .A2(n12872), .B1(n12877), .B2(n14607), .ZN(
        n12844) );
  NAND2_X1 U15194 ( .A1(n15025), .A2(n12871), .ZN(n12842) );
  NAND2_X1 U15195 ( .A1(n14607), .A2(n12872), .ZN(n12841) );
  NAND2_X1 U15196 ( .A1(n12842), .A2(n12841), .ZN(n12843) );
  XNOR2_X1 U15197 ( .A(n12843), .B(n12866), .ZN(n12846) );
  XOR2_X1 U15198 ( .A(n12844), .B(n12846), .Z(n14472) );
  INV_X1 U15199 ( .A(n12844), .ZN(n12845) );
  NAND2_X1 U15200 ( .A1(n14781), .A2(n12871), .ZN(n12848) );
  NAND2_X1 U15201 ( .A1(n14606), .A2(n12872), .ZN(n12847) );
  NAND2_X1 U15202 ( .A1(n12848), .A2(n12847), .ZN(n12849) );
  XNOR2_X1 U15203 ( .A(n12849), .B(n12866), .ZN(n12852) );
  AOI22_X1 U15204 ( .A1(n14781), .A2(n12872), .B1(n12877), .B2(n14606), .ZN(
        n12850) );
  XNOR2_X1 U15205 ( .A(n12852), .B(n12850), .ZN(n14536) );
  INV_X1 U15206 ( .A(n12850), .ZN(n12851) );
  NAND2_X1 U15207 ( .A1(n12854), .A2(n12853), .ZN(n14504) );
  OAI22_X1 U15208 ( .A1(n14768), .A2(n12857), .B1(n12856), .B2(n12855), .ZN(
        n12861) );
  NAND2_X1 U15209 ( .A1(n15012), .A2(n12871), .ZN(n12859) );
  NAND2_X1 U15210 ( .A1(n14605), .A2(n12872), .ZN(n12858) );
  NAND2_X1 U15211 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  XNOR2_X1 U15212 ( .A(n12860), .B(n12866), .ZN(n12862) );
  XOR2_X1 U15213 ( .A(n12861), .B(n12862), .Z(n14505) );
  OR2_X1 U15214 ( .A1(n12862), .A2(n12861), .ZN(n12863) );
  NAND2_X1 U15215 ( .A1(n14750), .A2(n12871), .ZN(n12865) );
  NAND2_X1 U15216 ( .A1(n14604), .A2(n12872), .ZN(n12864) );
  NAND2_X1 U15217 ( .A1(n12865), .A2(n12864), .ZN(n12867) );
  XNOR2_X1 U15218 ( .A(n12867), .B(n12866), .ZN(n12868) );
  AOI22_X1 U15219 ( .A1(n14750), .A2(n12872), .B1(n12877), .B2(n14604), .ZN(
        n12869) );
  XNOR2_X1 U15220 ( .A(n12868), .B(n12869), .ZN(n14583) );
  INV_X1 U15221 ( .A(n12868), .ZN(n12870) );
  NAND2_X1 U15222 ( .A1(n14737), .A2(n12871), .ZN(n12874) );
  NAND2_X1 U15223 ( .A1(n14603), .A2(n12872), .ZN(n12873) );
  NAND2_X1 U15224 ( .A1(n12874), .A2(n12873), .ZN(n12876) );
  XNOR2_X1 U15225 ( .A(n12876), .B(n12875), .ZN(n12881) );
  AND2_X1 U15226 ( .A1(n14603), .A2(n12877), .ZN(n12878) );
  AOI21_X1 U15227 ( .B1(n14737), .B2(n11176), .A(n12878), .ZN(n12880) );
  XNOR2_X1 U15228 ( .A(n12881), .B(n12880), .ZN(n14454) );
  INV_X1 U15229 ( .A(n14454), .ZN(n12879) );
  NAND2_X1 U15230 ( .A1(n12881), .A2(n12880), .ZN(n12884) );
  AOI22_X1 U15231 ( .A1(n12882), .A2(n14597), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12883) );
  OAI21_X1 U15232 ( .B1(n14992), .B2(n14595), .A(n12883), .ZN(n12887) );
  NOR3_X1 U15233 ( .A1(n12885), .A2(n15237), .A3(n12884), .ZN(n12886) );
  AOI211_X1 U15234 ( .C1(n14586), .C2(n14991), .A(n12887), .B(n12886), .ZN(
        n12888) );
  OAI211_X1 U15235 ( .C1(n12891), .C2(n12890), .A(n12889), .B(n12888), .ZN(
        P1_U3220) );
  INV_X1 U15236 ( .A(n12892), .ZN(n14448) );
  OAI222_X1 U15237 ( .A1(n15149), .A2(n12893), .B1(n15141), .B2(n14448), .C1(
        n10115), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U15238 ( .A(n12894), .ZN(n12936) );
  OAI222_X1 U15239 ( .A1(n12896), .A2(P1_U3086), .B1(n15141), .B2(n12936), 
        .C1(n12895), .C2(n15149), .ZN(P1_U3326) );
  XNOR2_X1 U15240 ( .A(n13350), .B(n6400), .ZN(n12904) );
  INV_X1 U15241 ( .A(n12904), .ZN(n12897) );
  NAND2_X1 U15242 ( .A1(n12897), .A2(n13095), .ZN(n12910) );
  INV_X1 U15243 ( .A(n12898), .ZN(n12899) );
  NAND4_X1 U15244 ( .A1(n12909), .A2(n13095), .A3(n12899), .A4(n12904), .ZN(
        n12908) );
  NAND2_X1 U15245 ( .A1(n13354), .A2(n13100), .ZN(n12901) );
  AOI22_X1 U15246 ( .A1(n13349), .A2(n13111), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12900) );
  OAI211_X1 U15247 ( .C1(n12902), .C2(n13098), .A(n12901), .B(n12900), .ZN(
        n12906) );
  NOR4_X1 U15248 ( .A1(n12904), .A2(n12903), .A3(n13115), .A4(n13379), .ZN(
        n12905) );
  AOI211_X1 U15249 ( .C1(n13112), .C2(n13548), .A(n12906), .B(n12905), .ZN(
        n12907) );
  OAI211_X1 U15250 ( .C1(n12910), .C2(n12909), .A(n12908), .B(n12907), .ZN(
        P3_U3160) );
  AND2_X1 U15251 ( .A1(n14398), .A2(n14050), .ZN(n12912) );
  XNOR2_X1 U15252 ( .A(n12915), .B(n12914), .ZN(n12921) );
  INV_X1 U15253 ( .A(n14050), .ZN(n12919) );
  NAND2_X1 U15254 ( .A1(n12916), .A2(P2_B_REG_SCAN_IN), .ZN(n12917) );
  NAND2_X1 U15255 ( .A1(n14082), .A2(n12917), .ZN(n12944) );
  OAI22_X1 U15256 ( .A1(n12919), .A2(n14197), .B1(n12918), .B2(n12944), .ZN(
        n12920) );
  AOI21_X2 U15257 ( .B1(n12921), .B2(n14252), .A(n12920), .ZN(n14294) );
  AOI21_X1 U15258 ( .B1(n14292), .B2(n12923), .A(n14363), .ZN(n12924) );
  AND2_X1 U15259 ( .A1(n14042), .A2(n12924), .ZN(n14291) );
  NAND2_X1 U15260 ( .A1(n14292), .A2(n14278), .ZN(n12926) );
  NAND2_X1 U15261 ( .A1(n14280), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n12925) );
  OAI211_X1 U15262 ( .C1(n14239), .C2(n12927), .A(n12926), .B(n12925), .ZN(
        n12928) );
  OAI21_X1 U15263 ( .B1(n14295), .B2(n14248), .A(n12931), .ZN(P2_U3236) );
  OAI222_X1 U15264 ( .A1(n15149), .A2(n12933), .B1(n15141), .B2(n12932), .C1(
        n10007), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI222_X1 U15265 ( .A1(n13707), .A2(n12935), .B1(n13705), .B2(n12934), .C1(
        P3_U3151), .C2(n13313), .ZN(P3_U3276) );
  OAI222_X1 U15266 ( .A1(n12742), .A2(n12938), .B1(P2_U3088), .B2(n12937), 
        .C1(n14447), .C2(n12936), .ZN(P2_U3298) );
  OAI222_X1 U15267 ( .A1(n15149), .A2(n12941), .B1(n15141), .B2(n12940), .C1(
        P1_U3086), .C2(n12939), .ZN(P1_U3334) );
  XNOR2_X1 U15268 ( .A(n14387), .B(n14040), .ZN(n12942) );
  INV_X1 U15269 ( .A(n13928), .ZN(n12943) );
  OR2_X1 U15270 ( .A1(n12944), .A2(n12943), .ZN(n14035) );
  XOR2_X1 U15271 ( .A(n12946), .B(n12945), .Z(n12952) );
  AND2_X1 U15272 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13218) );
  AOI21_X1 U15273 ( .B1(n13100), .B2(n13538), .A(n13218), .ZN(n12947) );
  OAI21_X1 U15274 ( .B1(n12948), .B2(n13098), .A(n12947), .ZN(n12950) );
  NOR2_X1 U15275 ( .A1(n13680), .A2(n13103), .ZN(n12949) );
  AOI211_X1 U15276 ( .C1(n13532), .C2(n13045), .A(n12950), .B(n12949), .ZN(
        n12951) );
  OAI21_X1 U15277 ( .B1(n12952), .B2(n13115), .A(n12951), .ZN(P3_U3155) );
  INV_X1 U15278 ( .A(n13630), .ZN(n12962) );
  OAI21_X1 U15279 ( .B1(n12954), .B2(n12953), .A(n12955), .ZN(n13064) );
  OAI21_X1 U15280 ( .B1(n6502), .B2(n13431), .A(n13023), .ZN(n12957) );
  NAND2_X1 U15281 ( .A1(n12957), .A2(n13095), .ZN(n12961) );
  AOI22_X1 U15282 ( .A1(n13440), .A2(n13107), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12958) );
  OAI21_X1 U15283 ( .B1(n13419), .B2(n13109), .A(n12958), .ZN(n12959) );
  AOI21_X1 U15284 ( .B1(n13415), .B2(n13111), .A(n12959), .ZN(n12960) );
  OAI211_X1 U15285 ( .C1(n12962), .C2(n13103), .A(n12961), .B(n12960), .ZN(
        P3_U3156) );
  XNOR2_X1 U15286 ( .A(n12964), .B(n12963), .ZN(n12969) );
  AND2_X1 U15287 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13316) );
  AOI21_X1 U15288 ( .B1(n13100), .B2(n13470), .A(n13316), .ZN(n12966) );
  NAND2_X1 U15289 ( .A1(n13045), .A2(n13475), .ZN(n12965) );
  OAI211_X1 U15290 ( .C1(n13501), .C2(n13098), .A(n12966), .B(n12965), .ZN(
        n12967) );
  AOI21_X1 U15291 ( .B1(n13651), .B2(n13112), .A(n12967), .ZN(n12968) );
  OAI21_X1 U15292 ( .B1(n12969), .B2(n13115), .A(n12968), .ZN(P3_U3159) );
  AOI21_X1 U15293 ( .B1(n12971), .B2(n12970), .A(n6520), .ZN(n12976) );
  AOI22_X1 U15294 ( .A1(n13107), .A2(n13470), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12973) );
  NAND2_X1 U15295 ( .A1(n13045), .A2(n13437), .ZN(n12972) );
  OAI211_X1 U15296 ( .C1(n13418), .C2(n13109), .A(n12973), .B(n12972), .ZN(
        n12974) );
  AOI21_X1 U15297 ( .B1(n13641), .B2(n13112), .A(n12974), .ZN(n12975) );
  OAI21_X1 U15298 ( .B1(n12976), .B2(n13115), .A(n12975), .ZN(P3_U3163) );
  INV_X1 U15299 ( .A(n12977), .ZN(n12979) );
  NOR2_X1 U15300 ( .A1(n12978), .A2(n12979), .ZN(n12980) );
  AOI21_X1 U15301 ( .B1(n12979), .B2(n12978), .A(n12980), .ZN(n13072) );
  NAND2_X1 U15302 ( .A1(n13072), .A2(n13073), .ZN(n13071) );
  INV_X1 U15303 ( .A(n12980), .ZN(n12981) );
  NAND2_X1 U15304 ( .A1(n13071), .A2(n12981), .ZN(n12984) );
  XNOR2_X1 U15305 ( .A(n12982), .B(n13076), .ZN(n12983) );
  XNOR2_X1 U15306 ( .A(n12984), .B(n12983), .ZN(n12991) );
  NAND2_X1 U15307 ( .A1(n13100), .A2(n13537), .ZN(n12985) );
  NAND2_X1 U15308 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13159)
         );
  OAI211_X1 U15309 ( .C1(n13073), .C2(n13098), .A(n12985), .B(n13159), .ZN(
        n12986) );
  AOI21_X1 U15310 ( .B1(n12987), .B2(n13111), .A(n12986), .ZN(n12990) );
  NAND2_X1 U15311 ( .A1(n13112), .A2(n12988), .ZN(n12989) );
  OAI211_X1 U15312 ( .C1(n12991), .C2(n13115), .A(n12990), .B(n12989), .ZN(
        P3_U3164) );
  INV_X1 U15313 ( .A(n12993), .ZN(n12997) );
  NOR3_X1 U15314 ( .A1(n13021), .A2(n12995), .A3(n12994), .ZN(n12996) );
  OAI21_X1 U15315 ( .B1(n12997), .B2(n12996), .A(n13095), .ZN(n13002) );
  INV_X1 U15316 ( .A(n13392), .ZN(n12999) );
  AOI22_X1 U15317 ( .A1(n13119), .A2(n13107), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12998) );
  OAI21_X1 U15318 ( .B1(n12999), .B2(n13088), .A(n12998), .ZN(n13000) );
  AOI21_X1 U15319 ( .B1(n13100), .B2(n13118), .A(n13000), .ZN(n13001) );
  OAI211_X1 U15320 ( .C1(n13622), .C2(n13103), .A(n13002), .B(n13001), .ZN(
        P3_U3165) );
  XNOR2_X1 U15321 ( .A(n13003), .B(n13498), .ZN(n13004) );
  XNOR2_X1 U15322 ( .A(n13005), .B(n13004), .ZN(n13010) );
  NAND2_X1 U15323 ( .A1(n13107), .A2(n13538), .ZN(n13006) );
  NAND2_X1 U15324 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13254)
         );
  OAI211_X1 U15325 ( .C1(n13511), .C2(n13109), .A(n13006), .B(n13254), .ZN(
        n13008) );
  INV_X1 U15326 ( .A(n13585), .ZN(n13514) );
  NOR2_X1 U15327 ( .A1(n13514), .A2(n13103), .ZN(n13007) );
  AOI211_X1 U15328 ( .C1(n13512), .C2(n13045), .A(n13008), .B(n13007), .ZN(
        n13009) );
  OAI21_X1 U15329 ( .B1(n13010), .B2(n13115), .A(n13009), .ZN(P3_U3166) );
  XNOR2_X1 U15330 ( .A(n13012), .B(n13011), .ZN(n13017) );
  NOR2_X1 U15331 ( .A1(n15627), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13278) );
  AOI21_X1 U15332 ( .B1(n13100), .B2(n13469), .A(n13278), .ZN(n13014) );
  NAND2_X1 U15333 ( .A1(n13045), .A2(n13494), .ZN(n13013) );
  OAI211_X1 U15334 ( .C1(n13525), .C2(n13098), .A(n13014), .B(n13013), .ZN(
        n13015) );
  AOI21_X1 U15335 ( .B1(n13660), .B2(n13112), .A(n13015), .ZN(n13016) );
  OAI21_X1 U15336 ( .B1(n13017), .B2(n13115), .A(n13016), .ZN(P3_U3168) );
  INV_X1 U15337 ( .A(n13018), .ZN(n13020) );
  NOR2_X1 U15338 ( .A1(n13020), .A2(n13019), .ZN(n13022) );
  AOI21_X1 U15339 ( .B1(n13023), .B2(n13022), .A(n13021), .ZN(n13028) );
  AOI22_X1 U15340 ( .A1(n13120), .A2(n13107), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13025) );
  NAND2_X1 U15341 ( .A1(n13408), .A2(n13111), .ZN(n13024) );
  OAI211_X1 U15342 ( .C1(n13404), .C2(n13109), .A(n13025), .B(n13024), .ZN(
        n13026) );
  AOI21_X1 U15343 ( .B1(n13565), .B2(n13112), .A(n13026), .ZN(n13027) );
  OAI21_X1 U15344 ( .B1(n13028), .B2(n13115), .A(n13027), .ZN(P3_U3169) );
  OAI21_X1 U15345 ( .B1(n13030), .B2(n13029), .A(n10549), .ZN(n13031) );
  NAND2_X1 U15346 ( .A1(n13031), .A2(n13095), .ZN(n13042) );
  OAI21_X1 U15347 ( .B1(n13109), .B2(n13033), .A(n13032), .ZN(n13036) );
  NOR2_X1 U15348 ( .A1(n13098), .A2(n13034), .ZN(n13035) );
  NOR2_X1 U15349 ( .A1(n13036), .A2(n13035), .ZN(n13041) );
  NAND2_X1 U15350 ( .A1(n13111), .A2(n13037), .ZN(n13040) );
  NAND2_X1 U15351 ( .A1(n13112), .A2(n13038), .ZN(n13039) );
  NAND4_X1 U15352 ( .A1(n13042), .A2(n13041), .A3(n13040), .A4(n13039), .ZN(
        P3_U3171) );
  XNOR2_X1 U15353 ( .A(n13044), .B(n13043), .ZN(n13050) );
  AOI22_X1 U15354 ( .A1(n13065), .A2(n13100), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13047) );
  NAND2_X1 U15355 ( .A1(n13045), .A2(n13448), .ZN(n13046) );
  OAI211_X1 U15356 ( .C1(n13085), .C2(n13098), .A(n13047), .B(n13046), .ZN(
        n13048) );
  AOI21_X1 U15357 ( .B1(n13646), .B2(n13112), .A(n13048), .ZN(n13049) );
  OAI21_X1 U15358 ( .B1(n13050), .B2(n13115), .A(n13049), .ZN(P3_U3173) );
  NAND2_X1 U15359 ( .A1(n13052), .A2(n13051), .ZN(n13054) );
  XOR2_X1 U15360 ( .A(n13054), .B(n13053), .Z(n13061) );
  NAND2_X1 U15361 ( .A1(n13107), .A2(n10479), .ZN(n13055) );
  NAND2_X1 U15362 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13192)
         );
  OAI211_X1 U15363 ( .C1(n13524), .C2(n13109), .A(n13055), .B(n13192), .ZN(
        n13056) );
  AOI21_X1 U15364 ( .B1(n13057), .B2(n13111), .A(n13056), .ZN(n13060) );
  NAND2_X1 U15365 ( .A1(n13058), .A2(n13112), .ZN(n13059) );
  OAI211_X1 U15366 ( .C1(n13061), .C2(n13115), .A(n13060), .B(n13059), .ZN(
        P3_U3174) );
  INV_X1 U15367 ( .A(n13062), .ZN(n13063) );
  AOI21_X1 U15368 ( .B1(n13440), .B2(n13064), .A(n13063), .ZN(n13070) );
  AOI22_X1 U15369 ( .A1(n13065), .A2(n13107), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13067) );
  NAND2_X1 U15370 ( .A1(n13427), .A2(n13111), .ZN(n13066) );
  OAI211_X1 U15371 ( .C1(n13431), .C2(n13109), .A(n13067), .B(n13066), .ZN(
        n13068) );
  AOI21_X1 U15372 ( .B1(n13635), .B2(n13112), .A(n13068), .ZN(n13069) );
  OAI21_X1 U15373 ( .B1(n13070), .B2(n13115), .A(n13069), .ZN(P3_U3175) );
  OAI21_X1 U15374 ( .B1(n13073), .B2(n13072), .A(n13071), .ZN(n13074) );
  NAND2_X1 U15375 ( .A1(n13074), .A2(n13095), .ZN(n13080) );
  NAND2_X1 U15376 ( .A1(n13107), .A2(n13122), .ZN(n13075) );
  NAND2_X1 U15377 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n13139)
         );
  OAI211_X1 U15378 ( .C1(n13076), .C2(n13109), .A(n13075), .B(n13139), .ZN(
        n13077) );
  AOI21_X1 U15379 ( .B1(n13078), .B2(n13111), .A(n13077), .ZN(n13079) );
  OAI211_X1 U15380 ( .C1(n13103), .C2(n13601), .A(n13080), .B(n13079), .ZN(
        P3_U3176) );
  XNOR2_X1 U15381 ( .A(n13081), .B(n13469), .ZN(n13082) );
  XNOR2_X1 U15382 ( .A(n13083), .B(n13082), .ZN(n13091) );
  INV_X1 U15383 ( .A(n13084), .ZN(n13479) );
  NAND2_X1 U15384 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13290)
         );
  OAI21_X1 U15385 ( .B1(n13085), .B2(n13109), .A(n13290), .ZN(n13086) );
  AOI21_X1 U15386 ( .B1(n13107), .B2(n13487), .A(n13086), .ZN(n13087) );
  OAI21_X1 U15387 ( .B1(n13479), .B2(n13088), .A(n13087), .ZN(n13089) );
  AOI21_X1 U15388 ( .B1(n13580), .B2(n13112), .A(n13089), .ZN(n13090) );
  OAI21_X1 U15389 ( .B1(n13091), .B2(n13115), .A(n13090), .ZN(P3_U3178) );
  INV_X1 U15390 ( .A(n13615), .ZN(n13104) );
  OAI21_X1 U15391 ( .B1(n13094), .B2(n13093), .A(n13092), .ZN(n13096) );
  NAND2_X1 U15392 ( .A1(n13096), .A2(n13095), .ZN(n13102) );
  AOI22_X1 U15393 ( .A1(n13375), .A2(n13111), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13097) );
  OAI21_X1 U15394 ( .B1(n13404), .B2(n13098), .A(n13097), .ZN(n13099) );
  AOI21_X1 U15395 ( .B1(n13379), .B2(n13100), .A(n13099), .ZN(n13101) );
  OAI211_X1 U15396 ( .C1(n13104), .C2(n13103), .A(n13102), .B(n13101), .ZN(
        P3_U3180) );
  XOR2_X1 U15397 ( .A(n13106), .B(n13105), .Z(n13116) );
  NAND2_X1 U15398 ( .A1(n13107), .A2(n13121), .ZN(n13108) );
  NAND2_X1 U15399 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13238)
         );
  OAI211_X1 U15400 ( .C1(n13525), .C2(n13109), .A(n13108), .B(n13238), .ZN(
        n13110) );
  AOI21_X1 U15401 ( .B1(n13518), .B2(n13111), .A(n13110), .ZN(n13114) );
  NAND2_X1 U15402 ( .A1(n13669), .A2(n13112), .ZN(n13113) );
  OAI211_X1 U15403 ( .C1(n13116), .C2(n13115), .A(n13114), .B(n13113), .ZN(
        P3_U3181) );
  MUX2_X1 U15404 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13117), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15405 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n13354), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15406 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13379), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15407 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13118), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15408 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13378), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15409 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13119), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15410 ( .A(n13120), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13130), .Z(
        P3_U3514) );
  MUX2_X1 U15411 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13440), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15412 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13470), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15413 ( .A(n13488), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13130), .Z(
        P3_U3510) );
  MUX2_X1 U15414 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13469), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15415 ( .A(n13487), .B(P3_DATAO_REG_17__SCAN_IN), .S(n13130), .Z(
        P3_U3508) );
  MUX2_X1 U15416 ( .A(n13498), .B(P3_DATAO_REG_16__SCAN_IN), .S(n13130), .Z(
        P3_U3507) );
  MUX2_X1 U15417 ( .A(n13538), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13130), .Z(
        P3_U3506) );
  MUX2_X1 U15418 ( .A(n13121), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13130), .Z(
        P3_U3505) );
  MUX2_X1 U15419 ( .A(n13537), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13130), .Z(
        P3_U3504) );
  MUX2_X1 U15420 ( .A(n10479), .B(P3_DATAO_REG_12__SCAN_IN), .S(n13130), .Z(
        P3_U3503) );
  MUX2_X1 U15421 ( .A(n13122), .B(P3_DATAO_REG_10__SCAN_IN), .S(n13130), .Z(
        P3_U3501) );
  MUX2_X1 U15422 ( .A(n13123), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13130), .Z(
        P3_U3500) );
  MUX2_X1 U15423 ( .A(n13124), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13130), .Z(
        P3_U3498) );
  MUX2_X1 U15424 ( .A(n13125), .B(P3_DATAO_REG_6__SCAN_IN), .S(n13130), .Z(
        P3_U3497) );
  MUX2_X1 U15425 ( .A(n13126), .B(P3_DATAO_REG_5__SCAN_IN), .S(n13130), .Z(
        P3_U3496) );
  MUX2_X1 U15426 ( .A(n13127), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13130), .Z(
        P3_U3495) );
  MUX2_X1 U15427 ( .A(n13128), .B(P3_DATAO_REG_3__SCAN_IN), .S(n13130), .Z(
        P3_U3494) );
  MUX2_X1 U15428 ( .A(n15536), .B(P3_DATAO_REG_2__SCAN_IN), .S(n13130), .Z(
        P3_U3493) );
  MUX2_X1 U15429 ( .A(n13129), .B(P3_DATAO_REG_1__SCAN_IN), .S(n13130), .Z(
        P3_U3492) );
  MUX2_X1 U15430 ( .A(n15534), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13130), .Z(
        P3_U3491) );
  NAND2_X1 U15431 ( .A1(n13132), .A2(n13131), .ZN(n13134) );
  NAND2_X1 U15432 ( .A1(n13140), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n13133) );
  NAND2_X1 U15433 ( .A1(n13134), .A2(n13133), .ZN(n13156) );
  INV_X1 U15434 ( .A(n13155), .ZN(n13170) );
  XNOR2_X1 U15435 ( .A(n13156), .B(n13170), .ZN(n13154) );
  XOR2_X1 U15436 ( .A(P3_REG1_REG_11__SCAN_IN), .B(n13154), .Z(n13152) );
  MUX2_X1 U15437 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13703), .Z(n13168) );
  XOR2_X1 U15438 ( .A(n13168), .B(n13155), .Z(n13171) );
  XNOR2_X1 U15439 ( .A(n13172), .B(n13171), .ZN(n13150) );
  NAND2_X1 U15440 ( .A1(n15503), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n13138) );
  OAI211_X1 U15441 ( .C1(n13314), .C2(n13155), .A(n13139), .B(n13138), .ZN(
        n13149) );
  INV_X1 U15442 ( .A(n13140), .ZN(n13143) );
  NAND2_X1 U15443 ( .A1(n13146), .A2(n13145), .ZN(n13147) );
  AOI21_X1 U15444 ( .B1(n13163), .B2(n13147), .A(n13164), .ZN(n13148) );
  AOI211_X1 U15445 ( .C1(n13329), .C2(n13150), .A(n13149), .B(n13148), .ZN(
        n13151) );
  OAI21_X1 U15446 ( .B1(n13152), .B2(n13283), .A(n13151), .ZN(P3_U3193) );
  XNOR2_X1 U15447 ( .A(n13180), .B(n13153), .ZN(n13178) );
  NAND2_X1 U15448 ( .A1(n13154), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n13158) );
  NAND2_X1 U15449 ( .A1(n13156), .A2(n13155), .ZN(n13157) );
  NAND2_X1 U15450 ( .A1(n13158), .A2(n13157), .ZN(n13179) );
  XOR2_X1 U15451 ( .A(n13178), .B(n13179), .Z(n13177) );
  OAI21_X1 U15452 ( .B1(n13291), .B2(n13160), .A(n13159), .ZN(n13167) );
  XNOR2_X1 U15453 ( .A(n13180), .B(P3_REG2_REG_12__SCAN_IN), .ZN(n13162) );
  NAND3_X1 U15454 ( .A1(n13163), .A2(n13162), .A3(n13161), .ZN(n13165) );
  AOI21_X1 U15455 ( .B1(n13182), .B2(n13165), .A(n13164), .ZN(n13166) );
  AOI211_X1 U15456 ( .C1(n13293), .C2(n13189), .A(n13167), .B(n13166), .ZN(
        n13176) );
  INV_X1 U15457 ( .A(n13168), .ZN(n13169) );
  MUX2_X1 U15458 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13703), .Z(n13186) );
  XNOR2_X1 U15459 ( .A(n13186), .B(n13189), .ZN(n13173) );
  OAI211_X1 U15460 ( .C1(n13174), .C2(n13173), .A(n13187), .B(n13329), .ZN(
        n13175) );
  OAI211_X1 U15461 ( .C1(n13177), .C2(n13283), .A(n13176), .B(n13175), .ZN(
        P3_U3194) );
  XOR2_X1 U15462 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n13202), .Z(n13199) );
  NAND2_X1 U15463 ( .A1(n13180), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13181) );
  OAI21_X1 U15464 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n13185), .A(n13208), 
        .ZN(n13197) );
  MUX2_X1 U15465 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13703), .Z(n13210) );
  XOR2_X1 U15466 ( .A(n13210), .B(n13213), .Z(n13191) );
  INV_X1 U15467 ( .A(n13186), .ZN(n13188) );
  OAI21_X1 U15468 ( .B1(n13189), .B2(n13188), .A(n13187), .ZN(n13190) );
  AOI21_X1 U15469 ( .B1(n13191), .B2(n13190), .A(n13211), .ZN(n13195) );
  INV_X1 U15470 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15161) );
  OAI21_X1 U15471 ( .B1(n13291), .B2(n15161), .A(n13192), .ZN(n13193) );
  AOI21_X1 U15472 ( .B1(n13213), .B2(n13293), .A(n13193), .ZN(n13194) );
  OAI21_X1 U15473 ( .B1(n13195), .B2(n13303), .A(n13194), .ZN(n13196) );
  AOI21_X1 U15474 ( .B1(n13197), .B2(n13311), .A(n13196), .ZN(n13198) );
  OAI21_X1 U15475 ( .B1(n13199), .B2(n13283), .A(n13198), .ZN(P3_U3195) );
  NOR2_X1 U15476 ( .A1(n13200), .A2(n13213), .ZN(n13201) );
  OR2_X1 U15477 ( .A1(n13221), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13203) );
  NAND2_X1 U15478 ( .A1(n13221), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13231) );
  AND2_X1 U15479 ( .A1(n13203), .A2(n13231), .ZN(n13226) );
  XNOR2_X1 U15480 ( .A(n13227), .B(n13226), .ZN(n13225) );
  NAND2_X1 U15481 ( .A1(n13208), .A2(n13206), .ZN(n13205) );
  OR2_X1 U15482 ( .A1(n13221), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13204) );
  NAND2_X1 U15483 ( .A1(n13221), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13232) );
  AND2_X1 U15484 ( .A1(n13204), .A2(n13232), .ZN(n13215) );
  NAND2_X1 U15485 ( .A1(n13205), .A2(n13215), .ZN(n13228) );
  INV_X1 U15486 ( .A(n13215), .ZN(n13207) );
  NAND3_X1 U15487 ( .A1(n13208), .A2(n13207), .A3(n13206), .ZN(n13209) );
  NAND2_X1 U15488 ( .A1(n13228), .A2(n13209), .ZN(n13223) );
  INV_X1 U15489 ( .A(n13210), .ZN(n13212) );
  MUX2_X1 U15490 ( .A(n13226), .B(n13215), .S(n13214), .Z(n13216) );
  OAI211_X1 U15491 ( .C1(n13217), .C2(n13216), .A(n13234), .B(n13329), .ZN(
        n13220) );
  AOI21_X1 U15492 ( .B1(n15503), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13218), 
        .ZN(n13219) );
  OAI211_X1 U15493 ( .C1(n13314), .C2(n13221), .A(n13220), .B(n13219), .ZN(
        n13222) );
  AOI21_X1 U15494 ( .B1(n13223), .B2(n13311), .A(n13222), .ZN(n13224) );
  OAI21_X1 U15495 ( .B1(n13283), .B2(n13225), .A(n13224), .ZN(P3_U3196) );
  XNOR2_X1 U15496 ( .A(n13248), .B(P3_REG1_REG_15__SCAN_IN), .ZN(n13243) );
  NAND2_X1 U15497 ( .A1(n13228), .A2(n13232), .ZN(n13229) );
  OAI21_X1 U15498 ( .B1(P3_REG2_REG_15__SCAN_IN), .B2(n13230), .A(n13250), 
        .ZN(n13241) );
  MUX2_X1 U15499 ( .A(n13232), .B(n13231), .S(n13703), .Z(n13233) );
  INV_X1 U15500 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15643) );
  INV_X1 U15501 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13247) );
  MUX2_X1 U15502 ( .A(n15643), .B(n13247), .S(n13703), .Z(n13235) );
  AOI211_X1 U15503 ( .C1(n13236), .C2(n13235), .A(n13303), .B(n13257), .ZN(
        n13240) );
  NAND2_X1 U15504 ( .A1(n15503), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n13237) );
  OAI211_X1 U15505 ( .C1(n13314), .C2(n7411), .A(n13238), .B(n13237), .ZN(
        n13239) );
  AOI211_X1 U15506 ( .C1(n13241), .C2(n13311), .A(n13240), .B(n13239), .ZN(
        n13242) );
  OAI21_X1 U15507 ( .B1(n13243), .B2(n13283), .A(n13242), .ZN(P3_U3197) );
  XNOR2_X1 U15508 ( .A(n13259), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13266) );
  INV_X1 U15509 ( .A(n13244), .ZN(n13245) );
  XOR2_X1 U15510 ( .A(n13266), .B(n13267), .Z(n13265) );
  INV_X1 U15511 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13249) );
  NOR2_X1 U15512 ( .A1(n13259), .A2(n13249), .ZN(n13268) );
  AOI21_X1 U15513 ( .B1(n13259), .B2(n13249), .A(n13268), .ZN(n13252) );
  NAND2_X1 U15514 ( .A1(n13251), .A2(n13252), .ZN(n13270) );
  OAI21_X1 U15515 ( .B1(n13252), .B2(n13251), .A(n13270), .ZN(n13256) );
  NAND2_X1 U15516 ( .A1(n15503), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n13253) );
  OAI211_X1 U15517 ( .C1(n13314), .C2(n13274), .A(n13254), .B(n13253), .ZN(
        n13255) );
  AOI21_X1 U15518 ( .B1(n13256), .B2(n13311), .A(n13255), .ZN(n13264) );
  MUX2_X1 U15519 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13703), .Z(n13275) );
  XNOR2_X1 U15520 ( .A(n13275), .B(n13259), .ZN(n13260) );
  OAI21_X1 U15521 ( .B1(n13261), .B2(n13260), .A(n13273), .ZN(n13262) );
  NAND2_X1 U15522 ( .A1(n13262), .A2(n13329), .ZN(n13263) );
  OAI211_X1 U15523 ( .C1(n13265), .C2(n13283), .A(n13264), .B(n13263), .ZN(
        P3_U3198) );
  XNOR2_X1 U15524 ( .A(n13294), .B(n13295), .ZN(n13296) );
  XNOR2_X1 U15525 ( .A(n13296), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n13284) );
  INV_X1 U15526 ( .A(n13268), .ZN(n13269) );
  INV_X1 U15527 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13503) );
  MUX2_X1 U15528 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13703), .Z(n13300) );
  XOR2_X1 U15529 ( .A(n13300), .B(n13295), .Z(n13277) );
  AOI211_X1 U15530 ( .C1(n13277), .C2(n13276), .A(n13303), .B(n13298), .ZN(
        n13281) );
  AOI21_X1 U15531 ( .B1(n15503), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13278), 
        .ZN(n13279) );
  OAI21_X1 U15532 ( .B1(n13314), .B2(n13299), .A(n13279), .ZN(n13280) );
  OAI21_X1 U15533 ( .B1(n13284), .B2(n13283), .A(n13282), .ZN(P3_U3199) );
  INV_X1 U15534 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13480) );
  OR2_X1 U15535 ( .A1(n13324), .A2(n13480), .ZN(n13308) );
  NAND2_X1 U15536 ( .A1(n13324), .A2(n13480), .ZN(n13285) );
  NAND2_X1 U15537 ( .A1(n13308), .A2(n13285), .ZN(n13286) );
  INV_X1 U15538 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15220) );
  OAI21_X1 U15539 ( .B1(n13291), .B2(n15220), .A(n13290), .ZN(n13292) );
  AOI21_X1 U15540 ( .B1(n13324), .B2(n13293), .A(n13292), .ZN(n13307) );
  INV_X1 U15541 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n15734) );
  XNOR2_X1 U15542 ( .A(n13324), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n13318) );
  XNOR2_X1 U15543 ( .A(n13319), .B(n13318), .ZN(n13297) );
  NAND2_X1 U15544 ( .A1(n13297), .A2(n13322), .ZN(n13306) );
  MUX2_X1 U15545 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13703), .Z(n13302) );
  XNOR2_X1 U15546 ( .A(n13325), .B(n13324), .ZN(n13301) );
  AOI21_X1 U15547 ( .B1(n13302), .B2(n13301), .A(n13323), .ZN(n13304) );
  OR2_X1 U15548 ( .A1(n13304), .A2(n13303), .ZN(n13305) );
  INV_X1 U15549 ( .A(n13308), .ZN(n13309) );
  NOR2_X1 U15550 ( .A1(n13314), .A2(n13313), .ZN(n13315) );
  AOI211_X1 U15551 ( .C1(P3_ADDR_REG_19__SCAN_IN), .C2(n15503), .A(n13316), 
        .B(n13315), .ZN(n13332) );
  XNOR2_X1 U15552 ( .A(n13321), .B(n13320), .ZN(n13326) );
  MUX2_X1 U15553 ( .A(n6624), .B(n13326), .S(n13703), .Z(n13327) );
  XNOR2_X1 U15554 ( .A(n13328), .B(n13327), .ZN(n13330) );
  NAND2_X1 U15555 ( .A1(n13330), .A2(n13329), .ZN(n13331) );
  NAND2_X1 U15556 ( .A1(n15549), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13337) );
  INV_X1 U15557 ( .A(n13333), .ZN(n13334) );
  NOR2_X1 U15558 ( .A1(n13336), .A2(n15509), .ZN(n13342) );
  OAI21_X1 U15559 ( .B1(n13602), .B2(n13342), .A(n15524), .ZN(n13338) );
  OAI211_X1 U15560 ( .C1(n13604), .C2(n13534), .A(n13337), .B(n13338), .ZN(
        P3_U3202) );
  NAND2_X1 U15561 ( .A1(n15549), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13339) );
  OAI211_X1 U15562 ( .C1(n13607), .C2(n13534), .A(n13339), .B(n13338), .ZN(
        P3_U3203) );
  NOR2_X1 U15563 ( .A1(n13340), .A2(n13534), .ZN(n13341) );
  AOI211_X1 U15564 ( .C1(n15549), .C2(P3_REG2_REG_29__SCAN_IN), .A(n13342), 
        .B(n13341), .ZN(n13345) );
  OR2_X1 U15565 ( .A1(n13343), .A2(n15549), .ZN(n13344) );
  OAI211_X1 U15566 ( .C1(n13346), .C2(n13529), .A(n13345), .B(n13344), .ZN(
        P3_U3204) );
  NAND2_X1 U15567 ( .A1(n6463), .A2(n13347), .ZN(n13348) );
  XNOR2_X1 U15568 ( .A(n13348), .B(n13350), .ZN(n13609) );
  AOI22_X1 U15569 ( .A1(n13548), .A2(n13519), .B1(n15544), .B2(n13349), .ZN(
        n13358) );
  OAI21_X1 U15570 ( .B1(n13351), .B2(n13350), .A(n15532), .ZN(n13353) );
  AOI22_X1 U15571 ( .A1(n13379), .A2(n15535), .B1(n13354), .B2(n15537), .ZN(
        n13355) );
  MUX2_X1 U15572 ( .A(n13610), .B(P3_REG2_REG_28__SCAN_IN), .S(n15549), .Z(
        n13356) );
  INV_X1 U15573 ( .A(n13356), .ZN(n13357) );
  OAI211_X1 U15574 ( .C1(n13609), .C2(n13529), .A(n13358), .B(n13357), .ZN(
        P3_U3205) );
  INV_X1 U15575 ( .A(n13359), .ZN(n13360) );
  OAI22_X1 U15576 ( .A1(n13362), .A2(n15513), .B1(n13387), .B2(n15516), .ZN(
        n13363) );
  AOI22_X1 U15577 ( .A1(n13364), .A2(n15544), .B1(n15549), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13365) );
  OAI21_X1 U15578 ( .B1(n13366), .B2(n13534), .A(n13365), .ZN(n13367) );
  AOI21_X1 U15579 ( .B1(n13551), .B2(n15545), .A(n13367), .ZN(n13368) );
  OAI21_X1 U15580 ( .B1(n13554), .B2(n15549), .A(n13368), .ZN(P3_U3206) );
  INV_X1 U15581 ( .A(n13369), .ZN(n13371) );
  OAI21_X1 U15582 ( .B1(n13414), .B2(n13371), .A(n13370), .ZN(n13373) );
  NAND2_X1 U15583 ( .A1(n13373), .A2(n13372), .ZN(n13374) );
  XNOR2_X1 U15584 ( .A(n13374), .B(n13376), .ZN(n13618) );
  AOI22_X1 U15585 ( .A1(n13615), .A2(n13519), .B1(n15544), .B2(n13375), .ZN(
        n13382) );
  INV_X1 U15586 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n13380) );
  MUX2_X1 U15587 ( .A(n13380), .B(n13613), .S(n15524), .Z(n13381) );
  OAI211_X1 U15588 ( .C1(n13618), .C2(n13529), .A(n13382), .B(n13381), .ZN(
        P3_U3207) );
  NAND3_X1 U15589 ( .A1(n13413), .A2(n13401), .A3(n13398), .ZN(n13397) );
  NAND2_X1 U15590 ( .A1(n13397), .A2(n13383), .ZN(n13384) );
  XNOR2_X1 U15591 ( .A(n13384), .B(n13386), .ZN(n13391) );
  XOR2_X1 U15592 ( .A(n13386), .B(n13385), .Z(n13389) );
  OAI22_X1 U15593 ( .A1(n13387), .A2(n15513), .B1(n13419), .B2(n15516), .ZN(
        n13388) );
  AOI21_X1 U15594 ( .B1(n13389), .B2(n15532), .A(n13388), .ZN(n13390) );
  INV_X1 U15595 ( .A(n13560), .ZN(n13396) );
  INV_X1 U15596 ( .A(n13391), .ZN(n13561) );
  AOI22_X1 U15597 ( .A1(n13392), .A2(n15544), .B1(n15549), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13393) );
  OAI21_X1 U15598 ( .B1(n13622), .B2(n13534), .A(n13393), .ZN(n13394) );
  AOI21_X1 U15599 ( .B1(n13561), .B2(n15545), .A(n13394), .ZN(n13395) );
  OAI21_X1 U15600 ( .B1(n13396), .B2(n15549), .A(n13395), .ZN(P3_U3208) );
  INV_X1 U15601 ( .A(n13397), .ZN(n13400) );
  AOI21_X1 U15602 ( .B1(n13413), .B2(n13398), .A(n13401), .ZN(n13399) );
  NOR2_X1 U15603 ( .A1(n13400), .A2(n13399), .ZN(n13626) );
  XNOR2_X1 U15604 ( .A(n13402), .B(n13401), .ZN(n13403) );
  NAND2_X1 U15605 ( .A1(n13403), .A2(n15532), .ZN(n13407) );
  OAI22_X1 U15606 ( .A1(n13404), .A2(n15513), .B1(n13431), .B2(n15516), .ZN(
        n13405) );
  INV_X1 U15607 ( .A(n13405), .ZN(n13406) );
  NAND2_X1 U15608 ( .A1(n13407), .A2(n13406), .ZN(n13564) );
  NAND2_X1 U15609 ( .A1(n13565), .A2(n13519), .ZN(n13410) );
  AOI22_X1 U15610 ( .A1(n13408), .A2(n15544), .B1(n15549), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13409) );
  NAND2_X1 U15611 ( .A1(n13410), .A2(n13409), .ZN(n13411) );
  AOI21_X1 U15612 ( .B1(n13564), .B2(n15524), .A(n13411), .ZN(n13412) );
  OAI21_X1 U15613 ( .B1(n13626), .B2(n13529), .A(n13412), .ZN(P3_U3209) );
  OAI21_X1 U15614 ( .B1(n13414), .B2(n13416), .A(n13413), .ZN(n13632) );
  AOI22_X1 U15615 ( .A1(n13630), .A2(n13519), .B1(n15544), .B2(n13415), .ZN(
        n13425) );
  INV_X1 U15616 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13423) );
  AOI21_X1 U15617 ( .B1(n13417), .B2(n13416), .A(n13522), .ZN(n13422) );
  OAI22_X1 U15618 ( .A1(n13419), .A2(n15513), .B1(n13418), .B2(n15516), .ZN(
        n13420) );
  AOI21_X1 U15619 ( .B1(n13422), .B2(n13421), .A(n13420), .ZN(n13627) );
  MUX2_X1 U15620 ( .A(n13423), .B(n13627), .S(n15524), .Z(n13424) );
  OAI211_X1 U15621 ( .C1(n13632), .C2(n13529), .A(n13425), .B(n13424), .ZN(
        P3_U3210) );
  XNOR2_X1 U15622 ( .A(n13426), .B(n13428), .ZN(n13637) );
  AOI22_X1 U15623 ( .A1(n13635), .A2(n13519), .B1(n15544), .B2(n13427), .ZN(
        n13435) );
  INV_X1 U15624 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13433) );
  XNOR2_X1 U15625 ( .A(n13429), .B(n13428), .ZN(n13430) );
  OAI222_X1 U15626 ( .A1(n15516), .A2(n13454), .B1(n15513), .B2(n13431), .C1(
        n13430), .C2(n13522), .ZN(n13633) );
  INV_X1 U15627 ( .A(n13633), .ZN(n13432) );
  MUX2_X1 U15628 ( .A(n13433), .B(n13432), .S(n15524), .Z(n13434) );
  OAI211_X1 U15629 ( .C1(n13637), .C2(n13529), .A(n13435), .B(n13434), .ZN(
        P3_U3211) );
  XNOR2_X1 U15630 ( .A(n13436), .B(n13438), .ZN(n13643) );
  AOI22_X1 U15631 ( .A1(n13641), .A2(n13519), .B1(n15544), .B2(n13437), .ZN(
        n13444) );
  INV_X1 U15632 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13442) );
  XNOR2_X1 U15633 ( .A(n13439), .B(n13438), .ZN(n13441) );
  AOI222_X1 U15634 ( .A1(n15532), .A2(n13441), .B1(n13440), .B2(n15537), .C1(
        n13470), .C2(n15535), .ZN(n13638) );
  MUX2_X1 U15635 ( .A(n13442), .B(n13638), .S(n15524), .Z(n13443) );
  OAI211_X1 U15636 ( .C1(n13643), .C2(n13529), .A(n13444), .B(n13443), .ZN(
        P3_U3212) );
  OAI21_X1 U15637 ( .B1(n13447), .B2(n13446), .A(n13445), .ZN(n13648) );
  AOI22_X1 U15638 ( .A1(n13646), .A2(n13519), .B1(n15544), .B2(n13448), .ZN(
        n13458) );
  INV_X1 U15639 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13456) );
  OAI211_X1 U15640 ( .C1(n13451), .C2(n13450), .A(n13449), .B(n15532), .ZN(
        n13453) );
  NAND2_X1 U15641 ( .A1(n13488), .A2(n15535), .ZN(n13452) );
  OAI211_X1 U15642 ( .C1(n13454), .C2(n15513), .A(n13453), .B(n13452), .ZN(
        n13644) );
  INV_X1 U15643 ( .A(n13644), .ZN(n13455) );
  MUX2_X1 U15644 ( .A(n13456), .B(n13455), .S(n15524), .Z(n13457) );
  OAI211_X1 U15645 ( .C1(n13648), .C2(n13529), .A(n13458), .B(n13457), .ZN(
        P3_U3213) );
  NAND2_X1 U15646 ( .A1(n6668), .A2(n13459), .ZN(n13461) );
  XNOR2_X1 U15647 ( .A(n13461), .B(n13460), .ZN(n13653) );
  NOR2_X1 U15648 ( .A1(n13462), .A2(n13534), .ZN(n13474) );
  INV_X1 U15649 ( .A(n13464), .ZN(n13466) );
  AOI21_X1 U15650 ( .B1(n13463), .B2(n13466), .A(n13465), .ZN(n13468) );
  XNOR2_X1 U15651 ( .A(n13468), .B(n13467), .ZN(n13472) );
  AOI22_X1 U15652 ( .A1(n13470), .A2(n15537), .B1(n15535), .B2(n13469), .ZN(
        n13471) );
  OAI21_X1 U15653 ( .B1(n13472), .B2(n13522), .A(n13471), .ZN(n13649) );
  MUX2_X1 U15654 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n13649), .S(n15524), .Z(
        n13473) );
  AOI211_X1 U15655 ( .C1(n15544), .C2(n13475), .A(n13474), .B(n13473), .ZN(
        n13476) );
  OAI21_X1 U15656 ( .B1(n13653), .B2(n13529), .A(n13476), .ZN(P3_U3214) );
  OAI21_X1 U15657 ( .B1(n13478), .B2(n13484), .A(n6668), .ZN(n13657) );
  OAI22_X1 U15658 ( .A1(n15524), .A2(n13480), .B1(n13479), .B2(n15509), .ZN(
        n13481) );
  AOI21_X1 U15659 ( .B1(n13580), .B2(n13519), .A(n13481), .ZN(n13492) );
  OR2_X1 U15660 ( .A1(n13463), .A2(n13482), .ZN(n13495) );
  NAND2_X1 U15661 ( .A1(n13495), .A2(n13483), .ZN(n13485) );
  XNOR2_X1 U15662 ( .A(n13485), .B(n13484), .ZN(n13486) );
  NAND2_X1 U15663 ( .A1(n13486), .A2(n15532), .ZN(n13490) );
  AOI22_X1 U15664 ( .A1(n13488), .A2(n15537), .B1(n15535), .B2(n13487), .ZN(
        n13489) );
  NAND2_X1 U15665 ( .A1(n13490), .A2(n13489), .ZN(n13579) );
  NAND2_X1 U15666 ( .A1(n13579), .A2(n15524), .ZN(n13491) );
  OAI211_X1 U15667 ( .C1(n13657), .C2(n13529), .A(n13492), .B(n13491), .ZN(
        P3_U3215) );
  XNOR2_X1 U15668 ( .A(n13493), .B(n13496), .ZN(n13662) );
  AOI22_X1 U15669 ( .A1(n13660), .A2(n13519), .B1(n15544), .B2(n13494), .ZN(
        n13505) );
  INV_X1 U15670 ( .A(n13463), .ZN(n13497) );
  OAI211_X1 U15671 ( .C1(n13497), .C2(n13496), .A(n15532), .B(n13495), .ZN(
        n13500) );
  NAND2_X1 U15672 ( .A1(n15535), .A2(n13498), .ZN(n13499) );
  OAI211_X1 U15673 ( .C1(n13501), .C2(n15513), .A(n13500), .B(n13499), .ZN(
        n13658) );
  INV_X1 U15674 ( .A(n13658), .ZN(n13502) );
  MUX2_X1 U15675 ( .A(n13503), .B(n13502), .S(n15524), .Z(n13504) );
  OAI211_X1 U15676 ( .C1(n13662), .C2(n13529), .A(n13505), .B(n13504), .ZN(
        P3_U3216) );
  XNOR2_X1 U15677 ( .A(n13506), .B(n7624), .ZN(n13666) );
  XNOR2_X1 U15678 ( .A(n13508), .B(n13507), .ZN(n13509) );
  OAI222_X1 U15679 ( .A1(n15513), .A2(n13511), .B1(n15516), .B2(n13510), .C1(
        n13522), .C2(n13509), .ZN(n13584) );
  AOI22_X1 U15680 ( .A1(n15549), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15544), 
        .B2(n13512), .ZN(n13513) );
  OAI21_X1 U15681 ( .B1(n13514), .B2(n13534), .A(n13513), .ZN(n13515) );
  AOI21_X1 U15682 ( .B1(n13584), .B2(n15524), .A(n13515), .ZN(n13516) );
  OAI21_X1 U15683 ( .B1(n13666), .B2(n13529), .A(n13516), .ZN(P3_U3217) );
  XNOR2_X1 U15684 ( .A(n13517), .B(n13520), .ZN(n13672) );
  AOI22_X1 U15685 ( .A1(n13519), .A2(n13669), .B1(n15544), .B2(n13518), .ZN(
        n13528) );
  XNOR2_X1 U15686 ( .A(n13521), .B(n13520), .ZN(n13523) );
  OAI222_X1 U15687 ( .A1(n15513), .A2(n13525), .B1(n15516), .B2(n13524), .C1(
        n13523), .C2(n13522), .ZN(n13667) );
  INV_X1 U15688 ( .A(n13667), .ZN(n13526) );
  MUX2_X1 U15689 ( .A(n15643), .B(n13526), .S(n15524), .Z(n13527) );
  OAI211_X1 U15690 ( .C1(n13672), .C2(n13529), .A(n13528), .B(n13527), .ZN(
        P3_U3218) );
  OAI21_X1 U15691 ( .B1(n13531), .B2(n13535), .A(n13530), .ZN(n13675) );
  INV_X1 U15692 ( .A(n13532), .ZN(n13533) );
  OAI22_X1 U15693 ( .A1(n13680), .A2(n13534), .B1(n13533), .B2(n15509), .ZN(
        n13542) );
  XNOR2_X1 U15694 ( .A(n13536), .B(n13535), .ZN(n13539) );
  AOI222_X1 U15695 ( .A1(n15532), .A2(n13539), .B1(n13538), .B2(n15537), .C1(
        n13537), .C2(n15535), .ZN(n13676) );
  INV_X1 U15696 ( .A(n13676), .ZN(n13540) );
  MUX2_X1 U15697 ( .A(P3_REG2_REG_14__SCAN_IN), .B(n13540), .S(n15524), .Z(
        n13541) );
  AOI211_X1 U15698 ( .C1(n13543), .C2(n13675), .A(n13542), .B(n13541), .ZN(
        n13544) );
  INV_X1 U15699 ( .A(n13544), .ZN(P3_U3219) );
  NAND2_X1 U15700 ( .A1(n15593), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13545) );
  NAND2_X1 U15701 ( .A1(n13602), .A2(n15595), .ZN(n13547) );
  OAI211_X1 U15702 ( .C1(n13604), .C2(n13597), .A(n13545), .B(n13547), .ZN(
        P3_U3490) );
  NAND2_X1 U15703 ( .A1(n15593), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13546) );
  OAI211_X1 U15704 ( .C1(n13607), .C2(n13597), .A(n13547), .B(n13546), .ZN(
        P3_U3489) );
  INV_X1 U15705 ( .A(n13548), .ZN(n13608) );
  OAI22_X1 U15706 ( .A1(n13609), .A2(n13592), .B1(n13608), .B2(n13597), .ZN(
        n13550) );
  MUX2_X1 U15707 ( .A(n13610), .B(P3_REG1_REG_28__SCAN_IN), .S(n15593), .Z(
        n13549) );
  OR2_X1 U15708 ( .A1(n13550), .A2(n13549), .ZN(P3_U3487) );
  INV_X1 U15709 ( .A(n13551), .ZN(n13556) );
  NAND2_X1 U15710 ( .A1(n13552), .A2(n13586), .ZN(n13553) );
  MUX2_X1 U15711 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13612), .S(n15595), .Z(
        P3_U3486) );
  MUX2_X1 U15712 ( .A(n13557), .B(n13613), .S(n15595), .Z(n13559) );
  NAND2_X1 U15713 ( .A1(n13615), .A2(n13590), .ZN(n13558) );
  OAI211_X1 U15714 ( .C1(n13618), .C2(n13592), .A(n13559), .B(n13558), .ZN(
        P3_U3485) );
  AOI21_X1 U15715 ( .B1(n15579), .B2(n13561), .A(n13560), .ZN(n13619) );
  MUX2_X1 U15716 ( .A(n13562), .B(n13619), .S(n15595), .Z(n13563) );
  INV_X1 U15717 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n15609) );
  AOI21_X1 U15718 ( .B1(n13586), .B2(n13565), .A(n13564), .ZN(n13623) );
  MUX2_X1 U15719 ( .A(n15609), .B(n13623), .S(n15595), .Z(n13566) );
  OAI21_X1 U15720 ( .B1(n13626), .B2(n13592), .A(n13566), .ZN(P3_U3483) );
  MUX2_X1 U15721 ( .A(n13567), .B(n13627), .S(n15595), .Z(n13569) );
  NAND2_X1 U15722 ( .A1(n13630), .A2(n13590), .ZN(n13568) );
  OAI211_X1 U15723 ( .C1(n13632), .C2(n13592), .A(n13569), .B(n13568), .ZN(
        P3_U3482) );
  MUX2_X1 U15724 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n13633), .S(n15595), .Z(
        n13570) );
  AOI21_X1 U15725 ( .B1(n13590), .B2(n13635), .A(n13570), .ZN(n13571) );
  OAI21_X1 U15726 ( .B1(n13637), .B2(n13592), .A(n13571), .ZN(P3_U3481) );
  MUX2_X1 U15727 ( .A(n13572), .B(n13638), .S(n15595), .Z(n13574) );
  NAND2_X1 U15728 ( .A1(n13641), .A2(n13590), .ZN(n13573) );
  OAI211_X1 U15729 ( .C1(n13643), .C2(n13592), .A(n13574), .B(n13573), .ZN(
        P3_U3480) );
  MUX2_X1 U15730 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13644), .S(n15595), .Z(
        n13575) );
  AOI21_X1 U15731 ( .B1(n13590), .B2(n13646), .A(n13575), .ZN(n13576) );
  OAI21_X1 U15732 ( .B1(n13648), .B2(n13592), .A(n13576), .ZN(P3_U3479) );
  MUX2_X1 U15733 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13649), .S(n15595), .Z(
        n13577) );
  AOI21_X1 U15734 ( .B1(n13590), .B2(n13651), .A(n13577), .ZN(n13578) );
  OAI21_X1 U15735 ( .B1(n13653), .B2(n13592), .A(n13578), .ZN(P3_U3478) );
  AOI21_X1 U15736 ( .B1(n13586), .B2(n13580), .A(n13579), .ZN(n13654) );
  MUX2_X1 U15737 ( .A(n7122), .B(n13654), .S(n15595), .Z(n13581) );
  OAI21_X1 U15738 ( .B1(n13657), .B2(n13592), .A(n13581), .ZN(P3_U3477) );
  MUX2_X1 U15739 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13658), .S(n15595), .Z(
        n13582) );
  AOI21_X1 U15740 ( .B1(n13590), .B2(n13660), .A(n13582), .ZN(n13583) );
  OAI21_X1 U15741 ( .B1(n13662), .B2(n13592), .A(n13583), .ZN(P3_U3476) );
  INV_X1 U15742 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13587) );
  AOI21_X1 U15743 ( .B1(n13586), .B2(n13585), .A(n13584), .ZN(n13663) );
  MUX2_X1 U15744 ( .A(n13587), .B(n13663), .S(n15595), .Z(n13588) );
  OAI21_X1 U15745 ( .B1(n13666), .B2(n13592), .A(n13588), .ZN(P3_U3475) );
  MUX2_X1 U15746 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13667), .S(n15595), .Z(
        n13589) );
  AOI21_X1 U15747 ( .B1(n13590), .B2(n13669), .A(n13589), .ZN(n13591) );
  OAI21_X1 U15748 ( .B1(n13672), .B2(n13592), .A(n13591), .ZN(P3_U3474) );
  INV_X1 U15749 ( .A(n13592), .ZN(n13593) );
  NAND2_X1 U15750 ( .A1(n13675), .A2(n13593), .ZN(n13596) );
  INV_X1 U15751 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13594) );
  MUX2_X1 U15752 ( .A(n13594), .B(n13676), .S(n15595), .Z(n13595) );
  OAI211_X1 U15753 ( .C1(n13597), .C2(n13680), .A(n13596), .B(n13595), .ZN(
        P3_U3473) );
  NAND2_X1 U15754 ( .A1(n13598), .A2(n15569), .ZN(n13600) );
  OAI211_X1 U15755 ( .C1(n13601), .C2(n15567), .A(n13600), .B(n13599), .ZN(
        n13682) );
  MUX2_X1 U15756 ( .A(P3_REG1_REG_11__SCAN_IN), .B(n13682), .S(n15595), .Z(
        P3_U3470) );
  NAND2_X1 U15757 ( .A1(n15583), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13603) );
  NAND2_X1 U15758 ( .A1(n13602), .A2(n15585), .ZN(n13606) );
  OAI211_X1 U15759 ( .C1(n13604), .C2(n13681), .A(n13603), .B(n13606), .ZN(
        P3_U3458) );
  NAND2_X1 U15760 ( .A1(n15583), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13605) );
  OAI211_X1 U15761 ( .C1(n13607), .C2(n13681), .A(n13606), .B(n13605), .ZN(
        P3_U3457) );
  OAI22_X1 U15762 ( .A1(n13609), .A2(n13673), .B1(n13608), .B2(n13681), .ZN(
        n13611) );
  MUX2_X1 U15763 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13612), .S(n15585), .Z(
        P3_U3454) );
  INV_X1 U15764 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13614) );
  MUX2_X1 U15765 ( .A(n13614), .B(n13613), .S(n15585), .Z(n13617) );
  NAND2_X1 U15766 ( .A1(n13615), .A2(n13670), .ZN(n13616) );
  OAI211_X1 U15767 ( .C1(n13618), .C2(n13673), .A(n13617), .B(n13616), .ZN(
        P3_U3453) );
  INV_X1 U15768 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13620) );
  MUX2_X1 U15769 ( .A(n13620), .B(n13619), .S(n15585), .Z(n13621) );
  OAI21_X1 U15770 ( .B1(n13622), .B2(n13681), .A(n13621), .ZN(P3_U3452) );
  INV_X1 U15771 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13624) );
  MUX2_X1 U15772 ( .A(n13624), .B(n13623), .S(n15585), .Z(n13625) );
  OAI21_X1 U15773 ( .B1(n13626), .B2(n13673), .A(n13625), .ZN(P3_U3451) );
  INV_X1 U15774 ( .A(n13627), .ZN(n13628) );
  MUX2_X1 U15775 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13628), .S(n15585), .Z(
        n13629) );
  AOI21_X1 U15776 ( .B1(n13670), .B2(n13630), .A(n13629), .ZN(n13631) );
  OAI21_X1 U15777 ( .B1(n13632), .B2(n13673), .A(n13631), .ZN(P3_U3450) );
  MUX2_X1 U15778 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n13633), .S(n15585), .Z(
        n13634) );
  AOI21_X1 U15779 ( .B1(n13670), .B2(n13635), .A(n13634), .ZN(n13636) );
  OAI21_X1 U15780 ( .B1(n13637), .B2(n13673), .A(n13636), .ZN(P3_U3449) );
  INV_X1 U15781 ( .A(n13638), .ZN(n13639) );
  MUX2_X1 U15782 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n13639), .S(n15585), .Z(
        n13640) );
  AOI21_X1 U15783 ( .B1(n13670), .B2(n13641), .A(n13640), .ZN(n13642) );
  OAI21_X1 U15784 ( .B1(n13643), .B2(n13673), .A(n13642), .ZN(P3_U3448) );
  MUX2_X1 U15785 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13644), .S(n15585), .Z(
        n13645) );
  AOI21_X1 U15786 ( .B1(n13670), .B2(n13646), .A(n13645), .ZN(n13647) );
  OAI21_X1 U15787 ( .B1(n13648), .B2(n13673), .A(n13647), .ZN(P3_U3447) );
  MUX2_X1 U15788 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13649), .S(n15585), .Z(
        n13650) );
  AOI21_X1 U15789 ( .B1(n13670), .B2(n13651), .A(n13650), .ZN(n13652) );
  OAI21_X1 U15790 ( .B1(n13653), .B2(n13673), .A(n13652), .ZN(P3_U3446) );
  INV_X1 U15791 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13655) );
  MUX2_X1 U15792 ( .A(n13655), .B(n13654), .S(n15585), .Z(n13656) );
  OAI21_X1 U15793 ( .B1(n13657), .B2(n13673), .A(n13656), .ZN(P3_U3444) );
  MUX2_X1 U15794 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13658), .S(n15585), .Z(
        n13659) );
  AOI21_X1 U15795 ( .B1(n13670), .B2(n13660), .A(n13659), .ZN(n13661) );
  OAI21_X1 U15796 ( .B1(n13662), .B2(n13673), .A(n13661), .ZN(P3_U3441) );
  INV_X1 U15797 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13664) );
  MUX2_X1 U15798 ( .A(n13664), .B(n13663), .S(n15585), .Z(n13665) );
  OAI21_X1 U15799 ( .B1(n13666), .B2(n13673), .A(n13665), .ZN(P3_U3438) );
  MUX2_X1 U15800 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13667), .S(n15585), .Z(
        n13668) );
  AOI21_X1 U15801 ( .B1(n13670), .B2(n13669), .A(n13668), .ZN(n13671) );
  OAI21_X1 U15802 ( .B1(n13672), .B2(n13673), .A(n13671), .ZN(P3_U3435) );
  INV_X1 U15803 ( .A(n13673), .ZN(n13674) );
  NAND2_X1 U15804 ( .A1(n13675), .A2(n13674), .ZN(n13679) );
  INV_X1 U15805 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13677) );
  MUX2_X1 U15806 ( .A(n13677), .B(n13676), .S(n15585), .Z(n13678) );
  OAI211_X1 U15807 ( .C1(n13681), .C2(n13680), .A(n13679), .B(n13678), .ZN(
        P3_U3432) );
  MUX2_X1 U15808 ( .A(P3_REG0_REG_11__SCAN_IN), .B(n13682), .S(n15585), .Z(
        P3_U3423) );
  MUX2_X1 U15809 ( .A(n13684), .B(P3_D_REG_1__SCAN_IN), .S(n13683), .Z(
        P3_U3377) );
  INV_X1 U15810 ( .A(n13685), .ZN(n13690) );
  NOR4_X1 U15811 ( .A1(n13687), .A2(P3_IR_REG_30__SCAN_IN), .A3(n13686), .A4(
        P3_U3151), .ZN(n13688) );
  AOI21_X1 U15812 ( .B1(n6622), .B2(SI_31_), .A(n13688), .ZN(n13689) );
  OAI21_X1 U15813 ( .B1(n13690), .B2(n13707), .A(n13689), .ZN(P3_U3264) );
  INV_X1 U15814 ( .A(n13691), .ZN(n13692) );
  OAI222_X1 U15815 ( .A1(n13694), .A2(P3_U3151), .B1(n13705), .B2(n13693), 
        .C1(n13707), .C2(n13692), .ZN(P3_U3265) );
  INV_X1 U15816 ( .A(n13695), .ZN(n13696) );
  OAI222_X1 U15817 ( .A1(n13705), .A2(n15690), .B1(P3_U3151), .B2(n13697), 
        .C1(n13707), .C2(n13696), .ZN(P3_U3266) );
  INV_X1 U15818 ( .A(n13698), .ZN(n13700) );
  OAI222_X1 U15819 ( .A1(P3_U3151), .A2(n13701), .B1(n13707), .B2(n13700), 
        .C1(n13699), .C2(n13705), .ZN(P3_U3267) );
  INV_X1 U15820 ( .A(n13702), .ZN(n13706) );
  OAI222_X1 U15821 ( .A1(n13707), .A2(n13706), .B1(n13705), .B2(n13704), .C1(
        P3_U3151), .C2(n13703), .ZN(P3_U3268) );
  NOR2_X1 U15822 ( .A1(n13710), .A2(n13709), .ZN(n13711) );
  XNOR2_X1 U15823 ( .A(n13712), .B(n13711), .ZN(n13718) );
  OAI22_X1 U15824 ( .A1(n14057), .A2(n13891), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13713), .ZN(n13715) );
  NOR2_X1 U15825 ( .A1(n13800), .A2(n13912), .ZN(n13714) );
  AOI211_X1 U15826 ( .C1(n13909), .C2(n14050), .A(n13715), .B(n13714), .ZN(
        n13717) );
  NAND2_X1 U15827 ( .A1(n14298), .A2(n13926), .ZN(n13716) );
  INV_X1 U15828 ( .A(n13722), .ZN(n13721) );
  NOR2_X1 U15829 ( .A1(n13721), .A2(n13720), .ZN(n13864) );
  NAND2_X1 U15830 ( .A1(n13719), .A2(n13864), .ZN(n13863) );
  NAND2_X1 U15831 ( .A1(n13863), .A2(n13722), .ZN(n13726) );
  XNOR2_X1 U15832 ( .A(n13724), .B(n13723), .ZN(n13725) );
  XNOR2_X1 U15833 ( .A(n13726), .B(n13725), .ZN(n13733) );
  NAND2_X1 U15834 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n15431)
         );
  OAI21_X1 U15835 ( .B1(n13891), .B2(n13727), .A(n15431), .ZN(n13728) );
  AOI21_X1 U15836 ( .B1(n13909), .B2(n13938), .A(n13728), .ZN(n13729) );
  OAI21_X1 U15837 ( .B1(n13730), .B2(n13912), .A(n13729), .ZN(n13731) );
  AOI21_X1 U15838 ( .B1(n14377), .B2(n13926), .A(n13731), .ZN(n13732) );
  OAI21_X1 U15839 ( .B1(n13733), .B2(n13921), .A(n13732), .ZN(P2_U3187) );
  INV_X1 U15840 ( .A(n14122), .ZN(n14320) );
  INV_X1 U15841 ( .A(n13875), .ZN(n13735) );
  NOR2_X1 U15842 ( .A1(n13735), .A2(n13734), .ZN(n13871) );
  NOR2_X1 U15843 ( .A1(n13871), .A2(n13736), .ZN(n13738) );
  XNOR2_X1 U15844 ( .A(n13738), .B(n13737), .ZN(n13740) );
  AOI21_X1 U15845 ( .B1(n13740), .B2(n13741), .A(n13921), .ZN(n13739) );
  OAI21_X1 U15846 ( .B1(n13741), .B2(n13740), .A(n13739), .ZN(n13746) );
  INV_X1 U15847 ( .A(n13912), .ZN(n13902) );
  INV_X1 U15848 ( .A(n13742), .ZN(n14121) );
  AOI22_X1 U15849 ( .A1(n13917), .A2(n14121), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13743) );
  OAI21_X1 U15850 ( .B1(n13900), .B2(n14114), .A(n13743), .ZN(n13744) );
  AOI21_X1 U15851 ( .B1(n13902), .B2(n13931), .A(n13744), .ZN(n13745) );
  OAI211_X1 U15852 ( .C1(n14320), .C2(n13905), .A(n13746), .B(n13745), .ZN(
        P2_U3188) );
  XNOR2_X1 U15853 ( .A(n13748), .B(n13747), .ZN(n13755) );
  NAND2_X1 U15854 ( .A1(n13888), .A2(n13749), .ZN(n13750) );
  NAND2_X1 U15855 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n15388)
         );
  OAI211_X1 U15856 ( .C1(n13891), .C2(n13751), .A(n13750), .B(n15388), .ZN(
        n13752) );
  AOI21_X1 U15857 ( .B1(n13753), .B2(n13926), .A(n13752), .ZN(n13754) );
  OAI21_X1 U15858 ( .B1(n13755), .B2(n13921), .A(n13754), .ZN(P2_U3189) );
  NAND2_X1 U15859 ( .A1(n13757), .A2(n13756), .ZN(n13759) );
  XOR2_X1 U15860 ( .A(n13759), .B(n7163), .Z(n13764) );
  AOI22_X1 U15861 ( .A1(n13935), .A2(n14097), .B1(n13933), .B2(n14082), .ZN(
        n14175) );
  NOR2_X1 U15862 ( .A1(n13760), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14033) );
  AOI21_X1 U15863 ( .B1(n13917), .B2(n14180), .A(n14033), .ZN(n13761) );
  OAI21_X1 U15864 ( .B1(n14175), .B2(n13919), .A(n13761), .ZN(n13762) );
  AOI21_X1 U15865 ( .B1(n14179), .B2(n13926), .A(n13762), .ZN(n13763) );
  OAI21_X1 U15866 ( .B1(n13764), .B2(n13921), .A(n13763), .ZN(P2_U3191) );
  INV_X1 U15867 ( .A(n13765), .ZN(n13766) );
  AOI21_X1 U15868 ( .B1(n13768), .B2(n13767), .A(n13766), .ZN(n13774) );
  NAND2_X1 U15869 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n13969) );
  OAI21_X1 U15870 ( .B1(n13891), .B2(n13769), .A(n13969), .ZN(n13771) );
  NOR2_X1 U15871 ( .A1(n13905), .A2(n10439), .ZN(n13770) );
  AOI211_X1 U15872 ( .C1(n13888), .C2(n13772), .A(n13771), .B(n13770), .ZN(
        n13773) );
  OAI21_X1 U15873 ( .B1(n13774), .B2(n13921), .A(n13773), .ZN(P2_U3193) );
  OAI211_X1 U15874 ( .C1(n13777), .C2(n13776), .A(n13775), .B(n13872), .ZN(
        n13783) );
  AOI22_X1 U15875 ( .A1(n13931), .A2(n14082), .B1(n14097), .B2(n13933), .ZN(
        n14146) );
  INV_X1 U15876 ( .A(n14146), .ZN(n13781) );
  INV_X1 U15877 ( .A(n14152), .ZN(n13779) );
  OAI22_X1 U15878 ( .A1(n13891), .A2(n13779), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13778), .ZN(n13780) );
  AOI21_X1 U15879 ( .B1(n13781), .B2(n13888), .A(n13780), .ZN(n13782) );
  OAI211_X1 U15880 ( .C1(n7435), .C2(n13905), .A(n13783), .B(n13782), .ZN(
        P2_U3195) );
  NAND2_X1 U15881 ( .A1(n13785), .A2(n13784), .ZN(n13787) );
  XOR2_X1 U15882 ( .A(n13787), .B(n13786), .Z(n13795) );
  NOR2_X1 U15883 ( .A1(n13919), .A2(n13788), .ZN(n13792) );
  OAI21_X1 U15884 ( .B1(n13891), .B2(n13790), .A(n13789), .ZN(n13791) );
  AOI211_X1 U15885 ( .C1(n13793), .C2(n13926), .A(n13792), .B(n13791), .ZN(
        n13794) );
  OAI21_X1 U15886 ( .B1(n13795), .B2(n13921), .A(n13794), .ZN(P2_U3196) );
  OAI211_X1 U15887 ( .C1(n13798), .C2(n13797), .A(n13796), .B(n13872), .ZN(
        n13803) );
  AOI22_X1 U15888 ( .A1(n14088), .A2(n13917), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13799) );
  OAI21_X1 U15889 ( .B1(n13800), .B2(n13900), .A(n13799), .ZN(n13801) );
  AOI21_X1 U15890 ( .B1(n13902), .B2(n14081), .A(n13801), .ZN(n13802) );
  OAI211_X1 U15891 ( .C1(n14404), .C2(n13905), .A(n13803), .B(n13802), .ZN(
        P2_U3197) );
  XNOR2_X1 U15892 ( .A(n13805), .B(n13804), .ZN(n13922) );
  NOR2_X1 U15893 ( .A1(n13922), .A2(n13923), .ZN(n13920) );
  AOI21_X1 U15894 ( .B1(n13805), .B2(n13804), .A(n13920), .ZN(n13809) );
  XOR2_X1 U15895 ( .A(n13807), .B(n13806), .Z(n13808) );
  NAND2_X1 U15896 ( .A1(n13809), .A2(n13808), .ZN(n13829) );
  OAI21_X1 U15897 ( .B1(n13809), .B2(n13808), .A(n13829), .ZN(n13810) );
  NAND2_X1 U15898 ( .A1(n13810), .A2(n13872), .ZN(n13814) );
  OAI22_X1 U15899 ( .A1(n14198), .A2(n14199), .B1(n13811), .B2(n14197), .ZN(
        n14235) );
  OAI22_X1 U15900 ( .A1(n13891), .A2(n14240), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15656), .ZN(n13812) );
  AOI21_X1 U15901 ( .B1(n13888), .B2(n14235), .A(n13812), .ZN(n13813) );
  OAI211_X1 U15902 ( .C1(n6838), .C2(n13905), .A(n13814), .B(n13813), .ZN(
        P2_U3198) );
  OAI21_X1 U15903 ( .B1(n13817), .B2(n13816), .A(n13815), .ZN(n13818) );
  NAND2_X1 U15904 ( .A1(n13818), .A2(n13872), .ZN(n13824) );
  AND2_X1 U15905 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n13960) );
  NOR2_X1 U15906 ( .A1(n13891), .A2(n13819), .ZN(n13820) );
  AOI211_X1 U15907 ( .C1(n13821), .C2(n13926), .A(n13960), .B(n13820), .ZN(
        n13823) );
  AOI22_X1 U15908 ( .A1(n13902), .A2(n13950), .B1(n13909), .B2(n13948), .ZN(
        n13822) );
  NAND3_X1 U15909 ( .A1(n13824), .A2(n13823), .A3(n13822), .ZN(P2_U3199) );
  AOI22_X1 U15910 ( .A1(n13935), .A2(n14082), .B1(n14097), .B2(n13937), .ZN(
        n14216) );
  INV_X1 U15911 ( .A(n13825), .ZN(n14223) );
  AOI22_X1 U15912 ( .A1(n13917), .A2(n14223), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13826) );
  OAI21_X1 U15913 ( .B1(n14216), .B2(n13919), .A(n13826), .ZN(n13833) );
  NAND3_X1 U15914 ( .A1(n13829), .A2(n13828), .A3(n13827), .ZN(n13831) );
  AOI21_X1 U15915 ( .B1(n13831), .B2(n13830), .A(n13921), .ZN(n13832) );
  AOI211_X1 U15916 ( .C1(n14222), .C2(n13926), .A(n13833), .B(n13832), .ZN(
        n13834) );
  INV_X1 U15917 ( .A(n13834), .ZN(P2_U3200) );
  OAI211_X1 U15918 ( .C1(n13837), .C2(n13836), .A(n13835), .B(n13872), .ZN(
        n13842) );
  OAI22_X1 U15919 ( .A1(n14104), .A2(n13891), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13838), .ZN(n13840) );
  NOR2_X1 U15920 ( .A1(n13877), .A2(n13912), .ZN(n13839) );
  AOI211_X1 U15921 ( .C1(n14096), .C2(n13909), .A(n13840), .B(n13839), .ZN(
        n13841) );
  OAI211_X1 U15922 ( .C1(n7432), .C2(n13905), .A(n13842), .B(n13841), .ZN(
        P2_U3201) );
  OAI21_X1 U15923 ( .B1(n13845), .B2(n13844), .A(n13843), .ZN(n13846) );
  NAND2_X1 U15924 ( .A1(n13846), .A2(n13872), .ZN(n13853) );
  OR2_X1 U15925 ( .A1(n13919), .A2(n13847), .ZN(n13848) );
  NAND2_X1 U15926 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n15385) );
  OAI211_X1 U15927 ( .C1(n13891), .C2(n13849), .A(n13848), .B(n15385), .ZN(
        n13850) );
  AOI21_X1 U15928 ( .B1(n13851), .B2(n13926), .A(n13850), .ZN(n13852) );
  NAND2_X1 U15929 ( .A1(n13853), .A2(n13852), .ZN(P2_U3203) );
  NAND2_X1 U15930 ( .A1(n13855), .A2(n13854), .ZN(n13857) );
  XOR2_X1 U15931 ( .A(n13857), .B(n13856), .Z(n13862) );
  AOI22_X1 U15932 ( .A1(n13932), .A2(n14082), .B1(n13934), .B2(n14097), .ZN(
        n14162) );
  INV_X1 U15933 ( .A(n14164), .ZN(n13858) );
  AOI22_X1 U15934 ( .A1(n13917), .A2(n13858), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13859) );
  OAI21_X1 U15935 ( .B1(n14162), .B2(n13919), .A(n13859), .ZN(n13860) );
  AOI21_X1 U15936 ( .B1(n14336), .B2(n13926), .A(n13860), .ZN(n13861) );
  OAI21_X1 U15937 ( .B1(n13862), .B2(n13921), .A(n13861), .ZN(P2_U3205) );
  OAI211_X1 U15938 ( .C1(n13719), .C2(n13864), .A(n13863), .B(n13872), .ZN(
        n13869) );
  NAND2_X1 U15939 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n15418)
         );
  OAI21_X1 U15940 ( .B1(n13891), .B2(n13865), .A(n15418), .ZN(n13866) );
  AOI21_X1 U15941 ( .B1(n13888), .B2(n13867), .A(n13866), .ZN(n13868) );
  OAI211_X1 U15942 ( .C1(n13870), .C2(n13905), .A(n13869), .B(n13868), .ZN(
        P2_U3206) );
  INV_X1 U15943 ( .A(n13871), .ZN(n13873) );
  OAI211_X1 U15944 ( .C1(n13875), .C2(n13874), .A(n13873), .B(n13872), .ZN(
        n13882) );
  OAI22_X1 U15945 ( .A1(n13877), .A2(n14199), .B1(n13876), .B2(n14197), .ZN(
        n14129) );
  INV_X1 U15946 ( .A(n14139), .ZN(n13879) );
  OAI22_X1 U15947 ( .A1(n13879), .A2(n13891), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13878), .ZN(n13880) );
  AOI21_X1 U15948 ( .B1(n14129), .B2(n13888), .A(n13880), .ZN(n13881) );
  OAI211_X1 U15949 ( .C1(n14411), .C2(n13905), .A(n13882), .B(n13881), .ZN(
        P2_U3207) );
  INV_X1 U15950 ( .A(n13883), .ZN(n13884) );
  AOI21_X1 U15951 ( .B1(n13886), .B2(n13885), .A(n13884), .ZN(n13894) );
  NAND2_X1 U15952 ( .A1(n13888), .A2(n13887), .ZN(n13889) );
  NAND2_X1 U15953 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n15416)
         );
  OAI211_X1 U15954 ( .C1(n13891), .C2(n13890), .A(n13889), .B(n15416), .ZN(
        n13892) );
  AOI21_X1 U15955 ( .B1(n14382), .B2(n13926), .A(n13892), .ZN(n13893) );
  OAI21_X1 U15956 ( .B1(n13894), .B2(n13921), .A(n13893), .ZN(P2_U3208) );
  AOI21_X1 U15957 ( .B1(n13896), .B2(n13895), .A(n13921), .ZN(n13898) );
  NAND2_X1 U15958 ( .A1(n13898), .A2(n13897), .ZN(n13904) );
  NAND2_X1 U15959 ( .A1(n13917), .A2(n14208), .ZN(n13899) );
  NAND2_X1 U15960 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14014)
         );
  OAI211_X1 U15961 ( .C1(n13900), .C2(n14200), .A(n13899), .B(n14014), .ZN(
        n13901) );
  AOI21_X1 U15962 ( .B1(n13902), .B2(n13936), .A(n13901), .ZN(n13903) );
  OAI211_X1 U15963 ( .C1(n14352), .C2(n13905), .A(n13904), .B(n13903), .ZN(
        P2_U3210) );
  AOI21_X1 U15964 ( .B1(n13908), .B2(n13907), .A(n13906), .ZN(n13916) );
  NAND2_X1 U15965 ( .A1(n14065), .A2(n13909), .ZN(n13911) );
  AOI22_X1 U15966 ( .A1(n14068), .A2(n13917), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13910) );
  OAI211_X1 U15967 ( .C1(n13913), .C2(n13912), .A(n13911), .B(n13910), .ZN(
        n13914) );
  AOI21_X1 U15968 ( .B1(n7254), .B2(n13926), .A(n13914), .ZN(n13915) );
  OAI21_X1 U15969 ( .B1(n13916), .B2(n13921), .A(n13915), .ZN(P2_U3212) );
  AOI22_X1 U15970 ( .A1(n13937), .A2(n14082), .B1(n13939), .B2(n14097), .ZN(
        n14254) );
  AOI22_X1 U15971 ( .A1(n13917), .A2(n14257), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13918) );
  OAI21_X1 U15972 ( .B1(n14254), .B2(n13919), .A(n13918), .ZN(n13925) );
  AOI211_X1 U15973 ( .C1(n13923), .C2(n13922), .A(n13921), .B(n13920), .ZN(
        n13924) );
  AOI211_X1 U15974 ( .C1(n14433), .C2(n13926), .A(n13925), .B(n13924), .ZN(
        n13927) );
  INV_X1 U15975 ( .A(n13927), .ZN(P2_U3213) );
  MUX2_X1 U15976 ( .A(n13928), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13945), .Z(
        P2_U3562) );
  MUX2_X1 U15977 ( .A(n13929), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13945), .Z(
        P2_U3561) );
  MUX2_X1 U15978 ( .A(n13930), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13945), .Z(
        P2_U3560) );
  MUX2_X1 U15979 ( .A(n14050), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13945), .Z(
        P2_U3559) );
  MUX2_X1 U15980 ( .A(n14065), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13945), .Z(
        P2_U3558) );
  MUX2_X1 U15981 ( .A(n14083), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13945), .Z(
        P2_U3557) );
  MUX2_X1 U15982 ( .A(n14096), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13945), .Z(
        P2_U3556) );
  MUX2_X1 U15983 ( .A(n14081), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13945), .Z(
        P2_U3555) );
  MUX2_X1 U15984 ( .A(n14098), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13945), .Z(
        P2_U3554) );
  MUX2_X1 U15985 ( .A(n13931), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13945), .Z(
        P2_U3553) );
  MUX2_X1 U15986 ( .A(n13932), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13945), .Z(
        P2_U3552) );
  MUX2_X1 U15987 ( .A(n13933), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13945), .Z(
        P2_U3551) );
  MUX2_X1 U15988 ( .A(n13934), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13945), .Z(
        P2_U3550) );
  MUX2_X1 U15989 ( .A(n13935), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13945), .Z(
        P2_U3549) );
  MUX2_X1 U15990 ( .A(n13936), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13945), .Z(
        P2_U3548) );
  MUX2_X1 U15991 ( .A(n13937), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13945), .Z(
        P2_U3547) );
  MUX2_X1 U15992 ( .A(n13938), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13945), .Z(
        P2_U3546) );
  MUX2_X1 U15993 ( .A(n13939), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13945), .Z(
        P2_U3545) );
  MUX2_X1 U15994 ( .A(n13940), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13945), .Z(
        P2_U3544) );
  MUX2_X1 U15995 ( .A(n13941), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13945), .Z(
        P2_U3543) );
  MUX2_X1 U15996 ( .A(n13942), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13945), .Z(
        P2_U3542) );
  MUX2_X1 U15997 ( .A(n13943), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13945), .Z(
        P2_U3541) );
  MUX2_X1 U15998 ( .A(n13944), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13945), .Z(
        P2_U3540) );
  MUX2_X1 U15999 ( .A(n13946), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13945), .Z(
        P2_U3539) );
  MUX2_X1 U16000 ( .A(n13947), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13945), .Z(
        P2_U3538) );
  MUX2_X1 U16001 ( .A(n13948), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13945), .Z(
        P2_U3537) );
  MUX2_X1 U16002 ( .A(n13949), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13945), .Z(
        P2_U3536) );
  MUX2_X1 U16003 ( .A(n13950), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13945), .Z(
        P2_U3535) );
  MUX2_X1 U16004 ( .A(n13951), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13945), .Z(
        P2_U3534) );
  MUX2_X1 U16005 ( .A(n13952), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13945), .Z(
        P2_U3533) );
  MUX2_X1 U16006 ( .A(n7158), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13945), .Z(
        P2_U3532) );
  MUX2_X1 U16007 ( .A(n13954), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13945), .Z(
        P2_U3531) );
  MUX2_X1 U16008 ( .A(n10885), .B(P2_REG2_REG_5__SCAN_IN), .S(n13964), .Z(
        n13955) );
  NAND3_X1 U16009 ( .A1(n13957), .A2(n13956), .A3(n13955), .ZN(n13958) );
  NAND3_X1 U16010 ( .A1(n15451), .A2(n13959), .A3(n13958), .ZN(n13968) );
  AOI21_X1 U16011 ( .B1(n15336), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n13960), .ZN(
        n13967) );
  OAI211_X1 U16012 ( .C1(n13963), .C2(n13962), .A(n15402), .B(n13961), .ZN(
        n13966) );
  NAND2_X1 U16013 ( .A1(n15450), .A2(n13964), .ZN(n13965) );
  NAND4_X1 U16014 ( .A1(n13968), .A2(n13967), .A3(n13966), .A4(n13965), .ZN(
        P2_U3219) );
  INV_X1 U16015 ( .A(n13969), .ZN(n13972) );
  NOR2_X1 U16016 ( .A1(n15457), .A2(n13970), .ZN(n13971) );
  AOI211_X1 U16017 ( .C1(n15450), .C2(n13975), .A(n13972), .B(n13971), .ZN(
        n13982) );
  OAI211_X1 U16018 ( .C1(n13974), .C2(n13973), .A(n15402), .B(n15378), .ZN(
        n13981) );
  MUX2_X1 U16019 ( .A(n12375), .B(P2_REG2_REG_8__SCAN_IN), .S(n13975), .Z(
        n13976) );
  NAND3_X1 U16020 ( .A1(n15370), .A2(n13977), .A3(n13976), .ZN(n13978) );
  NAND3_X1 U16021 ( .A1(n15451), .A2(n13979), .A3(n13978), .ZN(n13980) );
  NAND3_X1 U16022 ( .A1(n13982), .A2(n13981), .A3(n13980), .ZN(P2_U3222) );
  NAND2_X1 U16023 ( .A1(n13983), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n13986) );
  NAND2_X1 U16024 ( .A1(n13984), .A2(n13993), .ZN(n13985) );
  NAND2_X1 U16025 ( .A1(n13986), .A2(n13985), .ZN(n14001) );
  INV_X1 U16026 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13987) );
  XNOR2_X1 U16027 ( .A(n14011), .B(n13987), .ZN(n14000) );
  XNOR2_X1 U16028 ( .A(n14001), .B(n14000), .ZN(n13999) );
  NOR2_X1 U16029 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15656), .ZN(n13988) );
  AOI21_X1 U16030 ( .B1(n15336), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n13988), 
        .ZN(n13989) );
  INV_X1 U16031 ( .A(n13989), .ZN(n13997) );
  INV_X1 U16032 ( .A(n13990), .ZN(n13992) );
  XNOR2_X1 U16033 ( .A(n14011), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13994) );
  INV_X1 U16034 ( .A(n15402), .ZN(n15444) );
  NOR2_X1 U16035 ( .A1(n13995), .A2(n13994), .ZN(n14010) );
  AOI211_X1 U16036 ( .C1(n13995), .C2(n13994), .A(n15444), .B(n14010), .ZN(
        n13996) );
  AOI211_X1 U16037 ( .C1(n15450), .C2(n14011), .A(n13997), .B(n13996), .ZN(
        n13998) );
  OAI21_X1 U16038 ( .B1(n13999), .B2(n15411), .A(n13998), .ZN(P2_U3230) );
  NAND2_X1 U16039 ( .A1(n14001), .A2(n14000), .ZN(n14003) );
  NAND2_X1 U16040 ( .A1(n14011), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n14002) );
  NAND2_X1 U16041 ( .A1(n14003), .A2(n14002), .ZN(n15454) );
  INV_X1 U16042 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14004) );
  MUX2_X1 U16043 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n14004), .S(n15449), .Z(
        n15453) );
  NAND2_X1 U16044 ( .A1(n15454), .A2(n15453), .ZN(n15452) );
  NAND2_X1 U16045 ( .A1(n15449), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14005) );
  NAND2_X1 U16046 ( .A1(n15452), .A2(n14005), .ZN(n14006) );
  NAND2_X1 U16047 ( .A1(n14006), .A2(n14017), .ZN(n14007) );
  INV_X1 U16048 ( .A(n14026), .ZN(n14008) );
  AOI21_X1 U16049 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14009), .A(n14008), 
        .ZN(n14020) );
  XNOR2_X1 U16050 ( .A(n15449), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15445) );
  NOR2_X1 U16051 ( .A1(n15446), .A2(n15445), .ZN(n15443) );
  OAI211_X1 U16052 ( .C1(n14013), .C2(P2_REG1_REG_18__SCAN_IN), .A(n14023), 
        .B(n15402), .ZN(n14019) );
  INV_X1 U16053 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14015) );
  OAI21_X1 U16054 ( .B1(n15457), .B2(n14015), .A(n14014), .ZN(n14016) );
  AOI21_X1 U16055 ( .B1(n14017), .B2(n15450), .A(n14016), .ZN(n14018) );
  OAI211_X1 U16056 ( .C1(n14020), .C2(n15411), .A(n14019), .B(n14018), .ZN(
        P2_U3232) );
  INV_X1 U16057 ( .A(n14021), .ZN(n14022) );
  NAND2_X1 U16058 ( .A1(n14023), .A2(n14022), .ZN(n14024) );
  INV_X1 U16059 ( .A(n14030), .ZN(n14028) );
  NAND2_X1 U16060 ( .A1(n14026), .A2(n14025), .ZN(n14027) );
  XNOR2_X1 U16061 ( .A(n14027), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n14029) );
  INV_X1 U16062 ( .A(n14035), .ZN(n14287) );
  NAND2_X1 U16063 ( .A1(n14242), .A2(n14287), .ZN(n14043) );
  OAI21_X1 U16064 ( .B1(n14036), .B2(n14242), .A(n14043), .ZN(n14037) );
  AOI21_X1 U16065 ( .B1(n14387), .B2(n14278), .A(n14037), .ZN(n14038) );
  OAI21_X1 U16066 ( .B1(n14039), .B2(n14266), .A(n14038), .ZN(P2_U3234) );
  INV_X1 U16067 ( .A(n14040), .ZN(n14041) );
  AOI211_X1 U16068 ( .C1(n14042), .C2(n14286), .A(n14363), .B(n14041), .ZN(
        n14288) );
  INV_X1 U16069 ( .A(n14288), .ZN(n14047) );
  OAI21_X1 U16070 ( .B1(n14242), .B2(n14044), .A(n14043), .ZN(n14045) );
  AOI21_X1 U16071 ( .B1(n14286), .B2(n14278), .A(n14045), .ZN(n14046) );
  OAI21_X1 U16072 ( .B1(n14047), .B2(n14266), .A(n14046), .ZN(P2_U3235) );
  XNOR2_X1 U16073 ( .A(n14049), .B(n14048), .ZN(n14051) );
  AOI222_X1 U16074 ( .A1(n14252), .A2(n14051), .B1(n14050), .B2(n14082), .C1(
        n14083), .C2(n14097), .ZN(n14301) );
  AOI21_X1 U16075 ( .B1(n14066), .B2(n14298), .A(n14363), .ZN(n14053) );
  NAND2_X1 U16076 ( .A1(n14053), .A2(n14052), .ZN(n14300) );
  NAND3_X1 U16077 ( .A1(n14297), .A2(n14268), .A3(n14296), .ZN(n14060) );
  INV_X1 U16078 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n14056) );
  OAI22_X1 U16079 ( .A1(n14057), .A2(n14239), .B1(n14056), .B2(n14242), .ZN(
        n14058) );
  AOI21_X1 U16080 ( .B1(n14298), .B2(n14278), .A(n14058), .ZN(n14059) );
  OAI211_X1 U16081 ( .C1(n14300), .C2(n14266), .A(n14060), .B(n14059), .ZN(
        n14061) );
  INV_X1 U16082 ( .A(n14061), .ZN(n14062) );
  OAI21_X1 U16083 ( .B1(n14301), .B2(n14264), .A(n14062), .ZN(P2_U3238) );
  INV_X1 U16084 ( .A(n14086), .ZN(n14067) );
  AOI211_X1 U16085 ( .C1(n7254), .C2(n14067), .A(n14363), .B(n7428), .ZN(
        n14303) );
  AOI22_X1 U16086 ( .A1(n14068), .A2(n14276), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14264), .ZN(n14069) );
  OAI21_X1 U16087 ( .B1(n14070), .B2(n14226), .A(n14069), .ZN(n14074) );
  XNOR2_X1 U16088 ( .A(n14072), .B(n14071), .ZN(n14306) );
  NOR2_X1 U16089 ( .A1(n14306), .A2(n14248), .ZN(n14073) );
  AOI211_X1 U16090 ( .C1(n14303), .C2(n14273), .A(n14074), .B(n14073), .ZN(
        n14075) );
  OAI21_X1 U16091 ( .B1(n14305), .B2(n14264), .A(n14075), .ZN(P2_U3239) );
  OAI21_X1 U16092 ( .B1(n14080), .B2(n14079), .A(n14252), .ZN(n14085) );
  AOI22_X1 U16093 ( .A1(n14083), .A2(n14082), .B1(n14081), .B2(n14097), .ZN(
        n14084) );
  INV_X1 U16094 ( .A(n14308), .ZN(n14093) );
  OAI21_X1 U16095 ( .B1(n14103), .B2(n14404), .A(n14262), .ZN(n14087) );
  AOI22_X1 U16096 ( .A1(n14088), .A2(n14276), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14264), .ZN(n14091) );
  NAND2_X1 U16097 ( .A1(n14089), .A2(n14278), .ZN(n14090) );
  OAI211_X1 U16098 ( .C1(n14307), .C2(n14266), .A(n14091), .B(n14090), .ZN(
        n14092) );
  AOI21_X1 U16099 ( .B1(n14093), .B2(n14242), .A(n14092), .ZN(n14094) );
  OAI21_X1 U16100 ( .B1(n14309), .B2(n14248), .A(n14094), .ZN(P2_U3240) );
  OAI21_X1 U16101 ( .B1(n6500), .B2(n7791), .A(n14095), .ZN(n14099) );
  AOI222_X1 U16102 ( .A1(n14252), .A2(n14099), .B1(n14098), .B2(n14097), .C1(
        n14096), .C2(n14082), .ZN(n14318) );
  NAND2_X1 U16103 ( .A1(n14100), .A2(n7791), .ZN(n14313) );
  AND3_X1 U16104 ( .A1(n14314), .A2(n14313), .A3(n14268), .ZN(n14109) );
  NAND2_X1 U16105 ( .A1(n14119), .A2(n14312), .ZN(n14101) );
  NAND2_X1 U16106 ( .A1(n14101), .A2(n14262), .ZN(n14102) );
  OR2_X1 U16107 ( .A1(n14103), .A2(n14102), .ZN(n14315) );
  INV_X1 U16108 ( .A(n14104), .ZN(n14105) );
  AOI22_X1 U16109 ( .A1(n14105), .A2(n14276), .B1(n14264), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n14107) );
  NAND2_X1 U16110 ( .A1(n14312), .A2(n14278), .ZN(n14106) );
  OAI211_X1 U16111 ( .C1(n14315), .C2(n14266), .A(n14107), .B(n14106), .ZN(
        n14108) );
  NOR2_X1 U16112 ( .A1(n14109), .A2(n14108), .ZN(n14110) );
  OAI21_X1 U16113 ( .B1(n14318), .B2(n14264), .A(n14110), .ZN(P2_U3241) );
  INV_X1 U16114 ( .A(n14117), .ZN(n14111) );
  XNOR2_X1 U16115 ( .A(n14112), .B(n14111), .ZN(n14116) );
  OAI22_X1 U16116 ( .A1(n14114), .A2(n14199), .B1(n14113), .B2(n14197), .ZN(
        n14115) );
  AOI21_X1 U16117 ( .B1(n14116), .B2(n14252), .A(n14115), .ZN(n14324) );
  XNOR2_X1 U16118 ( .A(n14118), .B(n14117), .ZN(n14322) );
  AOI21_X1 U16119 ( .B1(n14135), .B2(n14122), .A(n14363), .ZN(n14120) );
  NAND2_X1 U16120 ( .A1(n14120), .A2(n14119), .ZN(n14319) );
  AOI22_X1 U16121 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(n14280), .B1(n14121), 
        .B2(n14276), .ZN(n14124) );
  NAND2_X1 U16122 ( .A1(n14122), .A2(n14278), .ZN(n14123) );
  OAI211_X1 U16123 ( .C1(n14319), .C2(n14266), .A(n14124), .B(n14123), .ZN(
        n14125) );
  AOI21_X1 U16124 ( .B1(n14322), .B2(n14268), .A(n14125), .ZN(n14126) );
  OAI21_X1 U16125 ( .B1(n14324), .B2(n14264), .A(n14126), .ZN(P2_U3242) );
  XNOR2_X1 U16126 ( .A(n14128), .B(n14127), .ZN(n14131) );
  INV_X1 U16127 ( .A(n14129), .ZN(n14130) );
  OAI21_X1 U16128 ( .B1(n14131), .B2(n14217), .A(n14130), .ZN(n14327) );
  INV_X1 U16129 ( .A(n14327), .ZN(n14144) );
  NAND2_X1 U16130 ( .A1(n14132), .A2(n6738), .ZN(n14133) );
  AND2_X1 U16131 ( .A1(n14134), .A2(n14133), .ZN(n14329) );
  INV_X1 U16132 ( .A(n14150), .ZN(n14137) );
  INV_X1 U16133 ( .A(n14135), .ZN(n14136) );
  AOI211_X1 U16134 ( .C1(n14138), .C2(n14137), .A(n14363), .B(n14136), .ZN(
        n14328) );
  NAND2_X1 U16135 ( .A1(n14328), .A2(n14273), .ZN(n14141) );
  AOI22_X1 U16136 ( .A1(n14280), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14276), 
        .B2(n14139), .ZN(n14140) );
  OAI211_X1 U16137 ( .C1(n14411), .C2(n14226), .A(n14141), .B(n14140), .ZN(
        n14142) );
  AOI21_X1 U16138 ( .B1(n14329), .B2(n14268), .A(n14142), .ZN(n14143) );
  OAI21_X1 U16139 ( .B1(n14144), .B2(n14280), .A(n14143), .ZN(P2_U3243) );
  XOR2_X1 U16140 ( .A(n14145), .B(n14148), .Z(n14147) );
  OAI21_X1 U16141 ( .B1(n14147), .B2(n14217), .A(n14146), .ZN(n14332) );
  INV_X1 U16142 ( .A(n14332), .ZN(n14157) );
  XNOR2_X1 U16143 ( .A(n14149), .B(n14148), .ZN(n14334) );
  AOI211_X1 U16144 ( .C1(n14151), .C2(n14166), .A(n14363), .B(n14150), .ZN(
        n14333) );
  NAND2_X1 U16145 ( .A1(n14333), .A2(n14273), .ZN(n14154) );
  AOI22_X1 U16146 ( .A1(n14280), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14276), 
        .B2(n14152), .ZN(n14153) );
  OAI211_X1 U16147 ( .C1(n7435), .C2(n14226), .A(n14154), .B(n14153), .ZN(
        n14155) );
  AOI21_X1 U16148 ( .B1(n14334), .B2(n14268), .A(n14155), .ZN(n14156) );
  OAI21_X1 U16149 ( .B1(n14157), .B2(n14280), .A(n14156), .ZN(P2_U3244) );
  XNOR2_X1 U16150 ( .A(n14158), .B(n14159), .ZN(n14339) );
  XNOR2_X1 U16151 ( .A(n14160), .B(n14159), .ZN(n14161) );
  NAND2_X1 U16152 ( .A1(n14161), .A2(n14252), .ZN(n14163) );
  NAND2_X1 U16153 ( .A1(n14163), .A2(n14162), .ZN(n14341) );
  NAND2_X1 U16154 ( .A1(n14341), .A2(n14242), .ZN(n14171) );
  INV_X1 U16155 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n14165) );
  OAI22_X1 U16156 ( .A1(n14242), .A2(n14165), .B1(n14164), .B2(n14239), .ZN(
        n14169) );
  AOI21_X1 U16157 ( .B1(n14177), .B2(n14336), .A(n14363), .ZN(n14167) );
  NAND2_X1 U16158 ( .A1(n14167), .A2(n14166), .ZN(n14338) );
  NOR2_X1 U16159 ( .A1(n14338), .A2(n14266), .ZN(n14168) );
  AOI211_X1 U16160 ( .C1(n14278), .C2(n14336), .A(n14169), .B(n14168), .ZN(
        n14170) );
  OAI211_X1 U16161 ( .C1(n14339), .C2(n14248), .A(n14171), .B(n14170), .ZN(
        P2_U3245) );
  XOR2_X1 U16162 ( .A(n14172), .B(n14173), .Z(n14346) );
  INV_X1 U16163 ( .A(n14346), .ZN(n14185) );
  XNOR2_X1 U16164 ( .A(n14174), .B(n14173), .ZN(n14176) );
  OAI21_X1 U16165 ( .B1(n14176), .B2(n14217), .A(n14175), .ZN(n14344) );
  NAND2_X1 U16166 ( .A1(n14344), .A2(n14242), .ZN(n14184) );
  INV_X1 U16167 ( .A(n14177), .ZN(n14178) );
  AOI211_X1 U16168 ( .C1(n14179), .C2(n14207), .A(n14363), .B(n14178), .ZN(
        n14345) );
  AOI22_X1 U16169 ( .A1(n14280), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14276), 
        .B2(n14180), .ZN(n14181) );
  OAI21_X1 U16170 ( .B1(n14421), .B2(n14226), .A(n14181), .ZN(n14182) );
  AOI21_X1 U16171 ( .B1(n14345), .B2(n14273), .A(n14182), .ZN(n14183) );
  OAI211_X1 U16172 ( .C1(n14248), .C2(n14185), .A(n14184), .B(n14183), .ZN(
        P2_U3246) );
  INV_X1 U16173 ( .A(n14186), .ZN(n14193) );
  XNOR2_X1 U16174 ( .A(n14187), .B(n14193), .ZN(n14188) );
  NAND2_X1 U16175 ( .A1(n14188), .A2(n14252), .ZN(n14204) );
  NAND2_X1 U16176 ( .A1(n14189), .A2(n14190), .ZN(n14219) );
  NAND2_X1 U16177 ( .A1(n14219), .A2(n14220), .ZN(n14192) );
  NAND2_X1 U16178 ( .A1(n14192), .A2(n14191), .ZN(n14194) );
  NAND2_X1 U16179 ( .A1(n14194), .A2(n14193), .ZN(n14196) );
  NAND2_X1 U16180 ( .A1(n14196), .A2(n14195), .ZN(n14349) );
  OAI22_X1 U16181 ( .A1(n14200), .A2(n14199), .B1(n14198), .B2(n14197), .ZN(
        n14201) );
  AOI21_X1 U16182 ( .B1(n14349), .B2(n14202), .A(n14201), .ZN(n14203) );
  NAND2_X1 U16183 ( .A1(n14204), .A2(n14203), .ZN(n14354) );
  INV_X1 U16184 ( .A(n14354), .ZN(n14214) );
  INV_X1 U16185 ( .A(n14221), .ZN(n14205) );
  NAND2_X1 U16186 ( .A1(n14205), .A2(n14209), .ZN(n14206) );
  NAND3_X1 U16187 ( .A1(n14207), .A2(n14206), .A3(n14262), .ZN(n14350) );
  AOI22_X1 U16188 ( .A1(n14280), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14276), 
        .B2(n14208), .ZN(n14211) );
  NAND2_X1 U16189 ( .A1(n14209), .A2(n14278), .ZN(n14210) );
  OAI211_X1 U16190 ( .C1(n14350), .C2(n14266), .A(n14211), .B(n14210), .ZN(
        n14212) );
  AOI21_X1 U16191 ( .B1(n14349), .B2(n14275), .A(n14212), .ZN(n14213) );
  OAI21_X1 U16192 ( .B1(n14214), .B2(n14280), .A(n14213), .ZN(P2_U3247) );
  XOR2_X1 U16193 ( .A(n14220), .B(n7138), .Z(n14218) );
  OAI21_X1 U16194 ( .B1(n14218), .B2(n14217), .A(n14216), .ZN(n14357) );
  INV_X1 U16195 ( .A(n14357), .ZN(n14229) );
  XOR2_X1 U16196 ( .A(n14220), .B(n14219), .Z(n14359) );
  AOI211_X1 U16197 ( .C1(n14222), .C2(n6840), .A(n14363), .B(n14221), .ZN(
        n14358) );
  NAND2_X1 U16198 ( .A1(n14358), .A2(n14273), .ZN(n14225) );
  AOI22_X1 U16199 ( .A1(n14280), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14276), 
        .B2(n14223), .ZN(n14224) );
  OAI211_X1 U16200 ( .C1(n14429), .C2(n14226), .A(n14225), .B(n14224), .ZN(
        n14227) );
  AOI21_X1 U16201 ( .B1(n14359), .B2(n14268), .A(n14227), .ZN(n14228) );
  OAI21_X1 U16202 ( .B1(n14229), .B2(n14280), .A(n14228), .ZN(P2_U3248) );
  INV_X1 U16203 ( .A(n14189), .ZN(n14230) );
  AOI21_X1 U16204 ( .B1(n14232), .B2(n14231), .A(n14230), .ZN(n14367) );
  INV_X1 U16205 ( .A(n14367), .ZN(n14249) );
  XNOR2_X1 U16206 ( .A(n14234), .B(n14233), .ZN(n14236) );
  AOI21_X1 U16207 ( .B1(n14236), .B2(n14252), .A(n14235), .ZN(n14368) );
  INV_X1 U16208 ( .A(n14368), .ZN(n14244) );
  AND2_X1 U16209 ( .A1(n14263), .A2(n14245), .ZN(n14238) );
  OR2_X1 U16210 ( .A1(n14238), .A2(n14237), .ZN(n14364) );
  OAI22_X1 U16211 ( .A1(n14364), .A2(n14241), .B1(n14240), .B2(n14239), .ZN(
        n14243) );
  OAI21_X1 U16212 ( .B1(n14244), .B2(n14243), .A(n14242), .ZN(n14247) );
  AOI22_X1 U16213 ( .A1(n14245), .A2(n14278), .B1(n14264), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n14246) );
  OAI211_X1 U16214 ( .C1(n14249), .C2(n14248), .A(n14247), .B(n14246), .ZN(
        P2_U3249) );
  NAND2_X1 U16215 ( .A1(n14250), .A2(n14258), .ZN(n14251) );
  NAND3_X1 U16216 ( .A1(n14253), .A2(n14252), .A3(n14251), .ZN(n14255) );
  INV_X1 U16217 ( .A(n14371), .ZN(n14256) );
  AOI21_X1 U16218 ( .B1(n14257), .B2(n14276), .A(n14256), .ZN(n14271) );
  XNOR2_X1 U16219 ( .A(n14259), .B(n14258), .ZN(n14372) );
  INV_X1 U16220 ( .A(n14372), .ZN(n14269) );
  NAND2_X1 U16221 ( .A1(n14260), .A2(n14433), .ZN(n14261) );
  NAND3_X1 U16222 ( .A1(n14263), .A2(n14262), .A3(n14261), .ZN(n14370) );
  AOI22_X1 U16223 ( .A1(n14433), .A2(n14278), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n14264), .ZN(n14265) );
  OAI21_X1 U16224 ( .B1(n14370), .B2(n14266), .A(n14265), .ZN(n14267) );
  AOI21_X1 U16225 ( .B1(n14269), .B2(n14268), .A(n14267), .ZN(n14270) );
  OAI21_X1 U16226 ( .B1(n14271), .B2(n14280), .A(n14270), .ZN(P2_U3250) );
  AOI22_X1 U16227 ( .A1(n14275), .A2(n14274), .B1(n14273), .B2(n14272), .ZN(
        n14285) );
  AOI22_X1 U16228 ( .A1(n14278), .A2(n14277), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n14276), .ZN(n14284) );
  INV_X1 U16229 ( .A(n14279), .ZN(n14282) );
  MUX2_X1 U16230 ( .A(n14282), .B(n14281), .S(n14280), .Z(n14283) );
  NAND3_X1 U16231 ( .A1(n14285), .A2(n14284), .A3(n14283), .ZN(P2_U3264) );
  NOR2_X1 U16232 ( .A1(n14288), .A2(n14287), .ZN(n14391) );
  MUX2_X1 U16233 ( .A(n14289), .B(n14391), .S(n15502), .Z(n14290) );
  OAI21_X1 U16234 ( .B1(n6841), .B2(n14362), .A(n14290), .ZN(P2_U3529) );
  AOI21_X1 U16235 ( .B1(n15479), .B2(n14292), .A(n14291), .ZN(n14293) );
  MUX2_X1 U16236 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14394), .S(n15502), .Z(
        P2_U3528) );
  NAND3_X1 U16237 ( .A1(n14297), .A2(n14366), .A3(n14296), .ZN(n14302) );
  NAND2_X1 U16238 ( .A1(n14298), .A2(n15479), .ZN(n14299) );
  NAND4_X1 U16239 ( .A1(n14302), .A2(n14301), .A3(n14300), .A4(n14299), .ZN(
        n14399) );
  MUX2_X1 U16240 ( .A(n14399), .B(P2_REG1_REG_27__SCAN_IN), .S(n15500), .Z(
        P2_U3526) );
  AOI21_X1 U16241 ( .B1(n15479), .B2(n7254), .A(n14303), .ZN(n14304) );
  OAI211_X1 U16242 ( .C1(n14386), .C2(n14306), .A(n14305), .B(n14304), .ZN(
        n14400) );
  MUX2_X1 U16243 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14400), .S(n15502), .Z(
        P2_U3525) );
  MUX2_X1 U16244 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14401), .S(n15502), .Z(
        n14310) );
  INV_X1 U16245 ( .A(n14310), .ZN(n14311) );
  OAI21_X1 U16246 ( .B1(n14404), .B2(n14362), .A(n14311), .ZN(P2_U3524) );
  NAND2_X1 U16247 ( .A1(n14312), .A2(n15479), .ZN(n14317) );
  NAND3_X1 U16248 ( .A1(n14314), .A2(n14313), .A3(n14366), .ZN(n14316) );
  NAND4_X1 U16249 ( .A1(n14318), .A2(n14317), .A3(n14316), .A4(n14315), .ZN(
        n14405) );
  MUX2_X1 U16250 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14405), .S(n15502), .Z(
        P2_U3523) );
  INV_X1 U16251 ( .A(n15479), .ZN(n15487) );
  OAI21_X1 U16252 ( .B1(n14320), .B2(n15487), .A(n14319), .ZN(n14321) );
  AOI21_X1 U16253 ( .B1(n14322), .B2(n14366), .A(n14321), .ZN(n14323) );
  AND2_X1 U16254 ( .A1(n14324), .A2(n14323), .ZN(n14406) );
  MUX2_X1 U16255 ( .A(n14325), .B(n14406), .S(n15502), .Z(n14326) );
  INV_X1 U16256 ( .A(n14326), .ZN(P2_U3522) );
  AOI211_X1 U16257 ( .C1(n14329), .C2(n14366), .A(n14328), .B(n14327), .ZN(
        n14408) );
  MUX2_X1 U16258 ( .A(n14330), .B(n14408), .S(n15502), .Z(n14331) );
  OAI21_X1 U16259 ( .B1(n14411), .B2(n14362), .A(n14331), .ZN(P2_U3521) );
  AOI211_X1 U16260 ( .C1(n14366), .C2(n14334), .A(n14333), .B(n14332), .ZN(
        n14412) );
  MUX2_X1 U16261 ( .A(n15668), .B(n14412), .S(n15502), .Z(n14335) );
  OAI21_X1 U16262 ( .B1(n7435), .B2(n14362), .A(n14335), .ZN(P2_U3520) );
  NAND2_X1 U16263 ( .A1(n14336), .A2(n15479), .ZN(n14337) );
  OAI211_X1 U16264 ( .C1(n14339), .C2(n14386), .A(n14338), .B(n14337), .ZN(
        n14340) );
  NOR2_X1 U16265 ( .A1(n14341), .A2(n14340), .ZN(n14415) );
  MUX2_X1 U16266 ( .A(n14342), .B(n14415), .S(n15502), .Z(n14343) );
  INV_X1 U16267 ( .A(n14343), .ZN(P2_U3519) );
  AOI211_X1 U16268 ( .C1(n14346), .C2(n14366), .A(n14345), .B(n14344), .ZN(
        n14418) );
  MUX2_X1 U16269 ( .A(n14347), .B(n14418), .S(n15502), .Z(n14348) );
  OAI21_X1 U16270 ( .B1(n14421), .B2(n14362), .A(n14348), .ZN(P2_U3518) );
  INV_X1 U16271 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14355) );
  NAND2_X1 U16272 ( .A1(n14349), .A2(n15476), .ZN(n14351) );
  OAI211_X1 U16273 ( .C1(n14352), .C2(n15487), .A(n14351), .B(n14350), .ZN(
        n14353) );
  NOR2_X1 U16274 ( .A1(n14354), .A2(n14353), .ZN(n14422) );
  MUX2_X1 U16275 ( .A(n14355), .B(n14422), .S(n15502), .Z(n14356) );
  INV_X1 U16276 ( .A(n14356), .ZN(P2_U3517) );
  INV_X1 U16277 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14360) );
  AOI211_X1 U16278 ( .C1(n14366), .C2(n14359), .A(n14358), .B(n14357), .ZN(
        n14425) );
  MUX2_X1 U16279 ( .A(n14360), .B(n14425), .S(n15502), .Z(n14361) );
  OAI21_X1 U16280 ( .B1(n14429), .B2(n14362), .A(n14361), .ZN(P2_U3516) );
  OAI22_X1 U16281 ( .A1(n14364), .A2(n14363), .B1(n6838), .B2(n15487), .ZN(
        n14365) );
  AOI21_X1 U16282 ( .B1(n14367), .B2(n14366), .A(n14365), .ZN(n14369) );
  NAND2_X1 U16283 ( .A1(n14369), .A2(n14368), .ZN(n14430) );
  MUX2_X1 U16284 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14430), .S(n15502), .Z(
        P2_U3515) );
  OAI211_X1 U16285 ( .C1(n14386), .C2(n14372), .A(n14371), .B(n14370), .ZN(
        n14431) );
  MUX2_X1 U16286 ( .A(n14431), .B(P2_REG1_REG_15__SCAN_IN), .S(n15500), .Z(
        n14373) );
  AOI21_X1 U16287 ( .B1(n14374), .B2(n14433), .A(n14373), .ZN(n14375) );
  INV_X1 U16288 ( .A(n14375), .ZN(P2_U3514) );
  AOI21_X1 U16289 ( .B1(n15479), .B2(n14377), .A(n14376), .ZN(n14378) );
  OAI211_X1 U16290 ( .C1(n14386), .C2(n14380), .A(n14379), .B(n14378), .ZN(
        n14436) );
  MUX2_X1 U16291 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14436), .S(n15502), .Z(
        P2_U3513) );
  AOI21_X1 U16292 ( .B1(n15479), .B2(n14382), .A(n14381), .ZN(n14383) );
  OAI211_X1 U16293 ( .C1(n14386), .C2(n14385), .A(n14384), .B(n14383), .ZN(
        n14437) );
  MUX2_X1 U16294 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14437), .S(n15502), .Z(
        P2_U3510) );
  INV_X1 U16295 ( .A(n14387), .ZN(n14390) );
  MUX2_X1 U16296 ( .A(n14392), .B(n14391), .S(n15494), .Z(n14393) );
  OAI21_X1 U16297 ( .B1(n6841), .B2(n14428), .A(n14393), .ZN(P2_U3497) );
  MUX2_X1 U16298 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14394), .S(n15494), .Z(
        P2_U3496) );
  OAI21_X1 U16299 ( .B1(n14398), .B2(n14428), .A(n14397), .ZN(P2_U3495) );
  MUX2_X1 U16300 ( .A(n14399), .B(P2_REG0_REG_27__SCAN_IN), .S(n15492), .Z(
        P2_U3494) );
  MUX2_X1 U16301 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14400), .S(n15494), .Z(
        P2_U3493) );
  MUX2_X1 U16302 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14401), .S(n15494), .Z(
        n14402) );
  INV_X1 U16303 ( .A(n14402), .ZN(n14403) );
  MUX2_X1 U16304 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14405), .S(n15494), .Z(
        P2_U3491) );
  INV_X1 U16305 ( .A(n14406), .ZN(n14407) );
  MUX2_X1 U16306 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14407), .S(n15494), .Z(
        P2_U3490) );
  INV_X1 U16307 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14409) );
  MUX2_X1 U16308 ( .A(n14409), .B(n14408), .S(n15494), .Z(n14410) );
  OAI21_X1 U16309 ( .B1(n14411), .B2(n14428), .A(n14410), .ZN(P2_U3489) );
  INV_X1 U16310 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14413) );
  MUX2_X1 U16311 ( .A(n14413), .B(n14412), .S(n15494), .Z(n14414) );
  OAI21_X1 U16312 ( .B1(n7435), .B2(n14428), .A(n14414), .ZN(P2_U3488) );
  INV_X1 U16313 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n14416) );
  MUX2_X1 U16314 ( .A(n14416), .B(n14415), .S(n15494), .Z(n14417) );
  INV_X1 U16315 ( .A(n14417), .ZN(P2_U3487) );
  INV_X1 U16316 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14419) );
  MUX2_X1 U16317 ( .A(n14419), .B(n14418), .S(n15494), .Z(n14420) );
  OAI21_X1 U16318 ( .B1(n14421), .B2(n14428), .A(n14420), .ZN(P2_U3486) );
  INV_X1 U16319 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14423) );
  MUX2_X1 U16320 ( .A(n14423), .B(n14422), .S(n15494), .Z(n14424) );
  INV_X1 U16321 ( .A(n14424), .ZN(P2_U3484) );
  INV_X1 U16322 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14426) );
  MUX2_X1 U16323 ( .A(n14426), .B(n14425), .S(n15494), .Z(n14427) );
  OAI21_X1 U16324 ( .B1(n14429), .B2(n14428), .A(n14427), .ZN(P2_U3481) );
  MUX2_X1 U16325 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14430), .S(n15494), .Z(
        P2_U3478) );
  MUX2_X1 U16326 ( .A(n14431), .B(P2_REG0_REG_15__SCAN_IN), .S(n15492), .Z(
        n14432) );
  AOI21_X1 U16327 ( .B1(n14434), .B2(n14433), .A(n14432), .ZN(n14435) );
  INV_X1 U16328 ( .A(n14435), .ZN(P2_U3475) );
  MUX2_X1 U16329 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14436), .S(n15494), .Z(
        P2_U3472) );
  MUX2_X1 U16330 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n14437), .S(n15494), .Z(
        P2_U3463) );
  INV_X1 U16331 ( .A(n14438), .ZN(n15142) );
  NOR4_X1 U16332 ( .A1(n14439), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14440), .A4(
        P2_U3088), .ZN(n14441) );
  AOI21_X1 U16333 ( .B1(n14445), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14441), 
        .ZN(n14442) );
  OAI21_X1 U16334 ( .B1(n15142), .B2(n14447), .A(n14442), .ZN(P2_U3296) );
  INV_X1 U16335 ( .A(n14443), .ZN(n15147) );
  AOI21_X1 U16336 ( .B1(n14445), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14444), 
        .ZN(n14446) );
  OAI21_X1 U16337 ( .B1(n15147), .B2(n14447), .A(n14446), .ZN(P2_U3299) );
  OAI222_X1 U16338 ( .A1(n12742), .A2(n14451), .B1(P2_U3088), .B2(n14449), 
        .C1(n14447), .C2(n14448), .ZN(P2_U3300) );
  INV_X1 U16339 ( .A(n14452), .ZN(n14453) );
  MUX2_X1 U16340 ( .A(n14453), .B(n15321), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  XNOR2_X1 U16341 ( .A(n14455), .B(n14454), .ZN(n14460) );
  AOI22_X1 U16342 ( .A1(n14604), .A2(n14560), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14457) );
  NAND2_X1 U16343 ( .A1(n14736), .A2(n14597), .ZN(n14456) );
  OAI211_X1 U16344 ( .C1(n14732), .C2(n14556), .A(n14457), .B(n14456), .ZN(
        n14458) );
  AOI21_X1 U16345 ( .B1(n14737), .B2(n14586), .A(n14458), .ZN(n14459) );
  OAI21_X1 U16346 ( .B1(n14460), .B2(n15237), .A(n14459), .ZN(P1_U3214) );
  INV_X1 U16347 ( .A(n14461), .ZN(n14462) );
  AOI21_X1 U16348 ( .B1(n14464), .B2(n14463), .A(n14462), .ZN(n14470) );
  OAI21_X1 U16349 ( .B1(n14556), .B2(n14917), .A(n14465), .ZN(n14466) );
  AOI21_X1 U16350 ( .B1(n14560), .B2(n14963), .A(n14466), .ZN(n14467) );
  OAI21_X1 U16351 ( .B1(n15246), .B2(n14947), .A(n14467), .ZN(n14468) );
  AOI21_X1 U16352 ( .B1(n15085), .B2(n14586), .A(n14468), .ZN(n14469) );
  OAI21_X1 U16353 ( .B1(n14470), .B2(n15237), .A(n14469), .ZN(P1_U3215) );
  XOR2_X1 U16354 ( .A(n14472), .B(n14471), .Z(n14477) );
  AOI22_X1 U16355 ( .A1(n14826), .A2(n14560), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14474) );
  NAND2_X1 U16356 ( .A1(n14796), .A2(n14597), .ZN(n14473) );
  OAI211_X1 U16357 ( .C1(n14798), .C2(n14556), .A(n14474), .B(n14473), .ZN(
        n14475) );
  AOI21_X1 U16358 ( .B1(n15025), .B2(n14586), .A(n14475), .ZN(n14476) );
  OAI21_X1 U16359 ( .B1(n14477), .B2(n15237), .A(n14476), .ZN(P1_U3216) );
  OAI211_X1 U16360 ( .C1(n14480), .C2(n14479), .A(n14478), .B(n14589), .ZN(
        n14484) );
  INV_X1 U16361 ( .A(n14858), .ZN(n14482) );
  AOI22_X1 U16362 ( .A1(n14825), .A2(n14960), .B1(n14962), .B2(n14889), .ZN(
        n15049) );
  NAND2_X1 U16363 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14691)
         );
  OAI21_X1 U16364 ( .B1(n15049), .B2(n14595), .A(n14691), .ZN(n14481) );
  AOI21_X1 U16365 ( .B1(n14482), .B2(n14597), .A(n14481), .ZN(n14483) );
  OAI211_X1 U16366 ( .C1(n7542), .C2(n14600), .A(n14484), .B(n14483), .ZN(
        P1_U3219) );
  AOI21_X1 U16367 ( .B1(n14487), .B2(n14486), .A(n14485), .ZN(n14493) );
  AOI22_X1 U16368 ( .A1(n14826), .A2(n14576), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14489) );
  NAND2_X1 U16369 ( .A1(n14597), .A2(n14831), .ZN(n14488) );
  OAI211_X1 U16370 ( .C1(n14490), .C2(n14579), .A(n14489), .B(n14488), .ZN(
        n14491) );
  AOI21_X1 U16371 ( .B1(n15036), .B2(n14586), .A(n14491), .ZN(n14492) );
  OAI21_X1 U16372 ( .B1(n14493), .B2(n15237), .A(n14492), .ZN(P1_U3223) );
  OAI211_X1 U16373 ( .C1(n6613), .C2(n14495), .A(n14494), .B(n14589), .ZN(
        n14502) );
  INV_X1 U16374 ( .A(n14496), .ZN(n14500) );
  OAI21_X1 U16375 ( .B1(n14595), .B2(n14498), .A(n14497), .ZN(n14499) );
  AOI21_X1 U16376 ( .B1(n14597), .B2(n14500), .A(n14499), .ZN(n14501) );
  OAI211_X1 U16377 ( .C1(n14503), .C2(n14600), .A(n14502), .B(n14501), .ZN(
        P1_U3224) );
  AOI22_X1 U16378 ( .A1(n14606), .A2(n14560), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14507) );
  NAND2_X1 U16379 ( .A1(n14764), .A2(n14597), .ZN(n14506) );
  OAI211_X1 U16380 ( .C1(n14765), .C2(n14556), .A(n14507), .B(n14506), .ZN(
        n14508) );
  AOI21_X1 U16381 ( .B1(n15012), .B2(n14586), .A(n14508), .ZN(n14509) );
  XNOR2_X1 U16382 ( .A(n14511), .B(n14510), .ZN(n14516) );
  XOR2_X1 U16383 ( .A(n14513), .B(n14514), .Z(n14592) );
  INV_X1 U16384 ( .A(n14512), .ZN(n14591) );
  NAND2_X1 U16385 ( .A1(n14592), .A2(n14591), .ZN(n14590) );
  OAI21_X1 U16386 ( .B1(n14514), .B2(n14513), .A(n14590), .ZN(n14515) );
  NOR2_X1 U16387 ( .A1(n14515), .A2(n14516), .ZN(n14526) );
  AOI21_X1 U16388 ( .B1(n14516), .B2(n14515), .A(n14526), .ZN(n14522) );
  NAND2_X1 U16389 ( .A1(n14597), .A2(n14919), .ZN(n14519) );
  AOI21_X1 U16390 ( .B1(n14576), .B2(n14610), .A(n14517), .ZN(n14518) );
  OAI211_X1 U16391 ( .C1(n14917), .C2(n14579), .A(n14519), .B(n14518), .ZN(
        n14520) );
  AOI21_X1 U16392 ( .B1(n15073), .B2(n14586), .A(n14520), .ZN(n14521) );
  OAI21_X1 U16393 ( .B1(n14522), .B2(n15237), .A(n14521), .ZN(P1_U3226) );
  INV_X1 U16394 ( .A(n14898), .ZN(n15066) );
  INV_X1 U16395 ( .A(n14523), .ZN(n14525) );
  NOR3_X1 U16396 ( .A1(n14526), .A2(n14525), .A3(n14524), .ZN(n14529) );
  INV_X1 U16397 ( .A(n14527), .ZN(n14528) );
  OAI21_X1 U16398 ( .B1(n14529), .B2(n14528), .A(n14589), .ZN(n14534) );
  NAND2_X1 U16399 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14664)
         );
  OAI21_X1 U16400 ( .B1(n14530), .B2(n14556), .A(n14664), .ZN(n14532) );
  NOR2_X1 U16401 ( .A1(n15246), .A2(n14891), .ZN(n14531) );
  AOI211_X1 U16402 ( .C1(n14560), .C2(n14887), .A(n14532), .B(n14531), .ZN(
        n14533) );
  OAI211_X1 U16403 ( .C1(n15066), .C2(n14600), .A(n14534), .B(n14533), .ZN(
        P1_U3228) );
  XOR2_X1 U16404 ( .A(n14536), .B(n14535), .Z(n14542) );
  NOR2_X1 U16405 ( .A1(n14784), .A2(n15065), .ZN(n15017) );
  AND2_X1 U16406 ( .A1(n14607), .A2(n14962), .ZN(n14537) );
  AOI21_X1 U16407 ( .B1(n14605), .B2(n14960), .A(n14537), .ZN(n14777) );
  INV_X1 U16408 ( .A(n14538), .ZN(n14782) );
  AOI22_X1 U16409 ( .A1(n14782), .A2(n14597), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14539) );
  OAI21_X1 U16410 ( .B1(n14777), .B2(n14595), .A(n14539), .ZN(n14540) );
  AOI21_X1 U16411 ( .B1(n15017), .B2(n15236), .A(n14540), .ZN(n14541) );
  OAI21_X1 U16412 ( .B1(n14542), .B2(n15237), .A(n14541), .ZN(P1_U3229) );
  OAI211_X1 U16413 ( .C1(n14545), .C2(n14544), .A(n14543), .B(n14589), .ZN(
        n14550) );
  INV_X1 U16414 ( .A(n14842), .ZN(n14548) );
  AOI22_X1 U16415 ( .A1(n14608), .A2(n14960), .B1(n14962), .B2(n14609), .ZN(
        n15041) );
  OAI22_X1 U16416 ( .A1(n15041), .A2(n14595), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14546), .ZN(n14547) );
  AOI21_X1 U16417 ( .B1(n14548), .B2(n14597), .A(n14547), .ZN(n14549) );
  OAI211_X1 U16418 ( .C1(n14846), .C2(n14600), .A(n14550), .B(n14549), .ZN(
        P1_U3233) );
  OAI211_X1 U16419 ( .C1(n14553), .C2(n14552), .A(n14551), .B(n14589), .ZN(
        n14562) );
  OAI21_X1 U16420 ( .B1(n14556), .B2(n14555), .A(n14554), .ZN(n14559) );
  NOR2_X1 U16421 ( .A1(n15246), .A2(n14557), .ZN(n14558) );
  AOI211_X1 U16422 ( .C1(n14560), .C2(n14613), .A(n14559), .B(n14558), .ZN(
        n14561) );
  OAI211_X1 U16423 ( .C1(n14563), .C2(n14600), .A(n14562), .B(n14561), .ZN(
        P1_U3234) );
  AOI21_X1 U16424 ( .B1(n14566), .B2(n14565), .A(n14564), .ZN(n14572) );
  OAI22_X1 U16425 ( .A1(n14568), .A2(n14916), .B1(n14567), .B2(n14918), .ZN(
        n14810) );
  AOI22_X1 U16426 ( .A1(n14810), .A2(n15241), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14569) );
  OAI21_X1 U16427 ( .B1(n15246), .B2(n14813), .A(n14569), .ZN(n14570) );
  AOI21_X1 U16428 ( .B1(n15030), .B2(n14586), .A(n14570), .ZN(n14571) );
  OAI21_X1 U16429 ( .B1(n14572), .B2(n15237), .A(n14571), .ZN(P1_U3235) );
  XOR2_X1 U16430 ( .A(n14573), .B(n14574), .Z(n14582) );
  NAND2_X1 U16431 ( .A1(n14597), .A2(n14875), .ZN(n14578) );
  NOR2_X1 U16432 ( .A1(n14575), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14674) );
  AOI21_X1 U16433 ( .B1(n14609), .B2(n14576), .A(n14674), .ZN(n14577) );
  OAI211_X1 U16434 ( .C1(n14915), .C2(n14579), .A(n14578), .B(n14577), .ZN(
        n14580) );
  AOI21_X1 U16435 ( .B1(n7159), .B2(n14586), .A(n14580), .ZN(n14581) );
  OAI21_X1 U16436 ( .B1(n14582), .B2(n15237), .A(n14581), .ZN(P1_U3238) );
  AOI22_X1 U16437 ( .A1(n14603), .A2(n14960), .B1(n14962), .B2(n14605), .ZN(
        n15001) );
  AOI22_X1 U16438 ( .A1(n14747), .A2(n14597), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14584) );
  OAI21_X1 U16439 ( .B1(n15001), .B2(n14595), .A(n14584), .ZN(n14585) );
  AOI21_X1 U16440 ( .B1(n14750), .B2(n14586), .A(n14585), .ZN(n14587) );
  OAI21_X1 U16441 ( .B1(n14588), .B2(n15237), .A(n14587), .ZN(P1_U3240) );
  OAI211_X1 U16442 ( .C1(n14592), .C2(n14591), .A(n14590), .B(n14589), .ZN(
        n14599) );
  INV_X1 U16443 ( .A(n14593), .ZN(n14935) );
  AND2_X1 U16444 ( .A1(n14612), .A2(n14962), .ZN(n14594) );
  AOI21_X1 U16445 ( .B1(n14887), .B2(n14960), .A(n14594), .ZN(n14933) );
  NAND2_X1 U16446 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15269)
         );
  OAI21_X1 U16447 ( .B1(n14933), .B2(n14595), .A(n15269), .ZN(n14596) );
  AOI21_X1 U16448 ( .B1(n14597), .B2(n14935), .A(n14596), .ZN(n14598) );
  OAI211_X1 U16449 ( .C1(n14938), .C2(n14600), .A(n14599), .B(n14598), .ZN(
        P1_U3241) );
  MUX2_X1 U16450 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14601), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16451 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14713), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16452 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14602), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16453 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14708), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16454 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14603), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16455 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14604), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16456 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14605), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16457 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14606), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16458 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14607), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16459 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14826), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16460 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14608), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16461 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14825), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16462 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14609), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16463 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14889), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16464 ( .A(n14610), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14611), .Z(
        P1_U3577) );
  MUX2_X1 U16465 ( .A(n14887), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14611), .Z(
        P1_U3576) );
  MUX2_X1 U16466 ( .A(n14961), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14611), .Z(
        P1_U3575) );
  MUX2_X1 U16467 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14612), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16468 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14963), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16469 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14613), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16470 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14614), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16471 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14615), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16472 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14616), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16473 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14617), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16474 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14618), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16475 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14619), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16476 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14620), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16477 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14621), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16478 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14622), .S(P1_U4016), .Z(
        P1_U3563) );
  INV_X1 U16479 ( .A(n14623), .ZN(n14624) );
  MUX2_X1 U16480 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14624), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16481 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14625), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16482 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14626), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16483 ( .C1(n14629), .C2(n14628), .A(n15266), .B(n14627), .ZN(
        n14638) );
  INV_X1 U16484 ( .A(n14630), .ZN(n14633) );
  OAI211_X1 U16485 ( .C1(n14633), .C2(n14632), .A(n15267), .B(n14631), .ZN(
        n14637) );
  AOI22_X1 U16486 ( .A1(n15255), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14636) );
  NAND2_X1 U16487 ( .A1(n15263), .A2(n14634), .ZN(n14635) );
  NAND4_X1 U16488 ( .A1(n14638), .A2(n14637), .A3(n14636), .A4(n14635), .ZN(
        P1_U3244) );
  AND2_X1 U16489 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14641) );
  NOR2_X1 U16490 ( .A1(n14686), .A2(n14639), .ZN(n14640) );
  AOI211_X1 U16491 ( .C1(n15255), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n14641), .B(
        n14640), .ZN(n14652) );
  OAI211_X1 U16492 ( .C1(n14644), .C2(n14643), .A(n15266), .B(n14642), .ZN(
        n14651) );
  OR3_X1 U16493 ( .A1(n14647), .A2(n14646), .A3(n14645), .ZN(n14648) );
  NAND3_X1 U16494 ( .A1(n15267), .A2(n14649), .A3(n14648), .ZN(n14650) );
  NAND3_X1 U16495 ( .A1(n14652), .A2(n14651), .A3(n14650), .ZN(P1_U3246) );
  AOI21_X1 U16496 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n14654), .A(n14653), 
        .ZN(n14656) );
  XNOR2_X1 U16497 ( .A(n14671), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14655) );
  NOR2_X1 U16498 ( .A1(n14656), .A2(n14655), .ZN(n14670) );
  AOI211_X1 U16499 ( .C1(n14656), .C2(n14655), .A(n14687), .B(n14670), .ZN(
        n14667) );
  NOR2_X1 U16500 ( .A1(n14657), .A2(n14908), .ZN(n14659) );
  MUX2_X1 U16501 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n14892), .S(n14671), .Z(
        n14658) );
  OAI21_X1 U16502 ( .B1(n14660), .B2(n14659), .A(n14658), .ZN(n14668) );
  INV_X1 U16503 ( .A(n14668), .ZN(n14662) );
  NOR3_X1 U16504 ( .A1(n14660), .A2(n14659), .A3(n14658), .ZN(n14661) );
  NOR3_X1 U16505 ( .A1(n14662), .A2(n14661), .A3(n14677), .ZN(n14666) );
  NAND2_X1 U16506 ( .A1(n15255), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n14663) );
  OAI211_X1 U16507 ( .C1(n14686), .C2(n14669), .A(n14664), .B(n14663), .ZN(
        n14665) );
  OR3_X1 U16508 ( .A1(n14667), .A2(n14666), .A3(n14665), .ZN(P1_U3260) );
  XNOR2_X1 U16509 ( .A(n14681), .B(n14876), .ZN(n14678) );
  NOR2_X1 U16510 ( .A1(n7292), .A2(n14672), .ZN(n14679) );
  OAI211_X1 U16511 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n6549), .A(n6442), .B(
        n15266), .ZN(n14676) );
  NOR2_X1 U16512 ( .A1(n14686), .A2(n14672), .ZN(n14673) );
  AOI211_X1 U16513 ( .C1(P1_ADDR_REG_18__SCAN_IN), .C2(n15255), .A(n14674), 
        .B(n14673), .ZN(n14675) );
  OAI211_X1 U16514 ( .C1(n14678), .C2(n14677), .A(n14676), .B(n14675), .ZN(
        P1_U3261) );
  XNOR2_X1 U16515 ( .A(n14680), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14689) );
  NAND2_X1 U16516 ( .A1(n14683), .A2(n14682), .ZN(n14684) );
  XOR2_X1 U16517 ( .A(n14685), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14688) );
  AOI22_X1 U16518 ( .A1(n14689), .A2(n15266), .B1(n15267), .B2(n14688), .ZN(
        n14690) );
  NAND2_X1 U16519 ( .A1(n14693), .A2(n14949), .ZN(n14971) );
  NOR2_X1 U16520 ( .A1(n14940), .A2(n14694), .ZN(n14698) );
  INV_X1 U16521 ( .A(P1_B_REG_SCAN_IN), .ZN(n14695) );
  NOR2_X1 U16522 ( .A1(n10115), .A2(n14695), .ZN(n14696) );
  OR2_X1 U16523 ( .A1(n14916), .A2(n14696), .ZN(n14714) );
  OR2_X1 U16524 ( .A1(n14714), .A2(n14697), .ZN(n14972) );
  NOR2_X1 U16525 ( .A1(n14920), .A2(n14972), .ZN(n14703) );
  AOI211_X1 U16526 ( .C1(n14699), .C2(n14956), .A(n14698), .B(n14703), .ZN(
        n14700) );
  OAI21_X1 U16527 ( .B1(n14971), .B2(n14953), .A(n14700), .ZN(P1_U3263) );
  OAI211_X1 U16528 ( .C1(n14712), .C2(n14974), .A(n14949), .B(n14701), .ZN(
        n14973) );
  NOR2_X1 U16529 ( .A1(n14940), .A2(n14702), .ZN(n14704) );
  AOI211_X1 U16530 ( .C1(n14705), .C2(n14956), .A(n14704), .B(n14703), .ZN(
        n14706) );
  OAI21_X1 U16531 ( .B1(n14973), .B2(n14953), .A(n14706), .ZN(P1_U3264) );
  OR2_X1 U16532 ( .A1(n14991), .A2(n14732), .ZN(n14977) );
  AND2_X1 U16533 ( .A1(n14991), .A2(n14732), .ZN(n14982) );
  AOI21_X1 U16534 ( .B1(n14976), .B2(n14977), .A(n14982), .ZN(n14707) );
  XNOR2_X1 U16535 ( .A(n14707), .B(n14980), .ZN(n14724) );
  XNOR2_X1 U16536 ( .A(n14711), .B(n14983), .ZN(n14984) );
  INV_X1 U16537 ( .A(n14713), .ZN(n14715) );
  OAI22_X1 U16538 ( .A1(n14732), .A2(n14918), .B1(n14715), .B2(n14714), .ZN(
        n14985) );
  AOI21_X1 U16539 ( .B1(n6433), .B2(n14716), .A(n14985), .ZN(n14721) );
  OAI22_X1 U16540 ( .A1(n14718), .A2(n14946), .B1(n14717), .B2(n14940), .ZN(
        n14719) );
  AOI21_X1 U16541 ( .B1(n14986), .B2(n14956), .A(n14719), .ZN(n14720) );
  OAI21_X1 U16542 ( .B1(n14721), .B2(n14920), .A(n14720), .ZN(n14722) );
  AOI21_X1 U16543 ( .B1(n14984), .B2(n14841), .A(n14722), .ZN(n14723) );
  OAI21_X1 U16544 ( .B1(n14724), .B2(n14754), .A(n14723), .ZN(P1_U3356) );
  OAI21_X1 U16545 ( .B1(n14726), .B2(n14728), .A(n14725), .ZN(n14727) );
  NAND2_X1 U16546 ( .A1(n14727), .A2(n15308), .ZN(n14734) );
  NAND2_X1 U16547 ( .A1(n14729), .A2(n14728), .ZN(n14730) );
  OAI22_X1 U16548 ( .A1(n14732), .A2(n14916), .B1(n14765), .B2(n14918), .ZN(
        n14733) );
  AOI21_X1 U16549 ( .B1(n14746), .B2(n14737), .A(n14893), .ZN(n14735) );
  NAND2_X1 U16550 ( .A1(n14735), .A2(n6413), .ZN(n14999) );
  AOI22_X1 U16551 ( .A1(n14736), .A2(n14934), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n14920), .ZN(n14739) );
  NAND2_X1 U16552 ( .A1(n14737), .A2(n14956), .ZN(n14738) );
  OAI211_X1 U16553 ( .C1(n14999), .C2(n14953), .A(n14739), .B(n14738), .ZN(
        n14740) );
  AOI21_X1 U16554 ( .B1(n14998), .B2(n14879), .A(n14740), .ZN(n14741) );
  OAI21_X1 U16555 ( .B1(n14742), .B2(n14920), .A(n14741), .ZN(P1_U3266) );
  XOR2_X1 U16556 ( .A(n14745), .B(n14743), .Z(n15008) );
  XOR2_X1 U16557 ( .A(n14745), .B(n14744), .Z(n15005) );
  OAI211_X1 U16558 ( .C1(n14762), .C2(n15003), .A(n14949), .B(n14746), .ZN(
        n15002) );
  AOI22_X1 U16559 ( .A1(n14747), .A2(n14934), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n14920), .ZN(n14748) );
  OAI21_X1 U16560 ( .B1(n15001), .B2(n14920), .A(n14748), .ZN(n14749) );
  AOI21_X1 U16561 ( .B1(n14750), .B2(n14956), .A(n14749), .ZN(n14751) );
  OAI21_X1 U16562 ( .B1(n15002), .B2(n14953), .A(n14751), .ZN(n14752) );
  AOI21_X1 U16563 ( .B1(n15005), .B2(n14841), .A(n14752), .ZN(n14753) );
  OAI21_X1 U16564 ( .B1(n15008), .B2(n14754), .A(n14753), .ZN(P1_U3267) );
  INV_X1 U16565 ( .A(n14755), .ZN(n14758) );
  INV_X1 U16566 ( .A(n14760), .ZN(n14757) );
  OAI21_X1 U16567 ( .B1(n14758), .B2(n14757), .A(n14756), .ZN(n15015) );
  OAI21_X1 U16568 ( .B1(n14761), .B2(n14760), .A(n14759), .ZN(n15009) );
  NAND2_X1 U16569 ( .A1(n15009), .A2(n14864), .ZN(n14771) );
  INV_X1 U16570 ( .A(n14779), .ZN(n14763) );
  AOI211_X1 U16571 ( .C1(n15012), .C2(n14763), .A(n14906), .B(n14762), .ZN(
        n15010) );
  AOI22_X1 U16572 ( .A1(n14764), .A2(n14934), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n14920), .ZN(n14767) );
  OAI22_X1 U16573 ( .A1(n14765), .A2(n14916), .B1(n14798), .B2(n14918), .ZN(
        n15011) );
  NAND2_X1 U16574 ( .A1(n15011), .A2(n14940), .ZN(n14766) );
  OAI211_X1 U16575 ( .C1(n14768), .C2(n14937), .A(n14767), .B(n14766), .ZN(
        n14769) );
  AOI21_X1 U16576 ( .B1(n15010), .B2(n14924), .A(n14769), .ZN(n14770) );
  OAI211_X1 U16577 ( .C1(n15015), .C2(n14969), .A(n14771), .B(n14770), .ZN(
        P1_U3268) );
  INV_X1 U16578 ( .A(n14772), .ZN(n14773) );
  AOI21_X1 U16579 ( .B1(n7849), .B2(n14774), .A(n14773), .ZN(n15021) );
  INV_X1 U16580 ( .A(n14775), .ZN(n14776) );
  OAI211_X1 U16581 ( .C1(n14776), .C2(n7849), .A(n15308), .B(n7851), .ZN(
        n15020) );
  INV_X1 U16582 ( .A(n15020), .ZN(n14778) );
  INV_X1 U16583 ( .A(n14777), .ZN(n15016) );
  OAI21_X1 U16584 ( .B1(n14778), .B2(n15016), .A(n14940), .ZN(n14787) );
  INV_X1 U16585 ( .A(n14795), .ZN(n14780) );
  AOI211_X1 U16586 ( .C1(n14781), .C2(n14780), .A(n14906), .B(n14779), .ZN(
        n15018) );
  AOI22_X1 U16587 ( .A1(n14782), .A2(n14934), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n14920), .ZN(n14783) );
  OAI21_X1 U16588 ( .B1(n14784), .B2(n14937), .A(n14783), .ZN(n14785) );
  AOI21_X1 U16589 ( .B1(n15018), .B2(n14924), .A(n14785), .ZN(n14786) );
  OAI211_X1 U16590 ( .C1(n15021), .C2(n14969), .A(n14787), .B(n14786), .ZN(
        P1_U3269) );
  OAI21_X1 U16591 ( .B1(n14788), .B2(n14805), .A(n14789), .ZN(n14791) );
  NAND2_X1 U16592 ( .A1(n14791), .A2(n14790), .ZN(n14792) );
  XNOR2_X1 U16593 ( .A(n14792), .B(n14793), .ZN(n15028) );
  XNOR2_X1 U16594 ( .A(n14794), .B(n14793), .ZN(n15022) );
  NAND2_X1 U16595 ( .A1(n15022), .A2(n14864), .ZN(n14803) );
  AOI211_X1 U16596 ( .C1(n15025), .C2(n6548), .A(n14893), .B(n14795), .ZN(
        n15023) );
  AOI22_X1 U16597 ( .A1(n14796), .A2(n14934), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n14920), .ZN(n14800) );
  OAI22_X1 U16598 ( .A1(n14798), .A2(n14916), .B1(n14797), .B2(n14918), .ZN(
        n15024) );
  NAND2_X1 U16599 ( .A1(n15024), .A2(n14940), .ZN(n14799) );
  OAI211_X1 U16600 ( .C1(n7554), .C2(n14937), .A(n14800), .B(n14799), .ZN(
        n14801) );
  AOI21_X1 U16601 ( .B1(n15023), .B2(n14924), .A(n14801), .ZN(n14802) );
  OAI211_X1 U16602 ( .C1(n15028), .C2(n14969), .A(n14803), .B(n14802), .ZN(
        P1_U3270) );
  NAND2_X1 U16603 ( .A1(n14788), .A2(n14804), .ZN(n14821) );
  NOR2_X1 U16604 ( .A1(n14821), .A2(n14824), .ZN(n14820) );
  NOR2_X1 U16605 ( .A1(n14820), .A2(n14805), .ZN(n14807) );
  XNOR2_X1 U16606 ( .A(n14807), .B(n14806), .ZN(n15033) );
  OAI21_X1 U16607 ( .B1(n14809), .B2(n6583), .A(n14808), .ZN(n14811) );
  AOI21_X1 U16608 ( .B1(n14811), .B2(n15308), .A(n14810), .ZN(n15032) );
  OAI22_X1 U16609 ( .A1(n14813), .A2(n14946), .B1(n14812), .B2(n14940), .ZN(
        n14814) );
  AOI21_X1 U16610 ( .B1(n15030), .B2(n14956), .A(n14814), .ZN(n14817) );
  AOI21_X1 U16611 ( .B1(n14829), .B2(n15030), .A(n14893), .ZN(n14815) );
  AND2_X1 U16612 ( .A1(n6548), .A2(n14815), .ZN(n15029) );
  NAND2_X1 U16613 ( .A1(n15029), .A2(n14924), .ZN(n14816) );
  OAI211_X1 U16614 ( .C1(n15032), .C2(n14920), .A(n14817), .B(n14816), .ZN(
        n14818) );
  INV_X1 U16615 ( .A(n14818), .ZN(n14819) );
  OAI21_X1 U16616 ( .B1(n15033), .B2(n14969), .A(n14819), .ZN(P1_U3271) );
  AOI21_X1 U16617 ( .B1(n14824), .B2(n14821), .A(n14820), .ZN(n15038) );
  OAI211_X1 U16618 ( .C1(n14824), .C2(n14823), .A(n14822), .B(n15308), .ZN(
        n14828) );
  AOI22_X1 U16619 ( .A1(n14826), .A2(n14960), .B1(n14962), .B2(n14825), .ZN(
        n14827) );
  NAND2_X1 U16620 ( .A1(n14828), .A2(n14827), .ZN(n15035) );
  INV_X1 U16621 ( .A(n15036), .ZN(n14834) );
  AOI21_X1 U16622 ( .B1(n14845), .B2(n15036), .A(n14893), .ZN(n14830) );
  AND2_X1 U16623 ( .A1(n14830), .A2(n14829), .ZN(n15034) );
  NAND2_X1 U16624 ( .A1(n15034), .A2(n14924), .ZN(n14833) );
  AOI22_X1 U16625 ( .A1(n14831), .A2(n14934), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n14920), .ZN(n14832) );
  OAI211_X1 U16626 ( .C1(n14834), .C2(n14937), .A(n14833), .B(n14832), .ZN(
        n14835) );
  AOI21_X1 U16627 ( .B1(n15035), .B2(n14940), .A(n14835), .ZN(n14836) );
  OAI21_X1 U16628 ( .B1(n15038), .B2(n14969), .A(n14836), .ZN(P1_U3272) );
  NAND2_X1 U16629 ( .A1(n14838), .A2(n14837), .ZN(n15039) );
  NAND3_X1 U16630 ( .A1(n15040), .A2(n15039), .A3(n14864), .ZN(n14850) );
  NAND2_X1 U16631 ( .A1(n14840), .A2(n14839), .ZN(n15044) );
  NAND3_X1 U16632 ( .A1(n14788), .A2(n14841), .A3(n15044), .ZN(n14849) );
  OAI22_X1 U16633 ( .A1(n15041), .A2(n14920), .B1(n14842), .B2(n14946), .ZN(
        n14844) );
  NOR2_X1 U16634 ( .A1(n14846), .A2(n14937), .ZN(n14843) );
  AOI211_X1 U16635 ( .C1(n14920), .C2(P1_REG2_REG_20__SCAN_IN), .A(n14844), 
        .B(n14843), .ZN(n14848) );
  OAI211_X1 U16636 ( .C1(n14855), .C2(n14846), .A(n14949), .B(n14845), .ZN(
        n15045) );
  OR2_X1 U16637 ( .A1(n15045), .A2(n14953), .ZN(n14847) );
  NAND4_X1 U16638 ( .A1(n14850), .A2(n14849), .A3(n14848), .A4(n14847), .ZN(
        P1_U3273) );
  XNOR2_X1 U16639 ( .A(n14851), .B(n14853), .ZN(n15054) );
  OAI21_X1 U16640 ( .B1(n14854), .B2(n14853), .A(n14852), .ZN(n15052) );
  INV_X1 U16641 ( .A(n14855), .ZN(n14856) );
  OAI211_X1 U16642 ( .C1(n7542), .C2(n6423), .A(n14856), .B(n14949), .ZN(
        n15050) );
  NOR2_X1 U16643 ( .A1(n14940), .A2(n14857), .ZN(n14860) );
  OAI22_X1 U16644 ( .A1(n15049), .A2(n14920), .B1(n14858), .B2(n14946), .ZN(
        n14859) );
  AOI211_X1 U16645 ( .C1(n6628), .C2(n14956), .A(n14860), .B(n14859), .ZN(
        n14862) );
  OAI21_X1 U16646 ( .B1(n15050), .B2(n14953), .A(n14862), .ZN(n14863) );
  AOI21_X1 U16647 ( .B1(n15052), .B2(n14864), .A(n14863), .ZN(n14865) );
  OAI21_X1 U16648 ( .B1(n15054), .B2(n14969), .A(n14865), .ZN(P1_U3274) );
  NOR2_X1 U16649 ( .A1(n14866), .A2(n14916), .ZN(n15057) );
  XNOR2_X1 U16650 ( .A(n14867), .B(n14870), .ZN(n15055) );
  NOR2_X1 U16651 ( .A1(n14885), .A2(n14886), .ZN(n14884) );
  NOR2_X1 U16652 ( .A1(n14884), .A2(n14868), .ZN(n14869) );
  XOR2_X1 U16653 ( .A(n14870), .B(n14869), .Z(n14871) );
  OAI22_X1 U16654 ( .A1(n14871), .A2(n15007), .B1(n14915), .B2(n14918), .ZN(
        n14872) );
  AOI21_X1 U16655 ( .B1(n14873), .B2(n15055), .A(n14872), .ZN(n15060) );
  INV_X1 U16656 ( .A(n15060), .ZN(n14874) );
  AOI211_X1 U16657 ( .C1(n14934), .C2(n14875), .A(n15057), .B(n14874), .ZN(
        n14882) );
  AOI211_X1 U16658 ( .C1(n7159), .C2(n14894), .A(n14893), .B(n6423), .ZN(
        n15056) );
  OAI22_X1 U16659 ( .A1(n14877), .A2(n14937), .B1(n14876), .B2(n14940), .ZN(
        n14878) );
  AOI21_X1 U16660 ( .B1(n15056), .B2(n14924), .A(n14878), .ZN(n14881) );
  NAND2_X1 U16661 ( .A1(n15055), .A2(n14879), .ZN(n14880) );
  OAI211_X1 U16662 ( .C1(n14882), .C2(n14920), .A(n14881), .B(n14880), .ZN(
        P1_U3275) );
  XNOR2_X1 U16663 ( .A(n14883), .B(n14886), .ZN(n15069) );
  INV_X1 U16664 ( .A(n15069), .ZN(n14901) );
  AOI211_X1 U16665 ( .C1(n14886), .C2(n14885), .A(n15007), .B(n14884), .ZN(
        n15067) );
  AND2_X1 U16666 ( .A1(n14887), .A2(n14962), .ZN(n14888) );
  AOI21_X1 U16667 ( .B1(n14889), .B2(n14960), .A(n14888), .ZN(n15063) );
  INV_X1 U16668 ( .A(n15063), .ZN(n14890) );
  OAI21_X1 U16669 ( .B1(n15067), .B2(n14890), .A(n14940), .ZN(n14900) );
  OAI22_X1 U16670 ( .A1(n14940), .A2(n14892), .B1(n14891), .B2(n14946), .ZN(
        n14897) );
  AOI21_X1 U16671 ( .B1(n14904), .B2(n14898), .A(n14893), .ZN(n14895) );
  NAND2_X1 U16672 ( .A1(n14895), .A2(n14894), .ZN(n15064) );
  NOR2_X1 U16673 ( .A1(n15064), .A2(n14953), .ZN(n14896) );
  AOI211_X1 U16674 ( .C1(n14956), .C2(n14898), .A(n14897), .B(n14896), .ZN(
        n14899) );
  OAI211_X1 U16675 ( .C1(n14901), .C2(n14969), .A(n14900), .B(n14899), .ZN(
        P1_U3276) );
  XNOR2_X1 U16676 ( .A(n14902), .B(n12689), .ZN(n15075) );
  INV_X1 U16677 ( .A(n14903), .ZN(n14907) );
  INV_X1 U16678 ( .A(n14904), .ZN(n14905) );
  AOI211_X1 U16679 ( .C1(n15073), .C2(n14907), .A(n14906), .B(n14905), .ZN(
        n15072) );
  OAI22_X1 U16680 ( .A1(n14909), .A2(n14937), .B1(n14940), .B2(n14908), .ZN(
        n14923) );
  INV_X1 U16681 ( .A(n14910), .ZN(n14911) );
  AOI21_X1 U16682 ( .B1(n14913), .B2(n14912), .A(n14911), .ZN(n14914) );
  OAI222_X1 U16683 ( .A1(n14918), .A2(n14917), .B1(n14916), .B2(n14915), .C1(
        n15007), .C2(n14914), .ZN(n15071) );
  AOI21_X1 U16684 ( .B1(n14919), .B2(n14934), .A(n15071), .ZN(n14921) );
  NOR2_X1 U16685 ( .A1(n14921), .A2(n14920), .ZN(n14922) );
  AOI211_X1 U16686 ( .C1(n15072), .C2(n14924), .A(n14923), .B(n14922), .ZN(
        n14925) );
  OAI21_X1 U16687 ( .B1(n14969), .B2(n15075), .A(n14925), .ZN(P1_U3277) );
  NOR2_X1 U16688 ( .A1(n14945), .A2(n14958), .ZN(n14944) );
  NOR2_X1 U16689 ( .A1(n14944), .A2(n14926), .ZN(n14928) );
  XNOR2_X1 U16690 ( .A(n14928), .B(n14927), .ZN(n15076) );
  INV_X1 U16691 ( .A(n15076), .ZN(n14943) );
  XNOR2_X1 U16692 ( .A(n14951), .B(n15078), .ZN(n14929) );
  NAND2_X1 U16693 ( .A1(n14929), .A2(n14949), .ZN(n15079) );
  OAI211_X1 U16694 ( .C1(n14932), .C2(n14931), .A(n14930), .B(n15308), .ZN(
        n15080) );
  INV_X1 U16695 ( .A(n14933), .ZN(n15077) );
  AOI21_X1 U16696 ( .B1(n14935), .B2(n14934), .A(n15077), .ZN(n14936) );
  OAI211_X1 U16697 ( .C1(n7274), .C2(n15079), .A(n15080), .B(n14936), .ZN(
        n14941) );
  OAI22_X1 U16698 ( .A1(n14938), .A2(n14937), .B1(n15260), .B2(n14940), .ZN(
        n14939) );
  AOI21_X1 U16699 ( .B1(n14941), .B2(n14940), .A(n14939), .ZN(n14942) );
  OAI21_X1 U16700 ( .B1(n14943), .B2(n14969), .A(n14942), .ZN(P1_U3278) );
  AOI21_X1 U16701 ( .B1(n14958), .B2(n14945), .A(n14944), .ZN(n15083) );
  INV_X1 U16702 ( .A(n15083), .ZN(n14970) );
  OAI22_X1 U16703 ( .A1(n14940), .A2(n12665), .B1(n14947), .B2(n14946), .ZN(
        n14955) );
  NAND2_X1 U16704 ( .A1(n14948), .A2(n15085), .ZN(n14950) );
  NAND2_X1 U16705 ( .A1(n14950), .A2(n14949), .ZN(n14952) );
  OR2_X1 U16706 ( .A1(n14952), .A2(n14951), .ZN(n15086) );
  NOR2_X1 U16707 ( .A1(n15086), .A2(n14953), .ZN(n14954) );
  AOI211_X1 U16708 ( .C1(n14956), .C2(n15085), .A(n14955), .B(n14954), .ZN(
        n14968) );
  OAI211_X1 U16709 ( .C1(n14959), .C2(n14958), .A(n14957), .B(n15308), .ZN(
        n15087) );
  INV_X1 U16710 ( .A(n15087), .ZN(n14966) );
  NAND2_X1 U16711 ( .A1(n14961), .A2(n14960), .ZN(n14965) );
  NAND2_X1 U16712 ( .A1(n14963), .A2(n14962), .ZN(n14964) );
  NAND2_X1 U16713 ( .A1(n14965), .A2(n14964), .ZN(n15084) );
  OAI21_X1 U16714 ( .B1(n14966), .B2(n15084), .A(n14940), .ZN(n14967) );
  OAI211_X1 U16715 ( .C1(n14970), .C2(n14969), .A(n14968), .B(n14967), .ZN(
        P1_U3279) );
  OAI211_X1 U16716 ( .C1(n6978), .C2(n15065), .A(n14971), .B(n14972), .ZN(
        n15113) );
  MUX2_X1 U16717 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15113), .S(n15316), .Z(
        P1_U3559) );
  OAI211_X1 U16718 ( .C1(n14974), .C2(n15065), .A(n14973), .B(n14972), .ZN(
        n15114) );
  MUX2_X1 U16719 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15114), .S(n15316), .Z(
        P1_U3558) );
  INV_X1 U16720 ( .A(n14982), .ZN(n14981) );
  INV_X1 U16721 ( .A(n14977), .ZN(n14978) );
  AOI21_X1 U16722 ( .B1(n14980), .B2(n14978), .A(n15007), .ZN(n14979) );
  NAND2_X1 U16723 ( .A1(n14984), .A2(n15297), .ZN(n14988) );
  OAI211_X1 U16724 ( .C1(n14990), .C2(n14989), .A(n14988), .B(n14987), .ZN(
        n15115) );
  MUX2_X1 U16725 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15115), .S(n15316), .Z(
        P1_U3557) );
  OAI21_X1 U16726 ( .B1(n6792), .B2(n15065), .A(n14992), .ZN(n14993) );
  AOI211_X1 U16727 ( .C1(n14995), .C2(n15297), .A(n14994), .B(n14993), .ZN(
        n14996) );
  OAI21_X1 U16728 ( .B1(n14997), .B2(n15007), .A(n14996), .ZN(n15116) );
  MUX2_X1 U16729 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15116), .S(n15316), .Z(
        P1_U3556) );
  MUX2_X1 U16730 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15117), .S(n15316), .Z(
        P1_U3555) );
  OAI211_X1 U16731 ( .C1(n15003), .C2(n15065), .A(n15002), .B(n15001), .ZN(
        n15004) );
  AOI21_X1 U16732 ( .B1(n15005), .B2(n15297), .A(n15004), .ZN(n15006) );
  OAI21_X1 U16733 ( .B1(n15008), .B2(n15007), .A(n15006), .ZN(n15118) );
  MUX2_X1 U16734 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15118), .S(n15316), .Z(
        P1_U3554) );
  NAND2_X1 U16735 ( .A1(n15009), .A2(n15308), .ZN(n15014) );
  AOI211_X1 U16736 ( .C1(n15302), .C2(n15012), .A(n15011), .B(n15010), .ZN(
        n15013) );
  OAI211_X1 U16737 ( .C1(n15304), .C2(n15015), .A(n15014), .B(n15013), .ZN(
        n15119) );
  MUX2_X1 U16738 ( .A(n15119), .B(P1_REG1_REG_25__SCAN_IN), .S(n15314), .Z(
        P1_U3553) );
  NOR3_X1 U16739 ( .A1(n15018), .A2(n15017), .A3(n15016), .ZN(n15019) );
  OAI211_X1 U16740 ( .C1(n15304), .C2(n15021), .A(n15020), .B(n15019), .ZN(
        n15120) );
  MUX2_X1 U16741 ( .A(n15120), .B(P1_REG1_REG_24__SCAN_IN), .S(n15314), .Z(
        P1_U3552) );
  NAND2_X1 U16742 ( .A1(n15022), .A2(n15308), .ZN(n15027) );
  AOI211_X1 U16743 ( .C1(n15302), .C2(n15025), .A(n15024), .B(n15023), .ZN(
        n15026) );
  OAI211_X1 U16744 ( .C1(n15304), .C2(n15028), .A(n15027), .B(n15026), .ZN(
        n15121) );
  MUX2_X1 U16745 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15121), .S(n15316), .Z(
        P1_U3551) );
  AOI21_X1 U16746 ( .B1(n15302), .B2(n15030), .A(n15029), .ZN(n15031) );
  OAI211_X1 U16747 ( .C1(n15033), .C2(n15304), .A(n15032), .B(n15031), .ZN(
        n15122) );
  MUX2_X1 U16748 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15122), .S(n15316), .Z(
        P1_U3550) );
  AOI211_X1 U16749 ( .C1(n15302), .C2(n15036), .A(n15035), .B(n15034), .ZN(
        n15037) );
  OAI21_X1 U16750 ( .B1(n15304), .B2(n15038), .A(n15037), .ZN(n15123) );
  MUX2_X1 U16751 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15123), .S(n15316), .Z(
        P1_U3549) );
  NAND3_X1 U16752 ( .A1(n15040), .A2(n15308), .A3(n15039), .ZN(n15048) );
  INV_X1 U16753 ( .A(n15041), .ZN(n15042) );
  AOI21_X1 U16754 ( .B1(n15043), .B2(n15302), .A(n15042), .ZN(n15047) );
  NAND3_X1 U16755 ( .A1(n14788), .A2(n15297), .A3(n15044), .ZN(n15046) );
  NAND4_X1 U16756 ( .A1(n15048), .A2(n15047), .A3(n15046), .A4(n15045), .ZN(
        n15124) );
  MUX2_X1 U16757 ( .A(n15124), .B(P1_REG1_REG_20__SCAN_IN), .S(n15314), .Z(
        P1_U3548) );
  OAI211_X1 U16758 ( .C1(n7542), .C2(n15065), .A(n15050), .B(n15049), .ZN(
        n15051) );
  AOI21_X1 U16759 ( .B1(n15052), .B2(n15308), .A(n15051), .ZN(n15053) );
  OAI21_X1 U16760 ( .B1(n15054), .B2(n15304), .A(n15053), .ZN(n15125) );
  MUX2_X1 U16761 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15125), .S(n15316), .Z(
        P1_U3547) );
  INV_X1 U16762 ( .A(n15055), .ZN(n15062) );
  AOI211_X1 U16763 ( .C1(n15302), .C2(n7159), .A(n15057), .B(n15056), .ZN(
        n15059) );
  OAI211_X1 U16764 ( .C1(n15062), .C2(n15061), .A(n15060), .B(n15059), .ZN(
        n15126) );
  MUX2_X1 U16765 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15126), .S(n15316), .Z(
        P1_U3546) );
  OAI211_X1 U16766 ( .C1(n15066), .C2(n15065), .A(n15064), .B(n15063), .ZN(
        n15068) );
  AOI211_X1 U16767 ( .C1(n15297), .C2(n15069), .A(n15068), .B(n15067), .ZN(
        n15070) );
  INV_X1 U16768 ( .A(n15070), .ZN(n15127) );
  MUX2_X1 U16769 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15127), .S(n15316), .Z(
        P1_U3545) );
  AOI211_X1 U16770 ( .C1(n15302), .C2(n15073), .A(n15072), .B(n15071), .ZN(
        n15074) );
  OAI21_X1 U16771 ( .B1(n15304), .B2(n15075), .A(n15074), .ZN(n15128) );
  MUX2_X1 U16772 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15128), .S(n15316), .Z(
        P1_U3544) );
  NAND2_X1 U16773 ( .A1(n15076), .A2(n15297), .ZN(n15082) );
  AOI21_X1 U16774 ( .B1(n15078), .B2(n15302), .A(n15077), .ZN(n15081) );
  NAND4_X1 U16775 ( .A1(n15082), .A2(n15081), .A3(n15080), .A4(n15079), .ZN(
        n15129) );
  MUX2_X1 U16776 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15129), .S(n15316), .Z(
        P1_U3543) );
  NAND2_X1 U16777 ( .A1(n15083), .A2(n15297), .ZN(n15089) );
  AOI21_X1 U16778 ( .B1(n15085), .B2(n15302), .A(n15084), .ZN(n15088) );
  NAND4_X1 U16779 ( .A1(n15089), .A2(n15088), .A3(n15087), .A4(n15086), .ZN(
        n15130) );
  MUX2_X1 U16780 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15130), .S(n15316), .Z(
        P1_U3542) );
  AOI211_X1 U16781 ( .C1(n15302), .C2(n15092), .A(n15091), .B(n15090), .ZN(
        n15093) );
  OAI21_X1 U16782 ( .B1(n15304), .B2(n15094), .A(n15093), .ZN(n15131) );
  MUX2_X1 U16783 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15131), .S(n15316), .Z(
        P1_U3541) );
  AOI211_X1 U16784 ( .C1(n15302), .C2(n15097), .A(n15096), .B(n15095), .ZN(
        n15098) );
  OAI21_X1 U16785 ( .B1(n15304), .B2(n15099), .A(n15098), .ZN(n15132) );
  MUX2_X1 U16786 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15132), .S(n15316), .Z(
        P1_U3540) );
  INV_X1 U16787 ( .A(n15100), .ZN(n15105) );
  NOR2_X1 U16788 ( .A1(n15102), .A2(n15101), .ZN(n15103) );
  OAI211_X1 U16789 ( .C1(n15304), .C2(n15105), .A(n15104), .B(n15103), .ZN(
        n15133) );
  MUX2_X1 U16790 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15133), .S(n15316), .Z(
        P1_U3539) );
  NOR4_X1 U16791 ( .A1(n15109), .A2(n15108), .A3(n15107), .A4(n15106), .ZN(
        n15110) );
  OAI21_X1 U16792 ( .B1(n15304), .B2(n15111), .A(n15110), .ZN(n15134) );
  MUX2_X1 U16793 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n15134), .S(n15316), .Z(
        P1_U3536) );
  MUX2_X1 U16794 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n15112), .S(n15316), .Z(
        P1_U3534) );
  MUX2_X1 U16795 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15113), .S(n15310), .Z(
        P1_U3527) );
  MUX2_X1 U16796 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15114), .S(n15310), .Z(
        P1_U3526) );
  MUX2_X1 U16797 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15115), .S(n15310), .Z(
        P1_U3525) );
  MUX2_X1 U16798 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15116), .S(n15310), .Z(
        P1_U3524) );
  MUX2_X1 U16799 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15117), .S(n15310), .Z(
        P1_U3523) );
  MUX2_X1 U16800 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15118), .S(n15310), .Z(
        P1_U3522) );
  MUX2_X1 U16801 ( .A(n15119), .B(P1_REG0_REG_25__SCAN_IN), .S(n15309), .Z(
        P1_U3521) );
  MUX2_X1 U16802 ( .A(n15120), .B(P1_REG0_REG_24__SCAN_IN), .S(n15309), .Z(
        P1_U3520) );
  MUX2_X1 U16803 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15121), .S(n15310), .Z(
        P1_U3519) );
  MUX2_X1 U16804 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15122), .S(n15310), .Z(
        P1_U3518) );
  MUX2_X1 U16805 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15123), .S(n15310), .Z(
        P1_U3517) );
  MUX2_X1 U16806 ( .A(n15124), .B(P1_REG0_REG_20__SCAN_IN), .S(n15309), .Z(
        P1_U3516) );
  MUX2_X1 U16807 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15125), .S(n15310), .Z(
        P1_U3515) );
  MUX2_X1 U16808 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15126), .S(n15310), .Z(
        P1_U3513) );
  MUX2_X1 U16809 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15127), .S(n15310), .Z(
        P1_U3510) );
  MUX2_X1 U16810 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15128), .S(n15310), .Z(
        P1_U3507) );
  MUX2_X1 U16811 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15129), .S(n15310), .Z(
        P1_U3504) );
  MUX2_X1 U16812 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15130), .S(n15310), .Z(
        P1_U3501) );
  MUX2_X1 U16813 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15131), .S(n15310), .Z(
        P1_U3498) );
  MUX2_X1 U16814 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15132), .S(n15310), .Z(
        P1_U3495) );
  MUX2_X1 U16815 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15133), .S(n15310), .Z(
        P1_U3492) );
  MUX2_X1 U16816 ( .A(P1_REG0_REG_8__SCAN_IN), .B(n15134), .S(n15310), .Z(
        P1_U3483) );
  NAND3_X1 U16817 ( .A1(n15135), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n15137) );
  OAI22_X1 U16818 ( .A1(n15138), .A2(n15137), .B1(n15136), .B2(n15149), .ZN(
        n15139) );
  INV_X1 U16819 ( .A(n15139), .ZN(n15140) );
  OAI21_X1 U16820 ( .B1(n15142), .B2(n15141), .A(n15140), .ZN(P1_U3324) );
  OAI222_X1 U16821 ( .A1(n15149), .A2(n15145), .B1(P1_U3086), .B2(n15144), 
        .C1(n15141), .C2(n15143), .ZN(P1_U3325) );
  OAI222_X1 U16822 ( .A1(n15149), .A2(n15148), .B1(n15141), .B2(n15147), .C1(
        P1_U3086), .C2(n15146), .ZN(P1_U3327) );
  MUX2_X1 U16823 ( .A(n15151), .B(n15150), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16824 ( .A(n15152), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U16825 ( .A(n15153), .B(n15154), .Z(SUB_1596_U59) );
  XOR2_X1 U16826 ( .A(n15155), .B(n15156), .Z(SUB_1596_U57) );
  XOR2_X1 U16827 ( .A(n15157), .B(n15158), .Z(SUB_1596_U56) );
  NAND2_X1 U16828 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15161), .ZN(n15162) );
  NAND2_X1 U16829 ( .A1(n15163), .A2(n15162), .ZN(n15166) );
  INV_X1 U16830 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15164) );
  NAND2_X1 U16831 ( .A1(n15164), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n15165) );
  NAND2_X1 U16832 ( .A1(n15166), .A2(n15165), .ZN(n15175) );
  INV_X1 U16833 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15167) );
  XNOR2_X1 U16834 ( .A(n15167), .B(P3_ADDR_REG_14__SCAN_IN), .ZN(n15174) );
  INV_X1 U16835 ( .A(n15174), .ZN(n15168) );
  XNOR2_X1 U16836 ( .A(n15175), .B(n15168), .ZN(n15169) );
  NAND2_X1 U16837 ( .A1(n15173), .A2(n15172), .ZN(n15171) );
  XNOR2_X1 U16838 ( .A(n15171), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  INV_X1 U16839 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15442) );
  INV_X1 U16840 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15176) );
  NAND2_X1 U16841 ( .A1(n15176), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U16842 ( .A1(n15178), .A2(n15177), .ZN(n15187) );
  XOR2_X1 U16843 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .Z(n15179) );
  XNOR2_X1 U16844 ( .A(n15187), .B(n15179), .ZN(n15180) );
  NAND2_X1 U16845 ( .A1(n15183), .A2(n15184), .ZN(n15181) );
  XNOR2_X1 U16846 ( .A(n15181), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  NAND2_X1 U16847 ( .A1(n15183), .A2(n15182), .ZN(n15185) );
  INV_X1 U16848 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15272) );
  NOR2_X1 U16849 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15272), .ZN(n15186) );
  NAND2_X1 U16850 ( .A1(n15272), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U16851 ( .A1(n15189), .A2(n15188), .ZN(n15202) );
  XOR2_X1 U16852 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(P3_ADDR_REG_16__SCAN_IN), 
        .Z(n15190) );
  XNOR2_X1 U16853 ( .A(n15202), .B(n15190), .ZN(n15191) );
  NAND2_X1 U16854 ( .A1(n15192), .A2(n15191), .ZN(n15198) );
  INV_X1 U16855 ( .A(n15198), .ZN(n15197) );
  INV_X1 U16856 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15193) );
  INV_X1 U16857 ( .A(n15194), .ZN(n15195) );
  OAI21_X1 U16858 ( .B1(n15195), .B2(n15197), .A(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n15196) );
  OAI21_X1 U16859 ( .B1(n15197), .B2(n15199), .A(n15196), .ZN(SUB_1596_U64) );
  INV_X1 U16860 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15200) );
  AND2_X1 U16861 ( .A1(n15200), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n15201) );
  OAI22_X1 U16862 ( .A1(n15202), .A2(n15201), .B1(P3_ADDR_REG_16__SCAN_IN), 
        .B2(n15200), .ZN(n15211) );
  XNOR2_X1 U16863 ( .A(n15211), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n15210) );
  XNOR2_X1 U16864 ( .A(n15210), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15203) );
  NAND2_X1 U16865 ( .A1(n15204), .A2(n15203), .ZN(n15208) );
  INV_X1 U16866 ( .A(n15208), .ZN(n15207) );
  OAI21_X1 U16867 ( .B1(n15205), .B2(n15207), .A(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n15206) );
  OAI21_X1 U16868 ( .B1(n15209), .B2(n15207), .A(n15206), .ZN(SUB_1596_U63) );
  INV_X1 U16869 ( .A(n15210), .ZN(n15213) );
  NOR2_X1 U16870 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15211), .ZN(n15212) );
  AOI21_X1 U16871 ( .B1(n15213), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n15212), 
        .ZN(n15222) );
  XNOR2_X1 U16872 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n15214) );
  XNOR2_X1 U16873 ( .A(n15222), .B(n15214), .ZN(n15215) );
  AOI21_X1 U16874 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15216), .A(n15219), 
        .ZN(n15217) );
  INV_X1 U16875 ( .A(n15217), .ZN(SUB_1596_U62) );
  AND2_X1 U16876 ( .A1(n15220), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n15221) );
  OAI22_X1 U16877 ( .A1(n15222), .A2(n15221), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n15220), .ZN(n15225) );
  XNOR2_X1 U16878 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P3_ADDR_REG_19__SCAN_IN), 
        .ZN(n15223) );
  XNOR2_X1 U16879 ( .A(n15223), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15224) );
  XNOR2_X1 U16880 ( .A(n15225), .B(n15224), .ZN(n15226) );
  XNOR2_X1 U16881 ( .A(n15227), .B(n15226), .ZN(SUB_1596_U4) );
  AOI21_X1 U16882 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15228) );
  OAI21_X1 U16883 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15228), 
        .ZN(U28) );
  AOI21_X1 U16884 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15229) );
  OAI21_X1 U16885 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15229), 
        .ZN(U29) );
  AND2_X1 U16886 ( .A1(n15231), .A2(n15230), .ZN(n15233) );
  XNOR2_X1 U16887 ( .A(n15233), .B(n15232), .ZN(SUB_1596_U61) );
  NAND2_X1 U16888 ( .A1(n15302), .A2(n15234), .ZN(n15277) );
  INV_X1 U16889 ( .A(n15277), .ZN(n15235) );
  AOI22_X1 U16890 ( .A1(n15236), .A2(n15235), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15245) );
  AOI21_X1 U16891 ( .B1(n15239), .B2(n15238), .A(n15237), .ZN(n15243) );
  AOI22_X1 U16892 ( .A1(n15243), .A2(n15242), .B1(n15241), .B2(n15240), .ZN(
        n15244) );
  OAI211_X1 U16893 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n15246), .A(n15245), .B(
        n15244), .ZN(P1_U3218) );
  NAND2_X1 U16894 ( .A1(n10115), .A2(n15247), .ZN(n15250) );
  NAND2_X1 U16895 ( .A1(n15248), .A2(n15250), .ZN(n15251) );
  MUX2_X1 U16896 ( .A(n15251), .B(n15250), .S(n15249), .Z(n15254) );
  INV_X1 U16897 ( .A(n15252), .ZN(n15253) );
  NAND2_X1 U16898 ( .A1(n15254), .A2(n15253), .ZN(n15257) );
  AOI22_X1 U16899 ( .A1(n15255), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15256) );
  OAI21_X1 U16900 ( .B1(n15258), .B2(n15257), .A(n15256), .ZN(P1_U3243) );
  OAI21_X1 U16901 ( .B1(n15261), .B2(n15260), .A(n15259), .ZN(n15268) );
  XNOR2_X1 U16902 ( .A(n15262), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n15265) );
  AOI222_X1 U16903 ( .A1(n15268), .A2(n15267), .B1(n15266), .B2(n15265), .C1(
        n15264), .C2(n15263), .ZN(n15270) );
  OAI211_X1 U16904 ( .C1(n15272), .C2(n15271), .A(n15270), .B(n15269), .ZN(
        P1_U3258) );
  AND2_X1 U16905 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15596), .ZN(P1_U3294) );
  AND2_X1 U16906 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15596), .ZN(P1_U3295) );
  AND2_X1 U16907 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15596), .ZN(P1_U3296) );
  INV_X1 U16908 ( .A(n15596), .ZN(n15273) );
  INV_X1 U16909 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15639) );
  NOR2_X1 U16910 ( .A1(n15273), .A2(n15639), .ZN(P1_U3297) );
  AND2_X1 U16911 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15596), .ZN(P1_U3298) );
  AND2_X1 U16912 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15596), .ZN(P1_U3299) );
  AND2_X1 U16913 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15596), .ZN(P1_U3300) );
  AND2_X1 U16914 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15596), .ZN(P1_U3301) );
  AND2_X1 U16915 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15596), .ZN(P1_U3302) );
  AND2_X1 U16916 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15596), .ZN(P1_U3303) );
  AND2_X1 U16917 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15596), .ZN(P1_U3304) );
  INV_X1 U16918 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15717) );
  NOR2_X1 U16919 ( .A1(n15273), .A2(n15717), .ZN(P1_U3305) );
  AND2_X1 U16920 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15596), .ZN(P1_U3306) );
  AND2_X1 U16921 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15596), .ZN(P1_U3307) );
  AND2_X1 U16922 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15596), .ZN(P1_U3308) );
  AND2_X1 U16923 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15596), .ZN(P1_U3309) );
  AND2_X1 U16924 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15596), .ZN(P1_U3310) );
  AND2_X1 U16925 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15596), .ZN(P1_U3311) );
  INV_X1 U16926 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15640) );
  NOR2_X1 U16927 ( .A1(n15273), .A2(n15640), .ZN(P1_U3312) );
  AND2_X1 U16928 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15596), .ZN(P1_U3313) );
  AND2_X1 U16929 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15596), .ZN(P1_U3314) );
  AND2_X1 U16930 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15596), .ZN(P1_U3315) );
  AND2_X1 U16931 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15596), .ZN(P1_U3316) );
  AND2_X1 U16932 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15596), .ZN(P1_U3317) );
  AND2_X1 U16933 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15596), .ZN(P1_U3318) );
  AND2_X1 U16934 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15596), .ZN(P1_U3319) );
  AND2_X1 U16935 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15596), .ZN(P1_U3321) );
  INV_X1 U16936 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15642) );
  NOR2_X1 U16937 ( .A1(n15273), .A2(n15642), .ZN(P1_U3322) );
  AND2_X1 U16938 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15596), .ZN(P1_U3323) );
  INV_X1 U16939 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15274) );
  AOI22_X1 U16940 ( .A1(n15310), .A2(n15275), .B1(n15274), .B2(n15309), .ZN(
        P1_U3459) );
  INV_X1 U16941 ( .A(n15276), .ZN(n15278) );
  NAND2_X1 U16942 ( .A1(n15278), .A2(n15277), .ZN(n15279) );
  AOI211_X1 U16943 ( .C1(n15282), .C2(n15281), .A(n15280), .B(n15279), .ZN(
        n15311) );
  INV_X1 U16944 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15283) );
  AOI22_X1 U16945 ( .A1(n15310), .A2(n15311), .B1(n15283), .B2(n15309), .ZN(
        P1_U3468) );
  INV_X1 U16946 ( .A(n15284), .ZN(n15286) );
  NAND4_X1 U16947 ( .A1(n15288), .A2(n15287), .A3(n15286), .A4(n15285), .ZN(
        n15289) );
  AOI21_X1 U16948 ( .B1(n15297), .B2(n15290), .A(n15289), .ZN(n15312) );
  INV_X1 U16949 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15729) );
  AOI22_X1 U16950 ( .A1(n15310), .A2(n15312), .B1(n15729), .B2(n15309), .ZN(
        P1_U3471) );
  OR3_X1 U16951 ( .A1(n15293), .A2(n15292), .A3(n15291), .ZN(n15295) );
  AOI211_X1 U16952 ( .C1(n15297), .C2(n15296), .A(n15295), .B(n15294), .ZN(
        n15313) );
  INV_X1 U16953 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15298) );
  AOI22_X1 U16954 ( .A1(n15310), .A2(n15313), .B1(n15298), .B2(n15309), .ZN(
        P1_U3474) );
  AOI211_X1 U16955 ( .C1(n15302), .C2(n15301), .A(n15300), .B(n15299), .ZN(
        n15303) );
  OAI21_X1 U16956 ( .B1(n15305), .B2(n15304), .A(n15303), .ZN(n15306) );
  AOI21_X1 U16957 ( .B1(n15308), .B2(n15307), .A(n15306), .ZN(n15315) );
  AOI22_X1 U16958 ( .A1(n15310), .A2(n15315), .B1(n9666), .B2(n15309), .ZN(
        P1_U3480) );
  AOI22_X1 U16959 ( .A1(n15316), .A2(n15311), .B1(n10694), .B2(n15314), .ZN(
        P1_U3531) );
  AOI22_X1 U16960 ( .A1(n15316), .A2(n15312), .B1(n9626), .B2(n15314), .ZN(
        P1_U3532) );
  AOI22_X1 U16961 ( .A1(n15316), .A2(n15313), .B1(n10695), .B2(n15314), .ZN(
        P1_U3533) );
  AOI22_X1 U16962 ( .A1(n15316), .A2(n15315), .B1(n10735), .B2(n15314), .ZN(
        P1_U3535) );
  NOR2_X1 U16963 ( .A1(n15336), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16964 ( .A1(n15451), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n15402), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15320) );
  AOI22_X1 U16965 ( .A1(n15336), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15319) );
  OAI22_X1 U16966 ( .A1(n15444), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n15411), .ZN(n15317) );
  OAI21_X1 U16967 ( .B1(n15450), .B2(n15317), .A(n15321), .ZN(n15318) );
  OAI211_X1 U16968 ( .C1(n15321), .C2(n15320), .A(n15319), .B(n15318), .ZN(
        P2_U3214) );
  OAI21_X1 U16969 ( .B1(n15323), .B2(n15322), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15324) );
  OAI21_X1 U16970 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15324), .ZN(n15335) );
  OAI211_X1 U16971 ( .C1(n15327), .C2(n15326), .A(n15402), .B(n15325), .ZN(
        n15328) );
  INV_X1 U16972 ( .A(n15328), .ZN(n15329) );
  AOI21_X1 U16973 ( .B1(n15336), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n15329), .ZN(
        n15334) );
  OAI211_X1 U16974 ( .C1(n15332), .C2(n15331), .A(n15451), .B(n15330), .ZN(
        n15333) );
  NAND3_X1 U16975 ( .A1(n15335), .A2(n15334), .A3(n15333), .ZN(P2_U3215) );
  AOI22_X1 U16976 ( .A1(n15336), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15348) );
  OAI211_X1 U16977 ( .C1(n15339), .C2(n15338), .A(n15402), .B(n15337), .ZN(
        n15340) );
  OAI21_X1 U16978 ( .B1(n15405), .B2(n15341), .A(n15340), .ZN(n15342) );
  INV_X1 U16979 ( .A(n15342), .ZN(n15347) );
  OAI211_X1 U16980 ( .C1(n15345), .C2(n15344), .A(n15451), .B(n15343), .ZN(
        n15346) );
  NAND3_X1 U16981 ( .A1(n15348), .A2(n15347), .A3(n15346), .ZN(P2_U3216) );
  INV_X1 U16982 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15362) );
  OAI211_X1 U16983 ( .C1(n15351), .C2(n15350), .A(n15402), .B(n15349), .ZN(
        n15356) );
  NAND2_X1 U16984 ( .A1(n15450), .A2(n15352), .ZN(n15355) );
  OR2_X1 U16985 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15353), .ZN(n15354) );
  AND3_X1 U16986 ( .A1(n15356), .A2(n15355), .A3(n15354), .ZN(n15361) );
  OAI211_X1 U16987 ( .C1(n15359), .C2(n15358), .A(n15451), .B(n15357), .ZN(
        n15360) );
  OAI211_X1 U16988 ( .C1(n15457), .C2(n15362), .A(n15361), .B(n15360), .ZN(
        P2_U3217) );
  OAI211_X1 U16989 ( .C1(n15365), .C2(n15364), .A(n15402), .B(n15363), .ZN(
        n15366) );
  OAI211_X1 U16990 ( .C1(n15405), .C2(n15368), .A(n15367), .B(n15366), .ZN(
        n15369) );
  INV_X1 U16991 ( .A(n15369), .ZN(n15374) );
  OAI211_X1 U16992 ( .C1(n15372), .C2(n15371), .A(n15451), .B(n15370), .ZN(
        n15373) );
  OAI211_X1 U16993 ( .C1(n15457), .C2(n11137), .A(n15374), .B(n15373), .ZN(
        P2_U3221) );
  INV_X1 U16994 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15387) );
  MUX2_X1 U16995 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n12221), .S(n15383), .Z(
        n15376) );
  OAI21_X1 U16996 ( .B1(n6461), .B2(n15376), .A(n15375), .ZN(n15384) );
  AND2_X1 U16997 ( .A1(n15378), .A2(n15377), .ZN(n15381) );
  OAI21_X1 U16998 ( .B1(n15381), .B2(n15380), .A(n15379), .ZN(n15382) );
  AOI222_X1 U16999 ( .A1(n15384), .A2(n15451), .B1(n15383), .B2(n15450), .C1(
        n15382), .C2(n15402), .ZN(n15386) );
  OAI211_X1 U17000 ( .C1(n15387), .C2(n15457), .A(n15386), .B(n15385), .ZN(
        P2_U3223) );
  INV_X1 U17001 ( .A(n15388), .ZN(n15394) );
  INV_X1 U17002 ( .A(n15389), .ZN(n15390) );
  AOI211_X1 U17003 ( .C1(n15392), .C2(n15391), .A(n15390), .B(n15444), .ZN(
        n15393) );
  AOI211_X1 U17004 ( .C1(n15450), .C2(n15395), .A(n15394), .B(n15393), .ZN(
        n15401) );
  AOI21_X1 U17005 ( .B1(n15397), .B2(n15396), .A(n15411), .ZN(n15399) );
  NAND2_X1 U17006 ( .A1(n15399), .A2(n15398), .ZN(n15400) );
  OAI211_X1 U17007 ( .C1(n15457), .C2(n6820), .A(n15401), .B(n15400), .ZN(
        P2_U3224) );
  OAI21_X1 U17008 ( .B1(n15404), .B2(n15403), .A(n15402), .ZN(n15408) );
  OAI22_X1 U17009 ( .A1(n15408), .A2(n15407), .B1(n15406), .B2(n15405), .ZN(
        n15415) );
  NAND2_X1 U17010 ( .A1(n15410), .A2(n15409), .ZN(n15412) );
  AOI21_X1 U17011 ( .B1(n15413), .B2(n15412), .A(n15411), .ZN(n15414) );
  NOR2_X1 U17012 ( .A1(n15415), .A2(n15414), .ZN(n15417) );
  OAI211_X1 U17013 ( .C1(n15607), .C2(n15457), .A(n15417), .B(n15416), .ZN(
        P2_U3225) );
  INV_X1 U17014 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15430) );
  INV_X1 U17015 ( .A(n15418), .ZN(n15423) );
  AOI211_X1 U17016 ( .C1(n15421), .C2(n15420), .A(n15444), .B(n15419), .ZN(
        n15422) );
  AOI211_X1 U17017 ( .C1(n15450), .C2(n15424), .A(n15423), .B(n15422), .ZN(
        n15429) );
  OAI211_X1 U17018 ( .C1(n15427), .C2(n15426), .A(n15425), .B(n15451), .ZN(
        n15428) );
  OAI211_X1 U17019 ( .C1(n15457), .C2(n15430), .A(n15429), .B(n15428), .ZN(
        P2_U3227) );
  INV_X1 U17020 ( .A(n15431), .ZN(n15436) );
  AOI211_X1 U17021 ( .C1(n15434), .C2(n15433), .A(n15444), .B(n15432), .ZN(
        n15435) );
  AOI211_X1 U17022 ( .C1(n15450), .C2(n15437), .A(n15436), .B(n15435), .ZN(
        n15441) );
  XOR2_X1 U17023 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n15438), .Z(n15439) );
  NAND2_X1 U17024 ( .A1(n15439), .A2(n15451), .ZN(n15440) );
  OAI211_X1 U17025 ( .C1(n15457), .C2(n15442), .A(n15441), .B(n15440), .ZN(
        P2_U3228) );
  AND2_X1 U17026 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15448) );
  AOI211_X1 U17027 ( .C1(n15446), .C2(n15445), .A(n15444), .B(n15443), .ZN(
        n15447) );
  AOI211_X1 U17028 ( .C1(n15450), .C2(n15449), .A(n15448), .B(n15447), .ZN(
        n15456) );
  OAI211_X1 U17029 ( .C1(n15454), .C2(n15453), .A(n15452), .B(n15451), .ZN(
        n15455) );
  OAI211_X1 U17030 ( .C1(n15457), .C2(n7151), .A(n15456), .B(n15455), .ZN(
        P2_U3231) );
  AND2_X1 U17031 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15460), .ZN(P2_U3266) );
  INV_X1 U17032 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15739) );
  NOR2_X1 U17033 ( .A1(n15459), .A2(n15739), .ZN(P2_U3267) );
  INV_X1 U17034 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15687) );
  NOR2_X1 U17035 ( .A1(n15459), .A2(n15687), .ZN(P2_U3268) );
  AND2_X1 U17036 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15460), .ZN(P2_U3269) );
  AND2_X1 U17037 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15460), .ZN(P2_U3270) );
  AND2_X1 U17038 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15460), .ZN(P2_U3271) );
  AND2_X1 U17039 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15460), .ZN(P2_U3272) );
  AND2_X1 U17040 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15460), .ZN(P2_U3273) );
  AND2_X1 U17041 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15460), .ZN(P2_U3274) );
  AND2_X1 U17042 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15460), .ZN(P2_U3275) );
  AND2_X1 U17043 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15460), .ZN(P2_U3276) );
  INV_X1 U17044 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15662) );
  NOR2_X1 U17045 ( .A1(n15459), .A2(n15662), .ZN(P2_U3277) );
  AND2_X1 U17046 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15460), .ZN(P2_U3278) );
  AND2_X1 U17047 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15460), .ZN(P2_U3279) );
  AND2_X1 U17048 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15460), .ZN(P2_U3280) );
  AND2_X1 U17049 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15460), .ZN(P2_U3281) );
  AND2_X1 U17050 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15460), .ZN(P2_U3282) );
  AND2_X1 U17051 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15460), .ZN(P2_U3283) );
  AND2_X1 U17052 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15460), .ZN(P2_U3284) );
  AND2_X1 U17053 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15460), .ZN(P2_U3285) );
  AND2_X1 U17054 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15460), .ZN(P2_U3286) );
  AND2_X1 U17055 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15460), .ZN(P2_U3287) );
  AND2_X1 U17056 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15460), .ZN(P2_U3288) );
  AND2_X1 U17057 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15460), .ZN(P2_U3289) );
  AND2_X1 U17058 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15460), .ZN(P2_U3290) );
  INV_X1 U17059 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15675) );
  NOR2_X1 U17060 ( .A1(n15459), .A2(n15675), .ZN(P2_U3291) );
  AND2_X1 U17061 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15460), .ZN(P2_U3292) );
  AND2_X1 U17062 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15460), .ZN(P2_U3293) );
  AND2_X1 U17063 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15460), .ZN(P2_U3294) );
  AND2_X1 U17064 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15460), .ZN(P2_U3295) );
  AOI22_X1 U17065 ( .A1(n15466), .A2(n15462), .B1(n15461), .B2(n15463), .ZN(
        P2_U3416) );
  AOI22_X1 U17066 ( .A1(n15466), .A2(n15465), .B1(n15464), .B2(n15463), .ZN(
        P2_U3417) );
  AOI211_X1 U17067 ( .C1(n15476), .C2(n15469), .A(n15468), .B(n15467), .ZN(
        n15496) );
  INV_X1 U17068 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15470) );
  AOI22_X1 U17069 ( .A1(n15494), .A2(n15496), .B1(n15470), .B2(n15492), .ZN(
        P2_U3430) );
  OAI21_X1 U17070 ( .B1(n15472), .B2(n15487), .A(n15471), .ZN(n15474) );
  AOI211_X1 U17071 ( .C1(n15476), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        n15498) );
  AOI22_X1 U17072 ( .A1(n15494), .A2(n15498), .B1(n8653), .B2(n15492), .ZN(
        P2_U3436) );
  AOI21_X1 U17073 ( .B1(n15479), .B2(n15478), .A(n15477), .ZN(n15480) );
  OAI211_X1 U17074 ( .C1(n15482), .C2(n15484), .A(n15481), .B(n15480), .ZN(
        n15483) );
  INV_X1 U17075 ( .A(n15483), .ZN(n15499) );
  AOI22_X1 U17076 ( .A1(n15494), .A2(n15499), .B1(n8707), .B2(n15492), .ZN(
        P2_U3442) );
  NOR2_X1 U17077 ( .A1(n15485), .A2(n15484), .ZN(n15490) );
  OAI21_X1 U17078 ( .B1(n15488), .B2(n15487), .A(n15486), .ZN(n15489) );
  NOR3_X1 U17079 ( .A1(n15491), .A2(n15490), .A3(n15489), .ZN(n15501) );
  INV_X1 U17080 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15493) );
  AOI22_X1 U17081 ( .A1(n15494), .A2(n15501), .B1(n15493), .B2(n15492), .ZN(
        P2_U3448) );
  INV_X1 U17082 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15495) );
  AOI22_X1 U17083 ( .A1(n15502), .A2(n15496), .B1(n15495), .B2(n15500), .ZN(
        P2_U3499) );
  AOI22_X1 U17084 ( .A1(n15502), .A2(n15498), .B1(n15497), .B2(n15500), .ZN(
        P2_U3501) );
  AOI22_X1 U17085 ( .A1(n15502), .A2(n15499), .B1(n8708), .B2(n15500), .ZN(
        P2_U3503) );
  AOI22_X1 U17086 ( .A1(n15502), .A2(n15501), .B1(n8760), .B2(n15500), .ZN(
        P2_U3505) );
  NOR2_X1 U17087 ( .A1(P3_U3897), .A2(n15503), .ZN(P3_U3150) );
  XNOR2_X1 U17088 ( .A(n15504), .B(n15511), .ZN(n15520) );
  INV_X1 U17089 ( .A(n15520), .ZN(n15557) );
  NOR2_X1 U17090 ( .A1(n15567), .A2(n15505), .ZN(n15556) );
  INV_X1 U17091 ( .A(n15556), .ZN(n15506) );
  OAI22_X1 U17092 ( .A1(n15509), .A2(n15508), .B1(n15507), .B2(n15506), .ZN(
        n15522) );
  OAI21_X1 U17093 ( .B1(n15512), .B2(n15511), .A(n15510), .ZN(n15518) );
  OAI22_X1 U17094 ( .A1(n15516), .A2(n15515), .B1(n15514), .B2(n15513), .ZN(
        n15517) );
  AOI21_X1 U17095 ( .B1(n15518), .B2(n15532), .A(n15517), .ZN(n15519) );
  OAI21_X1 U17096 ( .B1(n15521), .B2(n15520), .A(n15519), .ZN(n15555) );
  AOI211_X1 U17097 ( .C1(n15523), .C2(n15557), .A(n15522), .B(n15555), .ZN(
        n15525) );
  AOI22_X1 U17098 ( .A1(n15549), .A2(n6655), .B1(n15525), .B2(n15524), .ZN(
        P3_U3231) );
  NOR2_X1 U17099 ( .A1(n15567), .A2(n15526), .ZN(n15550) );
  XNOR2_X1 U17100 ( .A(n15527), .B(n15530), .ZN(n15551) );
  NAND2_X1 U17101 ( .A1(n15528), .A2(n15551), .ZN(n15541) );
  OAI21_X1 U17102 ( .B1(n15531), .B2(n15530), .A(n15529), .ZN(n15533) );
  NAND2_X1 U17103 ( .A1(n15533), .A2(n15532), .ZN(n15539) );
  AOI22_X1 U17104 ( .A1(n15537), .A2(n15536), .B1(n15535), .B2(n15534), .ZN(
        n15538) );
  AND2_X1 U17105 ( .A1(n15539), .A2(n15538), .ZN(n15540) );
  AND2_X1 U17106 ( .A1(n15541), .A2(n15540), .ZN(n15553) );
  INV_X1 U17107 ( .A(n15553), .ZN(n15542) );
  AOI21_X1 U17108 ( .B1(n15550), .B2(n15543), .A(n15542), .ZN(n15548) );
  AOI22_X1 U17109 ( .A1(n15545), .A2(n15551), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15544), .ZN(n15546) );
  OAI221_X1 U17110 ( .B1(n15549), .B2(n15548), .C1(n15524), .C2(n15547), .A(
        n15546), .ZN(P3_U3232) );
  AOI21_X1 U17111 ( .B1(n15551), .B2(n15579), .A(n15550), .ZN(n15552) );
  AND2_X1 U17112 ( .A1(n15553), .A2(n15552), .ZN(n15586) );
  INV_X1 U17113 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15554) );
  AOI22_X1 U17114 ( .A1(n15585), .A2(n15586), .B1(n15554), .B2(n15583), .ZN(
        P3_U3393) );
  AOI211_X1 U17115 ( .C1(n15557), .C2(n15579), .A(n15556), .B(n15555), .ZN(
        n15587) );
  INV_X1 U17116 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15558) );
  AOI22_X1 U17117 ( .A1(n15585), .A2(n15587), .B1(n15558), .B2(n15583), .ZN(
        P3_U3396) );
  INV_X1 U17118 ( .A(n15559), .ZN(n15560) );
  AOI211_X1 U17119 ( .C1(n15579), .C2(n15562), .A(n15561), .B(n15560), .ZN(
        n15589) );
  INV_X1 U17120 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15563) );
  AOI22_X1 U17121 ( .A1(n15585), .A2(n15589), .B1(n15563), .B2(n15583), .ZN(
        P3_U3399) );
  INV_X1 U17122 ( .A(n15564), .ZN(n15570) );
  OAI21_X1 U17123 ( .B1(n15567), .B2(n15566), .A(n15565), .ZN(n15568) );
  AOI21_X1 U17124 ( .B1(n15570), .B2(n15569), .A(n15568), .ZN(n15590) );
  INV_X1 U17125 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15571) );
  AOI22_X1 U17126 ( .A1(n15585), .A2(n15590), .B1(n15571), .B2(n15583), .ZN(
        P3_U3402) );
  INV_X1 U17127 ( .A(n15572), .ZN(n15575) );
  AND2_X1 U17128 ( .A1(n15573), .A2(n15579), .ZN(n15574) );
  NOR3_X1 U17129 ( .A1(n15576), .A2(n15575), .A3(n15574), .ZN(n15592) );
  INV_X1 U17130 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15577) );
  AOI22_X1 U17131 ( .A1(n15585), .A2(n15592), .B1(n15577), .B2(n15583), .ZN(
        P3_U3405) );
  AOI21_X1 U17132 ( .B1(n15580), .B2(n15579), .A(n15578), .ZN(n15581) );
  AND2_X1 U17133 ( .A1(n15582), .A2(n15581), .ZN(n15594) );
  INV_X1 U17134 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15584) );
  AOI22_X1 U17135 ( .A1(n15585), .A2(n15594), .B1(n15584), .B2(n15583), .ZN(
        P3_U3408) );
  AOI22_X1 U17136 ( .A1(n15595), .A2(n15586), .B1(n11117), .B2(n15593), .ZN(
        P3_U3460) );
  AOI22_X1 U17137 ( .A1(n15595), .A2(n15587), .B1(n11114), .B2(n15593), .ZN(
        P3_U3461) );
  INV_X1 U17138 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15588) );
  AOI22_X1 U17139 ( .A1(n15595), .A2(n15589), .B1(n15588), .B2(n15593), .ZN(
        P3_U3462) );
  AOI22_X1 U17140 ( .A1(n15595), .A2(n15590), .B1(n11245), .B2(n15593), .ZN(
        P3_U3463) );
  INV_X1 U17141 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15591) );
  AOI22_X1 U17142 ( .A1(n15595), .A2(n15592), .B1(n15591), .B2(n15593), .ZN(
        P3_U3464) );
  AOI22_X1 U17143 ( .A1(n15595), .A2(n15594), .B1(n11304), .B2(n15593), .ZN(
        P3_U3465) );
  NAND2_X1 U17144 ( .A1(n15596), .A2(P1_D_REG_5__SCAN_IN), .ZN(n15751) );
  AND4_X1 U17145 ( .A1(P3_REG0_REG_27__SCAN_IN), .A2(n15728), .A3(n15734), 
        .A4(n15729), .ZN(n15602) );
  NAND4_X1 U17146 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(P2_REG0_REG_4__SCAN_IN), 
        .A3(P1_REG0_REG_10__SCAN_IN), .A4(P3_DATAO_REG_8__SCAN_IN), .ZN(n15599) );
  INV_X1 U17147 ( .A(SI_4_), .ZN(n15597) );
  NAND3_X1 U17148 ( .A1(n15597), .A2(P2_IR_REG_30__SCAN_IN), .A3(
        P1_REG3_REG_12__SCAN_IN), .ZN(n15598) );
  NOR2_X1 U17149 ( .A1(n15599), .A2(n15598), .ZN(n15601) );
  AND4_X1 U17150 ( .A1(P2_REG1_REG_29__SCAN_IN), .A2(P3_REG3_REG_8__SCAN_IN), 
        .A3(P1_D_REG_20__SCAN_IN), .A4(n15714), .ZN(n15600) );
  AND4_X1 U17151 ( .A1(n15602), .A2(n15739), .A3(n15601), .A4(n15600), .ZN(
        n15749) );
  NAND4_X1 U17152 ( .A1(SI_17_), .A2(P1_IR_REG_30__SCAN_IN), .A3(
        P1_REG3_REG_17__SCAN_IN), .A4(n15627), .ZN(n15622) );
  NOR4_X1 U17153 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_5__SCAN_IN), .A4(n7149), .ZN(n15604) );
  NOR4_X1 U17154 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(SI_3_), .A3(n15639), .A4(
        n15624), .ZN(n15603) );
  NAND4_X1 U17155 ( .A1(n15606), .A2(n15605), .A3(n15604), .A4(n15603), .ZN(
        n15621) );
  INV_X1 U17156 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15672) );
  NOR4_X1 U17157 ( .A1(n15669), .A2(n15671), .A3(n15672), .A4(n15607), .ZN(
        n15613) );
  NOR4_X1 U17158 ( .A1(P3_D_REG_23__SCAN_IN), .A2(SI_11_), .A3(n15662), .A4(
        n15651), .ZN(n15612) );
  NOR4_X1 U17159 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(n15637), .A3(n15643), 
        .A4(n15655), .ZN(n15608) );
  NAND3_X1 U17160 ( .A1(n15674), .A2(P2_IR_REG_13__SCAN_IN), .A3(n15608), .ZN(
        n15610) );
  NOR3_X1 U17161 ( .A1(n15610), .A2(n15609), .A3(P2_IR_REG_4__SCAN_IN), .ZN(
        n15611) );
  NAND3_X1 U17162 ( .A1(n15613), .A2(n15612), .A3(n15611), .ZN(n15620) );
  NOR4_X1 U17163 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n12671), .A4(n15689), .ZN(n15618) );
  NOR4_X1 U17164 ( .A1(n10863), .A2(n10693), .A3(n15700), .A4(n15703), .ZN(
        n15615) );
  NOR4_X1 U17165 ( .A1(P3_REG2_REG_24__SCAN_IN), .A2(SI_29_), .A3(n15692), 
        .A4(n15702), .ZN(n15614) );
  NAND4_X1 U17166 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(n15615), .A3(n15614), 
        .A4(P1_REG3_REG_1__SCAN_IN), .ZN(n15616) );
  NOR3_X1 U17167 ( .A1(n15616), .A2(P2_REG1_REG_21__SCAN_IN), .A3(
        P3_DATAO_REG_28__SCAN_IN), .ZN(n15617) );
  NAND2_X1 U17168 ( .A1(n15618), .A2(n15617), .ZN(n15619) );
  NOR4_X1 U17169 ( .A1(n15622), .A2(n15621), .A3(n15620), .A4(n15619), .ZN(
        n15748) );
  AOI22_X1 U17170 ( .A1(n15624), .A2(keyinput50), .B1(keyinput34), .B2(n7149), 
        .ZN(n15623) );
  OAI221_X1 U17171 ( .B1(n15624), .B2(keyinput50), .C1(n7149), .C2(keyinput34), 
        .A(n15623), .ZN(n15634) );
  AOI22_X1 U17172 ( .A1(n15627), .A2(keyinput3), .B1(n15626), .B2(keyinput9), 
        .ZN(n15625) );
  OAI221_X1 U17173 ( .B1(n15627), .B2(keyinput3), .C1(n15626), .C2(keyinput9), 
        .A(n15625), .ZN(n15633) );
  XOR2_X1 U17174 ( .A(n15135), .B(keyinput40), .Z(n15631) );
  XNOR2_X1 U17175 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput23), .ZN(n15630) );
  XNOR2_X1 U17176 ( .A(P1_REG3_REG_17__SCAN_IN), .B(keyinput41), .ZN(n15629)
         );
  XNOR2_X1 U17177 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput28), .ZN(n15628)
         );
  NAND4_X1 U17178 ( .A1(n15631), .A2(n15630), .A3(n15629), .A4(n15628), .ZN(
        n15632) );
  NOR3_X1 U17179 ( .A1(n15634), .A2(n15633), .A3(n15632), .ZN(n15685) );
  AOI22_X1 U17180 ( .A1(n15637), .A2(keyinput57), .B1(keyinput59), .B2(n15636), 
        .ZN(n15635) );
  OAI221_X1 U17181 ( .B1(n15637), .B2(keyinput57), .C1(n15636), .C2(keyinput59), .A(n15635), .ZN(n15649) );
  AOI22_X1 U17182 ( .A1(n15640), .A2(keyinput21), .B1(keyinput33), .B2(n15639), 
        .ZN(n15638) );
  OAI221_X1 U17183 ( .B1(n15640), .B2(keyinput21), .C1(n15639), .C2(keyinput33), .A(n15638), .ZN(n15648) );
  AOI22_X1 U17184 ( .A1(n15643), .A2(keyinput47), .B1(keyinput36), .B2(n15642), 
        .ZN(n15641) );
  OAI221_X1 U17185 ( .B1(n15643), .B2(keyinput47), .C1(n15642), .C2(keyinput36), .A(n15641), .ZN(n15647) );
  XOR2_X1 U17186 ( .A(n7357), .B(keyinput8), .Z(n15645) );
  XNOR2_X1 U17187 ( .A(SI_3_), .B(keyinput54), .ZN(n15644) );
  NAND2_X1 U17188 ( .A1(n15645), .A2(n15644), .ZN(n15646) );
  NOR4_X1 U17189 ( .A1(n15649), .A2(n15648), .A3(n15647), .A4(n15646), .ZN(
        n15684) );
  AOI22_X1 U17190 ( .A1(n15652), .A2(keyinput19), .B1(keyinput12), .B2(n15651), 
        .ZN(n15650) );
  OAI221_X1 U17191 ( .B1(n15652), .B2(keyinput19), .C1(n15651), .C2(keyinput12), .A(n15650), .ZN(n15653) );
  INV_X1 U17192 ( .A(n15653), .ZN(n15666) );
  AOI22_X1 U17193 ( .A1(n15656), .A2(keyinput2), .B1(keyinput1), .B2(n15655), 
        .ZN(n15654) );
  OAI221_X1 U17194 ( .B1(n15656), .B2(keyinput2), .C1(n15655), .C2(keyinput1), 
        .A(n15654), .ZN(n15657) );
  INV_X1 U17195 ( .A(n15657), .ZN(n15665) );
  XNOR2_X1 U17196 ( .A(P3_REG1_REG_24__SCAN_IN), .B(keyinput6), .ZN(n15660) );
  XNOR2_X1 U17197 ( .A(SI_11_), .B(keyinput37), .ZN(n15659) );
  XNOR2_X1 U17198 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput51), .ZN(n15658) );
  AND3_X1 U17199 ( .A1(n15660), .A2(n15659), .A3(n15658), .ZN(n15664) );
  INV_X1 U17200 ( .A(keyinput10), .ZN(n15661) );
  XNOR2_X1 U17201 ( .A(n15662), .B(n15661), .ZN(n15663) );
  AND4_X1 U17202 ( .A1(n15666), .A2(n15665), .A3(n15664), .A4(n15663), .ZN(
        n15683) );
  AOI22_X1 U17203 ( .A1(n15669), .A2(keyinput35), .B1(n15668), .B2(keyinput25), 
        .ZN(n15667) );
  OAI221_X1 U17204 ( .B1(n15669), .B2(keyinput35), .C1(n15668), .C2(keyinput25), .A(n15667), .ZN(n15681) );
  AOI22_X1 U17205 ( .A1(n15672), .A2(keyinput5), .B1(n15671), .B2(keyinput20), 
        .ZN(n15670) );
  OAI221_X1 U17206 ( .B1(n15672), .B2(keyinput5), .C1(n15671), .C2(keyinput20), 
        .A(n15670), .ZN(n15680) );
  AOI22_X1 U17207 ( .A1(n15675), .A2(keyinput42), .B1(keyinput15), .B2(n15674), 
        .ZN(n15673) );
  OAI221_X1 U17208 ( .B1(n15675), .B2(keyinput42), .C1(n15674), .C2(keyinput15), .A(n15673), .ZN(n15679) );
  XNOR2_X1 U17209 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(keyinput55), .ZN(n15677)
         );
  XNOR2_X1 U17210 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput63), .ZN(n15676) );
  NAND2_X1 U17211 ( .A1(n15677), .A2(n15676), .ZN(n15678) );
  NOR4_X1 U17212 ( .A1(n15681), .A2(n15680), .A3(n15679), .A4(n15678), .ZN(
        n15682) );
  NAND4_X1 U17213 ( .A1(n15685), .A2(n15684), .A3(n15683), .A4(n15682), .ZN(
        n15747) );
  AOI22_X1 U17214 ( .A1(n15687), .A2(keyinput60), .B1(keyinput39), .B2(n12671), 
        .ZN(n15686) );
  OAI221_X1 U17215 ( .B1(n15687), .B2(keyinput60), .C1(n12671), .C2(keyinput39), .A(n15686), .ZN(n15698) );
  AOI22_X1 U17216 ( .A1(n15690), .A2(keyinput27), .B1(keyinput62), .B2(n15689), 
        .ZN(n15688) );
  OAI221_X1 U17217 ( .B1(n15690), .B2(keyinput27), .C1(n15689), .C2(keyinput62), .A(n15688), .ZN(n15697) );
  AOI22_X1 U17218 ( .A1(n8328), .A2(keyinput30), .B1(n15692), .B2(keyinput13), 
        .ZN(n15691) );
  OAI221_X1 U17219 ( .B1(n8328), .B2(keyinput30), .C1(n15692), .C2(keyinput13), 
        .A(n15691), .ZN(n15696) );
  XOR2_X1 U17220 ( .A(n9571), .B(keyinput49), .Z(n15694) );
  XNOR2_X1 U17221 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput11), .ZN(n15693) );
  NAND2_X1 U17222 ( .A1(n15694), .A2(n15693), .ZN(n15695) );
  NOR4_X1 U17223 ( .A1(n15698), .A2(n15697), .A3(n15696), .A4(n15695), .ZN(
        n15745) );
  AOI22_X1 U17224 ( .A1(n15700), .A2(keyinput32), .B1(n10693), .B2(keyinput45), 
        .ZN(n15699) );
  OAI221_X1 U17225 ( .B1(n15700), .B2(keyinput32), .C1(n10693), .C2(keyinput45), .A(n15699), .ZN(n15711) );
  AOI22_X1 U17226 ( .A1(n15703), .A2(keyinput16), .B1(n15702), .B2(keyinput44), 
        .ZN(n15701) );
  OAI221_X1 U17227 ( .B1(n15703), .B2(keyinput16), .C1(n15702), .C2(keyinput44), .A(n15701), .ZN(n15710) );
  AOI22_X1 U17228 ( .A1(n15705), .A2(keyinput48), .B1(n9577), .B2(keyinput14), 
        .ZN(n15704) );
  OAI221_X1 U17229 ( .B1(n15705), .B2(keyinput48), .C1(n9577), .C2(keyinput14), 
        .A(n15704), .ZN(n15709) );
  XNOR2_X1 U17230 ( .A(P1_REG3_REG_11__SCAN_IN), .B(keyinput43), .ZN(n15707)
         );
  XNOR2_X1 U17231 ( .A(keyinput29), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n15706) );
  NAND2_X1 U17232 ( .A1(n15707), .A2(n15706), .ZN(n15708) );
  NOR4_X1 U17233 ( .A1(n15711), .A2(n15710), .A3(n15709), .A4(n15708), .ZN(
        n15744) );
  INV_X1 U17234 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15713) );
  AOI22_X1 U17235 ( .A1(n15714), .A2(keyinput56), .B1(keyinput53), .B2(n15713), 
        .ZN(n15712) );
  OAI221_X1 U17236 ( .B1(n15714), .B2(keyinput56), .C1(n15713), .C2(keyinput53), .A(n15712), .ZN(n15726) );
  AOI22_X1 U17237 ( .A1(n15717), .A2(keyinput22), .B1(n15716), .B2(keyinput26), 
        .ZN(n15715) );
  OAI221_X1 U17238 ( .B1(n15717), .B2(keyinput22), .C1(n15716), .C2(keyinput26), .A(n15715), .ZN(n15725) );
  AOI22_X1 U17239 ( .A1(n15719), .A2(keyinput61), .B1(keyinput4), .B2(n8707), 
        .ZN(n15718) );
  OAI221_X1 U17240 ( .B1(n15719), .B2(keyinput61), .C1(n8707), .C2(keyinput4), 
        .A(n15718), .ZN(n15724) );
  AOI22_X1 U17241 ( .A1(n15722), .A2(keyinput52), .B1(keyinput31), .B2(n15721), 
        .ZN(n15720) );
  OAI221_X1 U17242 ( .B1(n15722), .B2(keyinput52), .C1(n15721), .C2(keyinput31), .A(n15720), .ZN(n15723) );
  NOR4_X1 U17243 ( .A1(n15726), .A2(n15725), .A3(n15724), .A4(n15723), .ZN(
        n15743) );
  AOI22_X1 U17244 ( .A1(n15729), .A2(keyinput24), .B1(n15728), .B2(keyinput0), 
        .ZN(n15727) );
  OAI221_X1 U17245 ( .B1(n15729), .B2(keyinput24), .C1(n15728), .C2(keyinput0), 
        .A(n15727), .ZN(n15738) );
  AOI22_X1 U17246 ( .A1(n8608), .A2(keyinput38), .B1(keyinput58), .B2(n15731), 
        .ZN(n15730) );
  OAI221_X1 U17247 ( .B1(n8608), .B2(keyinput38), .C1(n15731), .C2(keyinput58), 
        .A(n15730), .ZN(n15737) );
  AOI22_X1 U17248 ( .A1(n15734), .A2(keyinput7), .B1(n15733), .B2(keyinput46), 
        .ZN(n15732) );
  OAI221_X1 U17249 ( .B1(n15734), .B2(keyinput7), .C1(n15733), .C2(keyinput46), 
        .A(n15732), .ZN(n15736) );
  XOR2_X1 U17250 ( .A(SI_4_), .B(keyinput18), .Z(n15735) );
  NOR4_X1 U17251 ( .A1(n15738), .A2(n15737), .A3(n15736), .A4(n15735), .ZN(
        n15741) );
  XOR2_X1 U17252 ( .A(keyinput17), .B(n15739), .Z(n15740) );
  AND2_X1 U17253 ( .A1(n15741), .A2(n15740), .ZN(n15742) );
  NAND4_X1 U17254 ( .A1(n15745), .A2(n15744), .A3(n15743), .A4(n15742), .ZN(
        n15746) );
  AOI211_X1 U17255 ( .C1(n15749), .C2(n15748), .A(n15747), .B(n15746), .ZN(
        n15750) );
  XNOR2_X1 U17256 ( .A(n15751), .B(n15750), .ZN(P1_U3320) );
  XNOR2_X1 U17257 ( .A(n15753), .B(n15752), .ZN(n15754) );
  XNOR2_X1 U17258 ( .A(n15754), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U17259 ( .A(n15756), .B(n15755), .Z(SUB_1596_U5) );
  INV_X2 U7478 ( .A(n10015), .ZN(n9591) );
  BUF_X1 U7385 ( .A(n8675), .Z(n8950) );
  CLKBUF_X1 U7183 ( .A(n8965), .Z(n9244) );
  NOR2_X1 U7186 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n7884) );
  NAND2_X2 U7236 ( .A1(n6405), .A2(n10572), .ZN(n8070) );
  CLKBUF_X1 U7263 ( .A(n10459), .Z(n6400) );
  CLKBUF_X2 U7395 ( .A(n11096), .Z(n6405) );
  CLKBUF_X2 U7949 ( .A(n7991), .Z(n8363) );
  AND2_X1 U8036 ( .A1(n10436), .A2(n10435), .ZN(n12913) );
  CLKBUF_X1 U9305 ( .A(n10377), .Z(n7136) );
  CLKBUF_X1 U9563 ( .A(n9349), .Z(n14241) );
  XNOR2_X1 U9625 ( .A(n7999), .B(P3_IR_REG_2__SCAN_IN), .ZN(n11239) );
  CLKBUF_X1 U10261 ( .A(n13477), .Z(n6668) );
endmodule

