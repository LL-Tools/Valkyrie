

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n5011, n5012, n5013, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5737, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10983,
         n10984, n10985;

  OR2_X1 U5075 ( .A1(n7081), .A2(n7080), .ZN(n5109) );
  INV_X1 U5076 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n10983) );
  OR2_X1 U5077 ( .A1(n8211), .A2(n10753), .ZN(n7916) );
  INV_X1 U5079 ( .A(n6464), .ZN(n6499) );
  CLKBUF_X2 U5080 ( .A(n6179), .Z(n6352) );
  CLKBUF_X1 U5081 ( .A(n6357), .Z(n6284) );
  INV_X1 U5082 ( .A(n5824), .ZN(n5905) );
  INV_X2 U5083 ( .A(n7652), .ZN(n8732) );
  BUF_X1 U5085 ( .A(n5933), .Z(n8750) );
  INV_X1 U5086 ( .A(n10366), .ZN(n10740) );
  INV_X2 U5088 ( .A(n10985), .ZN(n5011) );
  INV_X1 U5090 ( .A(n10983), .ZN(n5012) );
  INV_X1 U5091 ( .A(n5012), .ZN(n5013) );
  INV_X1 U5092 ( .A(n5012), .ZN(P1_U3084) );
  AND2_X1 U5093 ( .A1(n5939), .A2(n5304), .ZN(n6464) );
  AOI21_X1 U5094 ( .B1(n10356), .B2(n10030), .A(n9975), .ZN(n10345) );
  INV_X1 U5095 ( .A(n6031), .ZN(n6254) );
  AND2_X1 U5096 ( .A1(n9548), .A2(n5225), .ZN(n5052) );
  NAND2_X1 U5097 ( .A1(n9550), .A2(n5484), .ZN(n9528) );
  INV_X1 U5098 ( .A(n7475), .ZN(n7279) );
  INV_X1 U5100 ( .A(n8823), .ZN(n6942) );
  INV_X1 U5101 ( .A(n6034), .ZN(n6311) );
  OAI21_X1 U5102 ( .B1(n8545), .B2(n5226), .A(n5052), .ZN(n6467) );
  INV_X1 U5103 ( .A(n10744), .ZN(n8014) );
  NAND2_X1 U5104 ( .A1(n5842), .A2(n5841), .ZN(n10753) );
  INV_X2 U5105 ( .A(n6575), .ZN(n5724) );
  AOI21_X1 U5106 ( .B1(n10353), .B2(n10357), .A(n8759), .ZN(n10340) );
  XNOR2_X2 U5107 ( .A(n5928), .B(n5927), .ZN(n6004) );
  XNOR2_X2 U5108 ( .A(n6549), .B(n6548), .ZN(n8794) );
  NAND2_X2 U5109 ( .A1(n6547), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6549) );
  NAND2_X2 U5110 ( .A1(n8559), .A2(n6431), .ZN(n8602) );
  XNOR2_X2 U5111 ( .A(n5770), .B(n5769), .ZN(n8545) );
  AOI21_X2 U5112 ( .B1(n6358), .B2(n6494), .A(n5475), .ZN(n6359) );
  OAI21_X2 U5113 ( .B1(n7764), .B2(n7765), .A(n6388), .ZN(n8205) );
  NAND2_X2 U5114 ( .A1(n6330), .A2(n6382), .ZN(n7764) );
  OAI21_X2 U5115 ( .B1(n6364), .B2(n6522), .A(n6495), .ZN(n6366) );
  AOI21_X2 U5116 ( .B1(n9755), .B2(n6360), .A(n6359), .ZN(n6364) );
  AOI21_X2 U5117 ( .B1(n5440), .B2(n5438), .A(n5437), .ZN(n5436) );
  OR2_X2 U5118 ( .A1(n5443), .A2(n5441), .ZN(n5440) );
  INV_X1 U5119 ( .A(n7912), .ZN(n8356) );
  OAI211_X2 U5120 ( .C1(n7475), .C2(n7521), .A(n5826), .B(n5825), .ZN(n7912)
         );
  XNOR2_X2 U5121 ( .A(n8455), .B(n10753), .ZN(n7954) );
  INV_X4 U5122 ( .A(n7009), .ZN(n6977) );
  NAND2_X2 U5123 ( .A1(n6708), .A2(n6585), .ZN(n7009) );
  OR2_X1 U5124 ( .A1(n6674), .A2(n6673), .ZN(n7945) );
  AND2_X1 U5125 ( .A1(n6402), .A2(n6398), .ZN(n8078) );
  NAND2_X1 U5126 ( .A1(n10064), .A2(n10037), .ZN(n10162) );
  INV_X1 U5127 ( .A(n10811), .ZN(n8304) );
  INV_X4 U5128 ( .A(n6764), .ZN(n7058) );
  NAND2_X2 U5129 ( .A1(n7160), .A2(n7843), .ZN(n6764) );
  OR2_X1 U5130 ( .A1(n9396), .A2(n8356), .ZN(n6388) );
  INV_X1 U5131 ( .A(n7903), .ZN(n7832) );
  CLKBUF_X1 U5132 ( .A(n7829), .Z(n10053) );
  NAND4_X1 U5133 ( .A1(n6622), .A2(n6621), .A3(n6620), .A4(n6619), .ZN(n10210)
         );
  INV_X1 U5134 ( .A(n7843), .ZN(n7123) );
  AOI21_X1 U5135 ( .B1(n5268), .B2(n9644), .A(n5266), .ZN(n9671) );
  OAI21_X1 U5136 ( .B1(n8840), .B2(n10178), .A(n8839), .ZN(n10460) );
  NAND2_X1 U5137 ( .A1(n8840), .A2(n10178), .ZN(n8839) );
  AND2_X1 U5138 ( .A1(n9314), .A2(n6265), .ZN(n9371) );
  OAI21_X1 U5139 ( .B1(n9292), .B2(n9291), .A(n5607), .ZN(n6252) );
  NAND2_X1 U5140 ( .A1(n6749), .A2(n5591), .ZN(n8328) );
  OAI21_X2 U5141 ( .B1(n8630), .B2(n5384), .A(n5382), .ZN(n8709) );
  NAND2_X1 U5142 ( .A1(n5224), .A2(n5771), .ZN(n9700) );
  INV_X1 U5143 ( .A(n5246), .ZN(n5245) );
  AND2_X1 U5144 ( .A1(n8224), .A2(n8330), .ZN(n5591) );
  NAND2_X1 U5145 ( .A1(n5775), .A2(n5774), .ZN(n9705) );
  NAND2_X1 U5146 ( .A1(n5779), .A2(n5778), .ZN(n9557) );
  AOI21_X1 U5147 ( .B1(n7945), .B2(n7944), .A(n6675), .ZN(n7940) );
  OR2_X1 U5148 ( .A1(n6292), .A2(n8934), .ZN(n8811) );
  OAI21_X1 U5149 ( .B1(n5777), .B2(n5682), .A(n5684), .ZN(n5773) );
  NAND2_X1 U5150 ( .A1(n6929), .A2(n6928), .ZN(n10426) );
  NOR2_X1 U5151 ( .A1(n10168), .A2(n5406), .ZN(n5405) );
  INV_X1 U5152 ( .A(n9512), .ZN(n9548) );
  NAND2_X1 U5153 ( .A1(n5808), .A2(n5807), .ZN(n9744) );
  OAI21_X1 U5154 ( .B1(n5902), .B2(n5669), .A(n5668), .ZN(n5789) );
  INV_X1 U5155 ( .A(n8078), .ZN(n5015) );
  NAND2_X1 U5156 ( .A1(n6774), .A2(n6773), .ZN(n10828) );
  INV_X2 U5157 ( .A(n10822), .ZN(n10969) );
  NAND2_X1 U5158 ( .A1(n5247), .A2(n5853), .ZN(n8463) );
  INV_X1 U5159 ( .A(n8146), .ZN(n5305) );
  NAND2_X2 U5160 ( .A1(n8252), .A2(n10819), .ZN(n10822) );
  NAND2_X1 U5161 ( .A1(n5525), .A2(n8034), .ZN(n6505) );
  NAND4_X2 U5162 ( .A1(n6051), .A2(n6050), .A3(n6049), .A4(n6048), .ZN(n8455)
         );
  NAND2_X1 U5163 ( .A1(n6640), .A2(n5599), .ZN(n10209) );
  OAI211_X1 U5164 ( .C1(n5623), .C2(n5215), .A(n5060), .B(n5214), .ZN(n5855)
         );
  NOR2_X1 U5165 ( .A1(n6159), .A2(n6158), .ZN(n5110) );
  NAND4_X2 U5166 ( .A1(n6011), .A2(n6010), .A3(n6009), .A4(n6008), .ZN(n7404)
         );
  INV_X2 U5167 ( .A(n6699), .ZN(n7810) );
  NAND2_X2 U5168 ( .A1(n7124), .A2(n7123), .ZN(n7652) );
  XNOR2_X1 U5169 ( .A(n6559), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7085) );
  OAI211_X1 U5170 ( .C1(n7140), .C2(n7373), .A(n6628), .B(n6627), .ZN(n7903)
         );
  NAND4_X1 U5171 ( .A1(n6608), .A2(n6607), .A3(n6606), .A4(n6605), .ZN(n7830)
         );
  NAND2_X1 U5172 ( .A1(n6576), .A2(n5398), .ZN(n7654) );
  NAND2_X1 U5173 ( .A1(n5138), .A2(n5620), .ZN(n5837) );
  INV_X1 U5174 ( .A(n7117), .ZN(n6656) );
  NAND2_X1 U5175 ( .A1(n6558), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6559) );
  AND2_X1 U5176 ( .A1(n10049), .A2(n8327), .ZN(n7843) );
  INV_X1 U5177 ( .A(n8240), .ZN(n8108) );
  NAND2_X1 U5178 ( .A1(n5139), .A2(n5617), .ZN(n5833) );
  NAND2_X1 U5179 ( .A1(n6563), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6560) );
  AND2_X1 U5180 ( .A1(n5039), .A2(n5126), .ZN(n8240) );
  NAND2_X2 U5181 ( .A1(n7155), .A2(n7126), .ZN(n7140) );
  CLKBUF_X2 U5182 ( .A(n5934), .Z(n8833) );
  AND2_X1 U5183 ( .A1(n5939), .A2(n8350), .ZN(n10702) );
  NAND2_X1 U5184 ( .A1(n5926), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5928) );
  XNOR2_X1 U5185 ( .A(n6570), .B(n6569), .ZN(n7126) );
  XNOR2_X1 U5186 ( .A(n5929), .B(n9789), .ZN(n5934) );
  NAND2_X1 U5187 ( .A1(n5615), .A2(n5614), .ZN(n5823) );
  XNOR2_X1 U5188 ( .A(n5923), .B(n5922), .ZN(n8350) );
  XNOR2_X1 U5189 ( .A(n5950), .B(n5949), .ZN(n5939) );
  NAND2_X1 U5190 ( .A1(n9792), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5929) );
  NAND2_X4 U5191 ( .A1(n5941), .A2(n5940), .ZN(n7475) );
  NAND2_X1 U5192 ( .A1(n5027), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U5193 ( .A1(n5920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5950) );
  OR2_X1 U5194 ( .A1(n5946), .A2(n5956), .ZN(n5742) );
  NAND2_X2 U5195 ( .A1(n5724), .A2(P2_U3152), .ZN(n8831) );
  OR2_X1 U5196 ( .A1(n5782), .A2(n5783), .ZN(n5017) );
  INV_X4 U5197 ( .A(n5608), .ZN(n6575) );
  NAND3_X1 U5198 ( .A1(n5734), .A2(n5829), .A3(n5735), .ZN(n5782) );
  AND2_X2 U5199 ( .A1(n5814), .A2(n5270), .ZN(n5829) );
  NOR2_X1 U5200 ( .A1(n6541), .A2(n6540), .ZN(n6542) );
  AND2_X1 U5201 ( .A1(n5271), .A2(n5810), .ZN(n5814) );
  AND4_X1 U5202 ( .A1(n5275), .A2(n5272), .A3(n5273), .A4(n5274), .ZN(n5734)
         );
  INV_X1 U5203 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9048) );
  NOR2_X1 U5204 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5270) );
  NOR2_X1 U5205 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6539) );
  INV_X1 U5206 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6903) );
  INV_X1 U5207 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6544) );
  NOR2_X1 U5208 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5273) );
  INV_X4 U5209 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U5210 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5272) );
  INV_X1 U5211 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U5212 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5274) );
  INV_X1 U5213 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9247) );
  INV_X1 U5214 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9266) );
  INV_X1 U5215 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6609) );
  INV_X1 U5216 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9246) );
  INV_X1 U5217 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6841) );
  NOR2_X1 U5218 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n6535) );
  NOR2_X1 U5219 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6536) );
  INV_X1 U5220 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6725) );
  INV_X2 U5221 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9251) );
  INV_X1 U5222 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5295) );
  INV_X1 U5223 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5804) );
  INV_X1 U5224 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5952) );
  INV_X1 U5225 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5895) );
  INV_X1 U5226 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5954) );
  INV_X1 U5227 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U5228 ( .A1(n6005), .A2(n7767), .ZN(n5016) );
  XNOR2_X2 U5229 ( .A(n5742), .B(n5743), .ZN(n5941) );
  NAND2_X4 U5230 ( .A1(n6551), .A2(n6552), .ZN(n7117) );
  OR2_X1 U5231 ( .A1(n8062), .A2(n8061), .ZN(n8064) );
  OAI211_X2 U5232 ( .C1(n7475), .C2(n7247), .A(n5819), .B(n5818), .ZN(n8061)
         );
  INV_X2 U5233 ( .A(n6298), .ZN(n6317) );
  NAND2_X1 U5234 ( .A1(n6462), .A2(n6463), .ZN(n5167) );
  MUX2_X1 U5235 ( .A(n6371), .B(n6370), .S(n6464), .Z(n6462) );
  AND2_X1 U5236 ( .A1(n6369), .A2(n6467), .ZN(n6370) );
  OR2_X1 U5237 ( .A1(n5167), .A2(n9536), .ZN(n5165) );
  INV_X1 U5238 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U5239 ( .A1(n8416), .A2(n8284), .ZN(n6415) );
  NAND2_X1 U5240 ( .A1(n5229), .A2(n5227), .ZN(n5902) );
  AOI21_X1 U5241 ( .B1(n5231), .B2(n5234), .A(n5228), .ZN(n5227) );
  INV_X1 U5242 ( .A(n5665), .ZN(n5228) );
  AND2_X1 U5243 ( .A1(n5184), .A2(n8563), .ZN(n5183) );
  AND2_X1 U5244 ( .A1(n5035), .A2(n5290), .ZN(n5184) );
  NAND2_X1 U5245 ( .A1(n5024), .A2(n5035), .ZN(n5185) );
  OAI21_X1 U5246 ( .B1(n6471), .B2(n6470), .A(n5222), .ZN(n5221) );
  AND2_X1 U5247 ( .A1(n9492), .A2(n6469), .ZN(n5222) );
  NOR2_X1 U5248 ( .A1(n8350), .A2(n9407), .ZN(n5304) );
  INV_X1 U5249 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5785) );
  AND2_X1 U5250 ( .A1(n10469), .A2(n10201), .ZN(n5366) );
  INV_X1 U5251 ( .A(n5378), .ZN(n5377) );
  OAI21_X1 U5252 ( .B1(n5379), .B2(n8755), .A(n5019), .ZN(n5378) );
  NOR2_X1 U5253 ( .A1(n5501), .A2(n5498), .ZN(n5497) );
  INV_X1 U5254 ( .A(n5637), .ZN(n5498) );
  INV_X1 U5255 ( .A(n5502), .ZN(n5501) );
  NAND2_X1 U5256 ( .A1(n5862), .A2(n5603), .ZN(n5638) );
  INV_X1 U5257 ( .A(n5627), .ZN(n5513) );
  INV_X1 U5258 ( .A(n5457), .ZN(n5455) );
  INV_X1 U5259 ( .A(n5933), .ZN(n5994) );
  NAND2_X1 U5260 ( .A1(n5161), .A2(n5159), .ZN(n5158) );
  INV_X1 U5261 ( .A(n5162), .ZN(n5159) );
  INV_X1 U5262 ( .A(n5533), .ZN(n5156) );
  AOI21_X1 U5263 ( .B1(n5534), .B2(n5536), .A(n5048), .ZN(n5533) );
  OR2_X1 U5264 ( .A1(n9679), .A2(n8807), .ZN(n6483) );
  OR2_X1 U5265 ( .A1(n9695), .A2(n9294), .ZN(n6469) );
  OR2_X1 U5266 ( .A1(n9588), .A2(n9361), .ZN(n6372) );
  AOI21_X1 U5267 ( .B1(n5258), .B2(n5255), .A(n5254), .ZN(n5253) );
  INV_X1 U5268 ( .A(n6441), .ZN(n5254) );
  INV_X1 U5269 ( .A(n5260), .ZN(n5255) );
  NOR2_X1 U5270 ( .A1(n8608), .A2(n8656), .ZN(n8609) );
  OR2_X1 U5271 ( .A1(n9716), .A2(n9563), .ZN(n6453) );
  AND4_X1 U5272 ( .A1(n5784), .A2(n5895), .A3(n5785), .A4(n5295), .ZN(n5739)
         );
  NAND2_X1 U5273 ( .A1(n5560), .A2(n7046), .ZN(n5556) );
  AND2_X1 U5274 ( .A1(n7160), .A2(n7123), .ZN(n6708) );
  NAND2_X1 U5275 ( .A1(n10002), .A2(n5594), .ZN(n10003) );
  NAND2_X1 U5276 ( .A1(n10006), .A2(n10100), .ZN(n10002) );
  NAND2_X1 U5277 ( .A1(n5520), .A2(n10007), .ZN(n5519) );
  INV_X1 U5278 ( .A(n5518), .ZN(n5517) );
  OAI21_X1 U5279 ( .B1(n10111), .B2(n10011), .A(n10143), .ZN(n5518) );
  OR2_X1 U5280 ( .A1(n8785), .A2(n8844), .ZN(n10005) );
  OR2_X1 U5281 ( .A1(n10474), .A2(n10315), .ZN(n10020) );
  NAND2_X1 U5282 ( .A1(n8784), .A2(n10302), .ZN(n5368) );
  NOR2_X1 U5283 ( .A1(n10484), .A2(n10491), .ZN(n5319) );
  NOR2_X1 U5284 ( .A1(n5380), .A2(n5419), .ZN(n5418) );
  INV_X1 U5285 ( .A(n10031), .ZN(n5419) );
  OR2_X1 U5286 ( .A1(n8473), .A2(n5389), .ZN(n5388) );
  INV_X1 U5287 ( .A(n8302), .ZN(n5389) );
  NAND2_X1 U5288 ( .A1(n8022), .A2(n10123), .ZN(n8135) );
  NAND2_X1 U5289 ( .A1(n8243), .A2(n8146), .ZN(n10126) );
  INV_X1 U5290 ( .A(n5415), .ZN(n5414) );
  AOI21_X1 U5291 ( .B1(n5413), .B2(n5415), .A(n5412), .ZN(n5411) );
  INV_X1 U5292 ( .A(n10037), .ZN(n5412) );
  NAND2_X1 U5293 ( .A1(n5719), .A2(n5718), .ZN(n5753) );
  INV_X1 U5294 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U5295 ( .A1(n5507), .A2(n5505), .ZN(n5916) );
  AOI21_X1 U5296 ( .B1(n5509), .B2(n5511), .A(n5506), .ZN(n5505) );
  NAND2_X1 U5297 ( .A1(n5912), .A2(n5509), .ZN(n5507) );
  INV_X1 U5298 ( .A(n5714), .ZN(n5506) );
  NAND3_X1 U5299 ( .A1(n6543), .A2(n5059), .A3(n6542), .ZN(n5309) );
  NOR2_X1 U5300 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6545) );
  INV_X1 U5301 ( .A(n5587), .ZN(n5585) );
  NOR2_X1 U5302 ( .A1(n5047), .A2(n5422), .ZN(n5421) );
  AND2_X1 U5303 ( .A1(n5714), .A2(n5713), .ZN(n5757) );
  NOR2_X1 U5304 ( .A1(n7100), .A2(n5422), .ZN(n6557) );
  NAND2_X1 U5305 ( .A1(n5240), .A2(n5490), .ZN(n5777) );
  AOI21_X1 U5306 ( .B1(n5494), .B2(n5492), .A(n5491), .ZN(n5490) );
  OR2_X1 U5307 ( .A1(n5781), .A2(n5493), .ZN(n5240) );
  INV_X1 U5308 ( .A(n5681), .ZN(n5491) );
  INV_X1 U5309 ( .A(SI_17_), .ZN(n5666) );
  AND2_X1 U5310 ( .A1(n5665), .A2(n5664), .ZN(n5793) );
  INV_X1 U5311 ( .A(n5893), .ZN(n5239) );
  NAND2_X1 U5312 ( .A1(n5655), .A2(n5654), .ZN(n5894) );
  INV_X1 U5313 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5211) );
  AND2_X1 U5314 ( .A1(n6002), .A2(n8350), .ZN(n6003) );
  INV_X1 U5315 ( .A(n5447), .ZN(n5135) );
  OAI21_X1 U5316 ( .B1(n5449), .B2(n5448), .A(n5061), .ZN(n5447) );
  INV_X1 U5317 ( .A(n8260), .ZN(n5448) );
  AOI21_X1 U5318 ( .B1(n8586), .B2(n6135), .A(n6146), .ZN(n5115) );
  INV_X1 U5319 ( .A(n8586), .ZN(n5116) );
  NAND2_X1 U5320 ( .A1(n8833), .A2(n8750), .ZN(n6163) );
  INV_X1 U5321 ( .A(n6025), .ZN(n6298) );
  INV_X1 U5322 ( .A(n7470), .ZN(n7281) );
  NAND2_X1 U5323 ( .A1(n7475), .A2(n5724), .ZN(n5824) );
  OR2_X1 U5324 ( .A1(n9695), .A2(n9530), .ZN(n5162) );
  OAI21_X1 U5325 ( .B1(n9527), .B2(n9548), .A(n9519), .ZN(n9505) );
  OR2_X1 U5326 ( .A1(n9705), .A2(n9564), .ZN(n6371) );
  INV_X1 U5327 ( .A(n5543), .ZN(n5538) );
  NOR2_X1 U5328 ( .A1(n5540), .A2(n5191), .ZN(n5189) );
  OR2_X1 U5329 ( .A1(n9596), .A2(n9716), .ZN(n9572) );
  NAND2_X1 U5330 ( .A1(n9587), .A2(n5190), .ZN(n9571) );
  NOR2_X1 U5331 ( .A1(n6337), .A2(n5486), .ZN(n5485) );
  INV_X1 U5332 ( .A(n6504), .ZN(n5486) );
  INV_X1 U5333 ( .A(n9619), .ZN(n9641) );
  NAND2_X1 U5334 ( .A1(n7475), .A2(n6575), .ZN(n5845) );
  OR2_X1 U5335 ( .A1(n10664), .A2(n5976), .ZN(n8038) );
  NOR2_X1 U5336 ( .A1(n5550), .A2(n5549), .ZN(n5548) );
  NAND2_X1 U5337 ( .A1(n5958), .A2(n5744), .ZN(n5549) );
  OR2_X1 U5338 ( .A1(n7155), .A2(n5397), .ZN(n5395) );
  OR2_X1 U5339 ( .A1(n8549), .A2(n5030), .ZN(n5584) );
  AOI21_X1 U5340 ( .B1(n10262), .B2(n10271), .A(n5598), .ZN(n8840) );
  OR2_X1 U5341 ( .A1(n10484), .A2(n10202), .ZN(n8762) );
  INV_X1 U5342 ( .A(n5372), .ZN(n5371) );
  OAI21_X1 U5343 ( .B1(n5374), .B2(n5373), .A(n10936), .ZN(n5372) );
  INV_X1 U5344 ( .A(n8751), .ZN(n5373) );
  OAI21_X1 U5345 ( .B1(n10869), .B2(n8622), .A(n10073), .ZN(n8623) );
  NAND2_X1 U5346 ( .A1(n8623), .A2(n10166), .ZN(n8675) );
  INV_X1 U5347 ( .A(n7140), .ZN(n7154) );
  NAND2_X1 U5348 ( .A1(n8149), .A2(n8016), .ZN(n8134) );
  AND2_X1 U5349 ( .A1(n5694), .A2(n5693), .ZN(n5769) );
  NAND2_X1 U5350 ( .A1(n5195), .A2(n5194), .ZN(n6412) );
  NAND2_X1 U5351 ( .A1(n6411), .A2(n6464), .ZN(n5195) );
  AND2_X1 U5352 ( .A1(n9646), .A2(n6440), .ZN(n5290) );
  AND2_X1 U5353 ( .A1(n9584), .A2(n5288), .ZN(n5287) );
  NAND2_X1 U5354 ( .A1(n5289), .A2(n9612), .ZN(n5288) );
  AND2_X1 U5355 ( .A1(n9492), .A2(n6468), .ZN(n5166) );
  NAND2_X1 U5356 ( .A1(n5018), .A2(n5167), .ZN(n5163) );
  OAI21_X1 U5357 ( .B1(n6481), .B2(n6474), .A(n5217), .ZN(n6475) );
  NOR2_X1 U5358 ( .A1(n5218), .A2(n6480), .ZN(n5217) );
  INV_X1 U5359 ( .A(n6482), .ZN(n5218) );
  AOI21_X1 U5360 ( .B1(n6481), .B2(n5299), .A(n5297), .ZN(n5296) );
  NAND2_X1 U5361 ( .A1(n5298), .A2(n6484), .ZN(n5297) );
  NAND2_X1 U5362 ( .A1(n5299), .A2(n5301), .ZN(n5298) );
  INV_X1 U5363 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8998) );
  INV_X1 U5364 ( .A(n5570), .ZN(n5567) );
  INV_X1 U5365 ( .A(n9882), .ZN(n5566) );
  NOR2_X1 U5366 ( .A1(n9882), .A2(n5569), .ZN(n5568) );
  INV_X1 U5367 ( .A(n5574), .ZN(n5569) );
  NOR2_X1 U5368 ( .A1(n8683), .A2(n10884), .ZN(n5324) );
  NOR2_X1 U5369 ( .A1(n9942), .A2(n9941), .ZN(n8305) );
  INV_X1 U5370 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9026) );
  NOR2_X1 U5371 ( .A1(n5645), .A2(n5503), .ZN(n5502) );
  INV_X1 U5372 ( .A(n5643), .ZN(n5503) );
  INV_X1 U5373 ( .A(n5601), .ZN(n5500) );
  AND2_X1 U5374 ( .A1(n8858), .A2(n5432), .ZN(n5431) );
  OR2_X1 U5375 ( .A1(n9370), .A2(n5022), .ZN(n5432) );
  NAND2_X1 U5376 ( .A1(n6217), .A2(n6216), .ZN(n5445) );
  NAND2_X1 U5377 ( .A1(n5133), .A2(n5137), .ZN(n5136) );
  NAND2_X1 U5378 ( .A1(n6367), .A2(n6485), .ZN(n5471) );
  INV_X1 U5379 ( .A(n5473), .ZN(n5472) );
  OAI21_X1 U5380 ( .B1(n9442), .B2(n5474), .A(n6486), .ZN(n5473) );
  NAND2_X1 U5381 ( .A1(n5172), .A2(n5171), .ZN(n5170) );
  INV_X1 U5382 ( .A(n6521), .ZN(n5171) );
  NOR2_X1 U5383 ( .A1(n5282), .A2(n5283), .ZN(n5281) );
  NOR2_X1 U5384 ( .A1(n6498), .A2(n6464), .ZN(n5169) );
  NAND2_X1 U5385 ( .A1(n5176), .A2(n6493), .ZN(n5175) );
  NAND2_X1 U5386 ( .A1(n5177), .A2(n6494), .ZN(n5176) );
  AND2_X1 U5387 ( .A1(n6004), .A2(n6001), .ZN(n6318) );
  INV_X1 U5388 ( .A(n5161), .ZN(n5160) );
  AOI21_X1 U5389 ( .B1(n9511), .B2(n5162), .A(n9492), .ZN(n5161) );
  NOR2_X1 U5390 ( .A1(n9700), .A2(n9705), .ZN(n5342) );
  INV_X1 U5391 ( .A(n6453), .ZN(n5481) );
  AND2_X1 U5392 ( .A1(n5348), .A2(n5347), .ZN(n5346) );
  INV_X1 U5393 ( .A(n5258), .ZN(n5256) );
  OR2_X1 U5394 ( .A1(n9627), .A2(n9639), .ZN(n8802) );
  NOR2_X1 U5395 ( .A1(n9627), .A2(n9656), .ZN(n5348) );
  NOR2_X1 U5396 ( .A1(n6341), .A2(n5261), .ZN(n5260) );
  INV_X1 U5397 ( .A(n6340), .ZN(n5261) );
  AOI21_X1 U5398 ( .B1(n5260), .B2(n8601), .A(n5259), .ZN(n5258) );
  INV_X1 U5399 ( .A(n6439), .ZN(n5259) );
  AND2_X1 U5400 ( .A1(n8660), .A2(n5153), .ZN(n5152) );
  NAND2_X1 U5401 ( .A1(n8658), .A2(n8657), .ZN(n5153) );
  OR2_X1 U5402 ( .A1(n9744), .A2(n9642), .ZN(n6438) );
  AND2_X1 U5403 ( .A1(n8390), .A2(n8386), .ZN(n5547) );
  NOR2_X1 U5404 ( .A1(n8385), .A2(n8281), .ZN(n5353) );
  OAI21_X1 U5405 ( .B1(n8078), .B2(n5529), .A(n8077), .ZN(n5528) );
  OR2_X1 U5406 ( .A1(n7957), .A2(n5530), .ZN(n5529) );
  INV_X1 U5407 ( .A(n7958), .ZN(n5530) );
  AND2_X1 U5408 ( .A1(n6407), .A2(n6408), .ZN(n8080) );
  NAND2_X1 U5409 ( .A1(n8205), .A2(n6331), .ZN(n5479) );
  NAND2_X1 U5410 ( .A1(n6329), .A2(n8108), .ZN(n5525) );
  NAND2_X1 U5411 ( .A1(n7404), .A2(n8240), .ZN(n7756) );
  NAND2_X1 U5412 ( .A1(n5743), .A2(n5551), .ZN(n5550) );
  AND2_X1 U5413 ( .A1(n5734), .A2(n5829), .ZN(n5883) );
  NAND2_X1 U5414 ( .A1(n8515), .A2(n5200), .ZN(n5199) );
  NAND2_X1 U5415 ( .A1(n5582), .A2(n5203), .ZN(n5202) );
  NAND2_X1 U5416 ( .A1(n5515), .A2(n10007), .ZN(n5514) );
  INV_X1 U5417 ( .A(n10143), .ZN(n5515) );
  INV_X1 U5418 ( .A(n8794), .ZN(n6552) );
  NOR2_X1 U5419 ( .A1(n5359), .A2(n5356), .ZN(n5355) );
  INV_X1 U5420 ( .A(n5360), .ZN(n5356) );
  INV_X1 U5421 ( .A(n5365), .ZN(n5359) );
  NOR2_X1 U5422 ( .A1(n10175), .A2(n5366), .ZN(n5365) );
  INV_X1 U5423 ( .A(n5366), .ZN(n5364) );
  NAND2_X1 U5424 ( .A1(n8765), .A2(n5367), .ZN(n5363) );
  NAND2_X1 U5425 ( .A1(n10117), .A2(n9983), .ZN(n5392) );
  AND2_X1 U5426 ( .A1(n10506), .A2(n10418), .ZN(n8757) );
  NOR2_X1 U5427 ( .A1(n10506), .A2(n10426), .ZN(n5313) );
  NOR2_X1 U5428 ( .A1(n5323), .A2(n9809), .ZN(n5322) );
  INV_X1 U5429 ( .A(n5324), .ZN(n5323) );
  NOR2_X1 U5430 ( .A1(n9964), .A2(n5375), .ZN(n5374) );
  INV_X1 U5431 ( .A(n8710), .ZN(n5375) );
  OR2_X1 U5432 ( .A1(n9809), .A2(n8719), .ZN(n10077) );
  INV_X1 U5433 ( .A(n10183), .ZN(n10049) );
  INV_X1 U5434 ( .A(n10496), .ZN(n5310) );
  NOR2_X1 U5435 ( .A1(n10162), .A2(n5416), .ZN(n5415) );
  INV_X1 U5436 ( .A(n10065), .ZN(n5416) );
  NAND2_X1 U5437 ( .A1(n8306), .A2(n8305), .ZN(n5417) );
  NAND2_X1 U5438 ( .A1(n5723), .A2(n5722), .ZN(n5749) );
  AND2_X1 U5439 ( .A1(n5709), .A2(n5708), .ZN(n5911) );
  NAND2_X1 U5440 ( .A1(n5705), .A2(n5704), .ZN(n5912) );
  INV_X1 U5441 ( .A(n5761), .ZN(n5524) );
  NAND2_X1 U5442 ( .A1(n6544), .A2(n5588), .ZN(n5587) );
  INV_X1 U5443 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U5444 ( .A1(n5673), .A2(n5672), .ZN(n5781) );
  NAND2_X1 U5445 ( .A1(n5789), .A2(n5670), .ZN(n5673) );
  OAI21_X1 U5446 ( .B1(n5882), .B2(n5881), .A(n5649), .ZN(n5889) );
  NAND2_X1 U5447 ( .A1(n5855), .A2(n5632), .ZN(n5862) );
  OAI21_X1 U5448 ( .B1(n6575), .B2(n5193), .A(n5192), .ZN(n5212) );
  NAND2_X1 U5449 ( .A1(n6575), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5192) );
  INV_X1 U5450 ( .A(n9315), .ZN(n5130) );
  AND2_X1 U5451 ( .A1(n9370), .A2(n6265), .ZN(n5132) );
  OAI211_X1 U5452 ( .C1(n9299), .C2(n5125), .A(n5434), .B(n5124), .ZN(n6241)
         );
  INV_X1 U5453 ( .A(n5436), .ZN(n5125) );
  AOI21_X1 U5454 ( .B1(n5436), .B2(n5439), .A(n6230), .ZN(n5434) );
  AND2_X1 U5455 ( .A1(n5431), .A2(n5433), .ZN(n5425) );
  NAND2_X1 U5456 ( .A1(n5430), .A2(n5428), .ZN(n5427) );
  OR2_X1 U5457 ( .A1(n5431), .A2(n5433), .ZN(n5428) );
  AOI21_X1 U5458 ( .B1(n5431), .B2(n5022), .A(n6291), .ZN(n5430) );
  XNOR2_X1 U5459 ( .A(n5016), .B(n8108), .ZN(n6012) );
  OR2_X1 U5460 ( .A1(n6208), .A2(n6207), .ZN(n5446) );
  AOI21_X1 U5461 ( .B1(n9332), .B2(n9333), .A(n6253), .ZN(n9316) );
  NAND2_X1 U5462 ( .A1(n8694), .A2(n8695), .ZN(n8693) );
  NAND2_X1 U5463 ( .A1(n8095), .A2(n8094), .ZN(n8093) );
  AND2_X1 U5464 ( .A1(n6318), .A2(n10702), .ZN(n6299) );
  INV_X1 U5465 ( .A(n5440), .ZN(n5439) );
  INV_X1 U5466 ( .A(n5442), .ZN(n5438) );
  INV_X1 U5467 ( .A(n9350), .ZN(n5437) );
  AND2_X1 U5468 ( .A1(n5446), .A2(n5445), .ZN(n5442) );
  INV_X1 U5469 ( .A(n5445), .ZN(n5441) );
  AOI21_X1 U5470 ( .B1(n9341), .B2(n5446), .A(n5444), .ZN(n5443) );
  INV_X1 U5471 ( .A(n9306), .ZN(n5444) );
  AOI21_X1 U5472 ( .B1(n5452), .B2(n5450), .A(n5054), .ZN(n5449) );
  INV_X1 U5473 ( .A(n8094), .ZN(n5450) );
  INV_X1 U5474 ( .A(n5136), .ZN(n8095) );
  NAND2_X1 U5475 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  AOI21_X1 U5476 ( .B1(n5460), .B2(n5458), .A(n5055), .ZN(n5457) );
  INV_X1 U5477 ( .A(n8695), .ZN(n5458) );
  AND2_X1 U5478 ( .A1(n6054), .A2(n6053), .ZN(n5465) );
  NAND2_X1 U5479 ( .A1(n9316), .A2(n9315), .ZN(n9314) );
  NAND2_X1 U5480 ( .A1(n5114), .A2(n5112), .ZN(n8638) );
  AOI21_X1 U5481 ( .B1(n5115), .B2(n5116), .A(n5113), .ZN(n5112) );
  INV_X1 U5482 ( .A(n8640), .ZN(n5113) );
  OR2_X1 U5483 ( .A1(n8038), .A2(n8036), .ZN(n6319) );
  NAND2_X1 U5484 ( .A1(n6506), .A2(n7760), .ZN(n7767) );
  NAND2_X1 U5485 ( .A1(n5995), .A2(n5994), .ZN(n6025) );
  NOR2_X1 U5486 ( .A1(n9668), .A2(n9436), .ZN(n9431) );
  NAND2_X1 U5487 ( .A1(n9441), .A2(n6485), .ZN(n5269) );
  NAND2_X1 U5488 ( .A1(n6367), .A2(n6486), .ZN(n8815) );
  NAND2_X1 U5489 ( .A1(n9443), .A2(n9442), .ZN(n9441) );
  OR2_X1 U5490 ( .A1(n9452), .A2(n9674), .ZN(n9436) );
  NOR2_X1 U5491 ( .A1(n9496), .A2(n9684), .ZN(n9480) );
  INV_X1 U5492 ( .A(n9477), .ZN(n5536) );
  AOI21_X1 U5493 ( .B1(n9477), .B2(n5535), .A(n5058), .ZN(n5534) );
  INV_X1 U5494 ( .A(n8805), .ZN(n5535) );
  OR2_X1 U5495 ( .A1(n9498), .A2(n6347), .ZN(n9474) );
  NAND2_X1 U5496 ( .A1(n5157), .A2(n5161), .ZN(n9487) );
  NAND2_X1 U5497 ( .A1(n9505), .A2(n5162), .ZN(n5157) );
  INV_X1 U5498 ( .A(n5771), .ZN(n5226) );
  NAND2_X1 U5499 ( .A1(n5771), .A2(n5845), .ZN(n5225) );
  AND2_X1 U5500 ( .A1(n9529), .A2(n6371), .ZN(n5484) );
  NAND2_X1 U5501 ( .A1(n6242), .A2(n6233), .ZN(n9524) );
  NAND2_X1 U5502 ( .A1(n5187), .A2(n5186), .ZN(n9519) );
  NOR2_X1 U5503 ( .A1(n5188), .A2(n9529), .ZN(n5186) );
  AND2_X1 U5504 ( .A1(n6503), .A2(n9577), .ZN(n5543) );
  NAND2_X1 U5505 ( .A1(n5064), .A2(n6503), .ZN(n5542) );
  AND2_X1 U5506 ( .A1(n6503), .A2(n6502), .ZN(n9560) );
  AND2_X1 U5507 ( .A1(n5243), .A2(n6372), .ZN(n5242) );
  NAND2_X1 U5508 ( .A1(n5245), .A2(n5028), .ZN(n5243) );
  NAND2_X1 U5509 ( .A1(n9611), .A2(n5084), .ZN(n9587) );
  OAI21_X1 U5510 ( .B1(n9624), .B2(n9623), .A(n8802), .ZN(n9613) );
  NAND2_X1 U5511 ( .A1(n9613), .A2(n9612), .ZN(n9611) );
  AND2_X1 U5512 ( .A1(n5545), .A2(n5149), .ZN(n5148) );
  NOR2_X1 U5513 ( .A1(n9646), .A2(n5546), .ZN(n5545) );
  NAND2_X1 U5514 ( .A1(n5152), .A2(n5150), .ZN(n5149) );
  INV_X1 U5515 ( .A(n8800), .ZN(n5546) );
  INV_X1 U5516 ( .A(n5152), .ZN(n5151) );
  NAND2_X1 U5517 ( .A1(n5147), .A2(n5152), .ZN(n8801) );
  NAND2_X1 U5518 ( .A1(n8659), .A2(n8657), .ZN(n5147) );
  NAND2_X1 U5519 ( .A1(n5900), .A2(n5899), .ZN(n8656) );
  OR2_X1 U5520 ( .A1(n8572), .A2(n8605), .ZN(n8608) );
  OR2_X1 U5521 ( .A1(n10852), .A2(n8506), .ZN(n8502) );
  AOI21_X1 U5522 ( .B1(n5142), .B2(n5144), .A(n5043), .ZN(n5141) );
  AND2_X1 U5523 ( .A1(n8090), .A2(n5349), .ZN(n8507) );
  NOR2_X1 U5524 ( .A1(n5351), .A2(n10852), .ZN(n5349) );
  NAND2_X1 U5525 ( .A1(n8387), .A2(n5547), .ZN(n8418) );
  NOR2_X1 U5526 ( .A1(n8390), .A2(n5489), .ZN(n5488) );
  INV_X1 U5527 ( .A(n6411), .ZN(n5489) );
  NAND2_X1 U5528 ( .A1(n8286), .A2(n6411), .ZN(n8391) );
  INV_X1 U5529 ( .A(n6402), .ZN(n8084) );
  AND2_X1 U5530 ( .A1(n8080), .A2(n6402), .ZN(n6334) );
  INV_X1 U5531 ( .A(n8080), .ZN(n8083) );
  NAND2_X1 U5532 ( .A1(n7960), .A2(n8078), .ZN(n8082) );
  OAI21_X1 U5533 ( .B1(n7264), .B2(n5845), .A(n5847), .ZN(n8450) );
  NAND2_X1 U5534 ( .A1(n7767), .A2(n7766), .ZN(n9644) );
  AND2_X1 U5535 ( .A1(n7281), .A2(n6320), .ZN(n9619) );
  NAND2_X1 U5536 ( .A1(n8240), .A2(n7754), .ZN(n8062) );
  NAND2_X1 U5537 ( .A1(n5747), .A2(n5746), .ZN(n6363) );
  NAND2_X1 U5538 ( .A1(n5760), .A2(n5759), .ZN(n9679) );
  NOR2_X1 U5539 ( .A1(n7257), .A2(n5724), .ZN(n5128) );
  NOR2_X1 U5540 ( .A1(n8704), .A2(n5964), .ZN(n10550) );
  XNOR2_X1 U5541 ( .A(n5932), .B(n5931), .ZN(n5933) );
  AND2_X1 U5542 ( .A1(n10984), .A2(n5551), .ZN(n5121) );
  INV_X1 U5543 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5924) );
  INV_X1 U5544 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U5545 ( .A1(n5468), .A2(n5467), .ZN(n5925) );
  AOI21_X1 U5546 ( .B1(n5469), .B2(n5956), .A(n5956), .ZN(n5467) );
  INV_X1 U5547 ( .A(n5470), .ZN(n5469) );
  NAND2_X1 U5548 ( .A1(n5782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U5549 ( .A1(n5557), .A2(n5554), .ZN(n7081) );
  INV_X1 U5550 ( .A(n5555), .ZN(n5554) );
  AOI21_X1 U5551 ( .B1(n9904), .B2(n5556), .A(n7062), .ZN(n5555) );
  NAND2_X1 U5552 ( .A1(n5576), .A2(n5082), .ZN(n5575) );
  INV_X1 U5553 ( .A(n9872), .ZN(n5576) );
  OR2_X2 U5554 ( .A1(n9824), .A2(n5079), .ZN(n6954) );
  OAI21_X1 U5555 ( .B1(n5327), .B2(n5021), .A(n7140), .ZN(n5326) );
  OR2_X1 U5556 ( .A1(n7140), .A2(n7252), .ZN(n5606) );
  INV_X1 U5557 ( .A(n6678), .ZN(n6699) );
  INV_X1 U5558 ( .A(n6655), .ZN(n6730) );
  OR2_X1 U5559 ( .A1(n7117), .A2(n7891), .ZN(n6639) );
  NAND2_X1 U5560 ( .A1(n6551), .A2(n8794), .ZN(n6604) );
  AND2_X1 U5561 ( .A1(n8836), .A2(n8794), .ZN(n6678) );
  NAND2_X1 U5562 ( .A1(n8768), .A2(n8767), .ZN(n8785) );
  NOR2_X1 U5563 ( .A1(n8841), .A2(n8776), .ZN(n8777) );
  NAND2_X1 U5564 ( .A1(n10004), .A2(n10103), .ZN(n10178) );
  INV_X1 U5565 ( .A(n5332), .ZN(n5330) );
  NOR2_X1 U5566 ( .A1(n10271), .A2(n10099), .ZN(n5410) );
  NAND2_X1 U5567 ( .A1(n10284), .A2(n10098), .ZN(n10270) );
  NAND2_X1 U5568 ( .A1(n10100), .A2(n10101), .ZN(n10271) );
  NOR2_X1 U5569 ( .A1(n10299), .A2(n8775), .ZN(n10285) );
  NAND2_X1 U5570 ( .A1(n10285), .A2(n10286), .ZN(n10284) );
  NAND2_X1 U5571 ( .A1(n10298), .A2(n10315), .ZN(n5367) );
  INV_X1 U5572 ( .A(n10201), .ZN(n10303) );
  NAND2_X1 U5573 ( .A1(n8763), .A2(n5360), .ZN(n5369) );
  INV_X1 U5574 ( .A(n10202), .ZN(n10348) );
  INV_X1 U5575 ( .A(n10288), .ZN(n10315) );
  NAND2_X1 U5576 ( .A1(n10345), .A2(n10090), .ZN(n10331) );
  NOR2_X1 U5577 ( .A1(n10354), .A2(n10491), .ZN(n10343) );
  NOR2_X1 U5578 ( .A1(n10396), .A2(n8774), .ZN(n10373) );
  OAI21_X1 U5579 ( .B1(n10415), .B2(n5404), .A(n5403), .ZN(n10396) );
  NAND2_X1 U5580 ( .A1(n10389), .A2(n10410), .ZN(n5404) );
  NAND2_X1 U5581 ( .A1(n10389), .A2(n8773), .ZN(n5403) );
  NOR2_X1 U5582 ( .A1(n10415), .A2(n10414), .ZN(n10417) );
  AND2_X1 U5583 ( .A1(n10081), .A2(n10036), .ZN(n9964) );
  NAND2_X1 U5584 ( .A1(n8711), .A2(n5374), .ZN(n8752) );
  AOI21_X1 U5585 ( .B1(n5383), .B2(n10868), .A(n5050), .ZN(n5382) );
  INV_X1 U5586 ( .A(n10041), .ZN(n5394) );
  NAND2_X1 U5587 ( .A1(n8630), .A2(n8629), .ZN(n10863) );
  INV_X1 U5588 ( .A(n5387), .ZN(n5386) );
  OAI21_X1 U5589 ( .B1(n5032), .B2(n5388), .A(n8472), .ZN(n5387) );
  OR2_X1 U5590 ( .A1(n8310), .A2(n8471), .ZN(n10803) );
  AOI21_X1 U5591 ( .B1(n8135), .B2(n10060), .A(n8024), .ZN(n8241) );
  NAND2_X1 U5592 ( .A1(n8241), .A2(n8242), .ZN(n8306) );
  INV_X1 U5593 ( .A(n10207), .ZN(n8243) );
  AND2_X1 U5594 ( .A1(n8015), .A2(n8012), .ZN(n5370) );
  INV_X1 U5595 ( .A(n10157), .ZN(n8015) );
  AND2_X1 U5596 ( .A1(n10125), .A2(n8023), .ZN(n10157) );
  INV_X1 U5597 ( .A(n10192), .ZN(n7845) );
  INV_X1 U5598 ( .A(n10403), .ZN(n10942) );
  INV_X1 U5599 ( .A(n10401), .ZN(n10944) );
  OR2_X1 U5600 ( .A1(n7127), .A2(n10018), .ZN(n10401) );
  NAND2_X1 U5601 ( .A1(n7127), .A2(n7387), .ZN(n10403) );
  NAND2_X1 U5602 ( .A1(n7064), .A2(n7063), .ZN(n10464) );
  INV_X1 U5603 ( .A(n8301), .ZN(n10776) );
  OR2_X1 U5604 ( .A1(n6626), .A2(n7255), .ZN(n6628) );
  OR2_X1 U5605 ( .A1(n7845), .A2(n7386), .ZN(n10970) );
  NOR2_X1 U5606 ( .A1(n7400), .A2(n7422), .ZN(n7409) );
  AND2_X1 U5607 ( .A1(n8538), .A2(n10183), .ZN(n7846) );
  AND2_X1 U5608 ( .A1(n7082), .A2(n7083), .ZN(n5196) );
  XNOR2_X1 U5609 ( .A(n6546), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U5610 ( .A1(n5590), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6546) );
  XNOR2_X1 U5611 ( .A(n5916), .B(n5915), .ZN(n8834) );
  INV_X1 U5612 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9271) );
  INV_X1 U5613 ( .A(n5421), .ZN(n5308) );
  XNOR2_X1 U5614 ( .A(n5912), .B(n5911), .ZN(n8702) );
  NAND2_X1 U5615 ( .A1(n5521), .A2(n5699), .ZN(n5762) );
  INV_X1 U5616 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9044) );
  INV_X1 U5617 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9262) );
  INV_X1 U5618 ( .A(n6582), .ZN(n5586) );
  NAND2_X1 U5619 ( .A1(n5230), .A2(n5235), .ZN(n5794) );
  NAND2_X1 U5620 ( .A1(n5894), .A2(n5237), .ZN(n5230) );
  NAND2_X1 U5621 ( .A1(n5504), .A2(n5643), .ZN(n5874) );
  NAND2_X1 U5622 ( .A1(n5867), .A2(n5601), .ZN(n5504) );
  OAI21_X1 U5623 ( .B1(n5512), .B2(n5038), .A(n5108), .ZN(n5854) );
  NOR2_X1 U5624 ( .A1(n5215), .A2(n5060), .ZN(n5108) );
  INV_X1 U5625 ( .A(n5623), .ZN(n5512) );
  XNOR2_X1 U5626 ( .A(n5248), .B(n5850), .ZN(n7269) );
  NAND2_X1 U5627 ( .A1(n5849), .A2(n5848), .ZN(n5248) );
  NAND2_X1 U5628 ( .A1(n5844), .A2(n5843), .ZN(n5849) );
  NAND2_X1 U5629 ( .A1(n5111), .A2(n6065), .ZN(n7872) );
  XNOR2_X1 U5630 ( .A(n6241), .B(n6240), .ZN(n9292) );
  AOI22_X1 U5631 ( .A1(n7403), .A2(n7402), .B1(n6024), .B2(n6023), .ZN(n7790)
         );
  NOR2_X1 U5632 ( .A1(n7380), .A2(n7379), .ZN(n7378) );
  NAND2_X1 U5633 ( .A1(n5768), .A2(n5767), .ZN(n9695) );
  NAND2_X1 U5634 ( .A1(n9299), .A2(n6198), .ZN(n9342) );
  NAND2_X1 U5635 ( .A1(n5099), .A2(n5910), .ZN(n9716) );
  NAND2_X1 U5636 ( .A1(n8325), .A2(n5856), .ZN(n5099) );
  INV_X1 U5637 ( .A(n9352), .ZN(n9381) );
  INV_X1 U5638 ( .A(n9294), .ZN(n9530) );
  OR2_X1 U5639 ( .A1(n6166), .A2(n6165), .ZN(n9618) );
  INV_X1 U5640 ( .A(n6363), .ZN(n9430) );
  NAND2_X1 U5641 ( .A1(n6999), .A2(n6998), .ZN(n10484) );
  INV_X1 U5642 ( .A(n5399), .ZN(n5398) );
  NAND2_X1 U5643 ( .A1(n8516), .A2(n8517), .ZN(n5204) );
  NAND2_X1 U5644 ( .A1(n6907), .A2(n6906), .ZN(n10516) );
  INV_X1 U5645 ( .A(n8538), .ZN(n10017) );
  AND2_X1 U5646 ( .A1(n8825), .A2(n8824), .ZN(n10011) );
  INV_X1 U5647 ( .A(n5303), .ZN(n6384) );
  OAI21_X1 U5648 ( .B1(n6392), .B2(n6508), .A(n6391), .ZN(n5280) );
  INV_X1 U5649 ( .A(n6430), .ZN(n5292) );
  NAND2_X1 U5650 ( .A1(n5182), .A2(n5180), .ZN(n6446) );
  AOI21_X1 U5651 ( .B1(n5025), .B2(n5290), .A(n5181), .ZN(n5180) );
  INV_X1 U5652 ( .A(n6443), .ZN(n5181) );
  NAND2_X1 U5653 ( .A1(n5284), .A2(n6455), .ZN(n6458) );
  NAND2_X1 U5654 ( .A1(n5302), .A2(n6482), .ZN(n5301) );
  INV_X1 U5655 ( .A(n5300), .ZN(n5299) );
  OAI21_X1 U5656 ( .B1(n5301), .B2(n6479), .A(n6483), .ZN(n5300) );
  NAND2_X1 U5657 ( .A1(n5223), .A2(n5219), .ZN(n6481) );
  NAND2_X1 U5658 ( .A1(n6473), .A2(n6464), .ZN(n5223) );
  NAND2_X1 U5659 ( .A1(n5220), .A2(n6499), .ZN(n5219) );
  INV_X1 U5660 ( .A(SI_16_), .ZN(n9096) );
  INV_X1 U5661 ( .A(SI_15_), .ZN(n8890) );
  INV_X1 U5662 ( .A(SI_13_), .ZN(n9094) );
  INV_X1 U5663 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9214) );
  INV_X1 U5664 ( .A(SI_12_), .ZN(n9101) );
  INV_X1 U5665 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9219) );
  INV_X1 U5666 ( .A(SI_9_), .ZN(n9109) );
  INV_X1 U5667 ( .A(SI_8_), .ZN(n9110) );
  INV_X1 U5668 ( .A(n6494), .ZN(n5282) );
  INV_X1 U5669 ( .A(n6496), .ZN(n5283) );
  NAND2_X1 U5670 ( .A1(n6490), .A2(n6499), .ZN(n5178) );
  INV_X1 U5671 ( .A(n6804), .ZN(n5203) );
  NOR2_X1 U5672 ( .A1(n5583), .A2(n5201), .ZN(n5200) );
  INV_X1 U5673 ( .A(n8517), .ZN(n5201) );
  AOI21_X1 U5674 ( .B1(n5582), .B2(n5030), .A(n5581), .ZN(n5580) );
  INV_X1 U5675 ( .A(n8667), .ZN(n5581) );
  OR2_X1 U5676 ( .A1(n10516), .A2(n8754), .ZN(n10024) );
  INV_X1 U5677 ( .A(n5510), .ZN(n5509) );
  OAI21_X1 U5678 ( .B1(n5911), .B2(n5511), .A(n5757), .ZN(n5510) );
  INV_X1 U5679 ( .A(n5709), .ZN(n5511) );
  INV_X1 U5680 ( .A(SI_21_), .ZN(n8881) );
  INV_X1 U5681 ( .A(n5494), .ZN(n5493) );
  AND2_X1 U5682 ( .A1(n5495), .A2(n5908), .ZN(n5494) );
  NAND2_X1 U5683 ( .A1(n5780), .A2(n5677), .ZN(n5495) );
  INV_X1 U5684 ( .A(n5677), .ZN(n5492) );
  AOI21_X1 U5685 ( .B1(n5235), .B2(n5233), .A(n5232), .ZN(n5231) );
  INV_X1 U5686 ( .A(n5793), .ZN(n5232) );
  INV_X1 U5687 ( .A(n5237), .ZN(n5233) );
  INV_X1 U5688 ( .A(n5235), .ZN(n5234) );
  INV_X1 U5689 ( .A(SI_14_), .ZN(n9095) );
  INV_X1 U5690 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5650) );
  INV_X1 U5691 ( .A(SI_10_), .ZN(n8898) );
  NAND2_X1 U5692 ( .A1(n5625), .A2(n5850), .ZN(n5216) );
  INV_X1 U5693 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5207) );
  INV_X1 U5694 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5210) );
  INV_X1 U5695 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5209) );
  OAI21_X1 U5696 ( .B1(n6515), .B2(n5028), .A(n9584), .ZN(n5246) );
  OR2_X1 U5697 ( .A1(n6199), .A2(n9343), .ZN(n6220) );
  NAND2_X1 U5698 ( .A1(n5253), .A2(n5256), .ZN(n5250) );
  INV_X1 U5699 ( .A(n8657), .ZN(n5150) );
  INV_X1 U5700 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6158) );
  INV_X1 U5701 ( .A(n5110), .ZN(n6171) );
  INV_X1 U5702 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8954) );
  OR2_X1 U5703 ( .A1(n6127), .A2(n8954), .ZN(n6138) );
  INV_X1 U5704 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8938) );
  INV_X1 U5705 ( .A(n5143), .ZN(n5142) );
  OAI21_X1 U5706 ( .B1(n5547), .B2(n5144), .A(n8499), .ZN(n5143) );
  INV_X1 U5707 ( .A(n8417), .ZN(n5144) );
  INV_X1 U5708 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9175) );
  NOR2_X1 U5709 ( .A1(n6055), .A2(n9175), .ZN(n6066) );
  AND2_X1 U5710 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6047) );
  NAND2_X1 U5711 ( .A1(n9556), .A2(n5338), .ZN(n9496) );
  NOR2_X1 U5712 ( .A1(n5340), .A2(n9498), .ZN(n5338) );
  INV_X1 U5713 ( .A(n5244), .ZN(n9590) );
  AOI21_X1 U5714 ( .B1(n9603), .B2(n6515), .A(n5028), .ZN(n5244) );
  OAI21_X1 U5715 ( .B1(n5784), .B2(n5956), .A(n5785), .ZN(n5470) );
  NOR2_X1 U5716 ( .A1(n7062), .A2(n5559), .ZN(n5558) );
  NAND2_X1 U5717 ( .A1(n7046), .A2(n9865), .ZN(n5559) );
  AND2_X1 U5718 ( .A1(n5565), .A2(n9880), .ZN(n5563) );
  NAND2_X1 U5719 ( .A1(n5567), .A2(n5566), .ZN(n5565) );
  NOR2_X1 U5720 ( .A1(n7251), .A2(n6575), .ZN(n5327) );
  NOR2_X1 U5721 ( .A1(n8785), .A2(n5332), .ZN(n5331) );
  OR2_X1 U5722 ( .A1(n10457), .A2(n10272), .ZN(n10004) );
  NAND2_X1 U5723 ( .A1(n10268), .A2(n5333), .ZN(n5332) );
  NAND2_X1 U5724 ( .A1(n5319), .A2(n8784), .ZN(n5318) );
  NOR2_X1 U5725 ( .A1(n8764), .A2(n5361), .ZN(n5360) );
  INV_X1 U5726 ( .A(n5597), .ZN(n5361) );
  INV_X1 U5727 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6538) );
  NOR2_X1 U5728 ( .A1(n10500), .A2(n5312), .ZN(n5311) );
  INV_X1 U5729 ( .A(n5313), .ZN(n5312) );
  NOR2_X1 U5730 ( .A1(n7993), .A2(n5401), .ZN(n5400) );
  INV_X1 U5731 ( .A(n10052), .ZN(n5401) );
  NAND2_X1 U5732 ( .A1(n7982), .A2(n7903), .ZN(n10119) );
  NAND2_X1 U5733 ( .A1(n7832), .A2(n10210), .ZN(n8021) );
  NAND2_X1 U5734 ( .A1(n10866), .A2(n5324), .ZN(n8678) );
  NAND2_X1 U5735 ( .A1(n10866), .A2(n10867), .ZN(n10865) );
  NAND2_X1 U5736 ( .A1(n5307), .A2(n8014), .ZN(n8153) );
  INV_X1 U5737 ( .A(n8152), .ZN(n5307) );
  OR2_X1 U5738 ( .A1(n7399), .A2(n7398), .ZN(n7422) );
  NAND2_X1 U5739 ( .A1(n5695), .A2(n5522), .ZN(n5521) );
  NOR2_X1 U5740 ( .A1(n5697), .A2(n5523), .ZN(n5522) );
  INV_X1 U5741 ( .A(n5694), .ZN(n5523) );
  NAND2_X1 U5742 ( .A1(n5770), .A2(n5769), .ZN(n5695) );
  NOR2_X1 U5743 ( .A1(n5800), .A2(n5238), .ZN(n5237) );
  INV_X1 U5744 ( .A(n5657), .ZN(n5238) );
  AOI21_X1 U5745 ( .B1(n5239), .B2(n5237), .A(n5236), .ZN(n5235) );
  INV_X1 U5746 ( .A(n5661), .ZN(n5236) );
  AOI21_X1 U5747 ( .B1(n5500), .B2(n5502), .A(n5057), .ZN(n5499) );
  NAND2_X1 U5748 ( .A1(n5638), .A2(n5637), .ZN(n5867) );
  NAND2_X1 U5749 ( .A1(n5212), .A2(SI_6_), .ZN(n5848) );
  OAI21_X1 U5750 ( .B1(n6575), .B2(n5107), .A(n5106), .ZN(n5616) );
  NAND2_X1 U5751 ( .A1(n6575), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5106) );
  OAI211_X1 U5752 ( .C1(n5608), .C2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n5262), .ZN(n5609) );
  INV_X1 U5753 ( .A(n5453), .ZN(n9301) );
  NAND2_X1 U5754 ( .A1(n5460), .A2(n9359), .ZN(n5456) );
  AOI21_X1 U5755 ( .B1(n5455), .B2(n9359), .A(n5034), .ZN(n5454) );
  INV_X1 U5756 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9144) );
  OR2_X1 U5757 ( .A1(n6242), .A2(n9157), .ZN(n6255) );
  NAND2_X1 U5758 ( .A1(n5173), .A2(n5168), .ZN(n6501) );
  NAND2_X1 U5759 ( .A1(n5175), .A2(n5174), .ZN(n5173) );
  NOR2_X1 U5760 ( .A1(n6492), .A2(n6499), .ZN(n5174) );
  OR2_X1 U5761 ( .A1(n5839), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5851) );
  AOI21_X1 U5762 ( .B1(n5037), .B2(n5160), .A(n5156), .ZN(n5155) );
  NAND2_X1 U5763 ( .A1(n9528), .A2(n5483), .ZN(n9510) );
  AND2_X1 U5764 ( .A1(n9511), .A2(n6467), .ZN(n5483) );
  NAND2_X1 U5765 ( .A1(n9556), .A2(n5342), .ZN(n9522) );
  NOR2_X1 U5766 ( .A1(n5481), .A2(n5033), .ZN(n5480) );
  NAND2_X1 U5767 ( .A1(n9556), .A2(n9544), .ZN(n9538) );
  NOR2_X1 U5768 ( .A1(n9557), .A2(n9572), .ZN(n9556) );
  NOR2_X1 U5769 ( .A1(n9588), .A2(n5345), .ZN(n5344) );
  INV_X1 U5770 ( .A(n5346), .ZN(n5345) );
  OR2_X1 U5771 ( .A1(n6177), .A2(n9174), .ZN(n6187) );
  NAND2_X1 U5772 ( .A1(n5110), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U5773 ( .A1(n5249), .A2(n5253), .ZN(n5478) );
  OR2_X1 U5774 ( .A1(n8602), .A2(n5256), .ZN(n5249) );
  NAND2_X1 U5775 ( .A1(n5146), .A2(n5145), .ZN(n9624) );
  AOI21_X1 U5776 ( .B1(n5148), .B2(n5151), .A(n5086), .ZN(n5145) );
  NAND2_X1 U5777 ( .A1(n9651), .A2(n5348), .ZN(n9625) );
  NAND2_X1 U5778 ( .A1(n8602), .A2(n5260), .ZN(n5252) );
  NAND2_X1 U5779 ( .A1(n9651), .A2(n9787), .ZN(n9650) );
  NAND2_X1 U5780 ( .A1(n6147), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6159) );
  AND2_X1 U5781 ( .A1(n8651), .A2(n8609), .ZN(n9651) );
  AND2_X1 U5782 ( .A1(n6425), .A2(n6426), .ZN(n8563) );
  NAND2_X1 U5783 ( .A1(n6105), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U5784 ( .A1(n8090), .A2(n5350), .ZN(n8423) );
  AND2_X1 U5785 ( .A1(n6097), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6105) );
  OR2_X1 U5786 ( .A1(n6076), .A2(n9144), .ZN(n6086) );
  NOR2_X1 U5787 ( .A1(n6086), .A2(n8946), .ZN(n6097) );
  INV_X1 U5788 ( .A(n8289), .ZN(n6335) );
  INV_X1 U5789 ( .A(n8288), .ZN(n6336) );
  OAI21_X1 U5790 ( .B1(n7960), .B2(n5265), .A(n5264), .ZN(n8288) );
  INV_X1 U5791 ( .A(n6334), .ZN(n5265) );
  AOI21_X1 U5792 ( .B1(n5015), .B2(n6334), .A(n5477), .ZN(n5264) );
  INV_X1 U5793 ( .A(n6408), .ZN(n5477) );
  INV_X1 U5794 ( .A(n5532), .ZN(n8081) );
  OAI21_X1 U5795 ( .B1(n8444), .B2(n5531), .A(n5527), .ZN(n5532) );
  NAND2_X1 U5796 ( .A1(n5015), .A2(n7958), .ZN(n5531) );
  INV_X1 U5797 ( .A(n5528), .ZN(n5527) );
  NAND2_X1 U5798 ( .A1(n8090), .A2(n8351), .ZN(n8295) );
  NOR2_X1 U5799 ( .A1(n7916), .A2(n8450), .ZN(n8445) );
  NAND2_X1 U5800 ( .A1(n8212), .A2(n7915), .ZN(n7953) );
  NOR2_X1 U5801 ( .A1(n8064), .A2(n7912), .ZN(n8209) );
  NAND2_X1 U5802 ( .A1(n6383), .A2(n6382), .ZN(n8052) );
  CLKBUF_X1 U5803 ( .A(n6377), .Z(n8051) );
  OR2_X1 U5804 ( .A1(n7755), .A2(n7754), .ZN(n7866) );
  NAND2_X1 U5805 ( .A1(n5525), .A2(n7756), .ZN(n7867) );
  NAND2_X1 U5806 ( .A1(n5756), .A2(n5755), .ZN(n9668) );
  NAND2_X1 U5807 ( .A1(n5482), .A2(n6453), .ZN(n9559) );
  AND2_X1 U5808 ( .A1(n5835), .A2(n5834), .ZN(n10731) );
  NAND2_X1 U5809 ( .A1(n7914), .A2(n7913), .ZN(n8214) );
  INV_X1 U5810 ( .A(n9746), .ZN(n10916) );
  INV_X1 U5811 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5931) );
  NOR2_X1 U5812 ( .A1(n5550), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5337) );
  AND2_X1 U5813 ( .A1(n5958), .A2(n5737), .ZN(n5335) );
  NOR2_X1 U5814 ( .A1(n5782), .A2(n5741), .ZN(n5957) );
  NAND2_X1 U5815 ( .A1(n5123), .A2(n5117), .ZN(n5741) );
  NAND2_X1 U5816 ( .A1(n5951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U5817 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  XNOR2_X1 U5818 ( .A(n5975), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6529) );
  INV_X1 U5819 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5949) );
  XNOR2_X1 U5820 ( .A(n5925), .B(n5924), .ZN(n6001) );
  NAND2_X1 U5821 ( .A1(n5784), .A2(n5295), .ZN(n5294) );
  INV_X1 U5822 ( .A(n5782), .ZN(n5885) );
  OR2_X1 U5823 ( .A1(n5863), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5864) );
  AND2_X1 U5824 ( .A1(n6769), .A2(n6785), .ZN(n5592) );
  NAND2_X1 U5825 ( .A1(n5205), .A2(n6786), .ZN(n8489) );
  NAND2_X1 U5826 ( .A1(n8328), .A2(n6769), .ZN(n5205) );
  NAND2_X1 U5827 ( .A1(n6575), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U5828 ( .A1(n6970), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6985) );
  AND2_X1 U5829 ( .A1(n6649), .A2(n6636), .ZN(n5578) );
  AND2_X1 U5830 ( .A1(n9831), .A2(n5576), .ZN(n5574) );
  AND2_X1 U5831 ( .A1(n5572), .A2(n5087), .ZN(n5570) );
  NAND2_X1 U5832 ( .A1(n5573), .A2(n9831), .ZN(n5572) );
  INV_X1 U5833 ( .A(n5575), .ZN(n5573) );
  XNOR2_X1 U5834 ( .A(n6612), .B(n7652), .ZN(n6614) );
  AND2_X1 U5835 ( .A1(n10053), .A2(n7058), .ZN(n6613) );
  NAND2_X1 U5836 ( .A1(n7044), .A2(n5561), .ZN(n5560) );
  OR2_X1 U5837 ( .A1(n9840), .A2(n7045), .ZN(n7044) );
  NAND2_X1 U5838 ( .A1(n9840), .A2(n7045), .ZN(n7046) );
  INV_X1 U5839 ( .A(n5069), .ZN(n5577) );
  NAND2_X1 U5840 ( .A1(n5516), .A2(n5045), .ZN(n10015) );
  OAI211_X1 U5841 ( .C1(n10009), .C2(n10007), .A(n5519), .B(n5517), .ZN(n5516)
         );
  NAND2_X1 U5842 ( .A1(n10182), .A2(n5097), .ZN(n5096) );
  NOR2_X1 U5843 ( .A1(n10016), .A2(n10017), .ZN(n5097) );
  AND3_X1 U5844 ( .A1(n10019), .A2(n7387), .A3(n5604), .ZN(n10190) );
  AND2_X1 U5845 ( .A1(n10279), .A2(n5328), .ZN(n10256) );
  AND2_X1 U5846 ( .A1(n5331), .A2(n5329), .ZN(n5328) );
  AOI21_X1 U5847 ( .B1(n5410), .B2(n10177), .A(n10001), .ZN(n5408) );
  INV_X1 U5848 ( .A(n5410), .ZN(n5409) );
  INV_X1 U5849 ( .A(n10287), .ZN(n8843) );
  AOI21_X1 U5850 ( .B1(n5365), .B2(n5358), .A(n5063), .ZN(n5357) );
  INV_X1 U5851 ( .A(n5368), .ZN(n5358) );
  OAI21_X1 U5852 ( .B1(n10345), .B2(n5391), .A(n5062), .ZN(n10301) );
  NAND2_X1 U5853 ( .A1(n10117), .A2(n9990), .ZN(n5391) );
  NOR2_X1 U5854 ( .A1(n10301), .A2(n10300), .ZN(n10299) );
  NOR2_X1 U5855 ( .A1(n10354), .A2(n5317), .ZN(n10324) );
  INV_X1 U5856 ( .A(n5319), .ZN(n5317) );
  INV_X1 U5857 ( .A(n6985), .ZN(n6986) );
  NAND2_X1 U5858 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n6986), .ZN(n7002) );
  OAI22_X1 U5859 ( .A1(n10371), .A2(n10372), .B1(n10402), .B2(n10383), .ZN(
        n10353) );
  NAND2_X1 U5860 ( .A1(n10422), .A2(n5311), .ZN(n10378) );
  OAI21_X1 U5861 ( .B1(n8756), .B2(n5380), .A(n5056), .ZN(n5379) );
  NAND2_X1 U5862 ( .A1(n10422), .A2(n8782), .ZN(n10424) );
  OR2_X1 U5863 ( .A1(n6910), .A2(n6909), .ZN(n6930) );
  NAND2_X1 U5864 ( .A1(n10939), .A2(n10031), .ZN(n10434) );
  NAND2_X1 U5865 ( .A1(n6888), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U5866 ( .A1(n10940), .A2(n10941), .ZN(n10939) );
  AND2_X1 U5867 ( .A1(n10866), .A2(n5320), .ZN(n10949) );
  NOR2_X1 U5868 ( .A1(n9929), .A2(n5321), .ZN(n5320) );
  INV_X1 U5869 ( .A(n5322), .ZN(n5321) );
  NOR2_X1 U5870 ( .A1(n6847), .A2(n7802), .ZN(n6871) );
  INV_X1 U5871 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7802) );
  INV_X1 U5872 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6825) );
  OR2_X1 U5873 ( .A1(n6826), .A2(n6825), .ZN(n6847) );
  NOR2_X1 U5874 ( .A1(n6791), .A2(n8518), .ZN(n6809) );
  AND2_X1 U5875 ( .A1(n10806), .A2(n10840), .ZN(n10866) );
  NAND2_X1 U5876 ( .A1(n10068), .A2(n10041), .ZN(n9948) );
  OR2_X1 U5877 ( .A1(n6755), .A2(n8332), .ZN(n6775) );
  OR2_X1 U5878 ( .A1(n6775), .A2(n8492), .ZN(n6791) );
  NOR2_X1 U5879 ( .A1(n10803), .A2(n10828), .ZN(n10806) );
  NAND2_X1 U5880 ( .A1(n8250), .A2(n10776), .ZN(n8310) );
  NAND2_X1 U5881 ( .A1(n5306), .A2(n5305), .ZN(n8251) );
  INV_X1 U5882 ( .A(n8153), .ZN(n5306) );
  NOR2_X1 U5883 ( .A1(n8251), .A2(n8408), .ZN(n8250) );
  INV_X1 U5884 ( .A(n10159), .ZN(n8017) );
  AND2_X1 U5885 ( .A1(n10126), .A2(n9935), .ZN(n10159) );
  AND2_X1 U5886 ( .A1(n7653), .A2(n7652), .ZN(n10737) );
  NOR2_X1 U5887 ( .A1(n7932), .A2(n7903), .ZN(n7988) );
  NAND2_X1 U5888 ( .A1(n5402), .A2(n10052), .ZN(n10124) );
  INV_X1 U5889 ( .A(n10011), .ZN(n10448) );
  INV_X1 U5890 ( .A(n10453), .ZN(n5104) );
  NAND2_X1 U5891 ( .A1(n6753), .A2(n6752), .ZN(n8471) );
  NAND2_X1 U5892 ( .A1(n5417), .A2(n5415), .ZN(n8478) );
  AND2_X1 U5893 ( .A1(n8848), .A2(n10520), .ZN(n10800) );
  OR2_X1 U5894 ( .A1(n10007), .A2(n10115), .ZN(n10520) );
  INV_X1 U5895 ( .A(n10970), .ZN(n10802) );
  INV_X1 U5896 ( .A(n7829), .ZN(n10708) );
  INV_X1 U5897 ( .A(n10973), .ZN(n10927) );
  INV_X1 U5898 ( .A(n7654), .ZN(n10047) );
  INV_X1 U5899 ( .A(n7408), .ZN(n7746) );
  OAI211_X1 U5900 ( .C1(P1_B_REG_SCAN_IN), .C2(n8583), .A(n7085), .B(n7084), 
        .ZN(n7393) );
  XNOR2_X1 U5901 ( .A(n5749), .B(n5748), .ZN(n8830) );
  AND2_X1 U5902 ( .A1(n9271), .A2(n6569), .ZN(n5589) );
  XNOR2_X1 U5903 ( .A(n5753), .B(n5752), .ZN(n8766) );
  OR2_X1 U5904 ( .A1(n6568), .A2(n6806), .ZN(n6570) );
  AND2_X1 U5905 ( .A1(n5421), .A2(n9271), .ZN(n5420) );
  XNOR2_X1 U5906 ( .A(n5758), .B(n5757), .ZN(n8707) );
  NAND2_X1 U5907 ( .A1(n5508), .A2(n5709), .ZN(n5758) );
  AND2_X1 U5908 ( .A1(n6564), .A2(n6563), .ZN(n7082) );
  NAND2_X1 U5909 ( .A1(n7099), .A2(n9048), .ZN(n6561) );
  XNOR2_X1 U5910 ( .A(n7101), .B(n9048), .ZN(n8546) );
  NAND2_X1 U5911 ( .A1(n9246), .A2(n6841), .ZN(n6864) );
  OAI21_X1 U5912 ( .B1(n5894), .B2(n5239), .A(n5657), .ZN(n5801) );
  CLKBUF_X1 U5913 ( .A(n6770), .Z(n6771) );
  XNOR2_X1 U5914 ( .A(n5867), .B(n5601), .ZN(n7293) );
  XNOR2_X1 U5915 ( .A(n5862), .B(n5603), .ZN(n7284) );
  OR2_X1 U5916 ( .A1(n6704), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6724) );
  XNOR2_X1 U5917 ( .A(n5212), .B(n5624), .ZN(n5843) );
  OAI21_X1 U5918 ( .B1(n9316), .B2(n5131), .A(n5129), .ZN(n8859) );
  INV_X1 U5919 ( .A(n5132), .ZN(n5131) );
  AOI21_X1 U5920 ( .B1(n5132), .B2(n5130), .A(n5022), .ZN(n5129) );
  NAND2_X1 U5921 ( .A1(n8585), .A2(n8586), .ZN(n8584) );
  NAND2_X1 U5922 ( .A1(n8525), .A2(n6136), .ZN(n8585) );
  NAND2_X1 U5923 ( .A1(n8545), .A2(n5856), .ZN(n5224) );
  NAND2_X1 U5924 ( .A1(n8093), .A2(n6096), .ZN(n8170) );
  AND2_X1 U5925 ( .A1(n6323), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9374) );
  NAND2_X1 U5926 ( .A1(n5918), .A2(n5917), .ZN(n9674) );
  NAND2_X1 U5927 ( .A1(n5430), .A2(n6301), .ZN(n5429) );
  OAI21_X1 U5928 ( .B1(n5433), .B2(n5430), .A(n5427), .ZN(n5426) );
  MUX2_X1 U5929 ( .A(n6006), .B(n6031), .S(n7754), .Z(n7380) );
  INV_X1 U5930 ( .A(n9531), .ZN(n9564) );
  OAI21_X1 U5931 ( .B1(n9342), .B2(n9341), .A(n5446), .ZN(n9307) );
  AND2_X1 U5932 ( .A1(n5135), .A2(n5134), .ZN(n8436) );
  NAND2_X1 U5933 ( .A1(n8693), .A2(n6170), .ZN(n9326) );
  NAND2_X1 U5934 ( .A1(n5907), .A2(n5906), .ZN(n9627) );
  OR2_X1 U5935 ( .A1(n7706), .A2(n7707), .ZN(n5466) );
  INV_X1 U5936 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9343) );
  INV_X1 U5937 ( .A(n9335), .ZN(n9365) );
  NAND2_X1 U5938 ( .A1(n5892), .A2(n5891), .ZN(n8605) );
  OAI21_X1 U5939 ( .B1(n9342), .B2(n5439), .A(n5436), .ZN(n9349) );
  NAND2_X1 U5940 ( .A1(n5435), .A2(n5440), .ZN(n9351) );
  NAND2_X1 U5941 ( .A1(n9342), .A2(n5442), .ZN(n5435) );
  OAI21_X1 U5942 ( .B1(n8095), .B2(n5451), .A(n5449), .ZN(n8261) );
  AND2_X1 U5943 ( .A1(n9373), .A2(n9619), .ZN(n9335) );
  INV_X1 U5944 ( .A(n9604), .ZN(n9361) );
  OAI21_X1 U5945 ( .B1(n8694), .B2(n5459), .A(n5457), .ZN(n9360) );
  OR2_X1 U5946 ( .A1(n5465), .A2(n7707), .ZN(n5463) );
  INV_X1 U5947 ( .A(n5465), .ZN(n5464) );
  OAI21_X1 U5948 ( .B1(n8525), .B2(n5116), .A(n5115), .ZN(n8639) );
  NOR2_X2 U5949 ( .A1(n6319), .A2(n6305), .ZN(n9352) );
  AND2_X1 U5950 ( .A1(n9373), .A2(n9638), .ZN(n9334) );
  INV_X1 U5951 ( .A(n5939), .ZN(n7761) );
  AND3_X1 U5952 ( .A1(n5938), .A2(n5937), .A3(n5936), .ZN(n7287) );
  OR2_X1 U5953 ( .A1(n9524), .A2(n6317), .ZN(n6239) );
  OR2_X1 U5954 ( .A1(n6357), .A2(n6007), .ZN(n6011) );
  AND2_X1 U5955 ( .A1(n7283), .A2(n7282), .ZN(n8373) );
  INV_X1 U5956 ( .A(n5267), .ZN(n5266) );
  XNOR2_X1 U5957 ( .A(n5269), .B(n8815), .ZN(n5268) );
  AOI22_X1 U5958 ( .A1(n9468), .A2(n9619), .B1(n8816), .B2(n9383), .ZN(n5267)
         );
  AND2_X1 U5959 ( .A1(n9447), .A2(n9446), .ZN(n9677) );
  OAI21_X1 U5960 ( .B1(n9487), .B2(n5536), .A(n5534), .ZN(n9451) );
  NAND2_X1 U5961 ( .A1(n9473), .A2(n9477), .ZN(n9472) );
  NAND2_X1 U5962 ( .A1(n9487), .A2(n8805), .ZN(n9473) );
  NAND2_X1 U5963 ( .A1(n5914), .A2(n5913), .ZN(n9684) );
  OAI21_X1 U5964 ( .B1(n9505), .B2(n9511), .A(n5162), .ZN(n9489) );
  AND2_X1 U5965 ( .A1(n5187), .A2(n5537), .ZN(n9521) );
  NAND2_X1 U5966 ( .A1(n5541), .A2(n5542), .ZN(n9537) );
  NAND2_X1 U5967 ( .A1(n9571), .A2(n5543), .ZN(n5541) );
  AND2_X1 U5968 ( .A1(n5544), .A2(n5040), .ZN(n9555) );
  NAND2_X1 U5969 ( .A1(n9571), .A2(n9577), .ZN(n5544) );
  NAND2_X1 U5970 ( .A1(n9611), .A2(n8803), .ZN(n9585) );
  NAND2_X1 U5971 ( .A1(n8801), .A2(n8800), .ZN(n9647) );
  NAND2_X1 U5972 ( .A1(n5257), .A2(n6340), .ZN(n8648) );
  OR2_X1 U5973 ( .A1(n8602), .A2(n8601), .ZN(n5257) );
  NAND2_X1 U5974 ( .A1(n8418), .A2(n8417), .ZN(n8500) );
  AND2_X1 U5975 ( .A1(n8387), .A2(n8386), .ZN(n8388) );
  NAND2_X1 U5976 ( .A1(n8082), .A2(n6334), .ZN(n8086) );
  NAND2_X1 U5977 ( .A1(n5526), .A2(n7958), .ZN(n8079) );
  NAND2_X1 U5978 ( .A1(n8444), .A2(n7957), .ZN(n5526) );
  NAND2_X1 U5979 ( .A1(n10856), .A2(n5600), .ZN(n9628) );
  OR2_X1 U5980 ( .A1(n8046), .A2(n6274), .ZN(n8615) );
  NAND2_X1 U5981 ( .A1(n10856), .A2(n10848), .ZN(n9602) );
  INV_X1 U5982 ( .A(n9628), .ZN(n9655) );
  INV_X1 U5983 ( .A(n8615), .ZN(n9610) );
  NAND2_X1 U5984 ( .A1(n7269), .A2(n5856), .ZN(n5247) );
  INV_X1 U5985 ( .A(n6362), .ZN(n9755) );
  NAND2_X1 U5986 ( .A1(n5880), .A2(n5879), .ZN(n10852) );
  OAI21_X1 U5987 ( .B1(n5127), .B2(n5128), .A(n7475), .ZN(n5126) );
  NOR2_X1 U5988 ( .A1(n6575), .A2(n7256), .ZN(n5127) );
  NOR2_X1 U5989 ( .A1(n6529), .A2(P2_U3152), .ZN(n10663) );
  INV_X1 U5990 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U5991 ( .A1(n5948), .A2(n5947), .ZN(n8704) );
  INV_X1 U5992 ( .A(n5946), .ZN(n5947) );
  XNOR2_X1 U5993 ( .A(n5955), .B(n5954), .ZN(n8580) );
  NAND2_X1 U5994 ( .A1(n5953), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U5995 ( .A1(n5975), .A2(n5952), .ZN(n5953) );
  INV_X1 U5996 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8540) );
  INV_X1 U5997 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8405) );
  CLKBUF_X1 U5998 ( .A(n6001), .Z(n9407) );
  INV_X1 U5999 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8165) );
  INV_X1 U6000 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7857) );
  INV_X1 U6001 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7377) );
  CLKBUF_X1 U6002 ( .A(n9798), .Z(n9799) );
  NAND2_X1 U6003 ( .A1(n6944), .A2(n6943), .ZN(n10506) );
  NAND2_X1 U6004 ( .A1(n7081), .A2(n7080), .ZN(n8748) );
  INV_X1 U6005 ( .A(n6600), .ZN(n7420) );
  NAND2_X1 U6006 ( .A1(n5571), .A2(n5575), .ZN(n9830) );
  NAND2_X1 U6007 ( .A1(n7029), .A2(n7028), .ZN(n10474) );
  CLKBUF_X1 U6008 ( .A(n9856), .Z(n9857) );
  NAND2_X1 U6009 ( .A1(n5579), .A2(n6636), .ZN(n7897) );
  INV_X1 U6010 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8332) );
  AND2_X1 U6011 ( .A1(n6749), .A2(n8224), .ZN(n8329) );
  NAND2_X1 U6012 ( .A1(n6955), .A2(n6954), .ZN(n9871) );
  AND2_X1 U6013 ( .A1(n5584), .A2(n5036), .ZN(n8664) );
  XNOR2_X1 U6014 ( .A(n6801), .B(n6802), .ZN(n8517) );
  CLKBUF_X1 U6015 ( .A(n8515), .Z(n8516) );
  INV_X1 U6016 ( .A(n9919), .ZN(n9906) );
  CLKBUF_X1 U6017 ( .A(n7940), .Z(n7941) );
  AND2_X1 U6018 ( .A1(n7104), .A2(n7102), .ZN(n9893) );
  OAI21_X1 U6019 ( .B1(n9864), .B2(n5560), .A(n5552), .ZN(n9905) );
  INV_X1 U6020 ( .A(n5553), .ZN(n5552) );
  OAI21_X1 U6021 ( .B1(n5560), .B2(n9865), .A(n7046), .ZN(n5553) );
  NAND2_X1 U6022 ( .A1(n7048), .A2(n7047), .ZN(n10469) );
  CLKBUF_X1 U6023 ( .A(n9912), .Z(n9913) );
  INV_X1 U6024 ( .A(n9903), .ZN(n9928) );
  INV_X1 U6025 ( .A(n9893), .ZN(n9931) );
  INV_X1 U6026 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5628) );
  OR2_X1 U6027 ( .A1(n6699), .A2(n6679), .ZN(n6680) );
  AND2_X1 U6028 ( .A1(n6639), .A2(n5041), .ZN(n5599) );
  AND3_X1 U6029 ( .A1(n6556), .A2(n6553), .A3(n6555), .ZN(n5101) );
  OR2_X1 U6030 ( .A1(n6604), .A2(n6550), .ZN(n6556) );
  OR2_X1 U6031 ( .A1(n5333), .A2(n10272), .ZN(n5595) );
  AND2_X1 U6032 ( .A1(n10284), .A2(n5410), .ZN(n10269) );
  INV_X1 U6033 ( .A(n10464), .ZN(n10268) );
  AOI21_X1 U6034 ( .B1(n10293), .B2(n10300), .A(n5362), .ZN(n10278) );
  INV_X1 U6035 ( .A(n5367), .ZN(n5362) );
  NAND2_X1 U6036 ( .A1(n10331), .A2(n10117), .ZN(n10311) );
  NAND2_X1 U6037 ( .A1(n8763), .A2(n5597), .ZN(n10309) );
  NAND2_X1 U6038 ( .A1(n6984), .A2(n6983), .ZN(n10491) );
  NAND2_X1 U6039 ( .A1(n6969), .A2(n6968), .ZN(n10496) );
  NOR2_X1 U6040 ( .A1(n10417), .A2(n8773), .ZN(n10398) );
  NOR2_X1 U6041 ( .A1(n10407), .A2(n8756), .ZN(n10412) );
  NAND2_X1 U6042 ( .A1(n6887), .A2(n6886), .ZN(n10960) );
  NAND2_X1 U6043 ( .A1(n8752), .A2(n8751), .ZN(n10937) );
  NAND2_X1 U6044 ( .A1(n8711), .A2(n8710), .ZN(n8713) );
  NAND2_X1 U6045 ( .A1(n8675), .A2(n10074), .ZN(n8714) );
  NAND2_X1 U6046 ( .A1(n6846), .A2(n6845), .ZN(n9809) );
  NAND2_X1 U6047 ( .A1(n6824), .A2(n6823), .ZN(n8683) );
  NAND2_X1 U6048 ( .A1(n10863), .A2(n5383), .ZN(n8684) );
  NAND2_X1 U6049 ( .A1(n6790), .A2(n6789), .ZN(n8626) );
  NAND2_X1 U6050 ( .A1(n8303), .A2(n8302), .ZN(n8474) );
  NAND2_X1 U6051 ( .A1(n6729), .A2(n6728), .ZN(n8301) );
  INV_X1 U6052 ( .A(n10792), .ZN(n10959) );
  NAND2_X1 U6053 ( .A1(n8013), .A2(n8012), .ZN(n8150) );
  NAND2_X1 U6054 ( .A1(n10822), .A2(n10743), .ZN(n10792) );
  OR2_X1 U6055 ( .A1(n7399), .A2(n7395), .ZN(n10819) );
  NAND2_X1 U6056 ( .A1(n5105), .A2(n5102), .ZN(n10523) );
  INV_X1 U6057 ( .A(n10454), .ZN(n5105) );
  INV_X1 U6058 ( .A(n5103), .ZN(n5102) );
  OAI21_X1 U6059 ( .B1(n10455), .B2(n10800), .A(n5104), .ZN(n5103) );
  NAND2_X1 U6060 ( .A1(n7409), .A2(n7746), .ZN(n10978) );
  XNOR2_X1 U6061 ( .A(n5733), .B(n5732), .ZN(n10537) );
  CLKBUF_X1 U6062 ( .A(n7126), .Z(n7127) );
  OR2_X1 U6063 ( .A1(n6571), .A2(n6806), .ZN(n5390) );
  INV_X1 U6064 ( .A(n7082), .ZN(n8583) );
  INV_X1 U6065 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8548) );
  AND2_X1 U6066 ( .A1(n5724), .A2(n5013), .ZN(n8544) );
  INV_X1 U6067 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8537) );
  XNOR2_X1 U6068 ( .A(n6581), .B(n9044), .ZN(n8538) );
  INV_X1 U6069 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8326) );
  NAND2_X1 U6070 ( .A1(n6567), .A2(n5027), .ZN(n8327) );
  INV_X1 U6071 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8987) );
  INV_X1 U6072 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9209) );
  INV_X1 U6073 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9007) );
  NOR2_X1 U6074 ( .A1(n5724), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10539) );
  NOR2_X1 U6075 ( .A1(n10610), .A2(n10609), .ZN(n10612) );
  NOR2_X1 U6076 ( .A1(n10608), .A2(n10607), .ZN(n10609) );
  OAI22_X1 U6077 ( .A1(n9430), .A2(n9742), .B1(n10923), .B2(n5980), .ZN(n5981)
         );
  OAI22_X1 U6078 ( .A1(n9430), .A2(n9786), .B1(n5011), .B2(n5990), .ZN(n5991)
         );
  INV_X1 U6079 ( .A(n5309), .ZN(n7099) );
  AND2_X1 U6080 ( .A1(n5165), .A2(n5077), .ZN(n5018) );
  OR2_X1 U6081 ( .A1(n10506), .A2(n10418), .ZN(n5019) );
  OR2_X1 U6082 ( .A1(n9668), .A2(n6351), .ZN(n6367) );
  INV_X1 U6083 ( .A(n10074), .ZN(n5406) );
  OR2_X1 U6084 ( .A1(n5513), .A2(n5843), .ZN(n5020) );
  NAND2_X1 U6085 ( .A1(n7013), .A2(n7012), .ZN(n10481) );
  NAND2_X1 U6086 ( .A1(n5764), .A2(n5763), .ZN(n9498) );
  NAND2_X1 U6087 ( .A1(n5586), .A2(n6544), .ZN(n6565) );
  AND2_X1 U6088 ( .A1(n10069), .A2(n10073), .ZN(n10868) );
  AND2_X1 U6089 ( .A1(n6575), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5021) );
  AND2_X1 U6090 ( .A1(n6278), .A2(n6277), .ZN(n5022) );
  AND2_X1 U6091 ( .A1(n10024), .A2(n10032), .ZN(n10171) );
  INV_X1 U6092 ( .A(n10171), .ZN(n5380) );
  NAND2_X1 U6093 ( .A1(n5216), .A2(n5020), .ZN(n5215) );
  INV_X1 U6094 ( .A(n5540), .ZN(n5539) );
  NAND2_X1 U6095 ( .A1(n5542), .A2(n9545), .ZN(n5540) );
  NAND3_X1 U6096 ( .A1(n5073), .A2(n10103), .A3(n10004), .ZN(n5023) );
  OR2_X1 U6097 ( .A1(n5292), .A2(n5291), .ZN(n5024) );
  NAND2_X1 U6098 ( .A1(n5078), .A2(n5185), .ZN(n5025) );
  AND2_X1 U6099 ( .A1(n5589), .A2(n6548), .ZN(n5026) );
  INV_X1 U6100 ( .A(n5384), .ZN(n5383) );
  NAND2_X1 U6101 ( .A1(n5385), .A2(n8631), .ZN(n5384) );
  NAND2_X2 U6102 ( .A1(n8538), .A2(n10366), .ZN(n10007) );
  NAND2_X1 U6103 ( .A1(n5872), .A2(n5871), .ZN(n8416) );
  INV_X1 U6104 ( .A(n8416), .ZN(n5352) );
  NAND2_X1 U6105 ( .A1(n8245), .A2(n5032), .ZN(n8303) );
  OR2_X1 U6106 ( .A1(n6582), .A2(n5587), .ZN(n5027) );
  NOR2_X1 U6107 ( .A1(n9727), .A2(n9593), .ZN(n5028) );
  NOR2_X1 U6108 ( .A1(n10413), .A2(n10412), .ZN(n5029) );
  AND2_X1 U6109 ( .A1(n8551), .A2(n8550), .ZN(n5030) );
  XNOR2_X1 U6111 ( .A(n5844), .B(n5843), .ZN(n7264) );
  NAND4_X1 U6112 ( .A1(n6590), .A2(n5593), .A3(n6589), .A4(n6588), .ZN(n7651)
         );
  AND2_X1 U6113 ( .A1(n10279), .A2(n5330), .ZN(n5031) );
  NOR2_X1 U6114 ( .A1(n10432), .A2(n10171), .ZN(n10407) );
  INV_X1 U6115 ( .A(n8755), .ZN(n8756) );
  OR2_X1 U6116 ( .A1(n10464), .A2(n8843), .ZN(n10100) );
  AND2_X1 U6117 ( .A1(n9942), .A2(n8020), .ZN(n5032) );
  NOR2_X1 U6118 ( .A1(n9557), .A2(n9547), .ZN(n5033) );
  AND2_X1 U6119 ( .A1(n6185), .A2(n6184), .ZN(n5034) );
  AND2_X1 U6120 ( .A1(n6433), .A2(n8658), .ZN(n5035) );
  NAND2_X1 U6121 ( .A1(n6820), .A2(n6819), .ZN(n5036) );
  NAND2_X1 U6122 ( .A1(n5369), .A2(n5368), .ZN(n10293) );
  AND2_X1 U6123 ( .A1(n5564), .A2(n5570), .ZN(n9879) );
  AND2_X1 U6124 ( .A1(n5158), .A2(n5534), .ZN(n5037) );
  NAND2_X1 U6125 ( .A1(n5627), .A2(n5622), .ZN(n5038) );
  NAND2_X1 U6126 ( .A1(n5799), .A2(n5798), .ZN(n9656) );
  NAND2_X1 U6127 ( .A1(n10020), .A2(n10105), .ZN(n10300) );
  OR2_X1 U6128 ( .A1(n7475), .A2(n7696), .ZN(n5039) );
  NAND2_X1 U6129 ( .A1(n9716), .A2(n9591), .ZN(n5040) );
  INV_X1 U6130 ( .A(n10418), .ZN(n9898) );
  INV_X2 U6131 ( .A(n6163), .ZN(n6179) );
  INV_X1 U6132 ( .A(n9488), .ZN(n9492) );
  AND2_X1 U6133 ( .A1(n6638), .A2(n6637), .ZN(n5041) );
  NAND2_X1 U6134 ( .A1(n6957), .A2(n6956), .ZN(n10500) );
  AND2_X1 U6135 ( .A1(n10021), .A2(n10098), .ZN(n10286) );
  NAND2_X1 U6136 ( .A1(n6808), .A2(n6807), .ZN(n10884) );
  INV_X1 U6137 ( .A(n10484), .ZN(n10329) );
  AND2_X1 U6138 ( .A1(n9998), .A2(n9997), .ZN(n5042) );
  INV_X1 U6139 ( .A(n9588), .ZN(n9777) );
  NAND2_X1 U6140 ( .A1(n5787), .A2(n5786), .ZN(n9588) );
  INV_X1 U6141 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5958) );
  AND2_X1 U6142 ( .A1(n10852), .A2(n9390), .ZN(n5043) );
  AND2_X1 U6143 ( .A1(n10138), .A2(n5392), .ZN(n5044) );
  INV_X1 U6144 ( .A(n6485), .ZN(n5474) );
  OR2_X1 U6145 ( .A1(n9674), .A2(n8862), .ZN(n6485) );
  AND2_X1 U6146 ( .A1(n10182), .A2(n5514), .ZN(n5045) );
  AND2_X1 U6147 ( .A1(n9544), .A2(n9564), .ZN(n5046) );
  NAND2_X1 U6148 ( .A1(n9266), .A2(n9053), .ZN(n5047) );
  INV_X1 U6149 ( .A(n10410), .ZN(n10414) );
  AND2_X1 U6150 ( .A1(n10025), .A2(n10034), .ZN(n10410) );
  AND2_X1 U6151 ( .A1(n6441), .A2(n6442), .ZN(n9646) );
  AND2_X1 U6152 ( .A1(n9679), .A2(n9444), .ZN(n5048) );
  NOR3_X1 U6153 ( .A1(n5017), .A2(n5294), .A3(n5049), .ZN(n5293) );
  INV_X1 U6154 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5744) );
  INV_X1 U6155 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6548) );
  INV_X1 U6156 ( .A(n5583), .ZN(n5582) );
  NAND2_X1 U6157 ( .A1(n8665), .A2(n5036), .ZN(n5583) );
  OR2_X1 U6158 ( .A1(n5919), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5049) );
  NOR2_X1 U6159 ( .A1(n8683), .A2(n10870), .ZN(n5050) );
  AND2_X1 U6160 ( .A1(n5541), .A2(n5539), .ZN(n5051) );
  INV_X1 U6161 ( .A(n5340), .ZN(n5339) );
  NAND2_X1 U6162 ( .A1(n5342), .A2(n5341), .ZN(n5340) );
  INV_X1 U6163 ( .A(n5351), .ZN(n5350) );
  NAND2_X1 U6164 ( .A1(n5353), .A2(n5352), .ZN(n5351) );
  OR2_X1 U6165 ( .A1(n5336), .A2(n5334), .ZN(n5053) );
  NOR2_X1 U6166 ( .A1(n6104), .A2(n6103), .ZN(n5054) );
  NOR2_X1 U6167 ( .A1(n6176), .A2(n6175), .ZN(n5055) );
  NAND2_X1 U6168 ( .A1(n10426), .A2(n10435), .ZN(n5056) );
  NAND2_X1 U6169 ( .A1(n6543), .A2(n6542), .ZN(n6582) );
  NAND2_X1 U6170 ( .A1(n9048), .A2(n5423), .ZN(n5422) );
  INV_X1 U6171 ( .A(n10117), .ZN(n5393) );
  AND2_X1 U6172 ( .A1(n5644), .A2(SI_11_), .ZN(n5057) );
  AND2_X1 U6173 ( .A1(n8806), .A2(n9459), .ZN(n5058) );
  INV_X1 U6174 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5735) );
  AND2_X1 U6175 ( .A1(n5585), .A2(n6545), .ZN(n5059) );
  INV_X1 U6176 ( .A(n5452), .ZN(n5451) );
  NOR2_X1 U6177 ( .A1(n8169), .A2(n6095), .ZN(n5452) );
  INV_X1 U6178 ( .A(n5460), .ZN(n5459) );
  NOR2_X1 U6179 ( .A1(n9325), .A2(n6169), .ZN(n5460) );
  AND2_X1 U6180 ( .A1(n5632), .A2(n5631), .ZN(n5060) );
  NAND2_X1 U6181 ( .A1(n6116), .A2(n6115), .ZN(n5061) );
  OR2_X1 U6182 ( .A1(n5044), .A2(n10023), .ZN(n5062) );
  AND2_X1 U6183 ( .A1(n5364), .A2(n5363), .ZN(n5063) );
  OR2_X1 U6184 ( .A1(n10448), .A2(n10012), .ZN(n10182) );
  NAND2_X1 U6185 ( .A1(n9560), .A2(n5040), .ZN(n5064) );
  INV_X1 U6186 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5784) );
  AND2_X1 U6187 ( .A1(n5452), .A2(n8260), .ZN(n5065) );
  AND2_X1 U6188 ( .A1(n9623), .A2(n6442), .ZN(n5066) );
  AND2_X1 U6189 ( .A1(n8289), .A2(n8282), .ZN(n5067) );
  AND2_X1 U6190 ( .A1(n5311), .A2(n5310), .ZN(n5068) );
  XNOR2_X1 U6191 ( .A(n8770), .B(n10151), .ZN(n10455) );
  XOR2_X1 U6192 ( .A(n6879), .B(n8732), .Z(n5069) );
  AND2_X1 U6193 ( .A1(n10941), .A2(n9966), .ZN(n5070) );
  AND2_X1 U6194 ( .A1(n5580), .A2(n5202), .ZN(n5071) );
  AND2_X1 U6195 ( .A1(n10389), .A2(n9970), .ZN(n5072) );
  NAND2_X1 U6196 ( .A1(n10000), .A2(n10007), .ZN(n5073) );
  AND2_X1 U6197 ( .A1(n9992), .A2(n10175), .ZN(n5074) );
  AND2_X1 U6198 ( .A1(n6371), .A2(n6369), .ZN(n9536) );
  AND2_X1 U6199 ( .A1(n9528), .A2(n6467), .ZN(n5075) );
  NAND2_X1 U6200 ( .A1(n10077), .A2(n10035), .ZN(n10168) );
  AND2_X1 U6201 ( .A1(n9550), .A2(n6371), .ZN(n5076) );
  INV_X1 U6202 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U6203 ( .A1(n6465), .A2(n6464), .ZN(n5077) );
  AND2_X1 U6204 ( .A1(n6437), .A2(n6436), .ZN(n5078) );
  INV_X1 U6205 ( .A(n6451), .ZN(n5289) );
  XNOR2_X1 U6206 ( .A(n7652), .B(n6951), .ZN(n5079) );
  INV_X1 U6207 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5193) );
  INV_X1 U6208 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6209 ( .A1(n8729), .A2(n8728), .ZN(n10457) );
  INV_X1 U6210 ( .A(n10457), .ZN(n5333) );
  NAND2_X1 U6211 ( .A1(n8821), .A2(n8820), .ZN(n10258) );
  INV_X1 U6212 ( .A(n10258), .ZN(n5329) );
  AND2_X1 U6213 ( .A1(n6432), .A2(n6431), .ZN(n8567) );
  INV_X1 U6214 ( .A(n8567), .ZN(n5291) );
  AND2_X1 U6215 ( .A1(n9651), .A2(n5346), .ZN(n5080) );
  AND2_X1 U6216 ( .A1(n10422), .A2(n5068), .ZN(n8783) );
  AND2_X1 U6217 ( .A1(n6372), .A2(n6373), .ZN(n9584) );
  INV_X1 U6218 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5107) );
  INV_X1 U6219 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6220 ( .A1(n5204), .A2(n6804), .ZN(n8549) );
  NAND2_X1 U6221 ( .A1(n5478), .A2(n6442), .ZN(n9616) );
  AND2_X1 U6222 ( .A1(n5252), .A2(n5258), .ZN(n5081) );
  AOI21_X1 U6223 ( .B1(n10432), .B2(n8755), .A(n5379), .ZN(n5376) );
  INV_X1 U6224 ( .A(n9695), .ZN(n5341) );
  OAI21_X1 U6225 ( .B1(n8711), .B2(n5373), .A(n5371), .ZN(n10935) );
  AND2_X1 U6226 ( .A1(n6967), .A2(n6966), .ZN(n5082) );
  NOR2_X1 U6227 ( .A1(n10948), .A2(n10516), .ZN(n10422) );
  NOR3_X1 U6228 ( .A1(n10354), .A2(n10474), .A3(n5318), .ZN(n5315) );
  NAND2_X1 U6229 ( .A1(n6870), .A2(n6869), .ZN(n9929) );
  AND2_X1 U6230 ( .A1(n10863), .A2(n8631), .ZN(n5083) );
  NAND2_X1 U6231 ( .A1(n9556), .A2(n5339), .ZN(n5343) );
  NAND2_X1 U6232 ( .A1(n10422), .A2(n5313), .ZN(n5314) );
  INV_X1 U6233 ( .A(n5316), .ZN(n10316) );
  NOR2_X1 U6234 ( .A1(n10354), .A2(n5318), .ZN(n5316) );
  AND2_X1 U6235 ( .A1(n9589), .A2(n8803), .ZN(n5084) );
  AND2_X1 U6236 ( .A1(n5584), .A2(n5582), .ZN(n5085) );
  INV_X1 U6237 ( .A(n5191), .ZN(n5190) );
  INV_X1 U6238 ( .A(n6301), .ZN(n5433) );
  AND2_X1 U6239 ( .A1(n9656), .A2(n9618), .ZN(n5086) );
  NAND2_X1 U6240 ( .A1(n10866), .A2(n5322), .ZN(n5325) );
  NAND2_X1 U6241 ( .A1(n6982), .A2(n6981), .ZN(n5087) );
  INV_X1 U6242 ( .A(n5537), .ZN(n5188) );
  AOI21_X1 U6243 ( .B1(n5539), .B2(n5538), .A(n5046), .ZN(n5537) );
  INV_X1 U6244 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6806) );
  AND2_X1 U6245 ( .A1(n5524), .A2(n5699), .ZN(n5088) );
  INV_X1 U6246 ( .A(n5596), .ZN(n5561) );
  OR2_X1 U6247 ( .A1(n5017), .A2(n5294), .ZN(n5089) );
  AND2_X1 U6248 ( .A1(n8090), .A2(n5353), .ZN(n5090) );
  NOR2_X1 U6249 ( .A1(n5120), .A2(n5122), .ZN(n5946) );
  NAND2_X1 U6250 ( .A1(n5792), .A2(n5791), .ZN(n9727) );
  INV_X1 U6251 ( .A(n9727), .ZN(n5347) );
  OAI21_X1 U6252 ( .B1(n8306), .B2(n5414), .A(n5411), .ZN(n10807) );
  NAND2_X1 U6253 ( .A1(n8328), .A2(n5592), .ZN(n8488) );
  NAND2_X1 U6254 ( .A1(n5479), .A2(n6332), .ZN(n7917) );
  AND2_X1 U6255 ( .A1(n5417), .A2(n10065), .ZN(n5091) );
  NAND2_X1 U6256 ( .A1(n6336), .A2(n6335), .ZN(n8286) );
  AND2_X1 U6257 ( .A1(n10076), .A2(n10074), .ZN(n10166) );
  INV_X1 U6258 ( .A(n10166), .ZN(n5385) );
  OR2_X1 U6259 ( .A1(n8389), .A2(n6337), .ZN(n5092) );
  AND2_X1 U6260 ( .A1(n5466), .A2(n6045), .ZN(n5093) );
  AND2_X1 U6261 ( .A1(n8245), .A2(n8020), .ZN(n5094) );
  AND2_X1 U6262 ( .A1(n8283), .A2(n8282), .ZN(n5095) );
  INV_X1 U6263 ( .A(n5487), .ZN(n8389) );
  NAND2_X1 U6264 ( .A1(n8286), .A2(n5488), .ZN(n5487) );
  INV_X1 U6265 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5213) );
  NOR2_X1 U6266 ( .A1(n10019), .A2(n5096), .ZN(n10191) );
  AOI21_X2 U6267 ( .B1(n9999), .B2(n5042), .A(n5023), .ZN(n10006) );
  OAI21_X1 U6268 ( .B1(n9972), .B2(n9971), .A(n5072), .ZN(n9974) );
  NAND2_X1 U6269 ( .A1(n5098), .A2(n5070), .ZN(n9968) );
  NAND3_X1 U6270 ( .A1(n9965), .A2(n9963), .A3(n9964), .ZN(n5098) );
  OAI21_X1 U6271 ( .B1(n9994), .B2(n9993), .A(n5074), .ZN(n9996) );
  OAI21_X2 U6272 ( .B1(n8155), .B2(n10127), .A(n10125), .ZN(n9934) );
  OR2_X1 U6273 ( .A1(n7836), .A2(n7654), .ZN(n7828) );
  INV_X1 U6274 ( .A(n10008), .ZN(n5520) );
  NAND2_X1 U6275 ( .A1(n5496), .A2(n5499), .ZN(n5882) );
  NAND2_X1 U6276 ( .A1(n5889), .A2(n5602), .ZN(n5655) );
  OAI211_X1 U6277 ( .C1(n9371), .C2(n5429), .A(n5426), .B(n5424), .ZN(n6306)
         );
  OAI21_X1 U6278 ( .B1(n5781), .B2(n5780), .A(n5677), .ZN(n5909) );
  INV_X1 U6279 ( .A(n5100), .ZN(n6537) );
  NAND4_X1 U6280 ( .A1(n6609), .A2(n6725), .A3(n9015), .A4(n6662), .ZN(n5100)
         );
  INV_X2 U6281 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6662) );
  OAI21_X2 U6282 ( .B1(n9814), .B2(n9815), .A(n9812), .ZN(n9864) );
  NAND2_X2 U6283 ( .A1(n6554), .A2(n5101), .ZN(n7836) );
  NOR2_X2 U6284 ( .A1(n6941), .A2(n6940), .ZN(n9890) );
  NAND2_X1 U6286 ( .A1(n8772), .A2(n10024), .ZN(n10415) );
  OAI21_X1 U6287 ( .B1(n8620), .B2(n5394), .A(n10068), .ZN(n10869) );
  NAND2_X1 U6288 ( .A1(n8489), .A2(n6787), .ZN(n8515) );
  NAND2_X1 U6289 ( .A1(n5199), .A2(n5071), .ZN(n6859) );
  NAND2_X1 U6290 ( .A1(n5578), .A2(n5579), .ZN(n7895) );
  XNOR2_X1 U6291 ( .A(n6614), .B(n6615), .ZN(n7446) );
  NAND2_X1 U6292 ( .A1(n10808), .A2(n10038), .ZN(n8620) );
  NAND2_X1 U6293 ( .A1(n8748), .A2(n5109), .ZN(n7103) );
  NAND2_X2 U6294 ( .A1(n6953), .A2(n6952), .ZN(n6955) );
  NAND2_X1 U6295 ( .A1(n7697), .A2(n7698), .ZN(n5579) );
  NAND2_X1 U6296 ( .A1(n6863), .A2(n9800), .ZN(n6882) );
  NAND2_X1 U6297 ( .A1(n5170), .A2(n5169), .ZN(n5168) );
  NAND2_X1 U6298 ( .A1(n6219), .A2(n6218), .ZN(n6232) );
  NAND2_X1 U6299 ( .A1(n6137), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U6300 ( .A1(n5177), .A2(n5281), .ZN(n5172) );
  NAND2_X1 U6301 ( .A1(n5221), .A2(n6472), .ZN(n5220) );
  INV_X1 U6302 ( .A(n6491), .ZN(n5179) );
  OAI21_X1 U6303 ( .B1(n7817), .B2(n7816), .A(n5111), .ZN(n7818) );
  NAND2_X1 U6304 ( .A1(n7816), .A2(n7817), .ZN(n5111) );
  NAND2_X1 U6305 ( .A1(n8525), .A2(n5115), .ZN(n5114) );
  AND2_X1 U6306 ( .A1(n5739), .A2(n10984), .ZN(n5123) );
  AND2_X1 U6307 ( .A1(n5740), .A2(n5737), .ZN(n5117) );
  NAND3_X1 U6308 ( .A1(n5119), .A2(n5123), .A3(n5118), .ZN(n5944) );
  AND2_X1 U6309 ( .A1(n5734), .A2(n5829), .ZN(n5118) );
  INV_X1 U6310 ( .A(n5122), .ZN(n5119) );
  NAND4_X1 U6311 ( .A1(n5121), .A2(n5739), .A3(n5829), .A4(n5734), .ZN(n5120)
         );
  NAND4_X1 U6312 ( .A1(n5740), .A2(n5958), .A3(n5735), .A4(n5737), .ZN(n5122)
         );
  NAND2_X1 U6313 ( .A1(n5436), .A2(n6197), .ZN(n5124) );
  NAND2_X1 U6314 ( .A1(n5065), .A2(n5136), .ZN(n5134) );
  NAND2_X1 U6315 ( .A1(n7885), .A2(n7884), .ZN(n5133) );
  NAND3_X1 U6316 ( .A1(n5135), .A2(n8437), .A3(n5134), .ZN(n8435) );
  NAND2_X1 U6317 ( .A1(n6085), .A2(n6084), .ZN(n5137) );
  NAND2_X1 U6318 ( .A1(n5833), .A2(n5832), .ZN(n5138) );
  NAND2_X1 U6319 ( .A1(n5822), .A2(n5823), .ZN(n5139) );
  NAND2_X1 U6320 ( .A1(n5140), .A2(n5141), .ZN(n8562) );
  NAND2_X1 U6321 ( .A1(n8387), .A2(n5142), .ZN(n5140) );
  NAND2_X1 U6322 ( .A1(n8659), .A2(n5148), .ZN(n5146) );
  OAI21_X1 U6323 ( .B1(n8659), .B2(n5151), .A(n5148), .ZN(n9649) );
  OAI21_X1 U6324 ( .B1(n8659), .B2(n8658), .A(n8657), .ZN(n8661) );
  NAND2_X1 U6325 ( .A1(n9505), .A2(n5037), .ZN(n5154) );
  NAND2_X1 U6326 ( .A1(n5154), .A2(n5155), .ZN(n8808) );
  NAND2_X1 U6327 ( .A1(n6461), .A2(n5018), .ZN(n5164) );
  NAND3_X1 U6328 ( .A1(n5164), .A2(n5166), .A3(n5163), .ZN(n6466) );
  OAI21_X1 U6329 ( .B1(n6461), .B2(n5167), .A(n5018), .ZN(n6471) );
  OAI21_X2 U6330 ( .B1(n5179), .B2(n6499), .A(n5178), .ZN(n5177) );
  NAND3_X1 U6331 ( .A1(n6422), .A2(n5183), .A3(n6423), .ZN(n5182) );
  NAND2_X1 U6332 ( .A1(n9587), .A2(n5189), .ZN(n5187) );
  NOR2_X1 U6333 ( .A1(n9777), .A2(n9361), .ZN(n5191) );
  MUX2_X1 U6334 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6575), .Z(n5626) );
  MUX2_X1 U6335 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n6575), .Z(n5619) );
  MUX2_X1 U6336 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6575), .Z(n5621) );
  MUX2_X1 U6337 ( .A(n9007), .B(n5628), .S(n6575), .Z(n5629) );
  MUX2_X1 U6338 ( .A(n7292), .B(n5633), .S(n6575), .Z(n5634) );
  MUX2_X1 U6339 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n6575), .Z(n5644) );
  MUX2_X1 U6340 ( .A(n9219), .B(n5639), .S(n6575), .Z(n5640) );
  MUX2_X1 U6341 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6575), .Z(n5656) );
  MUX2_X1 U6342 ( .A(n9210), .B(n7854), .S(n6575), .Z(n5658) );
  MUX2_X1 U6343 ( .A(n9214), .B(n7377), .S(n6575), .Z(n5646) );
  MUX2_X1 U6344 ( .A(n9209), .B(n7857), .S(n6575), .Z(n5662) );
  MUX2_X1 U6345 ( .A(n8998), .B(n5650), .S(n6575), .Z(n5651) );
  NAND2_X1 U6346 ( .A1(n5623), .A2(n5622), .ZN(n5844) );
  NAND3_X1 U6347 ( .A1(n6416), .A2(n6499), .A3(n6415), .ZN(n5194) );
  NAND2_X2 U6348 ( .A1(n7085), .A2(n5196), .ZN(n7160) );
  NAND2_X1 U6349 ( .A1(n6720), .A2(n5197), .ZN(n6716) );
  XNOR2_X1 U6350 ( .A(n8124), .B(n5197), .ZN(n8131) );
  XNOR2_X1 U6351 ( .A(n6714), .B(n5198), .ZN(n5197) );
  INV_X1 U6352 ( .A(n6713), .ZN(n5198) );
  NAND2_X2 U6353 ( .A1(n5208), .A2(n5206), .ZN(n5608) );
  NAND3_X1 U6354 ( .A1(n5207), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5206) );
  NAND3_X1 U6355 ( .A1(n5211), .A2(n5210), .A3(n5209), .ZN(n5208) );
  NAND3_X1 U6356 ( .A1(n5216), .A2(n5020), .A3(n5038), .ZN(n5214) );
  NAND2_X1 U6357 ( .A1(n5894), .A2(n5231), .ZN(n5229) );
  NAND2_X1 U6358 ( .A1(n9603), .A2(n5245), .ZN(n5241) );
  NAND2_X1 U6359 ( .A1(n5242), .A2(n5241), .ZN(n9578) );
  OR2_X2 U6360 ( .A1(n9546), .A2(n9545), .ZN(n9550) );
  NAND2_X1 U6361 ( .A1(n8602), .A2(n5253), .ZN(n5251) );
  NAND3_X1 U6362 ( .A1(n5251), .A2(n5066), .A3(n5250), .ZN(n6343) );
  NAND2_X1 U6363 ( .A1(n5812), .A2(n5811), .ZN(n5612) );
  XNOR2_X1 U6364 ( .A(n5609), .B(SI_1_), .ZN(n5812) );
  NAND2_X1 U6365 ( .A1(n5608), .A2(n5263), .ZN(n5262) );
  NOR2_X1 U6366 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5275) );
  NAND2_X1 U6367 ( .A1(n5276), .A2(n6396), .ZN(n6404) );
  NAND2_X1 U6368 ( .A1(n5277), .A2(n7954), .ZN(n5276) );
  NAND2_X1 U6369 ( .A1(n5280), .A2(n5278), .ZN(n5277) );
  NAND2_X1 U6370 ( .A1(n6392), .A2(n5279), .ZN(n5278) );
  INV_X1 U6371 ( .A(n7915), .ZN(n5279) );
  NAND2_X1 U6372 ( .A1(n5286), .A2(n5285), .ZN(n5284) );
  INV_X1 U6373 ( .A(n6456), .ZN(n5285) );
  OAI21_X1 U6374 ( .B1(n6452), .B2(n6451), .A(n5287), .ZN(n5286) );
  NAND2_X1 U6375 ( .A1(n6458), .A2(n8804), .ZN(n6459) );
  INV_X1 U6376 ( .A(n5293), .ZN(n5921) );
  NOR2_X1 U6377 ( .A1(n5017), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5903) );
  INV_X1 U6378 ( .A(n5296), .ZN(n6489) );
  NAND2_X1 U6379 ( .A1(n6480), .A2(n6479), .ZN(n5302) );
  MUX2_X1 U6380 ( .A(n6382), .B(n6383), .S(n6464), .Z(n5303) );
  NOR2_X2 U6381 ( .A1(n5309), .A2(n5308), .ZN(n6571) );
  INV_X1 U6382 ( .A(n5314), .ZN(n10390) );
  INV_X1 U6383 ( .A(n5315), .ZN(n10294) );
  INV_X1 U6384 ( .A(n5325), .ZN(n8721) );
  NAND2_X1 U6385 ( .A1(n5606), .A2(n5326), .ZN(n7829) );
  NAND2_X1 U6386 ( .A1(n7140), .A2(n5724), .ZN(n6626) );
  NAND2_X2 U6387 ( .A1(n7140), .A2(n6575), .ZN(n8823) );
  NAND2_X1 U6388 ( .A1(n10279), .A2(n5331), .ZN(n10257) );
  NAND2_X1 U6389 ( .A1(n10279), .A2(n10268), .ZN(n10263) );
  NAND4_X1 U6390 ( .A1(n5335), .A2(n5337), .A3(n10984), .A4(n5739), .ZN(n5334)
         );
  NAND3_X1 U6391 ( .A1(n5734), .A2(n5740), .A3(n5829), .ZN(n5336) );
  INV_X1 U6392 ( .A(n5343), .ZN(n9506) );
  NAND2_X1 U6393 ( .A1(n9651), .A2(n5344), .ZN(n9596) );
  NAND4_X1 U6394 ( .A1(n9246), .A2(n6841), .A3(n6903), .A4(n9247), .ZN(n6541)
         );
  NAND2_X1 U6395 ( .A1(n8763), .A2(n5355), .ZN(n5354) );
  NAND2_X1 U6396 ( .A1(n5354), .A2(n5357), .ZN(n10262) );
  NAND2_X1 U6397 ( .A1(n5370), .A2(n8013), .ZN(n8149) );
  OAI21_X1 U6398 ( .B1(n10432), .B2(n5379), .A(n5377), .ZN(n5381) );
  INV_X1 U6399 ( .A(n5381), .ZN(n8758) );
  OAI21_X1 U6400 ( .B1(n8245), .B2(n5388), .A(n5386), .ZN(n10799) );
  XNOR2_X2 U6401 ( .A(n5390), .B(n9271), .ZN(n7155) );
  AOI22_X1 U6402 ( .A1(n10340), .A2(n8761), .B1(n8760), .B2(n10362), .ZN(
        n10323) );
  NOR2_X2 U6403 ( .A1(n8758), .A2(n8757), .ZN(n10371) );
  NAND2_X1 U6404 ( .A1(n7986), .A2(n10155), .ZN(n8013) );
  AND2_X1 U6405 ( .A1(n9671), .A2(n9670), .ZN(n9672) );
  NAND2_X1 U6406 ( .A1(n8246), .A2(n10161), .ZN(n8245) );
  NAND2_X1 U6407 ( .A1(n7834), .A2(n7833), .ZN(n7984) );
  NAND2_X1 U6408 ( .A1(n8018), .A2(n8017), .ZN(n8132) );
  NAND2_X1 U6409 ( .A1(n7925), .A2(n7831), .ZN(n7834) );
  NAND2_X1 U6410 ( .A1(n8628), .A2(n8627), .ZN(n10862) );
  NAND2_X1 U6411 ( .A1(n10935), .A2(n8753), .ZN(n10432) );
  OAI211_X1 U6412 ( .C1(n7126), .C2(n5397), .A(n5396), .B(n5395), .ZN(n5399)
         );
  NAND3_X1 U6413 ( .A1(n7126), .A2(n7155), .A3(n10219), .ZN(n5396) );
  NAND2_X1 U6414 ( .A1(n7924), .A2(n7839), .ZN(n5402) );
  NAND2_X1 U6415 ( .A1(n5402), .A2(n5400), .ZN(n8022) );
  NAND2_X1 U6416 ( .A1(n8675), .A2(n5405), .ZN(n8715) );
  INV_X1 U6417 ( .A(n5407), .ZN(n8842) );
  OAI21_X1 U6418 ( .B1(n10285), .B2(n5409), .A(n5408), .ZN(n5407) );
  INV_X1 U6419 ( .A(n8305), .ZN(n5413) );
  NAND2_X1 U6420 ( .A1(n10939), .A2(n5418), .ZN(n8772) );
  AND2_X1 U6421 ( .A1(n7099), .A2(n5420), .ZN(n6568) );
  NAND2_X1 U6422 ( .A1(n9371), .A2(n5425), .ZN(n5424) );
  OAI21_X1 U6423 ( .B1(n8694), .B2(n5456), .A(n5454), .ZN(n5453) );
  NAND2_X1 U6424 ( .A1(n5461), .A2(n5464), .ZN(n5462) );
  NAND2_X1 U6425 ( .A1(n7731), .A2(n6045), .ZN(n5461) );
  OAI21_X1 U6426 ( .B1(n7706), .B2(n5463), .A(n5462), .ZN(n7816) );
  INV_X1 U6427 ( .A(n5466), .ZN(n7705) );
  NAND2_X1 U6428 ( .A1(n5903), .A2(n5469), .ZN(n5468) );
  NAND2_X1 U6429 ( .A1(n5089), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5790) );
  OAI22_X2 U6430 ( .A1(n9443), .A2(n5471), .B1(n5472), .B2(n6476), .ZN(n6358)
         );
  NOR2_X1 U6431 ( .A1(n5476), .A2(n8350), .ZN(n5475) );
  INV_X1 U6432 ( .A(n7287), .ZN(n5476) );
  NAND3_X1 U6433 ( .A1(n5479), .A2(n6332), .A3(n7954), .ZN(n7920) );
  NAND2_X1 U6434 ( .A1(n9578), .A2(n6344), .ZN(n5482) );
  NAND2_X1 U6435 ( .A1(n5482), .A2(n5480), .ZN(n6346) );
  NAND2_X1 U6436 ( .A1(n5487), .A2(n5485), .ZN(n8420) );
  NAND2_X1 U6437 ( .A1(n10457), .A2(n10272), .ZN(n10103) );
  NAND2_X1 U6438 ( .A1(n5638), .A2(n5497), .ZN(n5496) );
  NAND2_X1 U6439 ( .A1(n5912), .A2(n5911), .ZN(n5508) );
  NAND2_X1 U6440 ( .A1(n5521), .A2(n5088), .ZN(n5705) );
  NAND2_X1 U6441 ( .A1(n5695), .A2(n5694), .ZN(n5766) );
  NAND3_X1 U6442 ( .A1(n7914), .A2(n7913), .A3(n6509), .ZN(n8212) );
  NAND2_X1 U6443 ( .A1(n8283), .A2(n5067), .ZN(n8387) );
  AND2_X1 U6444 ( .A1(n5957), .A2(n5548), .ZN(n5930) );
  NAND2_X1 U6445 ( .A1(n9864), .A2(n5558), .ZN(n5557) );
  AOI21_X1 U6446 ( .B1(n9864), .B2(n9865), .A(n5596), .ZN(n9838) );
  NAND3_X1 U6447 ( .A1(n6955), .A2(n6954), .A3(n5568), .ZN(n5562) );
  NAND2_X1 U6448 ( .A1(n5562), .A2(n5563), .ZN(n7011) );
  NAND3_X1 U6449 ( .A1(n6955), .A2(n6954), .A3(n5574), .ZN(n5564) );
  NAND3_X1 U6450 ( .A1(n6955), .A2(n6954), .A3(n5576), .ZN(n5571) );
  NAND3_X1 U6451 ( .A1(n6863), .A2(n5577), .A3(n9800), .ZN(n9912) );
  NAND2_X1 U6452 ( .A1(n6571), .A2(n5589), .ZN(n6547) );
  NAND2_X1 U6453 ( .A1(n6571), .A2(n5026), .ZN(n5590) );
  INV_X1 U6454 ( .A(n10209), .ZN(n7985) );
  OR2_X1 U6455 ( .A1(n7117), .A2(n7106), .ZN(n7070) );
  OR2_X1 U6456 ( .A1(n7117), .A2(n10280), .ZN(n7054) );
  NAND2_X1 U6457 ( .A1(n10120), .A2(n10122), .ZN(n10155) );
  OR2_X1 U6458 ( .A1(n5930), .A2(n5956), .ZN(n5932) );
  INV_X1 U6459 ( .A(n5934), .ZN(n5995) );
  NAND2_X1 U6460 ( .A1(n6862), .A2(n6861), .ZN(n9800) );
  NAND2_X1 U6461 ( .A1(n6744), .A2(n6748), .ZN(n8224) );
  INV_X1 U6462 ( .A(n6859), .ZN(n6862) );
  AND2_X2 U6463 ( .A1(n8836), .A2(n6552), .ZN(n6655) );
  XNOR2_X1 U6464 ( .A(n6584), .B(n7652), .ZN(n6600) );
  OR2_X1 U6465 ( .A1(n6604), .A2(n10696), .ZN(n5593) );
  INV_X1 U6466 ( .A(n6604), .ZN(n6754) );
  AND2_X1 U6467 ( .A1(n10144), .A2(n10103), .ZN(n5594) );
  AND2_X1 U6468 ( .A1(n7027), .A2(n7026), .ZN(n5596) );
  OR2_X1 U6469 ( .A1(n10329), .A2(n10348), .ZN(n5597) );
  AND2_X1 U6470 ( .A1(n10268), .A2(n8843), .ZN(n5598) );
  NOR2_X1 U6471 ( .A1(n8045), .A2(n6004), .ZN(n5600) );
  AND2_X1 U6472 ( .A1(n5643), .A2(n5642), .ZN(n5601) );
  NAND2_X1 U6473 ( .A1(n7281), .A2(n5940), .ZN(n9565) );
  NAND2_X1 U6474 ( .A1(n10017), .A2(n10049), .ZN(n10018) );
  NAND2_X1 U6475 ( .A1(n5979), .A2(n10702), .ZN(n10914) );
  INV_X1 U6476 ( .A(n10914), .ZN(n9745) );
  AND2_X1 U6477 ( .A1(n5654), .A2(n5653), .ZN(n5602) );
  AND2_X1 U6478 ( .A1(n5637), .A2(n5636), .ZN(n5603) );
  INV_X1 U6479 ( .A(n7404), .ZN(n6329) );
  AND2_X1 U6480 ( .A1(n10115), .A2(n10366), .ZN(n5604) );
  AND3_X1 U6481 ( .A1(n6326), .A2(n6325), .A3(n6324), .ZN(n5605) );
  NAND2_X2 U6482 ( .A1(n8046), .A2(n10860), .ZN(n10856) );
  INV_X2 U6483 ( .A(n10856), .ZN(n10851) );
  AND2_X1 U6484 ( .A1(n7382), .A2(n6308), .ZN(n9379) );
  INV_X2 U6486 ( .A(n10922), .ZN(n10923) );
  INV_X1 U6487 ( .A(n9684), .ZN(n8806) );
  INV_X1 U6488 ( .A(n10426), .ZN(n8782) );
  OR2_X1 U6489 ( .A1(n6241), .A2(n6240), .ZN(n5607) );
  INV_X1 U6490 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9053) );
  INV_X1 U6491 ( .A(n6415), .ZN(n6337) );
  NAND2_X1 U6492 ( .A1(n6754), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6637) );
  INV_X1 U6493 ( .A(n6220), .ZN(n6219) );
  INV_X1 U6494 ( .A(n6138), .ZN(n6137) );
  INV_X1 U6495 ( .A(n6187), .ZN(n6186) );
  INV_X1 U6496 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8946) );
  INV_X1 U6497 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5743) );
  INV_X1 U6498 ( .A(n7898), .ZN(n6649) );
  INV_X1 U6499 ( .A(n9822), .ZN(n6952) );
  INV_X1 U6500 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8518) );
  INV_X1 U6501 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6695) );
  INV_X1 U6502 ( .A(n10868), .ZN(n8629) );
  NAND2_X1 U6503 ( .A1(n7985), .A2(n7991), .ZN(n10120) );
  INV_X1 U6504 ( .A(SI_22_), .ZN(n5685) );
  NOR2_X1 U6505 ( .A1(n10702), .A2(n6003), .ZN(n6005) );
  OR2_X1 U6506 ( .A1(n6255), .A2(n9320), .ZN(n6267) );
  NAND2_X1 U6507 ( .A1(n6231), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6242) );
  INV_X1 U6508 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9174) );
  OR2_X1 U6509 ( .A1(n6117), .A2(n8938), .ZN(n6127) );
  OR2_X1 U6510 ( .A1(n9498), .A2(n9513), .ZN(n8805) );
  NAND2_X1 U6511 ( .A1(n6186), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6199) );
  INV_X1 U6512 ( .A(n6318), .ZN(n5979) );
  INV_X1 U6513 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5956) );
  INV_X1 U6514 ( .A(n9850), .ZN(n6898) );
  AND2_X1 U6515 ( .A1(n6871), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6888) );
  OAI22_X1 U6516 ( .A1(n10272), .A2(n10401), .B1(n8826), .B2(n10109), .ZN(
        n8779) );
  AND2_X1 U6517 ( .A1(n6945), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6958) );
  INV_X1 U6518 ( .A(n10407), .ZN(n10408) );
  OR2_X1 U6519 ( .A1(n8471), .A2(n10811), .ZN(n8472) );
  NAND2_X1 U6520 ( .A1(n5916), .A2(n5915), .ZN(n5719) );
  OR2_X1 U6521 ( .A1(n6884), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6885) );
  INV_X1 U6522 ( .A(SI_11_), .ZN(n9102) );
  INV_X1 U6523 ( .A(n9374), .ZN(n9363) );
  INV_X1 U6524 ( .A(n8350), .ZN(n7760) );
  AND2_X1 U6525 ( .A1(n8811), .A2(n6293), .ZN(n9438) );
  OR2_X1 U6526 ( .A1(n6034), .A2(n8102), .ZN(n6009) );
  INV_X1 U6527 ( .A(n9480), .ZN(n9454) );
  AND2_X1 U6528 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  AND2_X1 U6529 ( .A1(n10702), .A2(n6004), .ZN(n9746) );
  INV_X1 U6530 ( .A(n9390), .ZN(n8506) );
  OAI21_X1 U6531 ( .B1(n5974), .B2(n5973), .A(n10550), .ZN(n6302) );
  INV_X1 U6532 ( .A(n9644), .ZN(n9561) );
  INV_X1 U6533 ( .A(n6764), .ZN(n6995) );
  AND3_X1 U6534 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6677) );
  NOR2_X1 U6535 ( .A1(n6930), .A2(n9896), .ZN(n6945) );
  OR2_X1 U6536 ( .A1(n6699), .A2(n7112), .ZN(n7121) );
  AND2_X1 U6537 ( .A1(n6958), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6970) );
  INV_X1 U6538 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8492) );
  INV_X1 U6539 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9896) );
  INV_X1 U6540 ( .A(n8779), .ZN(n8780) );
  AND2_X1 U6541 ( .A1(n10496), .A2(n10374), .ZN(n8759) );
  OR2_X1 U6542 ( .A1(n7393), .A2(P1_D_REG_0__SCAN_IN), .ZN(n7086) );
  INV_X1 U6543 ( .A(n8327), .ZN(n10115) );
  AND2_X1 U6544 ( .A1(n7655), .A2(n10016), .ZN(n10873) );
  AND2_X1 U6545 ( .A1(n8546), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7135) );
  AND2_X1 U6546 ( .A1(n5681), .A2(n5680), .ZN(n5908) );
  OR3_X1 U6547 ( .A1(n8580), .A2(n8704), .A3(n8689), .ZN(n7137) );
  NOR2_X1 U6548 ( .A1(n6319), .A2(n6530), .ZN(n9373) );
  AND2_X1 U6549 ( .A1(n6249), .A2(n6248), .ZN(n9294) );
  NAND2_X1 U6550 ( .A1(n6017), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6019) );
  INV_X1 U6551 ( .A(n9422), .ZN(n10684) );
  AND2_X1 U6552 ( .A1(n7494), .A2(n5940), .ZN(n10680) );
  INV_X1 U6553 ( .A(n8809), .ZN(n9442) );
  AND2_X1 U6554 ( .A1(n6469), .A2(n6468), .ZN(n9511) );
  INV_X1 U6555 ( .A(n9565), .ZN(n9638) );
  INV_X1 U6556 ( .A(n6307), .ZN(n8041) );
  NAND2_X1 U6557 ( .A1(n8040), .A2(n8039), .ZN(n8046) );
  INV_X1 U6558 ( .A(n9602), .ZN(n9660) );
  INV_X1 U6559 ( .A(n7754), .ZN(n10701) );
  AND2_X1 U6560 ( .A1(n8393), .A2(n8316), .ZN(n9750) );
  OR2_X1 U6561 ( .A1(n6303), .A2(n8041), .ZN(n5987) );
  INV_X1 U6562 ( .A(n9750), .ZN(n10921) );
  AND3_X1 U6563 ( .A1(n6004), .A2(n6002), .A3(n5939), .ZN(n10836) );
  AND2_X1 U6564 ( .A1(n7137), .A2(n10663), .ZN(n10552) );
  INV_X1 U6565 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5922) );
  OAI21_X1 U6566 ( .B1(n10268), .B2(n9903), .A(n7131), .ZN(n7132) );
  AND2_X1 U6567 ( .A1(n6941), .A2(n6940), .ZN(n9894) );
  AND4_X1 U6568 ( .A1(n7122), .A2(n7121), .A3(n7120), .A4(n7119), .ZN(n10272)
         );
  INV_X1 U6569 ( .A(n10651), .ZN(n10216) );
  OR2_X1 U6570 ( .A1(P1_U3083), .A2(n7161), .ZN(n7784) );
  INV_X1 U6571 ( .A(n7784), .ZN(n10648) );
  AND2_X1 U6572 ( .A1(n10822), .A2(n7847), .ZN(n10786) );
  INV_X1 U6573 ( .A(n10873), .ZN(n10947) );
  INV_X1 U6574 ( .A(n8848), .ZN(n10876) );
  AND2_X1 U6575 ( .A1(n7086), .A2(n10536), .ZN(n7408) );
  AND2_X1 U6576 ( .A1(n7846), .A2(n8327), .ZN(n10973) );
  INV_X1 U6577 ( .A(n10800), .ZN(n10952) );
  INV_X1 U6578 ( .A(n10520), .ZN(n10879) );
  NAND2_X1 U6579 ( .A1(n7160), .A2(n7135), .ZN(n7399) );
  NOR2_X1 U6580 ( .A1(n10576), .A2(n10575), .ZN(n10577) );
  NOR2_X1 U6581 ( .A1(n10604), .A2(n10603), .ZN(n10605) );
  NOR2_X1 U6582 ( .A1(n7137), .A2(P2_U3152), .ZN(n7471) );
  INV_X1 U6583 ( .A(n9334), .ZN(n9362) );
  INV_X1 U6584 ( .A(n9705), .ZN(n9544) );
  INV_X1 U6585 ( .A(n9379), .ZN(n9358) );
  NAND2_X1 U6586 ( .A1(n6288), .A2(n6287), .ZN(n9444) );
  INV_X1 U6587 ( .A(P2_U3966), .ZN(n9385) );
  INV_X1 U6588 ( .A(n10680), .ZN(n10668) );
  NAND2_X1 U6589 ( .A1(n7494), .A2(n7493), .ZN(n10689) );
  NAND2_X1 U6590 ( .A1(n10552), .A2(n8041), .ZN(n10860) );
  NAND2_X1 U6591 ( .A1(n10923), .A2(n9745), .ZN(n9742) );
  OR2_X1 U6592 ( .A1(n5987), .A2(n5978), .ZN(n10922) );
  INV_X1 U6593 ( .A(n9498), .ZN(n9765) );
  INV_X1 U6594 ( .A(n9656), .ZN(n9787) );
  NAND2_X1 U6595 ( .A1(n5011), .A2(n9745), .ZN(n9786) );
  NAND2_X1 U6596 ( .A1(n10552), .A2(n10551), .ZN(n10661) );
  INV_X1 U6597 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8543) );
  INV_X1 U6598 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7854) );
  INV_X1 U6599 ( .A(n7132), .ZN(n7133) );
  INV_X1 U6600 ( .A(n9900), .ZN(n9926) );
  AND2_X1 U6601 ( .A1(n7105), .A2(n10819), .ZN(n9903) );
  AND3_X1 U6602 ( .A1(n7299), .A2(n7298), .A3(n7297), .ZN(n10012) );
  OR2_X1 U6603 ( .A1(n6950), .A2(n6949), .ZN(n10418) );
  OR2_X2 U6604 ( .A1(n7160), .A2(n7136), .ZN(n10211) );
  INV_X1 U6605 ( .A(n10786), .ZN(n10429) );
  NAND2_X1 U6606 ( .A1(n10822), .A2(n10737), .ZN(n10406) );
  AND2_X2 U6607 ( .A1(n7409), .A2(n7408), .ZN(n10977) );
  INV_X1 U6608 ( .A(n10977), .ZN(n10975) );
  INV_X2 U6609 ( .A(n10978), .ZN(n10981) );
  OR2_X1 U6610 ( .A1(n7265), .A2(n7399), .ZN(n10549) );
  INV_X1 U6611 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9195) );
  INV_X1 U6612 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9210) );
  NOR2_X1 U6613 ( .A1(n10606), .A2(n10605), .ZN(n10608) );
  AND2_X2 U6614 ( .A1(n7471), .A2(n7138), .ZN(P2_U3966) );
  INV_X1 U6615 ( .A(n10211), .ZN(P1_U4006) );
  MUX2_X1 U6616 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5608), .Z(n5811) );
  INV_X1 U6617 ( .A(n5609), .ZN(n5610) );
  NAND2_X1 U6618 ( .A1(n5610), .A2(SI_1_), .ZN(n5611) );
  NAND2_X1 U6619 ( .A1(n5612), .A2(n5611), .ZN(n5817) );
  MUX2_X1 U6620 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5608), .Z(n5613) );
  INV_X1 U6621 ( .A(SI_2_), .ZN(n9120) );
  XNOR2_X1 U6622 ( .A(n5613), .B(n9120), .ZN(n5816) );
  NAND2_X1 U6623 ( .A1(n5817), .A2(n5816), .ZN(n5615) );
  NAND2_X1 U6624 ( .A1(n5613), .A2(SI_2_), .ZN(n5614) );
  INV_X1 U6625 ( .A(SI_3_), .ZN(n9119) );
  XNOR2_X1 U6626 ( .A(n5616), .B(n9119), .ZN(n5822) );
  NAND2_X1 U6627 ( .A1(n5616), .A2(SI_3_), .ZN(n5617) );
  INV_X1 U6628 ( .A(SI_4_), .ZN(n5618) );
  XNOR2_X1 U6629 ( .A(n5619), .B(n5618), .ZN(n5832) );
  NAND2_X1 U6630 ( .A1(n5619), .A2(SI_4_), .ZN(n5620) );
  INV_X1 U6631 ( .A(SI_5_), .ZN(n8909) );
  XNOR2_X1 U6632 ( .A(n5621), .B(n8909), .ZN(n5836) );
  NAND2_X1 U6633 ( .A1(n5837), .A2(n5836), .ZN(n5623) );
  NAND2_X1 U6634 ( .A1(n5621), .A2(SI_5_), .ZN(n5622) );
  INV_X1 U6635 ( .A(SI_6_), .ZN(n5624) );
  NAND2_X1 U6636 ( .A1(n5626), .A2(SI_7_), .ZN(n5625) );
  AND2_X1 U6637 ( .A1(n5848), .A2(n5625), .ZN(n5627) );
  XNOR2_X1 U6638 ( .A(n5626), .B(SI_7_), .ZN(n5850) );
  NAND2_X1 U6639 ( .A1(n5629), .A2(n9110), .ZN(n5632) );
  INV_X1 U6640 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U6641 ( .A1(n5630), .A2(SI_8_), .ZN(n5631) );
  INV_X1 U6642 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U6643 ( .A1(n5634), .A2(n9109), .ZN(n5637) );
  INV_X1 U6644 ( .A(n5634), .ZN(n5635) );
  NAND2_X1 U6645 ( .A1(n5635), .A2(SI_9_), .ZN(n5636) );
  INV_X1 U6646 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U6647 ( .A1(n5640), .A2(n8898), .ZN(n5643) );
  INV_X1 U6648 ( .A(n5640), .ZN(n5641) );
  NAND2_X1 U6649 ( .A1(n5641), .A2(SI_10_), .ZN(n5642) );
  XNOR2_X1 U6650 ( .A(n5644), .B(n9102), .ZN(n5873) );
  INV_X1 U6651 ( .A(n5873), .ZN(n5645) );
  NAND2_X1 U6652 ( .A1(n5646), .A2(n9101), .ZN(n5649) );
  INV_X1 U6653 ( .A(n5646), .ZN(n5647) );
  NAND2_X1 U6654 ( .A1(n5647), .A2(SI_12_), .ZN(n5648) );
  NAND2_X1 U6655 ( .A1(n5649), .A2(n5648), .ZN(n5881) );
  NAND2_X1 U6656 ( .A1(n5651), .A2(n9094), .ZN(n5654) );
  INV_X1 U6657 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U6658 ( .A1(n5652), .A2(SI_13_), .ZN(n5653) );
  XNOR2_X1 U6659 ( .A(n5656), .B(n9095), .ZN(n5893) );
  NAND2_X1 U6660 ( .A1(n5656), .A2(SI_14_), .ZN(n5657) );
  NAND2_X1 U6661 ( .A1(n5658), .A2(n8890), .ZN(n5661) );
  INV_X1 U6662 ( .A(n5658), .ZN(n5659) );
  NAND2_X1 U6663 ( .A1(n5659), .A2(SI_15_), .ZN(n5660) );
  NAND2_X1 U6664 ( .A1(n5661), .A2(n5660), .ZN(n5800) );
  NAND2_X1 U6665 ( .A1(n5662), .A2(n9096), .ZN(n5665) );
  INV_X1 U6666 ( .A(n5662), .ZN(n5663) );
  NAND2_X1 U6667 ( .A1(n5663), .A2(SI_16_), .ZN(n5664) );
  MUX2_X1 U6668 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5724), .Z(n5667) );
  XNOR2_X1 U6669 ( .A(n5667), .B(n5666), .ZN(n5901) );
  INV_X1 U6670 ( .A(n5901), .ZN(n5669) );
  NAND2_X1 U6671 ( .A1(n5667), .A2(SI_17_), .ZN(n5668) );
  MUX2_X1 U6672 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5724), .Z(n5671) );
  XNOR2_X1 U6673 ( .A(n5671), .B(SI_18_), .ZN(n5788) );
  INV_X1 U6674 ( .A(n5788), .ZN(n5670) );
  NAND2_X1 U6675 ( .A1(n5671), .A2(SI_18_), .ZN(n5672) );
  MUX2_X1 U6676 ( .A(n8165), .B(n8987), .S(n5724), .Z(n5674) );
  INV_X1 U6677 ( .A(SI_19_), .ZN(n8883) );
  NAND2_X1 U6678 ( .A1(n5674), .A2(n8883), .ZN(n5677) );
  INV_X1 U6679 ( .A(n5674), .ZN(n5675) );
  NAND2_X1 U6680 ( .A1(n5675), .A2(SI_19_), .ZN(n5676) );
  NAND2_X1 U6681 ( .A1(n5677), .A2(n5676), .ZN(n5780) );
  MUX2_X1 U6682 ( .A(n8405), .B(n8326), .S(n5724), .Z(n5678) );
  INV_X1 U6683 ( .A(SI_20_), .ZN(n8882) );
  NAND2_X1 U6684 ( .A1(n5678), .A2(n8882), .ZN(n5681) );
  INV_X1 U6685 ( .A(n5678), .ZN(n5679) );
  NAND2_X1 U6686 ( .A1(n5679), .A2(SI_20_), .ZN(n5680) );
  MUX2_X1 U6687 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5724), .Z(n5683) );
  XNOR2_X1 U6688 ( .A(n5683), .B(n8881), .ZN(n5776) );
  INV_X1 U6689 ( .A(n5776), .ZN(n5682) );
  NAND2_X1 U6690 ( .A1(n5683), .A2(SI_21_), .ZN(n5684) );
  MUX2_X1 U6691 ( .A(n8540), .B(n8537), .S(n5724), .Z(n5686) );
  NAND2_X1 U6692 ( .A1(n5686), .A2(n5685), .ZN(n5689) );
  INV_X1 U6693 ( .A(n5686), .ZN(n5687) );
  NAND2_X1 U6694 ( .A1(n5687), .A2(SI_22_), .ZN(n5688) );
  NAND2_X1 U6695 ( .A1(n5689), .A2(n5688), .ZN(n5772) );
  OAI21_X1 U6696 ( .B1(n5773), .B2(n5772), .A(n5689), .ZN(n5770) );
  MUX2_X1 U6697 ( .A(n8543), .B(n8548), .S(n5724), .Z(n5691) );
  INV_X1 U6698 ( .A(SI_23_), .ZN(n5690) );
  NAND2_X1 U6699 ( .A1(n5691), .A2(n5690), .ZN(n5694) );
  INV_X1 U6700 ( .A(n5691), .ZN(n5692) );
  NAND2_X1 U6701 ( .A1(n5692), .A2(SI_23_), .ZN(n5693) );
  MUX2_X1 U6702 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n5724), .Z(n5698) );
  INV_X1 U6703 ( .A(SI_24_), .ZN(n5696) );
  XNOR2_X1 U6704 ( .A(n5698), .B(n5696), .ZN(n5765) );
  INV_X1 U6705 ( .A(n5765), .ZN(n5697) );
  NAND2_X1 U6706 ( .A1(n5698), .A2(SI_24_), .ZN(n5699) );
  INV_X1 U6707 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8692) );
  MUX2_X1 U6708 ( .A(n8692), .B(n9195), .S(n5724), .Z(n5701) );
  INV_X1 U6709 ( .A(SI_25_), .ZN(n5700) );
  NAND2_X1 U6710 ( .A1(n5701), .A2(n5700), .ZN(n5704) );
  INV_X1 U6711 ( .A(n5701), .ZN(n5702) );
  NAND2_X1 U6712 ( .A1(n5702), .A2(SI_25_), .ZN(n5703) );
  NAND2_X1 U6713 ( .A1(n5704), .A2(n5703), .ZN(n5761) );
  INV_X1 U6714 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8703) );
  INV_X1 U6715 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9191) );
  MUX2_X1 U6716 ( .A(n8703), .B(n9191), .S(n5724), .Z(n5706) );
  INV_X1 U6717 ( .A(SI_26_), .ZN(n8872) );
  NAND2_X1 U6718 ( .A1(n5706), .A2(n8872), .ZN(n5709) );
  INV_X1 U6719 ( .A(n5706), .ZN(n5707) );
  NAND2_X1 U6720 ( .A1(n5707), .A2(SI_26_), .ZN(n5708) );
  INV_X1 U6721 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8708) );
  INV_X1 U6722 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9190) );
  MUX2_X1 U6723 ( .A(n8708), .B(n9190), .S(n5724), .Z(n5711) );
  INV_X1 U6724 ( .A(SI_27_), .ZN(n5710) );
  NAND2_X1 U6725 ( .A1(n5711), .A2(n5710), .ZN(n5714) );
  INV_X1 U6726 ( .A(n5711), .ZN(n5712) );
  NAND2_X1 U6727 ( .A1(n5712), .A2(SI_27_), .ZN(n5713) );
  MUX2_X1 U6728 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5724), .Z(n5715) );
  INV_X1 U6729 ( .A(SI_28_), .ZN(n5716) );
  XNOR2_X1 U6730 ( .A(n5715), .B(n5716), .ZN(n5915) );
  INV_X1 U6731 ( .A(n5715), .ZN(n5717) );
  NAND2_X1 U6732 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  MUX2_X1 U6733 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5724), .Z(n5720) );
  INV_X1 U6734 ( .A(SI_29_), .ZN(n9075) );
  XNOR2_X1 U6735 ( .A(n5720), .B(n9075), .ZN(n5752) );
  NAND2_X1 U6736 ( .A1(n5753), .A2(n5752), .ZN(n5723) );
  INV_X1 U6737 ( .A(n5720), .ZN(n5721) );
  NAND2_X1 U6738 ( .A1(n5721), .A2(n9075), .ZN(n5722) );
  MUX2_X1 U6739 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n5724), .Z(n5725) );
  INV_X1 U6740 ( .A(SI_30_), .ZN(n5726) );
  XNOR2_X1 U6741 ( .A(n5725), .B(n5726), .ZN(n5748) );
  NAND2_X1 U6742 ( .A1(n5749), .A2(n5748), .ZN(n5729) );
  INV_X1 U6743 ( .A(n5725), .ZN(n5727) );
  NAND2_X1 U6744 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  NAND2_X1 U6745 ( .A1(n5729), .A2(n5728), .ZN(n5733) );
  MUX2_X1 U6746 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n5724), .Z(n5731) );
  INV_X1 U6747 ( .A(SI_31_), .ZN(n5730) );
  XNOR2_X1 U6748 ( .A(n5731), .B(n5730), .ZN(n5732) );
  NAND2_X1 U6749 ( .A1(n5924), .A2(n5927), .ZN(n5919) );
  INV_X1 U6750 ( .A(n5919), .ZN(n5740) );
  NOR2_X1 U6753 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5737) );
  NAND2_X1 U6754 ( .A1(n5053), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5745) );
  XNOR2_X2 U6755 ( .A(n5745), .B(n5744), .ZN(n5940) );
  INV_X2 U6756 ( .A(n5845), .ZN(n5856) );
  NAND2_X1 U6757 ( .A1(n10537), .A2(n5856), .ZN(n5747) );
  INV_X1 U6758 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9790) );
  OR2_X1 U6759 ( .A1(n5824), .A2(n9790), .ZN(n5746) );
  NAND2_X1 U6760 ( .A1(n8830), .A2(n5856), .ZN(n5751) );
  INV_X1 U6761 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8832) );
  OR2_X1 U6762 ( .A1(n5824), .A2(n8832), .ZN(n5750) );
  NAND2_X1 U6763 ( .A1(n5751), .A2(n5750), .ZN(n6362) );
  NAND2_X1 U6764 ( .A1(n8766), .A2(n5856), .ZN(n5756) );
  INV_X1 U6765 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5754) );
  OR2_X1 U6766 ( .A1(n5824), .A2(n5754), .ZN(n5755) );
  NAND2_X1 U6767 ( .A1(n8707), .A2(n5856), .ZN(n5760) );
  OR2_X1 U6768 ( .A1(n5824), .A2(n8708), .ZN(n5759) );
  INV_X1 U6769 ( .A(n9679), .ZN(n9458) );
  XNOR2_X1 U6770 ( .A(n5762), .B(n5761), .ZN(n8687) );
  NAND2_X1 U6771 ( .A1(n8687), .A2(n5856), .ZN(n5764) );
  OR2_X1 U6772 ( .A1(n5824), .A2(n8692), .ZN(n5763) );
  XNOR2_X1 U6773 ( .A(n5766), .B(n5765), .ZN(n8578) );
  NAND2_X1 U6774 ( .A1(n8578), .A2(n5856), .ZN(n5768) );
  INV_X1 U6775 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8579) );
  OR2_X1 U6776 ( .A1(n5824), .A2(n8579), .ZN(n5767) );
  OR2_X1 U6777 ( .A1(n5824), .A2(n8543), .ZN(n5771) );
  XNOR2_X1 U6778 ( .A(n5773), .B(n5772), .ZN(n8536) );
  NAND2_X1 U6779 ( .A1(n8536), .A2(n5856), .ZN(n5775) );
  OR2_X1 U6780 ( .A1(n5824), .A2(n8540), .ZN(n5774) );
  XNOR2_X1 U6781 ( .A(n5777), .B(n5776), .ZN(n8348) );
  NAND2_X1 U6782 ( .A1(n8348), .A2(n5856), .ZN(n5779) );
  INV_X1 U6783 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8349) );
  OR2_X1 U6784 ( .A1(n5824), .A2(n8349), .ZN(n5778) );
  XNOR2_X1 U6785 ( .A(n5781), .B(n5780), .ZN(n8163) );
  NAND2_X1 U6786 ( .A1(n8163), .A2(n5856), .ZN(n5787) );
  NAND3_X1 U6787 ( .A1(n5802), .A2(n5895), .A3(n5804), .ZN(n5783) );
  AOI22_X1 U6788 ( .A1(n5905), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6002), .B2(
        n7279), .ZN(n5786) );
  XNOR2_X1 U6789 ( .A(n5789), .B(n5788), .ZN(n7965) );
  NAND2_X1 U6790 ( .A1(n7965), .A2(n5856), .ZN(n5792) );
  XNOR2_X1 U6791 ( .A(n5790), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9414) );
  AOI22_X1 U6792 ( .A1(n5905), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7279), .B2(
        n9414), .ZN(n5791) );
  XNOR2_X1 U6793 ( .A(n5794), .B(n5793), .ZN(n7856) );
  NAND2_X1 U6794 ( .A1(n7856), .A2(n5856), .ZN(n5799) );
  NAND2_X1 U6795 ( .A1(n5017), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5795) );
  MUX2_X1 U6796 ( .A(n5795), .B(P2_IR_REG_31__SCAN_IN), .S(n5295), .Z(n5797)
         );
  INV_X1 U6797 ( .A(n5903), .ZN(n5796) );
  NAND2_X1 U6798 ( .A1(n5797), .A2(n5796), .ZN(n8364) );
  INV_X1 U6799 ( .A(n8364), .ZN(n8377) );
  AOI22_X1 U6800 ( .A1(n5905), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7279), .B2(
        n8377), .ZN(n5798) );
  XNOR2_X1 U6801 ( .A(n5801), .B(n5800), .ZN(n7853) );
  NAND2_X1 U6802 ( .A1(n7853), .A2(n5856), .ZN(n5808) );
  NAND2_X1 U6803 ( .A1(n5890), .A2(n5802), .ZN(n5803) );
  NAND2_X1 U6804 ( .A1(n5803), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U6805 ( .A1(n5896), .A2(n5895), .ZN(n5898) );
  NAND2_X1 U6806 ( .A1(n5898), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5805) );
  XNOR2_X1 U6807 ( .A(n5805), .B(n5804), .ZN(n8185) );
  INV_X1 U6808 ( .A(n8185), .ZN(n5806) );
  AOI22_X1 U6809 ( .A1(n5905), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7279), .B2(
        n5806), .ZN(n5807) );
  INV_X1 U6810 ( .A(n9744), .ZN(n8651) );
  INV_X1 U6811 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U6812 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5809) );
  XNOR2_X1 U6813 ( .A(n5810), .B(n5809), .ZN(n7696) );
  XNOR2_X1 U6814 ( .A(n5812), .B(n5811), .ZN(n7257) );
  INV_X1 U6815 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7256) );
  INV_X1 U6816 ( .A(SI_0_), .ZN(n8906) );
  NOR2_X1 U6817 ( .A1(n5724), .A2(n8906), .ZN(n5813) );
  XNOR2_X1 U6818 ( .A(n5813), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9796) );
  MUX2_X1 U6819 ( .A(n5271), .B(n9796), .S(n7475), .Z(n7754) );
  OR2_X1 U6820 ( .A1(n5814), .A2(n5956), .ZN(n5815) );
  XNOR2_X1 U6821 ( .A(n5815), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10679) );
  INV_X1 U6822 ( .A(n10679), .ZN(n7247) );
  XNOR2_X1 U6823 ( .A(n5817), .B(n5816), .ZN(n7251) );
  OR2_X1 U6824 ( .A1(n5845), .A2(n7251), .ZN(n5819) );
  INV_X1 U6825 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7248) );
  OR2_X1 U6826 ( .A1(n5824), .A2(n7248), .ZN(n5818) );
  OR3_X1 U6827 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U6828 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5820), .ZN(n5821) );
  XNOR2_X1 U6829 ( .A(n5821), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7499) );
  INV_X1 U6830 ( .A(n7499), .ZN(n7521) );
  XNOR2_X1 U6831 ( .A(n5823), .B(n5822), .ZN(n7255) );
  OR2_X1 U6832 ( .A1(n7255), .A2(n5845), .ZN(n5826) );
  INV_X1 U6833 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7249) );
  OR2_X1 U6834 ( .A1(n5824), .A2(n7249), .ZN(n5825) );
  NOR2_X1 U6835 ( .A1(n5829), .A2(n5956), .ZN(n5827) );
  MUX2_X1 U6836 ( .A(n5956), .B(n5827), .S(P2_IR_REG_4__SCAN_IN), .Z(n5831) );
  INV_X1 U6837 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U6838 ( .A1(n5829), .A2(n5828), .ZN(n5839) );
  INV_X1 U6839 ( .A(n5839), .ZN(n5830) );
  NOR2_X1 U6840 ( .A1(n5831), .A2(n5830), .ZN(n7608) );
  AOI22_X1 U6841 ( .A1(n5905), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7279), .B2(
        n7608), .ZN(n5835) );
  XNOR2_X1 U6842 ( .A(n5833), .B(n5832), .ZN(n7259) );
  OR2_X1 U6843 ( .A1(n7259), .A2(n5845), .ZN(n5834) );
  NAND2_X1 U6844 ( .A1(n8209), .A2(n10731), .ZN(n8211) );
  XNOR2_X1 U6845 ( .A(n5837), .B(n5836), .ZN(n7262) );
  OR2_X1 U6846 ( .A1(n7262), .A2(n5845), .ZN(n5842) );
  NAND2_X1 U6847 ( .A1(n5839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5838) );
  MUX2_X1 U6848 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5838), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5840) );
  AND2_X1 U6849 ( .A1(n5840), .A2(n5851), .ZN(n7545) );
  AOI22_X1 U6850 ( .A1(n5905), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7279), .B2(
        n7545), .ZN(n5841) );
  NAND2_X1 U6851 ( .A1(n5851), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5846) );
  XNOR2_X1 U6852 ( .A(n5846), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7571) );
  AOI22_X1 U6853 ( .A1(n5905), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7279), .B2(
        n7571), .ZN(n5847) );
  NOR2_X1 U6854 ( .A1(n5851), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5858) );
  OR2_X1 U6855 ( .A1(n5858), .A2(n5956), .ZN(n5852) );
  XNOR2_X1 U6856 ( .A(n5852), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7583) );
  AOI22_X1 U6857 ( .A1(n5905), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7279), .B2(
        n7583), .ZN(n5853) );
  INV_X1 U6858 ( .A(n8463), .ZN(n8344) );
  AND2_X1 U6859 ( .A1(n8445), .A2(n8344), .ZN(n8090) );
  NAND2_X1 U6860 ( .A1(n5855), .A2(n5854), .ZN(n7273) );
  NAND2_X1 U6861 ( .A1(n7273), .A2(n5856), .ZN(n5861) );
  INV_X1 U6862 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U6863 ( .A1(n5858), .A2(n5857), .ZN(n5863) );
  NAND2_X1 U6864 ( .A1(n5863), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5859) );
  XNOR2_X1 U6865 ( .A(n5859), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7558) );
  AOI22_X1 U6866 ( .A1(n5905), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7279), .B2(
        n7558), .ZN(n5860) );
  NAND2_X1 U6867 ( .A1(n5861), .A2(n5860), .ZN(n8281) );
  INV_X1 U6868 ( .A(n8281), .ZN(n8351) );
  NAND2_X1 U6869 ( .A1(n7284), .A2(n5856), .ZN(n5866) );
  NAND2_X1 U6870 ( .A1(n5864), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5869) );
  XNOR2_X1 U6871 ( .A(n5869), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7596) );
  AOI22_X1 U6872 ( .A1(n5905), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7279), .B2(
        n7596), .ZN(n5865) );
  NAND2_X1 U6873 ( .A1(n5866), .A2(n5865), .ZN(n8385) );
  NAND2_X1 U6874 ( .A1(n7293), .A2(n5856), .ZN(n5872) );
  INV_X1 U6875 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U6876 ( .A1(n5869), .A2(n5868), .ZN(n5870) );
  NAND2_X1 U6877 ( .A1(n5870), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5876) );
  XNOR2_X1 U6878 ( .A(n5876), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7629) );
  AOI22_X1 U6879 ( .A1(n5905), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7279), .B2(
        n7629), .ZN(n5871) );
  XNOR2_X1 U6880 ( .A(n5874), .B(n5873), .ZN(n7329) );
  NAND2_X1 U6881 ( .A1(n7329), .A2(n5856), .ZN(n5880) );
  INV_X1 U6882 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U6883 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  NAND2_X1 U6884 ( .A1(n5877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5878) );
  XNOR2_X1 U6885 ( .A(n5878), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7630) );
  AOI22_X1 U6886 ( .A1(n5905), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7630), .B2(
        n7279), .ZN(n5879) );
  XNOR2_X1 U6887 ( .A(n5882), .B(n5881), .ZN(n7374) );
  NAND2_X1 U6888 ( .A1(n7374), .A2(n5856), .ZN(n5888) );
  NOR2_X1 U6889 ( .A1(n5883), .A2(n5956), .ZN(n5884) );
  MUX2_X1 U6890 ( .A(n5956), .B(n5884), .S(P2_IR_REG_12__SCAN_IN), .Z(n5886)
         );
  NOR2_X1 U6891 ( .A1(n5886), .A2(n5885), .ZN(n7625) );
  AOI22_X1 U6892 ( .A1(n5905), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7279), .B2(
        n7625), .ZN(n5887) );
  NAND2_X1 U6893 ( .A1(n5888), .A2(n5887), .ZN(n8564) );
  INV_X1 U6894 ( .A(n8564), .ZN(n10892) );
  NAND2_X1 U6895 ( .A1(n8507), .A2(n10892), .ZN(n8572) );
  XNOR2_X1 U6896 ( .A(n5889), .B(n5602), .ZN(n7428) );
  NAND2_X1 U6897 ( .A1(n7428), .A2(n5856), .ZN(n5892) );
  XNOR2_X1 U6898 ( .A(n5890), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7723) );
  AOI22_X1 U6899 ( .A1(n5905), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7279), .B2(
        n7723), .ZN(n5891) );
  XNOR2_X1 U6900 ( .A(n5894), .B(n5893), .ZN(n7468) );
  NAND2_X1 U6901 ( .A1(n7468), .A2(n5856), .ZN(n5900) );
  OR2_X1 U6902 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  AND2_X1 U6903 ( .A1(n5898), .A2(n5897), .ZN(n7972) );
  AOI22_X1 U6904 ( .A1(n5905), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7279), .B2(
        n7972), .ZN(n5899) );
  XNOR2_X1 U6905 ( .A(n5902), .B(n5901), .ZN(n7880) );
  NAND2_X1 U6906 ( .A1(n7880), .A2(n5856), .ZN(n5907) );
  OR2_X1 U6907 ( .A1(n5903), .A2(n5956), .ZN(n5904) );
  XNOR2_X1 U6908 ( .A(n5904), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9400) );
  AOI22_X1 U6909 ( .A1(n5905), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7279), .B2(
        n9400), .ZN(n5906) );
  XNOR2_X1 U6910 ( .A(n5909), .B(n5908), .ZN(n8325) );
  OR2_X1 U6911 ( .A1(n5824), .A2(n8405), .ZN(n5910) );
  NAND2_X1 U6912 ( .A1(n8702), .A2(n5856), .ZN(n5914) );
  OR2_X1 U6913 ( .A1(n5824), .A2(n8703), .ZN(n5913) );
  NAND2_X1 U6914 ( .A1(n9458), .A2(n9480), .ZN(n9452) );
  NAND2_X1 U6915 ( .A1(n8834), .A2(n5856), .ZN(n5918) );
  INV_X1 U6916 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8835) );
  OR2_X1 U6917 ( .A1(n5824), .A2(n8835), .ZN(n5917) );
  NAND2_X1 U6918 ( .A1(n9755), .A2(n9431), .ZN(n9663) );
  XOR2_X1 U6919 ( .A(n6363), .B(n9663), .Z(n9426) );
  NAND2_X1 U6920 ( .A1(n5293), .A2(n5922), .ZN(n5920) );
  NAND2_X1 U6921 ( .A1(n5921), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U6922 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  NAND2_X1 U6923 ( .A1(n5930), .A2(n5931), .ZN(n9792) );
  NAND2_X1 U6924 ( .A1(n6179), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5938) );
  NAND2_X4 U6925 ( .A1(n8833), .A2(n5994), .ZN(n6357) );
  INV_X1 U6926 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5980) );
  OR2_X1 U6927 ( .A1(n6357), .A2(n5980), .ZN(n5937) );
  NAND2_X4 U6928 ( .A1(n5995), .A2(n8750), .ZN(n6034) );
  INV_X1 U6929 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n5935) );
  OR2_X1 U6930 ( .A1(n6034), .A2(n5935), .ZN(n5936) );
  NAND2_X1 U6931 ( .A1(n7761), .A2(n7760), .ZN(n7470) );
  INV_X1 U6932 ( .A(P2_B_REG_SCAN_IN), .ZN(n5961) );
  OR2_X1 U6933 ( .A1(n5941), .A2(n5961), .ZN(n5942) );
  AND2_X1 U6934 ( .A1(n9638), .A2(n5942), .ZN(n8816) );
  INV_X1 U6935 ( .A(n8816), .ZN(n5943) );
  NOR2_X1 U6936 ( .A1(n7287), .A2(n5943), .ZN(n9427) );
  AOI21_X1 U6937 ( .B1(n9426), .B2(n9746), .A(n9427), .ZN(n5989) );
  INV_X1 U6938 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10553) );
  NAND2_X1 U6939 ( .A1(n5944), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5945) );
  MUX2_X1 U6940 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5945), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5948) );
  INV_X1 U6941 ( .A(n8580), .ZN(n5962) );
  OR2_X1 U6942 ( .A1(n5957), .A2(n5956), .ZN(n5959) );
  MUX2_X1 U6943 ( .A(n5959), .B(P2_IR_REG_31__SCAN_IN), .S(n5958), .Z(n5960)
         );
  NAND2_X1 U6944 ( .A1(n5960), .A2(n5944), .ZN(n8689) );
  OAI221_X1 U6945 ( .B1(P2_B_REG_SCAN_IN), .B2(n5962), .C1(n5961), .C2(n8580), 
        .A(n8689), .ZN(n5963) );
  INV_X1 U6946 ( .A(n5963), .ZN(n5964) );
  AND2_X1 U6947 ( .A1(n8689), .A2(n8704), .ZN(n10554) );
  AOI21_X1 U6948 ( .B1(n10553), .B2(n10550), .A(n10554), .ZN(n6303) );
  NAND2_X1 U6949 ( .A1(n10836), .A2(n8350), .ZN(n6307) );
  NOR4_X1 U6950 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5968) );
  NOR4_X1 U6951 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5967) );
  NOR4_X1 U6952 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5966) );
  NOR4_X1 U6953 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5965) );
  NAND4_X1 U6954 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(n5974)
         );
  NOR2_X1 U6955 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5972) );
  NOR4_X1 U6956 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5971) );
  NOR4_X1 U6957 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5970) );
  NOR4_X1 U6958 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5969) );
  NAND4_X1 U6959 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(n5973)
         );
  NAND2_X1 U6960 ( .A1(n5979), .A2(n7281), .ZN(n6321) );
  NAND2_X1 U6961 ( .A1(n10552), .A2(n6321), .ZN(n7381) );
  AND2_X1 U6962 ( .A1(n8580), .A2(n8704), .ZN(n10664) );
  INV_X1 U6963 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10662) );
  AND2_X1 U6964 ( .A1(n10550), .A2(n10662), .ZN(n5976) );
  NOR2_X1 U6965 ( .A1(n7381), .A2(n8038), .ZN(n5977) );
  NAND2_X1 U6966 ( .A1(n6302), .A2(n5977), .ZN(n5978) );
  OR2_X1 U6967 ( .A1(n5989), .A2(n10922), .ZN(n5983) );
  INV_X1 U6968 ( .A(n5981), .ZN(n5982) );
  NAND2_X1 U6969 ( .A1(n5983), .A2(n5982), .ZN(P2_U3551) );
  INV_X1 U6970 ( .A(n8038), .ZN(n5984) );
  NOR2_X1 U6971 ( .A1(n7381), .A2(n5984), .ZN(n5985) );
  NAND2_X1 U6972 ( .A1(n6302), .A2(n5985), .ZN(n5986) );
  OR2_X1 U6973 ( .A1(n5989), .A2(n10985), .ZN(n5993) );
  INV_X1 U6974 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n5990) );
  INV_X1 U6975 ( .A(n5991), .ZN(n5992) );
  NAND2_X1 U6976 ( .A1(n5993), .A2(n5992), .ZN(P2_U3519) );
  NAND2_X1 U6977 ( .A1(n6179), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6000) );
  INV_X1 U6978 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8043) );
  OR2_X1 U6979 ( .A1(n6025), .A2(n8043), .ZN(n5999) );
  NAND2_X1 U6980 ( .A1(n6017), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5998) );
  INV_X1 U6981 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5996) );
  OR2_X1 U6982 ( .A1(n6034), .A2(n5996), .ZN(n5997) );
  AND4_X2 U6983 ( .A1(n6000), .A2(n5999), .A3(n5998), .A4(n5997), .ZN(n7755)
         );
  NOR2_X1 U6984 ( .A1(n7755), .A2(n6299), .ZN(n6006) );
  INV_X1 U6985 ( .A(n6001), .ZN(n6002) );
  INV_X1 U6986 ( .A(n6004), .ZN(n6506) );
  NAND2_X2 U6987 ( .A1(n6005), .A2(n7767), .ZN(n6031) );
  INV_X1 U6988 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U6989 ( .A1(n6298), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6010) );
  INV_X1 U6990 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U6991 ( .A1(n6179), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6008) );
  INV_X2 U6992 ( .A(n6299), .ZN(n6274) );
  NAND2_X1 U6993 ( .A1(n7404), .A2(n6274), .ZN(n6013) );
  OAI21_X1 U6994 ( .B1(n6013), .B2(n6012), .A(n6014), .ZN(n7379) );
  INV_X1 U6995 ( .A(n6014), .ZN(n6015) );
  NOR2_X1 U6996 ( .A1(n7378), .A2(n6015), .ZN(n7403) );
  XOR2_X1 U6997 ( .A(n6031), .B(n8061), .Z(n6024) );
  NAND2_X1 U6998 ( .A1(n6179), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6021) );
  INV_X1 U6999 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7000 ( .A1(n6025), .A2(n6016), .ZN(n6020) );
  INV_X1 U7001 ( .A(n6357), .ZN(n6017) );
  INV_X1 U7002 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8067) );
  OR2_X1 U7003 ( .A1(n6034), .A2(n8067), .ZN(n6018) );
  NAND4_X1 U7004 ( .A1(n6021), .A2(n6020), .A3(n6019), .A4(n6018), .ZN(n9397)
         );
  NAND2_X1 U7005 ( .A1(n9397), .A2(n6274), .ZN(n6022) );
  XNOR2_X1 U7006 ( .A(n6024), .B(n6022), .ZN(n7402) );
  INV_X1 U7007 ( .A(n6022), .ZN(n6023) );
  OR2_X1 U7008 ( .A1(n6025), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7009 ( .A1(n6179), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6029) );
  INV_X1 U7010 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6026) );
  OR2_X1 U7011 ( .A1(n6357), .A2(n6026), .ZN(n6028) );
  INV_X1 U7012 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7520) );
  OR2_X1 U7013 ( .A1(n6034), .A2(n7520), .ZN(n6027) );
  NAND4_X1 U7014 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n9396)
         );
  NAND2_X1 U7015 ( .A1(n9396), .A2(n6274), .ZN(n6032) );
  XNOR2_X1 U7016 ( .A(n7912), .B(n6031), .ZN(n6033) );
  XNOR2_X1 U7017 ( .A(n6032), .B(n6033), .ZN(n7789) );
  OAI22_X1 U7018 ( .A1(n7790), .A2(n7789), .B1(n6033), .B2(n6032), .ZN(n7706)
         );
  XOR2_X1 U7019 ( .A(n10731), .B(n6031), .Z(n6044) );
  NAND2_X1 U7020 ( .A1(n6311), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6042) );
  INV_X1 U7021 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6035) );
  OR2_X1 U7022 ( .A1(n6163), .A2(n6035), .ZN(n6041) );
  INV_X1 U7023 ( .A(n6047), .ZN(n6037) );
  INV_X1 U7024 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9139) );
  INV_X1 U7025 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U7026 ( .A1(n9139), .A2(n9156), .ZN(n6036) );
  NAND2_X1 U7027 ( .A1(n6037), .A2(n6036), .ZN(n8216) );
  OR2_X1 U7028 ( .A1(n6317), .A2(n8216), .ZN(n6040) );
  INV_X1 U7029 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6038) );
  OR2_X1 U7030 ( .A1(n6357), .A2(n6038), .ZN(n6039) );
  NAND4_X1 U7031 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n9395)
         );
  NAND2_X1 U7032 ( .A1(n9395), .A2(n6274), .ZN(n6043) );
  NAND2_X1 U7033 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  OAI21_X1 U7034 ( .B1(n6044), .B2(n6043), .A(n6045), .ZN(n7707) );
  XNOR2_X1 U7035 ( .A(n10753), .B(n6254), .ZN(n6054) );
  NAND2_X1 U7036 ( .A1(n6352), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6051) );
  INV_X1 U7037 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6046) );
  OR2_X1 U7038 ( .A1(n6357), .A2(n6046), .ZN(n6050) );
  NAND2_X1 U7039 ( .A1(n6047), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6055) );
  OAI21_X1 U7040 ( .B1(n6047), .B2(P2_REG3_REG_5__SCAN_IN), .A(n6055), .ZN(
        n10752) );
  OR2_X1 U7041 ( .A1(n6317), .A2(n10752), .ZN(n6049) );
  INV_X1 U7042 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7525) );
  OR2_X1 U7043 ( .A1(n6034), .A2(n7525), .ZN(n6048) );
  NAND2_X1 U7044 ( .A1(n8455), .A2(n6274), .ZN(n6052) );
  XNOR2_X1 U7045 ( .A(n6054), .B(n6052), .ZN(n7731) );
  INV_X1 U7046 ( .A(n6052), .ZN(n6053) );
  XNOR2_X1 U7047 ( .A(n8450), .B(n6254), .ZN(n6063) );
  NAND2_X1 U7048 ( .A1(n6179), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6061) );
  INV_X1 U7049 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7526) );
  OR2_X1 U7050 ( .A1(n6034), .A2(n7526), .ZN(n6060) );
  AND2_X1 U7051 ( .A1(n6055), .A2(n9175), .ZN(n6056) );
  OR2_X1 U7052 ( .A1(n6056), .A2(n6066), .ZN(n8448) );
  OR2_X1 U7053 ( .A1(n6317), .A2(n8448), .ZN(n6059) );
  INV_X1 U7054 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6057) );
  OR2_X1 U7055 ( .A1(n6284), .A2(n6057), .ZN(n6058) );
  NAND4_X1 U7056 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n9394)
         );
  AND2_X1 U7057 ( .A1(n9394), .A2(n6274), .ZN(n6062) );
  NOR2_X1 U7058 ( .A1(n6063), .A2(n6062), .ZN(n6064) );
  AOI21_X1 U7059 ( .B1(n6063), .B2(n6062), .A(n6064), .ZN(n7817) );
  INV_X1 U7060 ( .A(n6064), .ZN(n6065) );
  XNOR2_X1 U7061 ( .A(n8463), .B(n6031), .ZN(n6074) );
  NAND2_X1 U7062 ( .A1(n6352), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6072) );
  INV_X1 U7063 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7529) );
  OR2_X1 U7064 ( .A1(n6034), .A2(n7529), .ZN(n6071) );
  NAND2_X1 U7065 ( .A1(n6066), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6076) );
  OR2_X1 U7066 ( .A1(n6066), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7067 ( .A1(n6076), .A2(n6067), .ZN(n8461) );
  OR2_X1 U7068 ( .A1(n6317), .A2(n8461), .ZN(n6070) );
  INV_X1 U7069 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6068) );
  OR2_X1 U7070 ( .A1(n6357), .A2(n6068), .ZN(n6069) );
  NAND4_X1 U7071 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n9393)
         );
  NAND2_X1 U7072 ( .A1(n9393), .A2(n6274), .ZN(n6073) );
  XNOR2_X1 U7073 ( .A(n6074), .B(n6073), .ZN(n7871) );
  OAI22_X2 U7074 ( .A1(n7872), .A2(n7871), .B1(n6074), .B2(n6073), .ZN(n7885)
         );
  XNOR2_X1 U7075 ( .A(n8281), .B(n6254), .ZN(n6085) );
  NAND2_X1 U7076 ( .A1(n6311), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6082) );
  INV_X1 U7077 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6075) );
  OR2_X1 U7078 ( .A1(n6163), .A2(n6075), .ZN(n6081) );
  NAND2_X1 U7079 ( .A1(n6076), .A2(n9144), .ZN(n6077) );
  NAND2_X1 U7080 ( .A1(n6086), .A2(n6077), .ZN(n8196) );
  OR2_X1 U7081 ( .A1(n6317), .A2(n8196), .ZN(n6080) );
  INV_X1 U7082 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6078) );
  OR2_X1 U7083 ( .A1(n6357), .A2(n6078), .ZN(n6079) );
  NAND4_X1 U7084 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(n9392)
         );
  NAND2_X1 U7085 ( .A1(n9392), .A2(n6274), .ZN(n6083) );
  XNOR2_X1 U7086 ( .A(n6085), .B(n6083), .ZN(n7884) );
  INV_X1 U7087 ( .A(n6083), .ZN(n6084) );
  XNOR2_X1 U7088 ( .A(n8385), .B(n6254), .ZN(n6094) );
  NAND2_X1 U7089 ( .A1(n6179), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6092) );
  INV_X1 U7090 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8294) );
  OR2_X1 U7091 ( .A1(n6034), .A2(n8294), .ZN(n6091) );
  AND2_X1 U7092 ( .A1(n6086), .A2(n8946), .ZN(n6087) );
  OR2_X1 U7093 ( .A1(n6087), .A2(n6097), .ZN(n8296) );
  OR2_X1 U7094 ( .A1(n6317), .A2(n8296), .ZN(n6090) );
  INV_X1 U7095 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6088) );
  OR2_X1 U7096 ( .A1(n6284), .A2(n6088), .ZN(n6089) );
  NAND4_X1 U7097 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n8394)
         );
  AND2_X1 U7098 ( .A1(n8394), .A2(n6274), .ZN(n6093) );
  NOR2_X1 U7099 ( .A1(n6094), .A2(n6093), .ZN(n6095) );
  AOI21_X1 U7100 ( .B1(n6094), .B2(n6093), .A(n6095), .ZN(n8094) );
  INV_X1 U7101 ( .A(n6095), .ZN(n6096) );
  XNOR2_X1 U7102 ( .A(n8416), .B(n6031), .ZN(n6104) );
  NAND2_X1 U7103 ( .A1(n6352), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6102) );
  INV_X1 U7104 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8399) );
  OR2_X1 U7105 ( .A1(n6034), .A2(n8399), .ZN(n6101) );
  NOR2_X1 U7106 ( .A1(n6097), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6098) );
  OR2_X1 U7107 ( .A1(n6105), .A2(n6098), .ZN(n8398) );
  OR2_X1 U7108 ( .A1(n6317), .A2(n8398), .ZN(n6100) );
  INV_X1 U7109 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7510) );
  OR2_X1 U7110 ( .A1(n6357), .A2(n7510), .ZN(n6099) );
  NAND4_X1 U7111 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(n9391)
         );
  NAND2_X1 U7112 ( .A1(n9391), .A2(n6274), .ZN(n6103) );
  XNOR2_X1 U7113 ( .A(n6104), .B(n6103), .ZN(n8169) );
  NAND2_X1 U7114 ( .A1(n6352), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6112) );
  INV_X1 U7115 ( .A(n6105), .ZN(n6106) );
  INV_X1 U7116 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U7117 ( .A1(n6106), .A2(n8959), .ZN(n6107) );
  NAND2_X1 U7118 ( .A1(n6117), .A2(n6107), .ZN(n10861) );
  OR2_X1 U7119 ( .A1(n6317), .A2(n10861), .ZN(n6111) );
  INV_X1 U7120 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7617) );
  OR2_X1 U7121 ( .A1(n6357), .A2(n7617), .ZN(n6110) );
  INV_X1 U7122 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6108) );
  OR2_X1 U7123 ( .A1(n6034), .A2(n6108), .ZN(n6109) );
  NAND4_X1 U7124 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n9390)
         );
  NAND2_X1 U7125 ( .A1(n9390), .A2(n6274), .ZN(n6114) );
  XNOR2_X1 U7126 ( .A(n10852), .B(n6031), .ZN(n6113) );
  XOR2_X1 U7127 ( .A(n6114), .B(n6113), .Z(n8260) );
  INV_X1 U7128 ( .A(n6113), .ZN(n6116) );
  INV_X1 U7129 ( .A(n6114), .ZN(n6115) );
  XNOR2_X1 U7130 ( .A(n8564), .B(n6254), .ZN(n6124) );
  NAND2_X1 U7131 ( .A1(n6352), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6122) );
  INV_X1 U7132 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7615) );
  OR2_X1 U7133 ( .A1(n6284), .A2(n7615), .ZN(n6121) );
  NAND2_X1 U7134 ( .A1(n6117), .A2(n8938), .ZN(n6118) );
  NAND2_X1 U7135 ( .A1(n6127), .A2(n6118), .ZN(n8508) );
  OR2_X1 U7136 ( .A1(n6317), .A2(n8508), .ZN(n6120) );
  INV_X1 U7137 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8509) );
  OR2_X1 U7138 ( .A1(n6034), .A2(n8509), .ZN(n6119) );
  NAND4_X1 U7139 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n9389)
         );
  AND2_X1 U7140 ( .A1(n9389), .A2(n6274), .ZN(n6123) );
  NOR2_X1 U7141 ( .A1(n6124), .A2(n6123), .ZN(n6125) );
  AOI21_X1 U7142 ( .B1(n6124), .B2(n6123), .A(n6125), .ZN(n8437) );
  INV_X1 U7143 ( .A(n6125), .ZN(n6126) );
  NAND2_X1 U7144 ( .A1(n8435), .A2(n6126), .ZN(n8526) );
  XNOR2_X1 U7145 ( .A(n8605), .B(n6254), .ZN(n6134) );
  NAND2_X1 U7146 ( .A1(n6179), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6132) );
  INV_X1 U7147 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8570) );
  OR2_X1 U7148 ( .A1(n6034), .A2(n8570), .ZN(n6131) );
  NAND2_X1 U7149 ( .A1(n6127), .A2(n8954), .ZN(n6128) );
  NAND2_X1 U7150 ( .A1(n6138), .A2(n6128), .ZN(n8569) );
  OR2_X1 U7151 ( .A1(n6317), .A2(n8569), .ZN(n6130) );
  INV_X1 U7152 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7614) );
  OR2_X1 U7153 ( .A1(n6357), .A2(n7614), .ZN(n6129) );
  NAND4_X1 U7154 ( .A1(n6132), .A2(n6131), .A3(n6130), .A4(n6129), .ZN(n9388)
         );
  AND2_X1 U7155 ( .A1(n9388), .A2(n6274), .ZN(n6133) );
  NOR2_X1 U7156 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  AOI21_X1 U7157 ( .B1(n6134), .B2(n6133), .A(n6135), .ZN(n8527) );
  NAND2_X1 U7158 ( .A1(n8526), .A2(n8527), .ZN(n8525) );
  INV_X1 U7159 ( .A(n6135), .ZN(n6136) );
  XNOR2_X1 U7160 ( .A(n8656), .B(n6254), .ZN(n6145) );
  NAND2_X1 U7161 ( .A1(n6352), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6143) );
  INV_X1 U7162 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8612) );
  OR2_X1 U7163 ( .A1(n6034), .A2(n8612), .ZN(n6142) );
  INV_X1 U7164 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9131) );
  NAND2_X1 U7165 ( .A1(n6138), .A2(n9131), .ZN(n6139) );
  NAND2_X1 U7166 ( .A1(n6148), .A2(n6139), .ZN(n8611) );
  OR2_X1 U7167 ( .A1(n6317), .A2(n8611), .ZN(n6141) );
  INV_X1 U7168 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7714) );
  OR2_X1 U7169 ( .A1(n6357), .A2(n7714), .ZN(n6140) );
  NAND4_X1 U7170 ( .A1(n6143), .A2(n6142), .A3(n6141), .A4(n6140), .ZN(n9387)
         );
  AND2_X1 U7171 ( .A1(n9387), .A2(n6274), .ZN(n6144) );
  NOR2_X1 U7172 ( .A1(n6145), .A2(n6144), .ZN(n6146) );
  AOI21_X1 U7173 ( .B1(n6145), .B2(n6144), .A(n6146), .ZN(n8586) );
  XNOR2_X1 U7174 ( .A(n9744), .B(n6254), .ZN(n6155) );
  NAND2_X1 U7175 ( .A1(n6352), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6153) );
  INV_X1 U7176 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8653) );
  OR2_X1 U7177 ( .A1(n6034), .A2(n8653), .ZN(n6152) );
  INV_X1 U7178 ( .A(n6148), .ZN(n6147) );
  INV_X1 U7179 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U7180 ( .A1(n6148), .A2(n9179), .ZN(n6149) );
  NAND2_X1 U7181 ( .A1(n6159), .A2(n6149), .ZN(n8652) );
  OR2_X1 U7182 ( .A1(n6317), .A2(n8652), .ZN(n6151) );
  INV_X1 U7183 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7973) );
  OR2_X1 U7184 ( .A1(n6284), .A2(n7973), .ZN(n6150) );
  NAND4_X1 U7185 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n9386)
         );
  AND2_X1 U7186 ( .A1(n9386), .A2(n6274), .ZN(n6154) );
  NOR2_X1 U7187 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  AOI21_X1 U7188 ( .B1(n6155), .B2(n6154), .A(n6156), .ZN(n8640) );
  INV_X1 U7189 ( .A(n6156), .ZN(n6157) );
  NAND2_X1 U7190 ( .A1(n8638), .A2(n6157), .ZN(n8694) );
  XNOR2_X1 U7191 ( .A(n9656), .B(n6254), .ZN(n6168) );
  NAND2_X1 U7192 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  NAND2_X1 U7193 ( .A1(n6171), .A2(n6160), .ZN(n9652) );
  INV_X1 U7194 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8363) );
  OR2_X1 U7195 ( .A1(n6357), .A2(n8363), .ZN(n6161) );
  OAI21_X1 U7196 ( .B1(n9652), .B2(n6317), .A(n6161), .ZN(n6166) );
  INV_X1 U7197 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9653) );
  INV_X1 U7198 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6162) );
  OR2_X1 U7199 ( .A1(n6163), .A2(n6162), .ZN(n6164) );
  OAI21_X1 U7200 ( .B1(n6034), .B2(n9653), .A(n6164), .ZN(n6165) );
  AND2_X1 U7201 ( .A1(n9618), .A2(n6274), .ZN(n6167) );
  NOR2_X1 U7202 ( .A1(n6168), .A2(n6167), .ZN(n6169) );
  AOI21_X1 U7203 ( .B1(n6168), .B2(n6167), .A(n6169), .ZN(n8695) );
  INV_X1 U7204 ( .A(n6169), .ZN(n6170) );
  XNOR2_X1 U7205 ( .A(n9627), .B(n6031), .ZN(n6176) );
  INV_X1 U7206 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9735) );
  INV_X1 U7207 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9155) );
  NAND2_X1 U7208 ( .A1(n6171), .A2(n9155), .ZN(n6172) );
  NAND2_X1 U7209 ( .A1(n6177), .A2(n6172), .ZN(n9629) );
  OR2_X1 U7210 ( .A1(n9629), .A2(n6317), .ZN(n6174) );
  AOI22_X1 U7211 ( .A1(n6311), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n6179), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n6173) );
  OAI211_X1 U7212 ( .C1(n6284), .C2(n9735), .A(n6174), .B(n6173), .ZN(n9639)
         );
  NAND2_X1 U7213 ( .A1(n9639), .A2(n6274), .ZN(n6175) );
  XNOR2_X1 U7214 ( .A(n6176), .B(n6175), .ZN(n9325) );
  NAND2_X1 U7215 ( .A1(n6177), .A2(n9174), .ZN(n6178) );
  NAND2_X1 U7216 ( .A1(n6187), .A2(n6178), .ZN(n9606) );
  AOI22_X1 U7217 ( .A1(n6311), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n6179), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7218 ( .A1(n6017), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6180) );
  OAI211_X1 U7219 ( .C1(n9606), .C2(n6317), .A(n6181), .B(n6180), .ZN(n9620)
         );
  NAND2_X1 U7220 ( .A1(n9620), .A2(n6274), .ZN(n6183) );
  XNOR2_X1 U7221 ( .A(n9727), .B(n6031), .ZN(n6182) );
  XOR2_X1 U7222 ( .A(n6183), .B(n6182), .Z(n9359) );
  INV_X1 U7223 ( .A(n6182), .ZN(n6185) );
  INV_X1 U7224 ( .A(n6183), .ZN(n6184) );
  XNOR2_X1 U7225 ( .A(n9588), .B(n6254), .ZN(n6196) );
  INV_X1 U7226 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U7227 ( .A1(n6187), .A2(n9140), .ZN(n6188) );
  NAND2_X1 U7228 ( .A1(n6199), .A2(n6188), .ZN(n9597) );
  OR2_X1 U7229 ( .A1(n9597), .A2(n6317), .ZN(n6194) );
  INV_X1 U7230 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7231 ( .A1(n6017), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7232 ( .A1(n6352), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6189) );
  OAI211_X1 U7233 ( .C1(n6034), .C2(n6191), .A(n6190), .B(n6189), .ZN(n6192)
         );
  INV_X1 U7234 ( .A(n6192), .ZN(n6193) );
  NAND2_X1 U7235 ( .A1(n6194), .A2(n6193), .ZN(n9604) );
  AND2_X1 U7236 ( .A1(n9604), .A2(n6274), .ZN(n6195) );
  NOR2_X1 U7237 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  AOI21_X1 U7238 ( .B1(n6196), .B2(n6195), .A(n6197), .ZN(n9300) );
  NAND2_X1 U7239 ( .A1(n9301), .A2(n9300), .ZN(n9299) );
  INV_X1 U7240 ( .A(n6197), .ZN(n6198) );
  XNOR2_X1 U7241 ( .A(n9716), .B(n6031), .ZN(n6208) );
  NAND2_X1 U7242 ( .A1(n6199), .A2(n9343), .ZN(n6200) );
  AND2_X1 U7243 ( .A1(n6220), .A2(n6200), .ZN(n9574) );
  NAND2_X1 U7244 ( .A1(n9574), .A2(n6298), .ZN(n6206) );
  INV_X1 U7245 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7246 ( .A1(n6352), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7247 ( .A1(n6311), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6201) );
  OAI211_X1 U7248 ( .C1(n6357), .C2(n6203), .A(n6202), .B(n6201), .ZN(n6204)
         );
  INV_X1 U7249 ( .A(n6204), .ZN(n6205) );
  NAND2_X1 U7250 ( .A1(n6206), .A2(n6205), .ZN(n9591) );
  NAND2_X1 U7251 ( .A1(n9591), .A2(n6274), .ZN(n6207) );
  XNOR2_X1 U7252 ( .A(n6208), .B(n6207), .ZN(n9341) );
  XNOR2_X1 U7253 ( .A(n6220), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U7254 ( .A1(n9566), .A2(n6298), .ZN(n6213) );
  INV_X1 U7255 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9714) );
  NAND2_X1 U7256 ( .A1(n6311), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7257 ( .A1(n6352), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6209) );
  OAI211_X1 U7258 ( .C1(n9714), .C2(n6284), .A(n6210), .B(n6209), .ZN(n6211)
         );
  INV_X1 U7259 ( .A(n6211), .ZN(n6212) );
  NAND2_X1 U7260 ( .A1(n6213), .A2(n6212), .ZN(n9579) );
  NAND2_X1 U7261 ( .A1(n9579), .A2(n6274), .ZN(n6215) );
  XNOR2_X1 U7262 ( .A(n9557), .B(n6031), .ZN(n6214) );
  XOR2_X1 U7263 ( .A(n6215), .B(n6214), .Z(n9306) );
  INV_X1 U7264 ( .A(n6214), .ZN(n6217) );
  INV_X1 U7265 ( .A(n6215), .ZN(n6216) );
  XNOR2_X1 U7266 ( .A(n9705), .B(n6254), .ZN(n6229) );
  AND2_X1 U7267 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n6218) );
  INV_X1 U7268 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9308) );
  INV_X1 U7269 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9165) );
  OAI21_X1 U7270 ( .B1(n6220), .B2(n9308), .A(n9165), .ZN(n6221) );
  NAND2_X1 U7271 ( .A1(n6232), .A2(n6221), .ZN(n9541) );
  OR2_X1 U7272 ( .A1(n9541), .A2(n6317), .ZN(n6227) );
  INV_X1 U7273 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7274 ( .A1(n6311), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7275 ( .A1(n6352), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6222) );
  OAI211_X1 U7276 ( .C1(n6224), .C2(n6357), .A(n6223), .B(n6222), .ZN(n6225)
         );
  INV_X1 U7277 ( .A(n6225), .ZN(n6226) );
  NAND2_X1 U7278 ( .A1(n6227), .A2(n6226), .ZN(n9531) );
  AND2_X1 U7279 ( .A1(n9531), .A2(n6274), .ZN(n6228) );
  NOR2_X1 U7280 ( .A1(n6229), .A2(n6228), .ZN(n6230) );
  AOI21_X1 U7281 ( .B1(n6229), .B2(n6228), .A(n6230), .ZN(n9350) );
  XNOR2_X1 U7282 ( .A(n9700), .B(n6031), .ZN(n6240) );
  INV_X1 U7283 ( .A(n6232), .ZN(n6231) );
  INV_X1 U7284 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U7285 ( .A1(n6232), .A2(n9293), .ZN(n6233) );
  INV_X1 U7286 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7287 ( .A1(n6352), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U7288 ( .A1(n6311), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6234) );
  OAI211_X1 U7289 ( .C1(n6236), .C2(n6357), .A(n6235), .B(n6234), .ZN(n6237)
         );
  INV_X1 U7290 ( .A(n6237), .ZN(n6238) );
  NAND2_X1 U7291 ( .A1(n6239), .A2(n6238), .ZN(n9512) );
  NAND2_X1 U7292 ( .A1(n9512), .A2(n6274), .ZN(n9291) );
  XNOR2_X1 U7293 ( .A(n9695), .B(n6031), .ZN(n6250) );
  XNOR2_X1 U7294 ( .A(n6252), .B(n6250), .ZN(n9332) );
  INV_X1 U7295 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U7296 ( .A1(n6242), .A2(n9157), .ZN(n6243) );
  NAND2_X1 U7297 ( .A1(n6255), .A2(n6243), .ZN(n9507) );
  OR2_X1 U7298 ( .A1(n9507), .A2(n6317), .ZN(n6249) );
  INV_X1 U7299 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7300 ( .A1(n6352), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7301 ( .A1(n6311), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6244) );
  OAI211_X1 U7302 ( .C1(n6246), .C2(n6284), .A(n6245), .B(n6244), .ZN(n6247)
         );
  INV_X1 U7303 ( .A(n6247), .ZN(n6248) );
  NOR2_X1 U7304 ( .A1(n9294), .A2(n6299), .ZN(n9333) );
  INV_X1 U7305 ( .A(n6250), .ZN(n6251) );
  AND2_X1 U7306 ( .A1(n6252), .A2(n6251), .ZN(n6253) );
  XNOR2_X1 U7307 ( .A(n9498), .B(n6254), .ZN(n6263) );
  INV_X1 U7308 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U7309 ( .A1(n6255), .A2(n9320), .ZN(n6256) );
  AND2_X1 U7310 ( .A1(n6267), .A2(n6256), .ZN(n9499) );
  NAND2_X1 U7311 ( .A1(n9499), .A2(n6298), .ZN(n6261) );
  INV_X1 U7312 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9693) );
  NAND2_X1 U7313 ( .A1(n6311), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7314 ( .A1(n6352), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6257) );
  OAI211_X1 U7315 ( .C1(n9693), .C2(n6357), .A(n6258), .B(n6257), .ZN(n6259)
         );
  INV_X1 U7316 ( .A(n6259), .ZN(n6260) );
  NAND2_X1 U7317 ( .A1(n6261), .A2(n6260), .ZN(n9513) );
  AND2_X1 U7318 ( .A1(n9513), .A2(n6274), .ZN(n6262) );
  NOR2_X1 U7319 ( .A1(n6263), .A2(n6262), .ZN(n6264) );
  AOI21_X1 U7320 ( .B1(n6263), .B2(n6262), .A(n6264), .ZN(n9315) );
  INV_X1 U7321 ( .A(n6264), .ZN(n6265) );
  XNOR2_X1 U7322 ( .A(n9684), .B(n6031), .ZN(n6275) );
  INV_X1 U7323 ( .A(n6267), .ZN(n6266) );
  NAND2_X1 U7324 ( .A1(n6266), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6280) );
  INV_X1 U7325 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8967) );
  NAND2_X1 U7326 ( .A1(n6267), .A2(n8967), .ZN(n6268) );
  NAND2_X1 U7327 ( .A1(n6280), .A2(n6268), .ZN(n9481) );
  OR2_X1 U7328 ( .A1(n9481), .A2(n6317), .ZN(n6273) );
  INV_X1 U7329 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U7330 ( .A1(n6311), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7331 ( .A1(n6352), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6269) );
  OAI211_X1 U7332 ( .C1(n9688), .C2(n6357), .A(n6270), .B(n6269), .ZN(n6271)
         );
  INV_X1 U7333 ( .A(n6271), .ZN(n6272) );
  NAND2_X1 U7334 ( .A1(n6273), .A2(n6272), .ZN(n9384) );
  NAND2_X1 U7335 ( .A1(n9384), .A2(n6274), .ZN(n6276) );
  XOR2_X1 U7336 ( .A(n6275), .B(n6276), .Z(n9370) );
  INV_X1 U7337 ( .A(n6275), .ZN(n6278) );
  INV_X1 U7338 ( .A(n6276), .ZN(n6277) );
  XNOR2_X1 U7339 ( .A(n9679), .B(n5016), .ZN(n6290) );
  INV_X1 U7340 ( .A(n6280), .ZN(n6279) );
  NAND2_X1 U7341 ( .A1(n6279), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6292) );
  INV_X1 U7342 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U7343 ( .A1(n6280), .A2(n8923), .ZN(n6281) );
  NAND2_X1 U7344 ( .A1(n6292), .A2(n6281), .ZN(n9455) );
  OR2_X1 U7345 ( .A1(n9455), .A2(n6317), .ZN(n6288) );
  INV_X1 U7346 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7347 ( .A1(n6311), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7348 ( .A1(n6352), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6282) );
  OAI211_X1 U7349 ( .C1(n6285), .C2(n6284), .A(n6283), .B(n6282), .ZN(n6286)
         );
  INV_X1 U7350 ( .A(n6286), .ZN(n6287) );
  NAND2_X1 U7351 ( .A1(n9444), .A2(n6274), .ZN(n6289) );
  NOR2_X1 U7352 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  AOI21_X1 U7353 ( .B1(n6290), .B2(n6289), .A(n6291), .ZN(n8858) );
  INV_X1 U7354 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U7355 ( .A1(n6292), .A2(n8934), .ZN(n6293) );
  INV_X1 U7356 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7357 ( .A1(n6311), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7358 ( .A1(n6352), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6294) );
  OAI211_X1 U7359 ( .C1(n6296), .C2(n6357), .A(n6295), .B(n6294), .ZN(n6297)
         );
  AOI21_X1 U7360 ( .B1(n9438), .B2(n6298), .A(n6297), .ZN(n8862) );
  NOR2_X1 U7361 ( .A1(n8862), .A2(n6299), .ZN(n6300) );
  MUX2_X1 U7362 ( .A(n8862), .B(n6300), .S(n6031), .Z(n6301) );
  NAND2_X1 U7363 ( .A1(n6303), .A2(n6302), .ZN(n8036) );
  AND2_X1 U7364 ( .A1(n10914), .A2(n7470), .ZN(n6304) );
  NAND2_X1 U7365 ( .A1(n10552), .A2(n6304), .ZN(n6305) );
  OR2_X1 U7366 ( .A1(n6306), .A2(n9381), .ZN(n6328) );
  NAND2_X1 U7367 ( .A1(n6306), .A2(n9352), .ZN(n6309) );
  NAND2_X1 U7368 ( .A1(n6319), .A2(n6307), .ZN(n7382) );
  AND2_X1 U7369 ( .A1(n10552), .A2(n9745), .ZN(n6308) );
  NAND2_X1 U7370 ( .A1(n6309), .A2(n9358), .ZN(n6310) );
  NAND2_X1 U7371 ( .A1(n6310), .A2(n9674), .ZN(n6327) );
  INV_X1 U7372 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U7373 ( .A1(n6311), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U7374 ( .A1(n6352), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6312) );
  OAI211_X1 U7375 ( .C1(n6314), .C2(n6357), .A(n6313), .B(n6312), .ZN(n6315)
         );
  INV_X1 U7376 ( .A(n6315), .ZN(n6316) );
  OAI21_X1 U7377 ( .B1(n8811), .B2(n6317), .A(n6316), .ZN(n9445) );
  NAND2_X1 U7378 ( .A1(n10552), .A2(n6318), .ZN(n6530) );
  NAND2_X1 U7379 ( .A1(n9445), .A2(n9334), .ZN(n6326) );
  INV_X1 U7380 ( .A(n5940), .ZN(n6320) );
  NAND2_X1 U7381 ( .A1(n9444), .A2(n9335), .ZN(n6325) );
  INV_X1 U7382 ( .A(n6529), .ZN(n7138) );
  AND3_X1 U7383 ( .A1(n7137), .A2(n7138), .A3(n6321), .ZN(n6322) );
  NAND2_X1 U7384 ( .A1(n7382), .A2(n6322), .ZN(n6323) );
  AOI22_X1 U7385 ( .A1(n9438), .A2(n9374), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6324) );
  OAI211_X1 U7386 ( .C1(n6328), .C2(n9674), .A(n6327), .B(n5605), .ZN(P2_U3222) );
  NAND2_X1 U7387 ( .A1(n7755), .A2(n10701), .ZN(n8034) );
  NAND2_X1 U7388 ( .A1(n6505), .A2(n7756), .ZN(n6377) );
  INV_X1 U7389 ( .A(n8061), .ZN(n10716) );
  OR2_X1 U7390 ( .A1(n9397), .A2(n10716), .ZN(n6383) );
  NAND2_X1 U7391 ( .A1(n6377), .A2(n6383), .ZN(n6330) );
  NAND2_X1 U7392 ( .A1(n9397), .A2(n10716), .ZN(n6382) );
  NAND2_X1 U7393 ( .A1(n9396), .A2(n8356), .ZN(n6387) );
  NAND2_X2 U7394 ( .A1(n6388), .A2(n6387), .ZN(n7765) );
  NAND2_X1 U7395 ( .A1(n9395), .A2(n10731), .ZN(n6331) );
  OR2_X1 U7396 ( .A1(n10731), .A2(n9395), .ZN(n6332) );
  INV_X1 U7397 ( .A(n7954), .ZN(n7918) );
  INV_X1 U7398 ( .A(n10753), .ZN(n8339) );
  NAND2_X1 U7399 ( .A1(n8339), .A2(n8455), .ZN(n6333) );
  NAND2_X1 U7400 ( .A1(n7920), .A2(n6333), .ZN(n8454) );
  INV_X1 U7401 ( .A(n9394), .ZN(n7874) );
  OR2_X1 U7402 ( .A1(n8450), .A2(n7874), .ZN(n6397) );
  NAND2_X1 U7403 ( .A1(n8450), .A2(n7874), .ZN(n6403) );
  NAND2_X1 U7404 ( .A1(n6397), .A2(n6403), .ZN(n7957) );
  INV_X1 U7405 ( .A(n7957), .ZN(n8453) );
  NAND2_X1 U7406 ( .A1(n8454), .A2(n8453), .ZN(n8452) );
  NAND2_X1 U7407 ( .A1(n8452), .A2(n6397), .ZN(n7960) );
  INV_X1 U7408 ( .A(n9393), .ZN(n7886) );
  OR2_X1 U7409 ( .A1(n8463), .A2(n7886), .ZN(n6402) );
  NAND2_X1 U7410 ( .A1(n8463), .A2(n7886), .ZN(n6398) );
  INV_X1 U7411 ( .A(n9392), .ZN(n8285) );
  OR2_X1 U7412 ( .A1(n8281), .A2(n8285), .ZN(n6407) );
  NAND2_X1 U7413 ( .A1(n8281), .A2(n8285), .ZN(n6408) );
  INV_X1 U7414 ( .A(n8394), .ZN(n8172) );
  OR2_X1 U7415 ( .A1(n8385), .A2(n8172), .ZN(n6411) );
  NAND2_X1 U7416 ( .A1(n8385), .A2(n8172), .ZN(n6416) );
  NAND2_X1 U7417 ( .A1(n6411), .A2(n6416), .ZN(n8289) );
  INV_X1 U7418 ( .A(n9391), .ZN(n8284) );
  OR2_X1 U7419 ( .A1(n8416), .A2(n8284), .ZN(n6418) );
  NAND2_X1 U7420 ( .A1(n6418), .A2(n6415), .ZN(n8390) );
  NAND2_X1 U7421 ( .A1(n10852), .A2(n8506), .ZN(n6504) );
  INV_X1 U7422 ( .A(n9389), .ZN(n8530) );
  OR2_X1 U7423 ( .A1(n8564), .A2(n8530), .ZN(n6425) );
  NAND2_X1 U7424 ( .A1(n8564), .A2(n8530), .ZN(n6426) );
  INV_X1 U7425 ( .A(n8563), .ZN(n6338) );
  INV_X1 U7426 ( .A(n8502), .ZN(n8422) );
  NOR2_X1 U7427 ( .A1(n6338), .A2(n8422), .ZN(n6339) );
  NAND2_X1 U7428 ( .A1(n8420), .A2(n6339), .ZN(n8501) );
  NAND2_X1 U7429 ( .A1(n8501), .A2(n6426), .ZN(n8560) );
  INV_X1 U7430 ( .A(n9388), .ZN(n8604) );
  OR2_X1 U7431 ( .A1(n8605), .A2(n8604), .ZN(n6432) );
  NAND2_X1 U7432 ( .A1(n8605), .A2(n8604), .ZN(n6431) );
  NAND2_X1 U7433 ( .A1(n8560), .A2(n8567), .ZN(n8559) );
  XNOR2_X1 U7434 ( .A(n8656), .B(n9387), .ZN(n8658) );
  INV_X1 U7435 ( .A(n8658), .ZN(n8601) );
  INV_X1 U7436 ( .A(n9387), .ZN(n8643) );
  OR2_X1 U7437 ( .A1(n8656), .A2(n8643), .ZN(n6340) );
  INV_X1 U7438 ( .A(n9386), .ZN(n9642) );
  INV_X1 U7439 ( .A(n6438), .ZN(n6341) );
  NAND2_X1 U7440 ( .A1(n9744), .A2(n9642), .ZN(n6439) );
  INV_X1 U7441 ( .A(n9618), .ZN(n9327) );
  OR2_X1 U7442 ( .A1(n9656), .A2(n9327), .ZN(n6441) );
  NAND2_X1 U7443 ( .A1(n9656), .A2(n9327), .ZN(n6442) );
  NAND2_X1 U7444 ( .A1(n9627), .A2(n9639), .ZN(n6445) );
  NAND2_X1 U7445 ( .A1(n8802), .A2(n6445), .ZN(n9623) );
  INV_X1 U7446 ( .A(n9639), .ZN(n9364) );
  OR2_X1 U7447 ( .A1(n9627), .A2(n9364), .ZN(n6342) );
  NAND2_X1 U7448 ( .A1(n6343), .A2(n6342), .ZN(n9603) );
  INV_X1 U7449 ( .A(n9620), .ZN(n9593) );
  XNOR2_X1 U7450 ( .A(n9727), .B(n9593), .ZN(n9612) );
  INV_X1 U7451 ( .A(n9612), .ZN(n6515) );
  NAND2_X1 U7452 ( .A1(n9588), .A2(n9361), .ZN(n6373) );
  INV_X1 U7453 ( .A(n9591), .ZN(n9563) );
  NAND2_X1 U7454 ( .A1(n9716), .A2(n9563), .ZN(n6454) );
  NAND2_X1 U7455 ( .A1(n6453), .A2(n6454), .ZN(n9577) );
  INV_X1 U7456 ( .A(n9577), .ZN(n6344) );
  INV_X1 U7457 ( .A(n9579), .ZN(n9547) );
  NAND2_X1 U7458 ( .A1(n9557), .A2(n9547), .ZN(n6345) );
  NAND2_X1 U7459 ( .A1(n6346), .A2(n6345), .ZN(n9546) );
  NAND2_X1 U7460 ( .A1(n9705), .A2(n9564), .ZN(n6369) );
  INV_X1 U7461 ( .A(n9536), .ZN(n9545) );
  OR2_X1 U7462 ( .A1(n9700), .A2(n9548), .ZN(n6463) );
  NAND2_X1 U7463 ( .A1(n6463), .A2(n6467), .ZN(n9520) );
  INV_X1 U7464 ( .A(n9520), .ZN(n9529) );
  NAND2_X1 U7465 ( .A1(n9695), .A2(n9294), .ZN(n6468) );
  NAND2_X1 U7466 ( .A1(n9510), .A2(n6469), .ZN(n9491) );
  INV_X1 U7467 ( .A(n9513), .ZN(n6347) );
  NAND2_X1 U7468 ( .A1(n9498), .A2(n6347), .ZN(n6472) );
  NAND2_X1 U7469 ( .A1(n9474), .A2(n6472), .ZN(n9488) );
  NAND2_X1 U7470 ( .A1(n9491), .A2(n9492), .ZN(n9490) );
  INV_X1 U7471 ( .A(n9384), .ZN(n9459) );
  OR2_X1 U7472 ( .A1(n9684), .A2(n9459), .ZN(n6479) );
  NAND2_X1 U7473 ( .A1(n9684), .A2(n9459), .ZN(n9461) );
  NAND2_X1 U7474 ( .A1(n6479), .A2(n9461), .ZN(n9477) );
  INV_X1 U7475 ( .A(n9474), .ZN(n6348) );
  NOR2_X1 U7476 ( .A1(n9477), .A2(n6348), .ZN(n6349) );
  NAND2_X1 U7477 ( .A1(n9490), .A2(n6349), .ZN(n9460) );
  INV_X1 U7478 ( .A(n9444), .ZN(n8807) );
  NAND2_X1 U7479 ( .A1(n9679), .A2(n8807), .ZN(n6482) );
  NAND2_X1 U7480 ( .A1(n6483), .A2(n6482), .ZN(n9465) );
  INV_X1 U7481 ( .A(n9461), .ZN(n6480) );
  NOR2_X1 U7482 ( .A1(n9465), .A2(n6480), .ZN(n6350) );
  NAND2_X1 U7483 ( .A1(n9460), .A2(n6350), .ZN(n9462) );
  NAND2_X1 U7484 ( .A1(n9462), .A2(n6483), .ZN(n9443) );
  NAND2_X1 U7485 ( .A1(n9674), .A2(n8862), .ZN(n6484) );
  NAND2_X1 U7486 ( .A1(n6485), .A2(n6484), .ZN(n8809) );
  INV_X1 U7487 ( .A(n9445), .ZN(n6351) );
  NAND2_X1 U7488 ( .A1(n9668), .A2(n6351), .ZN(n6486) );
  INV_X1 U7489 ( .A(n6367), .ZN(n6476) );
  INV_X1 U7490 ( .A(n6358), .ZN(n6360) );
  INV_X1 U7491 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U7492 ( .A1(n6352), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6355) );
  INV_X1 U7493 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6353) );
  OR2_X1 U7494 ( .A1(n6034), .A2(n6353), .ZN(n6354) );
  OAI211_X1 U7495 ( .C1(n6357), .C2(n6356), .A(n6355), .B(n6354), .ZN(n9383)
         );
  INV_X1 U7496 ( .A(n9383), .ZN(n6361) );
  OR2_X1 U7497 ( .A1(n6362), .A2(n6361), .ZN(n6494) );
  OR2_X1 U7498 ( .A1(n6363), .A2(n7287), .ZN(n6497) );
  NAND2_X1 U7499 ( .A1(n6362), .A2(n6361), .ZN(n6496) );
  NAND2_X1 U7500 ( .A1(n6497), .A2(n6496), .ZN(n6522) );
  NAND2_X1 U7501 ( .A1(n6363), .A2(n7287), .ZN(n6495) );
  XNOR2_X1 U7502 ( .A(n6366), .B(n9407), .ZN(n6365) );
  OAI22_X1 U7503 ( .A1(n6274), .A2(n6366), .B1(n6365), .B2(n7767), .ZN(n6528)
         );
  INV_X1 U7504 ( .A(n6484), .ZN(n6368) );
  NOR2_X1 U7505 ( .A1(n8815), .A2(n6368), .ZN(n6478) );
  NAND2_X1 U7506 ( .A1(n6453), .A2(n6372), .ZN(n6375) );
  NAND2_X1 U7507 ( .A1(n6454), .A2(n6373), .ZN(n6374) );
  MUX2_X1 U7508 ( .A(n6375), .B(n6374), .S(n6499), .Z(n6456) );
  INV_X1 U7509 ( .A(n7756), .ZN(n6376) );
  OR2_X1 U7510 ( .A1(n6505), .A2(n6376), .ZN(n7863) );
  NOR2_X1 U7511 ( .A1(n7755), .A2(n10701), .ZN(n7414) );
  OAI21_X1 U7512 ( .B1(n7863), .B2(n7414), .A(n8051), .ZN(n6380) );
  INV_X1 U7513 ( .A(n7414), .ZN(n8035) );
  AND2_X1 U7514 ( .A1(n8035), .A2(n7760), .ZN(n6378) );
  OAI21_X1 U7515 ( .B1(n6378), .B2(n6505), .A(n7756), .ZN(n6379) );
  MUX2_X1 U7516 ( .A(n6380), .B(n6379), .S(n6499), .Z(n6381) );
  INV_X1 U7517 ( .A(n8052), .ZN(n8050) );
  NAND2_X1 U7518 ( .A1(n6381), .A2(n8050), .ZN(n6386) );
  NOR2_X1 U7519 ( .A1(n6384), .A2(n7765), .ZN(n6385) );
  NAND2_X1 U7520 ( .A1(n6386), .A2(n6385), .ZN(n6390) );
  MUX2_X1 U7521 ( .A(n6388), .B(n6387), .S(n6464), .Z(n6389) );
  NAND2_X1 U7522 ( .A1(n6390), .A2(n6389), .ZN(n6392) );
  INV_X1 U7523 ( .A(n10731), .ZN(n8218) );
  NAND2_X1 U7524 ( .A1(n9395), .A2(n8218), .ZN(n7915) );
  OR2_X1 U7525 ( .A1(n8218), .A2(n9395), .ZN(n6508) );
  INV_X1 U7526 ( .A(n9395), .ZN(n7791) );
  MUX2_X1 U7527 ( .A(n10731), .B(n7791), .S(n6499), .Z(n6391) );
  AND2_X1 U7528 ( .A1(n10753), .A2(n6499), .ZN(n6394) );
  NOR2_X1 U7529 ( .A1(n10753), .A2(n6499), .ZN(n6393) );
  MUX2_X1 U7530 ( .A(n6394), .B(n6393), .S(n8455), .Z(n6395) );
  NOR2_X1 U7531 ( .A1(n7957), .A2(n6395), .ZN(n6396) );
  AND2_X1 U7532 ( .A1(n8078), .A2(n6397), .ZN(n6400) );
  INV_X1 U7533 ( .A(n6398), .ZN(n6399) );
  AOI21_X1 U7534 ( .B1(n6404), .B2(n6400), .A(n6399), .ZN(n6401) );
  MUX2_X1 U7535 ( .A(n6402), .B(n6401), .S(n6499), .Z(n6406) );
  NAND4_X1 U7536 ( .A1(n6404), .A2(n6464), .A3(n8078), .A4(n6403), .ZN(n6405)
         );
  NAND3_X1 U7537 ( .A1(n6406), .A2(n8080), .A3(n6405), .ZN(n6410) );
  MUX2_X1 U7538 ( .A(n6408), .B(n6407), .S(n6499), .Z(n6409) );
  NAND3_X1 U7539 ( .A1(n6410), .A2(n6411), .A3(n6409), .ZN(n6413) );
  AND2_X1 U7540 ( .A1(n6412), .A2(n6418), .ZN(n6414) );
  NAND2_X1 U7541 ( .A1(n6413), .A2(n6414), .ZN(n6423) );
  INV_X1 U7542 ( .A(n6414), .ZN(n6417) );
  OAI211_X1 U7543 ( .C1(n6417), .C2(n6416), .A(n6415), .B(n6504), .ZN(n6420)
         );
  NAND2_X1 U7544 ( .A1(n8502), .A2(n6418), .ZN(n6419) );
  MUX2_X1 U7545 ( .A(n6420), .B(n6419), .S(n6499), .Z(n6421) );
  INV_X1 U7546 ( .A(n6421), .ZN(n6422) );
  NAND2_X1 U7547 ( .A1(n6426), .A2(n6504), .ZN(n6424) );
  NAND2_X1 U7548 ( .A1(n6424), .A2(n6425), .ZN(n6429) );
  NAND2_X1 U7549 ( .A1(n6425), .A2(n8502), .ZN(n6427) );
  NAND2_X1 U7550 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  MUX2_X1 U7551 ( .A(n6429), .B(n6428), .S(n6464), .Z(n6430) );
  MUX2_X1 U7552 ( .A(n6432), .B(n6431), .S(n6464), .Z(n6433) );
  NAND2_X1 U7553 ( .A1(n6438), .A2(n6439), .ZN(n8660) );
  INV_X1 U7554 ( .A(n8660), .ZN(n6437) );
  NAND2_X1 U7555 ( .A1(n9387), .A2(n6464), .ZN(n6435) );
  OR2_X1 U7556 ( .A1(n9387), .A2(n6464), .ZN(n6434) );
  MUX2_X1 U7557 ( .A(n6435), .B(n6434), .S(n8656), .Z(n6436) );
  MUX2_X1 U7558 ( .A(n6439), .B(n6438), .S(n6499), .Z(n6440) );
  MUX2_X1 U7559 ( .A(n6442), .B(n6441), .S(n6464), .Z(n6443) );
  INV_X1 U7560 ( .A(n6446), .ZN(n6448) );
  MUX2_X1 U7561 ( .A(n9639), .B(n9627), .S(n6499), .Z(n6444) );
  OAI21_X1 U7562 ( .B1(n6446), .B2(n6445), .A(n6444), .ZN(n6447) );
  OAI21_X1 U7563 ( .B1(n6448), .B2(n8802), .A(n6447), .ZN(n6452) );
  AND2_X1 U7564 ( .A1(n9620), .A2(n6464), .ZN(n6450) );
  NOR2_X1 U7565 ( .A1(n9620), .A2(n6464), .ZN(n6449) );
  MUX2_X1 U7566 ( .A(n6450), .B(n6449), .S(n9727), .Z(n6451) );
  INV_X1 U7567 ( .A(n9584), .ZN(n9589) );
  MUX2_X1 U7568 ( .A(n6454), .B(n6453), .S(n6499), .Z(n6455) );
  NAND2_X1 U7569 ( .A1(n9557), .A2(n9579), .ZN(n6502) );
  MUX2_X1 U7570 ( .A(n9579), .B(n9557), .S(n6464), .Z(n6457) );
  OAI21_X1 U7571 ( .B1(n6458), .B2(n6502), .A(n6457), .ZN(n6460) );
  OR2_X1 U7572 ( .A1(n9557), .A2(n9579), .ZN(n6503) );
  INV_X1 U7573 ( .A(n6503), .ZN(n8804) );
  NAND2_X1 U7574 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  NAND2_X1 U7575 ( .A1(n6469), .A2(n6463), .ZN(n6465) );
  NAND2_X1 U7576 ( .A1(n6466), .A2(n9474), .ZN(n6473) );
  NAND2_X1 U7577 ( .A1(n6468), .A2(n6467), .ZN(n6470) );
  INV_X1 U7578 ( .A(n6479), .ZN(n6474) );
  NAND3_X1 U7579 ( .A1(n6475), .A2(n6483), .A3(n6485), .ZN(n6477) );
  AOI21_X1 U7580 ( .B1(n6478), .B2(n6477), .A(n6476), .ZN(n6491) );
  NOR2_X1 U7581 ( .A1(n8815), .A2(n5474), .ZN(n6488) );
  INV_X1 U7582 ( .A(n6486), .ZN(n6487) );
  AOI21_X1 U7583 ( .B1(n6489), .B2(n6488), .A(n6487), .ZN(n6490) );
  INV_X1 U7584 ( .A(n6522), .ZN(n6493) );
  INV_X1 U7585 ( .A(n6495), .ZN(n6492) );
  NAND2_X1 U7586 ( .A1(n6495), .A2(n6494), .ZN(n6521) );
  INV_X1 U7587 ( .A(n6497), .ZN(n6498) );
  OR2_X1 U7588 ( .A1(n5939), .A2(n9407), .ZN(n7766) );
  XNOR2_X1 U7589 ( .A(n6501), .B(n7766), .ZN(n6500) );
  NOR3_X1 U7590 ( .A1(n6500), .A2(n6506), .A3(n10702), .ZN(n6527) );
  INV_X1 U7591 ( .A(n6501), .ZN(n6525) );
  INV_X1 U7592 ( .A(n9646), .ZN(n9637) );
  NAND2_X1 U7593 ( .A1(n8502), .A2(n6504), .ZN(n8499) );
  INV_X1 U7594 ( .A(n8499), .ZN(n8419) );
  INV_X1 U7595 ( .A(n6505), .ZN(n6507) );
  NAND4_X1 U7596 ( .A1(n6507), .A2(n6506), .A3(n7756), .A4(n8035), .ZN(n6510)
         );
  NAND2_X1 U7597 ( .A1(n6508), .A2(n7915), .ZN(n8215) );
  INV_X1 U7598 ( .A(n8215), .ZN(n6509) );
  NOR4_X1 U7599 ( .A1(n6510), .A2(n6509), .A3(n7765), .A4(n8052), .ZN(n6511)
         );
  NAND4_X1 U7600 ( .A1(n8080), .A2(n8453), .A3(n6511), .A4(n7954), .ZN(n6512)
         );
  NOR4_X1 U7601 ( .A1(n8390), .A2(n6512), .A3(n8289), .A4(n5015), .ZN(n6513)
         );
  NAND4_X1 U7602 ( .A1(n8567), .A2(n8563), .A3(n8419), .A4(n6513), .ZN(n6514)
         );
  NOR4_X1 U7603 ( .A1(n9637), .A2(n8601), .A3(n8660), .A4(n6514), .ZN(n6516)
         );
  NAND4_X1 U7604 ( .A1(n9584), .A2(n6516), .A3(n9623), .A4(n6515), .ZN(n6517)
         );
  NOR4_X1 U7605 ( .A1(n9545), .A2(n9560), .A3(n9577), .A4(n6517), .ZN(n6518)
         );
  NAND4_X1 U7606 ( .A1(n9492), .A2(n9511), .A3(n9529), .A4(n6518), .ZN(n6519)
         );
  OR4_X1 U7607 ( .A1(n8809), .A2(n9465), .A3(n9477), .A4(n6519), .ZN(n6520) );
  NOR4_X1 U7608 ( .A1(n6522), .A2(n6521), .A3(n8815), .A4(n6520), .ZN(n6523)
         );
  XNOR2_X1 U7609 ( .A(n6523), .B(n6002), .ZN(n6524) );
  AOI211_X1 U7610 ( .C1(n6525), .C2(n6004), .A(n7760), .B(n6524), .ZN(n6526)
         );
  NOR3_X1 U7611 ( .A1(n6528), .A2(n6527), .A3(n6526), .ZN(n6534) );
  NAND2_X1 U7612 ( .A1(n6529), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8541) );
  NOR3_X1 U7613 ( .A1(n6530), .A2(n5941), .A3(n9641), .ZN(n6532) );
  OAI21_X1 U7614 ( .B1(n8541), .B2(n7761), .A(P2_B_REG_SCAN_IN), .ZN(n6531) );
  OR2_X1 U7615 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  OAI21_X1 U7616 ( .B1(n6534), .B2(n8541), .A(n6533), .ZN(P2_U3244) );
  INV_X2 U7617 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9015) );
  NOR2_X2 U7618 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6686) );
  NAND4_X1 U7619 ( .A1(n6537), .A2(n6536), .A3(n6535), .A4(n6686), .ZN(n6770)
         );
  INV_X1 U7620 ( .A(n6770), .ZN(n6543) );
  NAND4_X1 U7621 ( .A1(n6539), .A2(n6538), .A3(n9251), .A4(n6924), .ZN(n6540)
         );
  INV_X1 U7622 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6550) );
  INV_X1 U7623 ( .A(n6551), .ZN(n8836) );
  NAND2_X1 U7624 ( .A1(n6678), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7625 ( .A1(n6656), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U7626 ( .A1(n6655), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6553) );
  INV_X1 U7627 ( .A(n6557), .ZN(n6563) );
  NAND2_X1 U7628 ( .A1(n6560), .A2(n9266), .ZN(n6558) );
  XNOR2_X1 U7629 ( .A(n6560), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U7630 ( .A1(n6561), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6562) );
  MUX2_X1 U7631 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6562), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6564) );
  XNOR2_X2 U7632 ( .A(n6579), .B(n9262), .ZN(n10183) );
  NAND2_X1 U7633 ( .A1(n6565), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6566) );
  MUX2_X1 U7634 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6566), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6567) );
  NAND2_X1 U7635 ( .A1(n7836), .A2(n7058), .ZN(n6578) );
  NAND2_X1 U7636 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6572) );
  MUX2_X1 U7637 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6572), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n6574) );
  INV_X1 U7638 ( .A(n6686), .ZN(n6573) );
  NAND2_X1 U7639 ( .A1(n6574), .A2(n6573), .ZN(n7253) );
  INV_X1 U7640 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7254) );
  OR2_X1 U7641 ( .A1(n6626), .A2(n7257), .ZN(n6576) );
  NAND2_X1 U7642 ( .A1(n7654), .A2(n7030), .ZN(n6577) );
  NAND2_X1 U7643 ( .A1(n6578), .A2(n6577), .ZN(n6584) );
  NAND2_X1 U7644 ( .A1(n6579), .A2(n9262), .ZN(n6580) );
  NAND2_X1 U7645 ( .A1(n6580), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U7646 ( .A1(n6582), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6583) );
  XNOR2_X2 U7647 ( .A(n6583), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10366) );
  NAND2_X1 U7648 ( .A1(n10017), .A2(n10740), .ZN(n7124) );
  NAND2_X1 U7649 ( .A1(n8327), .A2(n10740), .ZN(n10192) );
  NAND2_X1 U7650 ( .A1(n8538), .A2(n7845), .ZN(n6585) );
  NAND2_X1 U7651 ( .A1(n7836), .A2(n6977), .ZN(n6587) );
  NAND2_X1 U7652 ( .A1(n7654), .A2(n7058), .ZN(n6586) );
  NAND2_X1 U7653 ( .A1(n6587), .A2(n6586), .ZN(n6601) );
  NAND2_X1 U7654 ( .A1(n6600), .A2(n6601), .ZN(n6599) );
  NAND2_X1 U7655 ( .A1(n6655), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6590) );
  INV_X1 U7656 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10696) );
  NAND2_X1 U7657 ( .A1(n6656), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6589) );
  NAND2_X1 U7658 ( .A1(n6678), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6588) );
  INV_X1 U7659 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10637) );
  NAND2_X1 U7660 ( .A1(n5724), .A2(SI_0_), .ZN(n6591) );
  XNOR2_X1 U7661 ( .A(n6591), .B(n5263), .ZN(n10543) );
  MUX2_X1 U7662 ( .A(n10637), .B(n10543), .S(n7140), .Z(n8799) );
  OAI22_X1 U7663 ( .A1(n8799), .A2(n6764), .B1(n7160), .B2(n10637), .ZN(n6593)
         );
  AOI21_X1 U7664 ( .B1(n7651), .B2(n6977), .A(n6593), .ZN(n7188) );
  NAND2_X1 U7665 ( .A1(n7651), .A2(n7058), .ZN(n6596) );
  INV_X1 U7666 ( .A(n8799), .ZN(n10694) );
  INV_X1 U7667 ( .A(n7160), .ZN(n6594) );
  AOI22_X1 U7668 ( .A1(n10694), .A2(n6708), .B1(n6594), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U7669 ( .A1(n6596), .A2(n6595), .ZN(n7187) );
  NAND2_X1 U7670 ( .A1(n7188), .A2(n7187), .ZN(n7186) );
  INV_X1 U7671 ( .A(n7187), .ZN(n6597) );
  NAND2_X1 U7672 ( .A1(n6597), .A2(n7652), .ZN(n6598) );
  NAND2_X1 U7673 ( .A1(n7186), .A2(n6598), .ZN(n7419) );
  NAND2_X1 U7674 ( .A1(n6599), .A2(n7419), .ZN(n6603) );
  INV_X1 U7675 ( .A(n6601), .ZN(n7418) );
  NAND2_X1 U7676 ( .A1(n7420), .A2(n7418), .ZN(n6602) );
  NAND2_X1 U7677 ( .A1(n6603), .A2(n6602), .ZN(n7445) );
  NAND2_X1 U7678 ( .A1(n6655), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U7679 ( .A1(n6678), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6607) );
  INV_X1 U7680 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7933) );
  OR2_X1 U7681 ( .A1(n7117), .A2(n7933), .ZN(n6606) );
  NAND2_X1 U7682 ( .A1(n6754), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U7683 ( .A1(n7830), .A2(n7058), .ZN(n6611) );
  INV_X1 U7684 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7250) );
  OR2_X1 U7685 ( .A1(n6686), .A2(n6806), .ZN(n6642) );
  NAND2_X1 U7686 ( .A1(n6642), .A2(n6609), .ZN(n6623) );
  OAI21_X1 U7687 ( .B1(n6642), .B2(n6609), .A(n6623), .ZN(n7252) );
  NAND2_X1 U7688 ( .A1(n10053), .A2(n7030), .ZN(n6610) );
  NAND2_X1 U7689 ( .A1(n6611), .A2(n6610), .ZN(n6612) );
  AOI21_X1 U7690 ( .B1(n7830), .B2(n6977), .A(n6613), .ZN(n6615) );
  NAND2_X1 U7691 ( .A1(n7445), .A2(n7446), .ZN(n6618) );
  INV_X1 U7692 ( .A(n6614), .ZN(n6616) );
  NAND2_X1 U7693 ( .A1(n6616), .A2(n6615), .ZN(n6617) );
  NAND2_X1 U7694 ( .A1(n6618), .A2(n6617), .ZN(n7697) );
  NAND2_X1 U7695 ( .A1(n6754), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U7696 ( .A1(n6678), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6621) );
  OR2_X1 U7697 ( .A1(n7117), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U7698 ( .A1(n6655), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U7699 ( .A1(n10210), .A2(n7058), .ZN(n6630) );
  NAND2_X1 U7700 ( .A1(n6623), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6625) );
  INV_X1 U7701 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6624) );
  XNOR2_X1 U7702 ( .A(n6625), .B(n6624), .ZN(n7373) );
  OR2_X1 U7703 ( .A1(n8823), .A2(n5107), .ZN(n6627) );
  NAND2_X1 U7704 ( .A1(n7903), .A2(n7030), .ZN(n6629) );
  NAND2_X1 U7705 ( .A1(n6630), .A2(n6629), .ZN(n6631) );
  XNOR2_X1 U7706 ( .A(n6631), .B(n7652), .ZN(n6633) );
  AND2_X1 U7707 ( .A1(n7903), .A2(n7058), .ZN(n6632) );
  AOI21_X1 U7708 ( .B1(n10210), .B2(n6977), .A(n6632), .ZN(n6634) );
  XNOR2_X1 U7709 ( .A(n6633), .B(n6634), .ZN(n7698) );
  INV_X1 U7710 ( .A(n6633), .ZN(n6635) );
  NAND2_X1 U7711 ( .A1(n6635), .A2(n6634), .ZN(n6636) );
  INV_X1 U7712 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7147) );
  OR2_X1 U7713 ( .A1(n6730), .A2(n7147), .ZN(n6640) );
  XNOR2_X1 U7714 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7891) );
  NAND2_X1 U7715 ( .A1(n6678), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U7716 ( .A1(n10209), .A2(n7058), .ZN(n6646) );
  OAI21_X1 U7717 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7718 ( .A1(n6642), .A2(n6641), .ZN(n6663) );
  XNOR2_X1 U7719 ( .A(n6663), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7643) );
  OR2_X1 U7720 ( .A1(n6626), .A2(n7259), .ZN(n6644) );
  INV_X1 U7721 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7258) );
  OR2_X1 U7722 ( .A1(n8823), .A2(n7258), .ZN(n6643) );
  OAI211_X1 U7723 ( .C1(n7643), .C2(n7140), .A(n6644), .B(n6643), .ZN(n7991)
         );
  NAND2_X1 U7724 ( .A1(n7991), .A2(n7030), .ZN(n6645) );
  NAND2_X1 U7725 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  XNOR2_X1 U7726 ( .A(n6647), .B(n8732), .ZN(n6650) );
  AND2_X1 U7727 ( .A1(n7991), .A2(n7058), .ZN(n6648) );
  AOI21_X1 U7728 ( .B1(n10209), .B2(n6977), .A(n6648), .ZN(n6651) );
  XNOR2_X1 U7729 ( .A(n6650), .B(n6651), .ZN(n7898) );
  INV_X1 U7730 ( .A(n6650), .ZN(n6653) );
  INV_X1 U7731 ( .A(n6651), .ZN(n6652) );
  NAND2_X1 U7732 ( .A1(n6653), .A2(n6652), .ZN(n6654) );
  NAND2_X1 U7733 ( .A1(n7895), .A2(n6654), .ZN(n6674) );
  INV_X1 U7734 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7173) );
  OR2_X1 U7735 ( .A1(n6604), .A2(n7173), .ZN(n6661) );
  NAND2_X1 U7736 ( .A1(n6655), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6660) );
  AOI21_X1 U7737 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6657) );
  NOR2_X1 U7738 ( .A1(n6657), .A2(n6677), .ZN(n10742) );
  NAND2_X1 U7739 ( .A1(n6656), .A2(n10742), .ZN(n6659) );
  NAND2_X1 U7740 ( .A1(n6678), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6658) );
  NAND4_X1 U7741 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .ZN(n10208)
         );
  NAND2_X1 U7742 ( .A1(n10208), .A2(n7058), .ZN(n6669) );
  OAI21_X1 U7743 ( .B1(n6663), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6664) );
  XNOR2_X1 U7744 ( .A(n6662), .B(n6664), .ZN(n7311) );
  INV_X1 U7745 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6665) );
  OR2_X1 U7746 ( .A1(n8823), .A2(n6665), .ZN(n6667) );
  OR2_X1 U7747 ( .A1(n6626), .A2(n7262), .ZN(n6666) );
  OAI211_X1 U7748 ( .C1(n7140), .C2(n7311), .A(n6667), .B(n6666), .ZN(n10744)
         );
  NAND2_X1 U7749 ( .A1(n10744), .A2(n7030), .ZN(n6668) );
  NAND2_X1 U7750 ( .A1(n6669), .A2(n6668), .ZN(n6670) );
  XNOR2_X1 U7751 ( .A(n6670), .B(n7652), .ZN(n6673) );
  NAND2_X1 U7752 ( .A1(n10208), .A2(n6977), .ZN(n6672) );
  NAND2_X1 U7753 ( .A1(n10744), .A2(n7058), .ZN(n6671) );
  NAND2_X1 U7754 ( .A1(n6672), .A2(n6671), .ZN(n7944) );
  NAND2_X1 U7755 ( .A1(n6674), .A2(n6673), .ZN(n7942) );
  INV_X1 U7756 ( .A(n7942), .ZN(n6675) );
  INV_X1 U7757 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6676) );
  OR2_X1 U7758 ( .A1(n6730), .A2(n6676), .ZN(n6683) );
  INV_X1 U7759 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8142) );
  OR2_X1 U7760 ( .A1(n6604), .A2(n8142), .ZN(n6682) );
  NAND2_X1 U7761 ( .A1(n6677), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6696) );
  OAI21_X1 U7762 ( .B1(n6677), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6696), .ZN(
        n8141) );
  OR2_X1 U7763 ( .A1(n7117), .A2(n8141), .ZN(n6681) );
  INV_X1 U7764 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6679) );
  NAND4_X1 U7765 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n10207)
         );
  NAND2_X1 U7766 ( .A1(n10207), .A2(n7058), .ZN(n6691) );
  NOR2_X1 U7767 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n6685) );
  NOR2_X1 U7768 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6684) );
  NAND3_X1 U7769 ( .A1(n6686), .A2(n6685), .A3(n6684), .ZN(n6704) );
  NAND2_X1 U7770 ( .A1(n6704), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6687) );
  XNOR2_X1 U7771 ( .A(n6687), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7226) );
  INV_X1 U7772 ( .A(n7226), .ZN(n7263) );
  OR2_X1 U7773 ( .A1(n7264), .A2(n6626), .ZN(n6689) );
  OR2_X1 U7774 ( .A1(n8823), .A2(n5193), .ZN(n6688) );
  OAI211_X1 U7775 ( .C1(n7140), .C2(n7263), .A(n6689), .B(n6688), .ZN(n8146)
         );
  NAND2_X1 U7776 ( .A1(n8146), .A2(n7030), .ZN(n6690) );
  NAND2_X1 U7777 ( .A1(n6691), .A2(n6690), .ZN(n6692) );
  XNOR2_X1 U7778 ( .A(n6692), .B(n7652), .ZN(n6717) );
  AND2_X1 U7779 ( .A1(n8146), .A2(n7058), .ZN(n6693) );
  AOI21_X1 U7780 ( .B1(n10207), .B2(n6977), .A(n6693), .ZN(n6718) );
  XNOR2_X1 U7781 ( .A(n6717), .B(n6718), .ZN(n8002) );
  INV_X1 U7782 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6694) );
  OR2_X1 U7783 ( .A1(n6604), .A2(n6694), .ZN(n6703) );
  AND2_X1 U7784 ( .A1(n6696), .A2(n6695), .ZN(n6697) );
  NOR2_X1 U7785 ( .A1(n6696), .A2(n6695), .ZN(n6732) );
  OR2_X1 U7786 ( .A1(n6697), .A2(n6732), .ZN(n8125) );
  OR2_X1 U7787 ( .A1(n7117), .A2(n8125), .ZN(n6702) );
  INV_X1 U7788 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6698) );
  OR2_X1 U7789 ( .A1(n6730), .A2(n6698), .ZN(n6701) );
  NAND2_X1 U7790 ( .A1(n7810), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6700) );
  NAND4_X1 U7791 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n10206)
         );
  NAND2_X1 U7792 ( .A1(n10206), .A2(n6995), .ZN(n6710) );
  INV_X2 U7793 ( .A(n6626), .ZN(n6723) );
  NAND2_X1 U7794 ( .A1(n7269), .A2(n6723), .ZN(n6707) );
  NAND2_X1 U7795 ( .A1(n6724), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6705) );
  XNOR2_X1 U7796 ( .A(n6705), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7326) );
  AOI22_X1 U7797 ( .A1(n6942), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7154), .B2(
        n7326), .ZN(n6706) );
  NAND2_X1 U7798 ( .A1(n6707), .A2(n6706), .ZN(n8408) );
  NAND2_X1 U7799 ( .A1(n8408), .A2(n8735), .ZN(n6709) );
  NAND2_X1 U7800 ( .A1(n6710), .A2(n6709), .ZN(n6711) );
  XNOR2_X1 U7801 ( .A(n6711), .B(n7652), .ZN(n6714) );
  INV_X1 U7802 ( .A(n6714), .ZN(n6712) );
  AOI22_X1 U7803 ( .A1(n10206), .A2(n6977), .B1(n7058), .B2(n8408), .ZN(n6713)
         );
  NAND2_X1 U7804 ( .A1(n6712), .A2(n6713), .ZN(n6720) );
  AND2_X1 U7805 ( .A1(n8002), .A2(n6716), .ZN(n6715) );
  NAND2_X1 U7806 ( .A1(n7940), .A2(n6715), .ZN(n6744) );
  INV_X1 U7807 ( .A(n6716), .ZN(n6722) );
  INV_X1 U7808 ( .A(n6717), .ZN(n6719) );
  NAND2_X1 U7809 ( .A1(n6719), .A2(n6718), .ZN(n8122) );
  AND2_X1 U7810 ( .A1(n8122), .A2(n6720), .ZN(n6721) );
  OR2_X1 U7811 ( .A1(n6722), .A2(n6721), .ZN(n6746) );
  NAND2_X1 U7812 ( .A1(n6744), .A2(n6746), .ZN(n6740) );
  NAND2_X1 U7813 ( .A1(n7273), .A2(n6723), .ZN(n6729) );
  INV_X1 U7814 ( .A(n6724), .ZN(n6726) );
  NAND2_X1 U7815 ( .A1(n6726), .A2(n6725), .ZN(n6750) );
  NAND2_X1 U7816 ( .A1(n6750), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6727) );
  XNOR2_X1 U7817 ( .A(n6727), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7228) );
  AOI22_X1 U7818 ( .A1(n6942), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7154), .B2(
        n7228), .ZN(n6728) );
  NAND2_X1 U7819 ( .A1(n8301), .A2(n7058), .ZN(n6739) );
  INV_X1 U7820 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6731) );
  OR2_X1 U7821 ( .A1(n6730), .A2(n6731), .ZN(n6737) );
  INV_X1 U7822 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8027) );
  OR2_X1 U7823 ( .A1(n6604), .A2(n8027), .ZN(n6736) );
  NAND2_X1 U7824 ( .A1(n6732), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6755) );
  OR2_X1 U7825 ( .A1(n6732), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U7826 ( .A1(n6755), .A2(n6733), .ZN(n8227) );
  OR2_X1 U7827 ( .A1(n7117), .A2(n8227), .ZN(n6735) );
  NAND2_X1 U7828 ( .A1(n7810), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6734) );
  NAND4_X1 U7829 ( .A1(n6737), .A2(n6736), .A3(n6735), .A4(n6734), .ZN(n8335)
         );
  NAND2_X1 U7830 ( .A1(n8335), .A2(n6977), .ZN(n6738) );
  AND2_X1 U7831 ( .A1(n6739), .A2(n6738), .ZN(n6745) );
  NAND2_X1 U7832 ( .A1(n6740), .A2(n6745), .ZN(n8223) );
  NAND2_X1 U7833 ( .A1(n8301), .A2(n7030), .ZN(n6742) );
  NAND2_X1 U7834 ( .A1(n8335), .A2(n7058), .ZN(n6741) );
  NAND2_X1 U7835 ( .A1(n6742), .A2(n6741), .ZN(n6743) );
  XNOR2_X1 U7836 ( .A(n6743), .B(n7652), .ZN(n8226) );
  NAND2_X1 U7837 ( .A1(n8223), .A2(n8226), .ZN(n6749) );
  INV_X1 U7838 ( .A(n6745), .ZN(n6747) );
  AND2_X1 U7839 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  NAND2_X1 U7840 ( .A1(n7284), .A2(n6723), .ZN(n6753) );
  OAI21_X1 U7841 ( .B1(n6750), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6751) );
  XNOR2_X1 U7842 ( .A(n6751), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7290) );
  AOI22_X1 U7843 ( .A1(n6942), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7154), .B2(
        n7290), .ZN(n6752) );
  NAND2_X1 U7844 ( .A1(n8471), .A2(n7030), .ZN(n6762) );
  INV_X1 U7845 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7209) );
  OR2_X1 U7846 ( .A1(n6730), .A2(n7209), .ZN(n6760) );
  NAND2_X1 U7847 ( .A1(n7809), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U7848 ( .A1(n6755), .A2(n8332), .ZN(n6756) );
  NAND2_X1 U7849 ( .A1(n6775), .A2(n6756), .ZN(n10788) );
  OR2_X1 U7850 ( .A1(n7117), .A2(n10788), .ZN(n6758) );
  NAND2_X1 U7851 ( .A1(n7810), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6757) );
  NAND4_X1 U7852 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n10811)
         );
  NAND2_X1 U7853 ( .A1(n10811), .A2(n7058), .ZN(n6761) );
  NAND2_X1 U7854 ( .A1(n6762), .A2(n6761), .ZN(n6763) );
  XNOR2_X1 U7855 ( .A(n6763), .B(n7652), .ZN(n6766) );
  AND2_X1 U7856 ( .A1(n10811), .A2(n6977), .ZN(n6765) );
  AOI21_X1 U7857 ( .B1(n8471), .B2(n6995), .A(n6765), .ZN(n6767) );
  XNOR2_X1 U7858 ( .A(n6766), .B(n6767), .ZN(n8330) );
  INV_X1 U7859 ( .A(n6766), .ZN(n6768) );
  NAND2_X1 U7860 ( .A1(n6768), .A2(n6767), .ZN(n6769) );
  NAND2_X1 U7861 ( .A1(n7293), .A2(n6723), .ZN(n6774) );
  NAND2_X1 U7862 ( .A1(n6771), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6772) );
  XNOR2_X1 U7863 ( .A(n6772), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U7864 ( .A1(n6942), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7154), .B2(
        n10228), .ZN(n6773) );
  NAND2_X1 U7865 ( .A1(n10828), .A2(n7030), .ZN(n6782) );
  INV_X1 U7866 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7208) );
  OR2_X1 U7867 ( .A1(n6730), .A2(n7208), .ZN(n6780) );
  NAND2_X1 U7868 ( .A1(n7809), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U7869 ( .A1(n6775), .A2(n8492), .ZN(n6776) );
  NAND2_X1 U7870 ( .A1(n6791), .A2(n6776), .ZN(n10820) );
  OR2_X1 U7871 ( .A1(n7117), .A2(n10820), .ZN(n6778) );
  NAND2_X1 U7872 ( .A1(n7810), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6777) );
  NAND4_X1 U7873 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n10205)
         );
  NAND2_X1 U7874 ( .A1(n10205), .A2(n7058), .ZN(n6781) );
  NAND2_X1 U7875 ( .A1(n6782), .A2(n6781), .ZN(n6783) );
  XNOR2_X1 U7876 ( .A(n6783), .B(n7652), .ZN(n6785) );
  AND2_X1 U7877 ( .A1(n10205), .A2(n6977), .ZN(n6784) );
  AOI21_X1 U7878 ( .B1(n10828), .B2(n6995), .A(n6784), .ZN(n8490) );
  NAND2_X1 U7879 ( .A1(n8488), .A2(n8490), .ZN(n6787) );
  INV_X1 U7880 ( .A(n6785), .ZN(n6786) );
  NAND2_X1 U7881 ( .A1(n7329), .A2(n6723), .ZN(n6790) );
  NOR2_X1 U7882 ( .A1(n6771), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6805) );
  OR2_X1 U7883 ( .A1(n6805), .A2(n6806), .ZN(n6788) );
  XNOR2_X1 U7884 ( .A(n6788), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7454) );
  AOI22_X1 U7885 ( .A1(n6942), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7154), .B2(
        n7454), .ZN(n6789) );
  NAND2_X1 U7886 ( .A1(n8626), .A2(n7030), .ZN(n6798) );
  INV_X1 U7887 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8483) );
  OR2_X1 U7888 ( .A1(n6604), .A2(n8483), .ZN(n6796) );
  AND2_X1 U7889 ( .A1(n6791), .A2(n8518), .ZN(n6792) );
  OR2_X1 U7890 ( .A1(n6792), .A2(n6809), .ZN(n8521) );
  OR2_X1 U7891 ( .A1(n7117), .A2(n8521), .ZN(n6795) );
  INV_X1 U7892 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7207) );
  OR2_X1 U7893 ( .A1(n6730), .A2(n7207), .ZN(n6794) );
  NAND2_X1 U7894 ( .A1(n7810), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6793) );
  NAND4_X1 U7895 ( .A1(n6796), .A2(n6795), .A3(n6794), .A4(n6793), .ZN(n10871)
         );
  NAND2_X1 U7896 ( .A1(n10871), .A2(n6995), .ZN(n6797) );
  NAND2_X1 U7897 ( .A1(n6798), .A2(n6797), .ZN(n6799) );
  XNOR2_X1 U7898 ( .A(n6799), .B(n7652), .ZN(n6801) );
  AND2_X1 U7899 ( .A1(n10871), .A2(n6977), .ZN(n6800) );
  AOI21_X1 U7900 ( .B1(n8626), .B2(n6995), .A(n6800), .ZN(n6802) );
  INV_X1 U7901 ( .A(n6801), .ZN(n6803) );
  NAND2_X1 U7902 ( .A1(n6803), .A2(n6802), .ZN(n6804) );
  NAND2_X1 U7903 ( .A1(n7374), .A2(n6723), .ZN(n6808) );
  AND2_X1 U7904 ( .A1(n6805), .A2(n9026), .ZN(n6866) );
  OR2_X1 U7905 ( .A1(n6866), .A2(n6806), .ZN(n6821) );
  XNOR2_X1 U7906 ( .A(n6821), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7432) );
  AOI22_X1 U7907 ( .A1(n6942), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7154), .B2(
        n7432), .ZN(n6807) );
  NAND2_X1 U7908 ( .A1(n10884), .A2(n8735), .ZN(n6816) );
  NAND2_X1 U7909 ( .A1(n7809), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6814) );
  INV_X1 U7910 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7206) );
  OR2_X1 U7911 ( .A1(n6730), .A2(n7206), .ZN(n6813) );
  NAND2_X1 U7912 ( .A1(n6809), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6826) );
  OR2_X1 U7913 ( .A1(n6809), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U7914 ( .A1(n6826), .A2(n6810), .ZN(n10882) );
  OR2_X1 U7915 ( .A1(n7117), .A2(n10882), .ZN(n6812) );
  NAND2_X1 U7916 ( .A1(n7810), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6811) );
  NAND4_X1 U7917 ( .A1(n6814), .A2(n6813), .A3(n6812), .A4(n6811), .ZN(n10204)
         );
  NAND2_X1 U7918 ( .A1(n10204), .A2(n6995), .ZN(n6815) );
  NAND2_X1 U7919 ( .A1(n6816), .A2(n6815), .ZN(n6817) );
  XNOR2_X1 U7920 ( .A(n6817), .B(n8732), .ZN(n8551) );
  AND2_X1 U7921 ( .A1(n10204), .A2(n6977), .ZN(n6818) );
  AOI21_X1 U7922 ( .B1(n10884), .B2(n6995), .A(n6818), .ZN(n8550) );
  INV_X1 U7923 ( .A(n8551), .ZN(n6820) );
  INV_X1 U7924 ( .A(n8550), .ZN(n6819) );
  NAND2_X1 U7925 ( .A1(n7428), .A2(n6723), .ZN(n6824) );
  NAND2_X1 U7926 ( .A1(n6821), .A2(n9246), .ZN(n6822) );
  NAND2_X1 U7927 ( .A1(n6822), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6842) );
  XNOR2_X1 U7928 ( .A(n6842), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7780) );
  AOI22_X1 U7929 ( .A1(n6942), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7154), .B2(
        n7780), .ZN(n6823) );
  NAND2_X1 U7930 ( .A1(n8683), .A2(n8735), .ZN(n6833) );
  INV_X1 U7931 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8632) );
  OR2_X1 U7932 ( .A1(n6604), .A2(n8632), .ZN(n6831) );
  NAND2_X1 U7933 ( .A1(n6826), .A2(n6825), .ZN(n6827) );
  NAND2_X1 U7934 ( .A1(n6847), .A2(n6827), .ZN(n8671) );
  OR2_X1 U7935 ( .A1(n7117), .A2(n8671), .ZN(n6830) );
  INV_X1 U7936 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7205) );
  OR2_X1 U7937 ( .A1(n6730), .A2(n7205), .ZN(n6829) );
  NAND2_X1 U7938 ( .A1(n7810), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6828) );
  NAND4_X1 U7939 ( .A1(n6831), .A2(n6830), .A3(n6829), .A4(n6828), .ZN(n10870)
         );
  NAND2_X1 U7940 ( .A1(n10870), .A2(n6995), .ZN(n6832) );
  NAND2_X1 U7941 ( .A1(n6833), .A2(n6832), .ZN(n6834) );
  XNOR2_X1 U7942 ( .A(n6834), .B(n7652), .ZN(n6837) );
  NAND2_X1 U7943 ( .A1(n8683), .A2(n6995), .ZN(n6836) );
  NAND2_X1 U7944 ( .A1(n10870), .A2(n6977), .ZN(n6835) );
  NAND2_X1 U7945 ( .A1(n6836), .A2(n6835), .ZN(n6838) );
  NAND2_X1 U7946 ( .A1(n6837), .A2(n6838), .ZN(n8665) );
  INV_X1 U7947 ( .A(n6837), .ZN(n6840) );
  INV_X1 U7948 ( .A(n6838), .ZN(n6839) );
  NAND2_X1 U7949 ( .A1(n6840), .A2(n6839), .ZN(n8667) );
  NAND2_X1 U7950 ( .A1(n7468), .A2(n6723), .ZN(n6846) );
  NAND2_X1 U7951 ( .A1(n6842), .A2(n6841), .ZN(n6843) );
  NAND2_X1 U7952 ( .A1(n6843), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6844) );
  XNOR2_X1 U7953 ( .A(n6844), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7235) );
  AOI22_X1 U7954 ( .A1(n6942), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7154), .B2(
        n7235), .ZN(n6845) );
  NAND2_X1 U7955 ( .A1(n9809), .A2(n8735), .ZN(n6855) );
  INV_X1 U7956 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8677) );
  OR2_X1 U7957 ( .A1(n6604), .A2(n8677), .ZN(n6853) );
  AND2_X1 U7958 ( .A1(n6847), .A2(n7802), .ZN(n6848) );
  OR2_X1 U7959 ( .A1(n6848), .A2(n6871), .ZN(n9807) );
  OR2_X1 U7960 ( .A1(n7117), .A2(n9807), .ZN(n6852) );
  INV_X1 U7961 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6849) );
  OR2_X1 U7962 ( .A1(n6730), .A2(n6849), .ZN(n6851) );
  NAND2_X1 U7963 ( .A1(n7810), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6850) );
  NAND4_X1 U7964 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n10203)
         );
  NAND2_X1 U7965 ( .A1(n10203), .A2(n6995), .ZN(n6854) );
  NAND2_X1 U7966 ( .A1(n6855), .A2(n6854), .ZN(n6856) );
  XNOR2_X1 U7967 ( .A(n6856), .B(n8732), .ZN(n6860) );
  NAND2_X1 U7968 ( .A1(n6859), .A2(n6860), .ZN(n9798) );
  NAND2_X1 U7969 ( .A1(n9809), .A2(n6995), .ZN(n6858) );
  NAND2_X1 U7970 ( .A1(n10203), .A2(n6977), .ZN(n6857) );
  NAND2_X1 U7971 ( .A1(n6858), .A2(n6857), .ZN(n9802) );
  NAND2_X1 U7972 ( .A1(n9798), .A2(n9802), .ZN(n6863) );
  INV_X1 U7973 ( .A(n6860), .ZN(n6861) );
  NAND2_X1 U7974 ( .A1(n7853), .A2(n6723), .ZN(n6870) );
  NOR2_X1 U7975 ( .A1(n6864), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U7976 ( .A1(n6866), .A2(n6865), .ZN(n6884) );
  NAND2_X1 U7977 ( .A1(n6884), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6867) );
  XNOR2_X1 U7978 ( .A(n6867), .B(n9251), .ZN(n8118) );
  INV_X1 U7979 ( .A(n8118), .ZN(n6868) );
  AOI22_X1 U7980 ( .A1(n6942), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7154), .B2(
        n6868), .ZN(n6869) );
  NAND2_X1 U7981 ( .A1(n9929), .A2(n8735), .ZN(n6878) );
  NAND2_X1 U7982 ( .A1(n6655), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U7983 ( .A1(n7809), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6875) );
  NOR2_X1 U7984 ( .A1(n6871), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6872) );
  OR2_X1 U7985 ( .A1(n6888), .A2(n6872), .ZN(n9925) );
  OR2_X1 U7986 ( .A1(n7117), .A2(n9925), .ZN(n6874) );
  NAND2_X1 U7987 ( .A1(n7810), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6873) );
  NAND4_X1 U7988 ( .A1(n6876), .A2(n6875), .A3(n6874), .A4(n6873), .ZN(n10945)
         );
  NAND2_X1 U7989 ( .A1(n10945), .A2(n6995), .ZN(n6877) );
  NAND2_X1 U7990 ( .A1(n6878), .A2(n6877), .ZN(n6879) );
  NAND2_X1 U7991 ( .A1(n9929), .A2(n6995), .ZN(n6881) );
  NAND2_X1 U7992 ( .A1(n10945), .A2(n6977), .ZN(n6880) );
  NAND2_X1 U7993 ( .A1(n6881), .A2(n6880), .ZN(n9916) );
  NAND2_X1 U7994 ( .A1(n9912), .A2(n9916), .ZN(n6883) );
  NAND2_X1 U7995 ( .A1(n6882), .A2(n5069), .ZN(n9914) );
  NAND2_X1 U7996 ( .A1(n6883), .A2(n9914), .ZN(n9847) );
  INV_X1 U7997 ( .A(n9847), .ZN(n6899) );
  NAND2_X1 U7998 ( .A1(n7856), .A2(n6723), .ZN(n6887) );
  NAND2_X1 U7999 ( .A1(n6885), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6904) );
  XNOR2_X1 U8000 ( .A(n6904), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7858) );
  AOI22_X1 U8001 ( .A1(n6942), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7154), .B2(
        n7858), .ZN(n6886) );
  NAND2_X1 U8002 ( .A1(n10960), .A2(n8735), .ZN(n6895) );
  NAND2_X1 U8003 ( .A1(n6655), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6893) );
  NAND2_X1 U8004 ( .A1(n7809), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6892) );
  OR2_X1 U8005 ( .A1(n6888), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U8006 ( .A1(n6910), .A2(n6889), .ZN(n10956) );
  OR2_X1 U8007 ( .A1(n7117), .A2(n10956), .ZN(n6891) );
  NAND2_X1 U8008 ( .A1(n7810), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6890) );
  NAND4_X1 U8009 ( .A1(n6893), .A2(n6892), .A3(n6891), .A4(n6890), .ZN(n10436)
         );
  NAND2_X1 U8010 ( .A1(n10436), .A2(n6995), .ZN(n6894) );
  NAND2_X1 U8011 ( .A1(n6895), .A2(n6894), .ZN(n6896) );
  XNOR2_X1 U8012 ( .A(n6896), .B(n8732), .ZN(n6901) );
  AND2_X1 U8013 ( .A1(n10436), .A2(n6977), .ZN(n6897) );
  AOI21_X1 U8014 ( .B1(n10960), .B2(n6995), .A(n6897), .ZN(n6900) );
  XNOR2_X1 U8015 ( .A(n6901), .B(n6900), .ZN(n9850) );
  NAND2_X1 U8016 ( .A1(n6899), .A2(n6898), .ZN(n9848) );
  NAND2_X1 U8017 ( .A1(n6901), .A2(n6900), .ZN(n6902) );
  NAND2_X1 U8018 ( .A1(n9848), .A2(n6902), .ZN(n9856) );
  NAND2_X1 U8019 ( .A1(n7880), .A2(n6723), .ZN(n6907) );
  NAND2_X1 U8020 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  NAND2_X1 U8021 ( .A1(n6905), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6925) );
  XNOR2_X1 U8022 ( .A(n6925), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U8023 ( .A1(n6942), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7154), .B2(
        n10245), .ZN(n6906) );
  NAND2_X1 U8024 ( .A1(n10516), .A2(n8735), .ZN(n6917) );
  NAND2_X1 U8025 ( .A1(n7809), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6915) );
  INV_X1 U8026 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6908) );
  OR2_X1 U8027 ( .A1(n6730), .A2(n6908), .ZN(n6914) );
  INV_X1 U8028 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U8029 ( .A1(n6910), .A2(n6909), .ZN(n6911) );
  NAND2_X1 U8030 ( .A1(n6930), .A2(n6911), .ZN(n10442) );
  OR2_X1 U8031 ( .A1(n7117), .A2(n10442), .ZN(n6913) );
  NAND2_X1 U8032 ( .A1(n7810), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6912) );
  NAND4_X1 U8033 ( .A1(n6915), .A2(n6914), .A3(n6913), .A4(n6912), .ZN(n10943)
         );
  NAND2_X1 U8034 ( .A1(n10943), .A2(n6995), .ZN(n6916) );
  NAND2_X1 U8035 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  XNOR2_X1 U8036 ( .A(n6918), .B(n7652), .ZN(n6920) );
  AND2_X1 U8037 ( .A1(n10943), .A2(n6977), .ZN(n6919) );
  AOI21_X1 U8038 ( .B1(n10516), .B2(n6995), .A(n6919), .ZN(n6921) );
  XNOR2_X1 U8039 ( .A(n6920), .B(n6921), .ZN(n9858) );
  INV_X1 U8040 ( .A(n6920), .ZN(n6922) );
  AND2_X1 U8041 ( .A1(n6922), .A2(n6921), .ZN(n6923) );
  AOI21_X1 U8042 ( .B1(n9856), .B2(n9858), .A(n6923), .ZN(n6941) );
  NAND2_X1 U8043 ( .A1(n7965), .A2(n6723), .ZN(n6929) );
  NAND2_X1 U8044 ( .A1(n6925), .A2(n6924), .ZN(n6926) );
  NAND2_X1 U8045 ( .A1(n6926), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6927) );
  XNOR2_X1 U8046 ( .A(n6927), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U8047 ( .A1(n6942), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7154), .B2(
        n10658), .ZN(n6928) );
  NAND2_X1 U8048 ( .A1(n10426), .A2(n8735), .ZN(n6937) );
  NAND2_X1 U8049 ( .A1(n7809), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6935) );
  AND2_X1 U8050 ( .A1(n6930), .A2(n9896), .ZN(n6931) );
  NOR2_X1 U8051 ( .A1(n6945), .A2(n6931), .ZN(n10425) );
  NAND2_X1 U8052 ( .A1(n10425), .A2(n6656), .ZN(n6934) );
  INV_X1 U8053 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10240) );
  OR2_X1 U8054 ( .A1(n6730), .A2(n10240), .ZN(n6933) );
  NAND2_X1 U8055 ( .A1(n7810), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6932) );
  NAND4_X1 U8056 ( .A1(n6935), .A2(n6934), .A3(n6933), .A4(n6932), .ZN(n10435)
         );
  NAND2_X1 U8057 ( .A1(n10435), .A2(n6995), .ZN(n6936) );
  NAND2_X1 U8058 ( .A1(n6937), .A2(n6936), .ZN(n6938) );
  XNOR2_X1 U8059 ( .A(n6938), .B(n7652), .ZN(n6940) );
  AND2_X1 U8060 ( .A1(n10435), .A2(n6977), .ZN(n6939) );
  AOI21_X1 U8061 ( .B1(n10426), .B2(n6995), .A(n6939), .ZN(n9891) );
  NOR2_X1 U8062 ( .A1(n9890), .A2(n9891), .ZN(n9889) );
  NOR2_X2 U8063 ( .A1(n9889), .A2(n9894), .ZN(n9824) );
  NAND2_X1 U8064 ( .A1(n8163), .A2(n6723), .ZN(n6944) );
  AOI22_X1 U8065 ( .A1(n6942), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10366), 
        .B2(n7154), .ZN(n6943) );
  NOR2_X1 U8066 ( .A1(n6945), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6946) );
  OR2_X1 U8067 ( .A1(n6958), .A2(n6946), .ZN(n10392) );
  INV_X1 U8068 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6947) );
  OAI22_X1 U8069 ( .A1(n10392), .A2(n7117), .B1(n6730), .B2(n6947), .ZN(n6950)
         );
  INV_X1 U8070 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U8071 ( .A1(n7810), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6948) );
  OAI21_X1 U8072 ( .B1(n10393), .B2(n6604), .A(n6948), .ZN(n6949) );
  AOI22_X1 U8073 ( .A1(n10506), .A2(n8735), .B1(n7058), .B2(n10418), .ZN(n6951) );
  NAND2_X1 U8074 ( .A1(n9824), .A2(n5079), .ZN(n6953) );
  AOI22_X1 U8075 ( .A1(n10506), .A2(n7058), .B1(n6977), .B2(n10418), .ZN(n9822) );
  NAND2_X1 U8076 ( .A1(n8325), .A2(n6723), .ZN(n6957) );
  OR2_X1 U8077 ( .A1(n8823), .A2(n8326), .ZN(n6956) );
  NAND2_X1 U8078 ( .A1(n10500), .A2(n8735), .ZN(n6963) );
  NOR2_X1 U8079 ( .A1(n6958), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6959) );
  OR2_X1 U8080 ( .A1(n6970), .A2(n6959), .ZN(n10380) );
  AOI22_X1 U8081 ( .A1(n7809), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n6655), .B2(
        P1_REG1_REG_20__SCAN_IN), .ZN(n6961) );
  NAND2_X1 U8082 ( .A1(n7810), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6960) );
  OAI211_X1 U8083 ( .C1(n10380), .C2(n7117), .A(n6961), .B(n6960), .ZN(n10359)
         );
  NAND2_X1 U8084 ( .A1(n10359), .A2(n6995), .ZN(n6962) );
  NAND2_X1 U8085 ( .A1(n6963), .A2(n6962), .ZN(n6964) );
  XNOR2_X1 U8086 ( .A(n6964), .B(n8732), .ZN(n6967) );
  AND2_X1 U8087 ( .A1(n10359), .A2(n6977), .ZN(n6965) );
  AOI21_X1 U8088 ( .B1(n10500), .B2(n7058), .A(n6965), .ZN(n6966) );
  NOR2_X1 U8089 ( .A1(n6967), .A2(n6966), .ZN(n9872) );
  NAND2_X1 U8090 ( .A1(n8348), .A2(n6723), .ZN(n6969) );
  INV_X1 U8091 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8383) );
  OR2_X1 U8092 ( .A1(n8823), .A2(n8383), .ZN(n6968) );
  NAND2_X1 U8093 ( .A1(n10496), .A2(n7030), .ZN(n6975) );
  OR2_X1 U8094 ( .A1(n6970), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U8095 ( .A1(n6971), .A2(n6985), .ZN(n10361) );
  AOI22_X1 U8096 ( .A1(n7809), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n7810), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6973) );
  NAND2_X1 U8097 ( .A1(n6655), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6972) );
  OAI211_X1 U8098 ( .C1(n10361), .C2(n7117), .A(n6973), .B(n6972), .ZN(n10374)
         );
  NAND2_X1 U8099 ( .A1(n10374), .A2(n6995), .ZN(n6974) );
  NAND2_X1 U8100 ( .A1(n6975), .A2(n6974), .ZN(n6976) );
  XNOR2_X1 U8101 ( .A(n6976), .B(n8732), .ZN(n6982) );
  INV_X1 U8102 ( .A(n6982), .ZN(n6980) );
  AND2_X1 U8103 ( .A1(n10374), .A2(n6977), .ZN(n6978) );
  AOI21_X1 U8104 ( .B1(n10496), .B2(n6995), .A(n6978), .ZN(n6981) );
  INV_X1 U8105 ( .A(n6981), .ZN(n6979) );
  NAND2_X1 U8106 ( .A1(n6980), .A2(n6979), .ZN(n9831) );
  NAND2_X1 U8107 ( .A1(n8536), .A2(n6723), .ZN(n6984) );
  OR2_X1 U8108 ( .A1(n8823), .A2(n8537), .ZN(n6983) );
  NAND2_X1 U8109 ( .A1(n10491), .A2(n8735), .ZN(n6992) );
  NAND2_X1 U8110 ( .A1(n6655), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U8111 ( .A1(n7809), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6989) );
  OAI21_X1 U8112 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n6986), .A(n7002), .ZN(
        n10341) );
  OR2_X1 U8113 ( .A1(n7117), .A2(n10341), .ZN(n6988) );
  NAND2_X1 U8114 ( .A1(n7810), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6987) );
  NAND4_X1 U8115 ( .A1(n6990), .A2(n6989), .A3(n6988), .A4(n6987), .ZN(n10335)
         );
  NAND2_X1 U8116 ( .A1(n10335), .A2(n6995), .ZN(n6991) );
  NAND2_X1 U8117 ( .A1(n6992), .A2(n6991), .ZN(n6993) );
  XNOR2_X1 U8118 ( .A(n6993), .B(n8732), .ZN(n6997) );
  AND2_X1 U8119 ( .A1(n10335), .A2(n6977), .ZN(n6994) );
  AOI21_X1 U8120 ( .B1(n10491), .B2(n6995), .A(n6994), .ZN(n6996) );
  NOR2_X1 U8121 ( .A1(n6997), .A2(n6996), .ZN(n9882) );
  NAND2_X1 U8122 ( .A1(n6997), .A2(n6996), .ZN(n9880) );
  NAND2_X1 U8123 ( .A1(n8545), .A2(n6723), .ZN(n6999) );
  OR2_X1 U8124 ( .A1(n8823), .A2(n8548), .ZN(n6998) );
  NAND2_X1 U8125 ( .A1(n7809), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7007) );
  NAND2_X1 U8126 ( .A1(n7810), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7006) );
  INV_X1 U8127 ( .A(n7002), .ZN(n7000) );
  NAND2_X1 U8128 ( .A1(n7000), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7016) );
  INV_X1 U8129 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7001) );
  NAND2_X1 U8130 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  NAND2_X1 U8131 ( .A1(n7016), .A2(n7003), .ZN(n10326) );
  OR2_X1 U8132 ( .A1(n7117), .A2(n10326), .ZN(n7005) );
  NAND2_X1 U8133 ( .A1(n6655), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7004) );
  NAND4_X1 U8134 ( .A1(n7007), .A2(n7006), .A3(n7005), .A4(n7004), .ZN(n10202)
         );
  AOI22_X1 U8135 ( .A1(n10484), .A2(n8735), .B1(n7058), .B2(n10202), .ZN(n7008) );
  XNOR2_X1 U8136 ( .A(n7008), .B(n7652), .ZN(n7010) );
  NOR2_X1 U8137 ( .A1(n7011), .A2(n7010), .ZN(n9814) );
  OAI22_X1 U8138 ( .A1(n10329), .A2(n6764), .B1(n10348), .B2(n7009), .ZN(n9815) );
  NAND2_X1 U8139 ( .A1(n7011), .A2(n7010), .ZN(n9812) );
  NAND2_X1 U8140 ( .A1(n8578), .A2(n6723), .ZN(n7013) );
  INV_X1 U8141 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8581) );
  OR2_X1 U8142 ( .A1(n8823), .A2(n8581), .ZN(n7012) );
  NAND2_X1 U8143 ( .A1(n10481), .A2(n8735), .ZN(n7023) );
  NAND2_X1 U8144 ( .A1(n7809), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U8145 ( .A1(n6655), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n7020) );
  INV_X1 U8146 ( .A(n7016), .ZN(n7014) );
  NAND2_X1 U8147 ( .A1(n7014), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7033) );
  INV_X1 U8148 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n7015) );
  NAND2_X1 U8149 ( .A1(n7016), .A2(n7015), .ZN(n7017) );
  NAND2_X1 U8150 ( .A1(n7033), .A2(n7017), .ZN(n10318) );
  OR2_X1 U8151 ( .A1(n7117), .A2(n10318), .ZN(n7019) );
  NAND2_X1 U8152 ( .A1(n7810), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7018) );
  NAND4_X1 U8153 ( .A1(n7021), .A2(n7020), .A3(n7019), .A4(n7018), .ZN(n10334)
         );
  NAND2_X1 U8154 ( .A1(n10334), .A2(n7058), .ZN(n7022) );
  NAND2_X1 U8155 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  XNOR2_X1 U8156 ( .A(n7024), .B(n7652), .ZN(n7025) );
  AOI22_X1 U8157 ( .A1(n10481), .A2(n7058), .B1(n6977), .B2(n10334), .ZN(n7026) );
  XNOR2_X1 U8158 ( .A(n7025), .B(n7026), .ZN(n9865) );
  INV_X1 U8159 ( .A(n7025), .ZN(n7027) );
  NAND2_X1 U8160 ( .A1(n8687), .A2(n6723), .ZN(n7029) );
  OR2_X1 U8161 ( .A1(n8823), .A2(n9195), .ZN(n7028) );
  NAND2_X1 U8162 ( .A1(n10474), .A2(n7030), .ZN(n7040) );
  NAND2_X1 U8163 ( .A1(n7809), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7038) );
  NAND2_X1 U8164 ( .A1(n6655), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7037) );
  INV_X1 U8165 ( .A(n7033), .ZN(n7031) );
  NAND2_X1 U8166 ( .A1(n7031), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7051) );
  INV_X1 U8167 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7032) );
  NAND2_X1 U8168 ( .A1(n7033), .A2(n7032), .ZN(n7034) );
  NAND2_X1 U8169 ( .A1(n7051), .A2(n7034), .ZN(n10295) );
  OR2_X1 U8170 ( .A1(n7117), .A2(n10295), .ZN(n7036) );
  NAND2_X1 U8171 ( .A1(n7810), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7035) );
  NAND4_X1 U8172 ( .A1(n7038), .A2(n7037), .A3(n7036), .A4(n7035), .ZN(n10288)
         );
  NAND2_X1 U8173 ( .A1(n10288), .A2(n7058), .ZN(n7039) );
  NAND2_X1 U8174 ( .A1(n7040), .A2(n7039), .ZN(n7041) );
  XNOR2_X1 U8175 ( .A(n7041), .B(n7652), .ZN(n9840) );
  NAND2_X1 U8176 ( .A1(n10474), .A2(n7058), .ZN(n7043) );
  NAND2_X1 U8177 ( .A1(n10288), .A2(n6977), .ZN(n7042) );
  NAND2_X1 U8178 ( .A1(n7043), .A2(n7042), .ZN(n7045) );
  INV_X1 U8179 ( .A(n7045), .ZN(n9839) );
  NAND2_X1 U8180 ( .A1(n8702), .A2(n6723), .ZN(n7048) );
  OR2_X1 U8181 ( .A1(n8823), .A2(n9191), .ZN(n7047) );
  NAND2_X1 U8182 ( .A1(n7809), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7056) );
  NAND2_X1 U8183 ( .A1(n6655), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n7055) );
  INV_X1 U8184 ( .A(n7051), .ZN(n7049) );
  NAND2_X1 U8185 ( .A1(n7049), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7067) );
  INV_X1 U8186 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U8187 ( .A1(n7051), .A2(n7050), .ZN(n7052) );
  NAND2_X1 U8188 ( .A1(n7067), .A2(n7052), .ZN(n10280) );
  NAND2_X1 U8189 ( .A1(n7810), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7053) );
  NAND4_X1 U8190 ( .A1(n7056), .A2(n7055), .A3(n7054), .A4(n7053), .ZN(n10201)
         );
  AND2_X1 U8191 ( .A1(n10201), .A2(n6977), .ZN(n7057) );
  AOI21_X1 U8192 ( .B1(n10469), .B2(n7058), .A(n7057), .ZN(n7060) );
  AOI22_X1 U8193 ( .A1(n10469), .A2(n8735), .B1(n7058), .B2(n10201), .ZN(n7059) );
  XNOR2_X1 U8194 ( .A(n7059), .B(n7652), .ZN(n7061) );
  XOR2_X1 U8195 ( .A(n7060), .B(n7061), .Z(n9904) );
  NOR2_X1 U8196 ( .A1(n7061), .A2(n7060), .ZN(n7062) );
  NAND2_X1 U8197 ( .A1(n8707), .A2(n6723), .ZN(n7064) );
  OR2_X1 U8198 ( .A1(n8823), .A2(n9190), .ZN(n7063) );
  NAND2_X1 U8199 ( .A1(n10464), .A2(n8735), .ZN(n7074) );
  NAND2_X1 U8200 ( .A1(n7809), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7072) );
  NAND2_X1 U8201 ( .A1(n6655), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7071) );
  INV_X1 U8202 ( .A(n7067), .ZN(n7065) );
  NAND2_X1 U8203 ( .A1(n7065), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n7115) );
  INV_X1 U8204 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7066) );
  NAND2_X1 U8205 ( .A1(n7067), .A2(n7066), .ZN(n7068) );
  NAND2_X1 U8206 ( .A1(n7115), .A2(n7068), .ZN(n7106) );
  NAND2_X1 U8207 ( .A1(n7810), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7069) );
  NAND4_X1 U8208 ( .A1(n7072), .A2(n7071), .A3(n7070), .A4(n7069), .ZN(n10287)
         );
  NAND2_X1 U8209 ( .A1(n10287), .A2(n7058), .ZN(n7073) );
  NAND2_X1 U8210 ( .A1(n7074), .A2(n7073), .ZN(n7075) );
  XNOR2_X1 U8211 ( .A(n7075), .B(n7652), .ZN(n7079) );
  NAND2_X1 U8212 ( .A1(n10464), .A2(n7058), .ZN(n7077) );
  NAND2_X1 U8213 ( .A1(n10287), .A2(n6977), .ZN(n7076) );
  NAND2_X1 U8214 ( .A1(n7077), .A2(n7076), .ZN(n7078) );
  NOR2_X1 U8215 ( .A1(n7079), .A2(n7078), .ZN(n8739) );
  AOI21_X1 U8216 ( .B1(n7079), .B2(n7078), .A(n8739), .ZN(n7080) );
  INV_X1 U8217 ( .A(n7083), .ZN(n8688) );
  NAND3_X1 U8218 ( .A1(n8688), .A2(P1_B_REG_SCAN_IN), .A3(n8583), .ZN(n7084)
         );
  INV_X1 U8219 ( .A(n7085), .ZN(n8706) );
  NAND2_X1 U8220 ( .A1(n8706), .A2(n8583), .ZN(n10536) );
  NOR4_X1 U8221 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n7090) );
  NOR4_X1 U8222 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n7089) );
  NOR4_X1 U8223 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n7088) );
  NOR4_X1 U8224 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n7087) );
  AND4_X1 U8225 ( .A1(n7090), .A2(n7089), .A3(n7088), .A4(n7087), .ZN(n7096)
         );
  NOR2_X1 U8226 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n7094) );
  NOR4_X1 U8227 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n7093) );
  NOR4_X1 U8228 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n7092) );
  NOR4_X1 U8229 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n7091) );
  AND4_X1 U8230 ( .A1(n7094), .A2(n7093), .A3(n7092), .A4(n7091), .ZN(n7095)
         );
  NAND2_X1 U8231 ( .A1(n7096), .A2(n7095), .ZN(n7391) );
  INV_X1 U8232 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7268) );
  NOR2_X1 U8233 ( .A1(n7391), .A2(n7268), .ZN(n7097) );
  OR2_X1 U8234 ( .A1(n7393), .A2(n7097), .ZN(n7098) );
  NAND2_X1 U8235 ( .A1(n8706), .A2(n8688), .ZN(n7390) );
  AND2_X1 U8236 ( .A1(n7098), .A2(n7390), .ZN(n7745) );
  NAND2_X1 U8237 ( .A1(n7408), .A2(n7745), .ZN(n7125) );
  INV_X1 U8238 ( .A(n7099), .ZN(n7100) );
  NAND2_X1 U8239 ( .A1(n7100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7101) );
  NOR2_X1 U8240 ( .A1(n7125), .A2(n7399), .ZN(n7104) );
  INV_X1 U8241 ( .A(n7846), .ZN(n7386) );
  AND2_X1 U8242 ( .A1(n10970), .A2(n10018), .ZN(n7102) );
  NAND2_X1 U8243 ( .A1(n7103), .A2(n9893), .ZN(n7134) );
  NAND2_X1 U8244 ( .A1(n7846), .A2(n10115), .ZN(n7109) );
  INV_X1 U8245 ( .A(n7109), .ZN(n10743) );
  NAND2_X1 U8246 ( .A1(n7104), .A2(n10743), .ZN(n7105) );
  NAND2_X1 U8247 ( .A1(n10973), .A2(n10366), .ZN(n7395) );
  INV_X1 U8248 ( .A(n7106), .ZN(n10266) );
  OR2_X1 U8249 ( .A1(n7845), .A2(n10018), .ZN(n7397) );
  AND3_X1 U8250 ( .A1(n7160), .A2(n8546), .A3(n7397), .ZN(n7107) );
  NAND2_X1 U8251 ( .A1(n7125), .A2(n10970), .ZN(n7423) );
  NAND2_X1 U8252 ( .A1(n7107), .A2(n7423), .ZN(n7108) );
  NAND2_X1 U8253 ( .A1(n7108), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7111) );
  NOR2_X1 U8254 ( .A1(n7109), .A2(n7399), .ZN(n7110) );
  NAND2_X1 U8255 ( .A1(n7125), .A2(n7110), .ZN(n7424) );
  NAND2_X1 U8256 ( .A1(n7111), .A2(n7424), .ZN(n9900) );
  NAND2_X1 U8257 ( .A1(n7809), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7122) );
  INV_X1 U8258 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7112) );
  INV_X1 U8259 ( .A(n7115), .ZN(n7113) );
  NAND2_X1 U8260 ( .A1(n7113), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8786) );
  INV_X1 U8261 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7114) );
  NAND2_X1 U8262 ( .A1(n7115), .A2(n7114), .ZN(n7116) );
  NAND2_X1 U8263 ( .A1(n8786), .A2(n7116), .ZN(n8849) );
  OR2_X1 U8264 ( .A1(n7117), .A2(n8849), .ZN(n7120) );
  INV_X1 U8265 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7118) );
  OR2_X1 U8266 ( .A1(n6730), .A2(n7118), .ZN(n7119) );
  OR2_X1 U8267 ( .A1(n7124), .A2(n7123), .ZN(n7653) );
  OR2_X1 U8268 ( .A1(n7399), .A2(n7653), .ZN(n9933) );
  NOR2_X1 U8269 ( .A1(n7125), .A2(n9933), .ZN(n7128) );
  NAND2_X1 U8270 ( .A1(n7128), .A2(n7127), .ZN(n9919) );
  INV_X1 U8271 ( .A(n7127), .ZN(n7179) );
  AND2_X2 U8272 ( .A1(n7128), .A2(n7179), .ZN(n9923) );
  AOI22_X1 U8273 ( .A1(n10201), .A2(n9923), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n7129) );
  OAI21_X1 U8274 ( .B1(n10272), .B2(n9919), .A(n7129), .ZN(n7130) );
  AOI21_X1 U8275 ( .B1(n10266), .B2(n9900), .A(n7130), .ZN(n7131) );
  NAND2_X1 U8276 ( .A1(n7134), .A2(n7133), .ZN(P1_U3212) );
  INV_X1 U8277 ( .A(n7135), .ZN(n7136) );
  NAND2_X1 U8278 ( .A1(n7160), .A2(n10018), .ZN(n7139) );
  NAND2_X1 U8279 ( .A1(n7139), .A2(n8546), .ZN(n7153) );
  NAND2_X1 U8280 ( .A1(n7153), .A2(n7140), .ZN(n7141) );
  NAND2_X1 U8281 ( .A1(n7141), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8282 ( .A(n7311), .ZN(n7151) );
  XNOR2_X1 U8283 ( .A(n7253), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n10214) );
  AND2_X1 U8284 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n10213) );
  NAND2_X1 U8285 ( .A1(n10214), .A2(n10213), .ZN(n10212) );
  INV_X1 U8286 ( .A(n7253), .ZN(n10219) );
  NAND2_X1 U8287 ( .A1(n10219), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7142) );
  NAND2_X1 U8288 ( .A1(n10212), .A2(n7142), .ZN(n7192) );
  XNOR2_X1 U8289 ( .A(n7252), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n7193) );
  AND2_X1 U8290 ( .A1(n7192), .A2(n7193), .ZN(n7194) );
  INV_X1 U8291 ( .A(n7194), .ZN(n7144) );
  INV_X1 U8292 ( .A(n7252), .ZN(n7166) );
  NAND2_X1 U8293 ( .A1(n7166), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7143) );
  NAND2_X1 U8294 ( .A1(n7144), .A2(n7143), .ZN(n7362) );
  XNOR2_X1 U8295 ( .A(n7373), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n7363) );
  NAND2_X1 U8296 ( .A1(n7362), .A2(n7363), .ZN(n7361) );
  INV_X1 U8297 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7145) );
  OR2_X1 U8298 ( .A1(n7373), .A2(n7145), .ZN(n7146) );
  NAND2_X1 U8299 ( .A1(n7361), .A2(n7146), .ZN(n7644) );
  MUX2_X1 U8300 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7147), .S(n7643), .Z(n7645)
         );
  OR2_X1 U8301 ( .A1(n7644), .A2(n7645), .ZN(n7149) );
  NAND2_X1 U8302 ( .A1(n7643), .A2(n7147), .ZN(n7148) );
  NAND2_X1 U8303 ( .A1(n7149), .A2(n7148), .ZN(n7306) );
  INV_X1 U8304 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7150) );
  XNOR2_X1 U8305 ( .A(n7311), .B(n7150), .ZN(n7307) );
  NOR2_X1 U8306 ( .A1(n7306), .A2(n7307), .ZN(n7305) );
  AOI21_X1 U8307 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n7151), .A(n7305), .ZN(
        n7158) );
  NAND2_X1 U8308 ( .A1(n7226), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7152) );
  OAI21_X1 U8309 ( .B1(n7226), .B2(P1_REG1_REG_6__SCAN_IN), .A(n7152), .ZN(
        n7157) );
  NOR2_X1 U8310 ( .A1(n7158), .A2(n7157), .ZN(n7210) );
  NAND2_X1 U8311 ( .A1(n7153), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7178) );
  OR2_X1 U8312 ( .A1(n7178), .A2(n7154), .ZN(n10644) );
  INV_X1 U8313 ( .A(n10644), .ZN(n7156) );
  NAND2_X1 U8314 ( .A1(n7156), .A2(n7155), .ZN(n10254) );
  AOI211_X1 U8315 ( .C1(n7158), .C2(n7157), .A(n7210), .B(n10254), .ZN(n7185)
         );
  INV_X1 U8316 ( .A(n8546), .ZN(n7159) );
  NOR2_X1 U8317 ( .A1(n7160), .A2(n7159), .ZN(n7161) );
  INV_X1 U8318 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7164) );
  INV_X1 U8319 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7162) );
  NOR2_X1 U8320 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7162), .ZN(n8003) );
  INV_X1 U8321 ( .A(n8003), .ZN(n7163) );
  OAI21_X1 U8322 ( .B1(n7784), .B2(n7164), .A(n7163), .ZN(n7184) );
  XNOR2_X1 U8323 ( .A(n7253), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n10218) );
  AND2_X1 U8324 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n10217) );
  NAND2_X1 U8325 ( .A1(n10218), .A2(n10217), .ZN(n10215) );
  NAND2_X1 U8326 ( .A1(n10219), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7165) );
  NAND2_X1 U8327 ( .A1(n10215), .A2(n7165), .ZN(n7198) );
  XNOR2_X1 U8328 ( .A(n7252), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n7199) );
  NAND2_X1 U8329 ( .A1(n7198), .A2(n7199), .ZN(n7197) );
  NAND2_X1 U8330 ( .A1(n7166), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7167) );
  NAND2_X1 U8331 ( .A1(n7197), .A2(n7167), .ZN(n7369) );
  XNOR2_X1 U8332 ( .A(n7373), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n7370) );
  NAND2_X1 U8333 ( .A1(n7369), .A2(n7370), .ZN(n7368) );
  INV_X1 U8334 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7168) );
  OR2_X1 U8335 ( .A1(n7373), .A2(n7168), .ZN(n7169) );
  NAND2_X1 U8336 ( .A1(n7368), .A2(n7169), .ZN(n7640) );
  INV_X1 U8337 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7170) );
  MUX2_X1 U8338 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7170), .S(n7643), .Z(n7641)
         );
  NOR2_X1 U8339 ( .A1(n7640), .A2(n7641), .ZN(n7639) );
  AND2_X1 U8340 ( .A1(n7643), .A2(n7170), .ZN(n7171) );
  NOR2_X1 U8341 ( .A1(n7639), .A2(n7171), .ZN(n7309) );
  XNOR2_X1 U8342 ( .A(n7311), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n7308) );
  INV_X1 U8343 ( .A(n7308), .ZN(n7172) );
  OR2_X1 U8344 ( .A1(n7309), .A2(n7172), .ZN(n7175) );
  NAND2_X1 U8345 ( .A1(n7311), .A2(n7173), .ZN(n7174) );
  NAND2_X1 U8346 ( .A1(n7175), .A2(n7174), .ZN(n7181) );
  OR2_X1 U8347 ( .A1(n7226), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7177) );
  NAND2_X1 U8348 ( .A1(n7226), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7176) );
  NAND2_X1 U8349 ( .A1(n7177), .A2(n7176), .ZN(n7180) );
  NOR2_X1 U8350 ( .A1(n7181), .A2(n7180), .ZN(n7225) );
  NOR2_X1 U8351 ( .A1(n7178), .A2(n7155), .ZN(n7453) );
  NAND2_X1 U8352 ( .A1(n7453), .A2(n7179), .ZN(n10651) );
  AOI211_X1 U8353 ( .C1(n7181), .C2(n7180), .A(n7225), .B(n10651), .ZN(n7183)
         );
  NAND2_X1 U8354 ( .A1(n7453), .A2(n7127), .ZN(n10249) );
  NOR2_X1 U8355 ( .A1(n10249), .A2(n7263), .ZN(n7182) );
  OR4_X1 U8356 ( .A1(n7185), .A2(n7184), .A3(n7183), .A4(n7182), .ZN(P1_U3247)
         );
  OAI21_X1 U8357 ( .B1(n7188), .B2(n7187), .A(n7186), .ZN(n8795) );
  MUX2_X1 U8358 ( .A(n10637), .B(n8795), .S(n7155), .Z(n7190) );
  NOR2_X1 U8359 ( .A1(n7155), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7189) );
  OR2_X1 U8360 ( .A1(n7189), .A2(n7127), .ZN(n10634) );
  NAND2_X1 U8361 ( .A1(n10634), .A2(n10637), .ZN(n10640) );
  OAI211_X1 U8362 ( .C1(n7190), .C2(n10634), .A(P1_U4006), .B(n10640), .ZN(
        n7191) );
  INV_X1 U8363 ( .A(n7191), .ZN(n7650) );
  INV_X1 U8364 ( .A(n7192), .ZN(n7196) );
  INV_X1 U8365 ( .A(n7193), .ZN(n7195) );
  AOI211_X1 U8366 ( .C1(n7196), .C2(n7195), .A(n7194), .B(n10254), .ZN(n7204)
         );
  OAI211_X1 U8367 ( .C1(n7199), .C2(n7198), .A(n10216), .B(n7197), .ZN(n7200)
         );
  OAI21_X1 U8368 ( .B1(n10249), .B2(n7252), .A(n7200), .ZN(n7203) );
  INV_X1 U8369 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7201) );
  OAI22_X1 U8370 ( .A1(n7784), .A2(n7201), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7933), .ZN(n7202) );
  OR4_X1 U8371 ( .A1(n7650), .A2(n7204), .A3(n7203), .A4(n7202), .ZN(P1_U3243)
         );
  INV_X1 U8372 ( .A(n7235), .ZN(n7804) );
  AOI22_X1 U8373 ( .A1(n7235), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n6849), .B2(
        n7804), .ZN(n7801) );
  MUX2_X1 U8374 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7205), .S(n7780), .Z(n7779)
         );
  MUX2_X1 U8375 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7206), .S(n7432), .Z(n7435)
         );
  MUX2_X1 U8376 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7207), .S(n7454), .Z(n7452)
         );
  OR2_X1 U8377 ( .A1(n10228), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7212) );
  MUX2_X1 U8378 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7208), .S(n10228), .Z(
        n10231) );
  MUX2_X1 U8379 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7209), .S(n7290), .Z(n7334)
         );
  INV_X1 U8380 ( .A(n7228), .ZN(n7357) );
  AOI22_X1 U8381 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n7228), .B1(n7357), .B2(
        n6731), .ZN(n7349) );
  AOI21_X1 U8382 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n7226), .A(n7210), .ZN(
        n7318) );
  NOR2_X1 U8383 ( .A1(n7326), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7211) );
  AOI21_X1 U8384 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n7326), .A(n7211), .ZN(
        n7317) );
  NAND2_X1 U8385 ( .A1(n7318), .A2(n7317), .ZN(n7316) );
  OAI21_X1 U8386 ( .B1(n7326), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7316), .ZN(
        n7348) );
  NAND2_X1 U8387 ( .A1(n7349), .A2(n7348), .ZN(n7347) );
  OAI21_X1 U8388 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7228), .A(n7347), .ZN(
        n7335) );
  NAND2_X1 U8389 ( .A1(n7334), .A2(n7335), .ZN(n7333) );
  OAI21_X1 U8390 ( .B1(n7290), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7333), .ZN(
        n10232) );
  NAND2_X1 U8391 ( .A1(n10231), .A2(n10232), .ZN(n10230) );
  NAND2_X1 U8392 ( .A1(n7212), .A2(n10230), .ZN(n7451) );
  NAND2_X1 U8393 ( .A1(n7452), .A2(n7451), .ZN(n7450) );
  OAI21_X1 U8394 ( .B1(n7454), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7450), .ZN(
        n7434) );
  NAND2_X1 U8395 ( .A1(n7435), .A2(n7434), .ZN(n7433) );
  OAI21_X1 U8396 ( .B1(n7432), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7433), .ZN(
        n7778) );
  NAND2_X1 U8397 ( .A1(n7779), .A2(n7778), .ZN(n7777) );
  OAI21_X1 U8398 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7780), .A(n7777), .ZN(
        n7800) );
  NAND2_X1 U8399 ( .A1(n7801), .A2(n7800), .ZN(n7799) );
  OAI21_X1 U8400 ( .B1(n7235), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7799), .ZN(
        n7213) );
  NOR2_X1 U8401 ( .A1(n8118), .A2(n7213), .ZN(n7214) );
  INV_X1 U8402 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10932) );
  XNOR2_X1 U8403 ( .A(n7213), .B(n8118), .ZN(n8113) );
  NOR2_X1 U8404 ( .A1(n10932), .A2(n8113), .ZN(n8112) );
  NOR2_X1 U8405 ( .A1(n7214), .A2(n8112), .ZN(n8274) );
  INV_X1 U8406 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10953) );
  NOR2_X1 U8407 ( .A1(n7858), .A2(n10953), .ZN(n7215) );
  AOI21_X1 U8408 ( .B1(n7858), .B2(n10953), .A(n7215), .ZN(n8273) );
  NOR2_X1 U8409 ( .A1(n8274), .A2(n8273), .ZN(n8272) );
  AOI21_X1 U8410 ( .B1(n7858), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8272), .ZN(
        n7217) );
  XNOR2_X1 U8411 ( .A(n10245), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7216) );
  NOR2_X1 U8412 ( .A1(n7217), .A2(n7216), .ZN(n10238) );
  AOI211_X1 U8413 ( .C1(n7217), .C2(n7216), .A(n10238), .B(n10254), .ZN(n7246)
         );
  INV_X1 U8414 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7219) );
  NAND2_X1 U8415 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(n5013), .ZN(n7218) );
  OAI21_X1 U8416 ( .B1(n7784), .B2(n7219), .A(n7218), .ZN(n7245) );
  NOR2_X1 U8417 ( .A1(n7804), .A2(n8677), .ZN(n7796) );
  NAND2_X1 U8418 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7780), .ZN(n7234) );
  MUX2_X1 U8419 ( .A(n8632), .B(P1_REG2_REG_13__SCAN_IN), .S(n7780), .Z(n7220)
         );
  INV_X1 U8420 ( .A(n7220), .ZN(n7775) );
  NAND2_X1 U8421 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7432), .ZN(n7233) );
  INV_X1 U8422 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7221) );
  MUX2_X1 U8423 ( .A(n7221), .B(P1_REG2_REG_12__SCAN_IN), .S(n7432), .Z(n7222)
         );
  INV_X1 U8424 ( .A(n7222), .ZN(n7441) );
  INV_X1 U8425 ( .A(n7454), .ZN(n7223) );
  NAND2_X1 U8426 ( .A1(n7223), .A2(n8483), .ZN(n7459) );
  NAND2_X1 U8427 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n10228), .ZN(n7230) );
  NAND2_X1 U8428 ( .A1(n7290), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7224) );
  OAI21_X1 U8429 ( .B1(n7290), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7224), .ZN(
        n7340) );
  AOI22_X1 U8430 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7228), .B1(n7357), .B2(
        n8027), .ZN(n7352) );
  AOI21_X1 U8431 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n7226), .A(n7225), .ZN(
        n7321) );
  NOR2_X1 U8432 ( .A1(n7326), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7227) );
  AOI21_X1 U8433 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7326), .A(n7227), .ZN(
        n7320) );
  NAND2_X1 U8434 ( .A1(n7321), .A2(n7320), .ZN(n7319) );
  OAI21_X1 U8435 ( .B1(n7326), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7319), .ZN(
        n7351) );
  NAND2_X1 U8436 ( .A1(n7352), .A2(n7351), .ZN(n7350) );
  OAI21_X1 U8437 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7228), .A(n7350), .ZN(
        n7341) );
  NOR2_X1 U8438 ( .A1(n7340), .A2(n7341), .ZN(n7339) );
  AOI21_X1 U8439 ( .B1(n7290), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7339), .ZN(
        n10226) );
  OAI21_X1 U8440 ( .B1(n10228), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7230), .ZN(
        n10225) );
  NOR2_X1 U8441 ( .A1(n10226), .A2(n10225), .ZN(n10224) );
  INV_X1 U8442 ( .A(n10224), .ZN(n7229) );
  NAND2_X1 U8443 ( .A1(n7230), .A2(n7229), .ZN(n7460) );
  NAND2_X1 U8444 ( .A1(n7459), .A2(n7460), .ZN(n7232) );
  NAND2_X1 U8445 ( .A1(n7454), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7231) );
  NAND2_X1 U8446 ( .A1(n7232), .A2(n7231), .ZN(n7461) );
  NAND2_X1 U8447 ( .A1(n7441), .A2(n7461), .ZN(n7440) );
  NAND2_X1 U8448 ( .A1(n7233), .A2(n7440), .ZN(n7776) );
  NAND2_X1 U8449 ( .A1(n7775), .A2(n7776), .ZN(n7774) );
  NAND2_X1 U8450 ( .A1(n7234), .A2(n7774), .ZN(n7797) );
  OAI22_X1 U8451 ( .A1(n7796), .A2(n7797), .B1(n7235), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n7236) );
  NOR2_X1 U8452 ( .A1(n8118), .A2(n7236), .ZN(n7237) );
  INV_X1 U8453 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8115) );
  XNOR2_X1 U8454 ( .A(n7236), .B(n8118), .ZN(n8116) );
  NOR2_X1 U8455 ( .A1(n8115), .A2(n8116), .ZN(n8114) );
  NOR2_X1 U8456 ( .A1(n7237), .A2(n8114), .ZN(n8271) );
  NAND2_X1 U8457 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7858), .ZN(n7238) );
  OAI21_X1 U8458 ( .B1(n7858), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7238), .ZN(
        n8270) );
  NOR2_X1 U8459 ( .A1(n8271), .A2(n8270), .ZN(n8269) );
  AOI21_X1 U8460 ( .B1(n7858), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8269), .ZN(
        n7241) );
  NAND2_X1 U8461 ( .A1(n10245), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7239) );
  OAI21_X1 U8462 ( .B1(n10245), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7239), .ZN(
        n7240) );
  NOR2_X1 U8463 ( .A1(n7241), .A2(n7240), .ZN(n10244) );
  AOI211_X1 U8464 ( .C1(n7241), .C2(n7240), .A(n10244), .B(n10651), .ZN(n7244)
         );
  INV_X1 U8465 ( .A(n10245), .ZN(n7242) );
  NOR2_X1 U8466 ( .A1(n10249), .A2(n7242), .ZN(n7243) );
  OR4_X1 U8467 ( .A1(n7246), .A2(n7245), .A3(n7244), .A4(n7243), .ZN(P1_U3258)
         );
  NOR2_X1 U8468 ( .A1(n5724), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9794) );
  INV_X2 U8469 ( .A(n9794), .ZN(n8691) );
  OAI222_X1 U8470 ( .A1(n8831), .A2(n7248), .B1(n8691), .B2(n7251), .C1(
        P2_U3152), .C2(n7247), .ZN(P2_U3356) );
  OAI222_X1 U8471 ( .A1(n8831), .A2(n7249), .B1(n8691), .B2(n7255), .C1(
        P2_U3152), .C2(n7521), .ZN(P2_U3355) );
  INV_X2 U8472 ( .A(n8544), .ZN(n10541) );
  INV_X1 U8473 ( .A(n10539), .ZN(n8855) );
  OAI222_X1 U8474 ( .A1(n7252), .A2(P1_U3084), .B1(n10541), .B2(n7251), .C1(
        n7250), .C2(n8855), .ZN(P1_U3351) );
  OAI222_X1 U8475 ( .A1(n8855), .A2(n7254), .B1(n10541), .B2(n7257), .C1(
        P1_U3084), .C2(n7253), .ZN(P1_U3352) );
  OAI222_X1 U8476 ( .A1(n7373), .A2(n5013), .B1(n10541), .B2(n7255), .C1(n5107), .C2(n8855), .ZN(P1_U3350) );
  OAI222_X1 U8477 ( .A1(n8691), .A2(n7257), .B1(n7696), .B2(P2_U3152), .C1(
        n7256), .C2(n8831), .ZN(P2_U3357) );
  OAI222_X1 U8478 ( .A1(n8855), .A2(n7258), .B1(n10541), .B2(n7259), .C1(n5013), .C2(n7643), .ZN(P1_U3349) );
  INV_X1 U8479 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7260) );
  INV_X1 U8480 ( .A(n7608), .ZN(n7523) );
  OAI222_X1 U8481 ( .A1(n8831), .A2(n7260), .B1(n8691), .B2(n7259), .C1(
        P2_U3152), .C2(n7523), .ZN(P2_U3354) );
  INV_X1 U8482 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7261) );
  INV_X1 U8483 ( .A(n7545), .ZN(n7524) );
  OAI222_X1 U8484 ( .A1(n8831), .A2(n7261), .B1(n8691), .B2(n7262), .C1(
        P2_U3152), .C2(n7524), .ZN(P2_U3353) );
  OAI222_X1 U8485 ( .A1(n7311), .A2(P1_U3084), .B1(n10541), .B2(n7262), .C1(
        n8855), .C2(n6665), .ZN(P1_U3348) );
  OAI222_X1 U8486 ( .A1(n8855), .A2(n5193), .B1(n10541), .B2(n7264), .C1(n7263), .C2(n5013), .ZN(P1_U3347) );
  INV_X1 U8487 ( .A(n7571), .ZN(n7527) );
  OAI222_X1 U8488 ( .A1(n8831), .A2(n5213), .B1(n8691), .B2(n7264), .C1(
        P2_U3152), .C2(n7527), .ZN(P2_U3352) );
  INV_X1 U8489 ( .A(n7393), .ZN(n7265) );
  INV_X1 U8490 ( .A(n7399), .ZN(n7267) );
  INV_X1 U8491 ( .A(n7390), .ZN(n7266) );
  AOI22_X1 U8492 ( .A1(n10549), .A2(n7268), .B1(n7267), .B2(n7266), .ZN(
        P1_U3441) );
  INV_X1 U8493 ( .A(n7269), .ZN(n7271) );
  AOI22_X1 U8494 ( .A1(n7326), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10539), .ZN(n7270) );
  OAI21_X1 U8495 ( .B1(n7271), .B2(n10541), .A(n7270), .ZN(P1_U3346) );
  INV_X1 U8496 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7272) );
  INV_X1 U8497 ( .A(n7583), .ZN(n7528) );
  OAI222_X1 U8498 ( .A1(n8831), .A2(n7272), .B1(n8691), .B2(n7271), .C1(
        P2_U3152), .C2(n7528), .ZN(P2_U3351) );
  INV_X1 U8499 ( .A(n7558), .ZN(n7530) );
  INV_X1 U8500 ( .A(n7273), .ZN(n7274) );
  OAI222_X1 U8501 ( .A1(n7530), .A2(P2_U3152), .B1(n8691), .B2(n7274), .C1(
        n8831), .C2(n5628), .ZN(P2_U3350) );
  OAI222_X1 U8502 ( .A1(n7357), .A2(n5013), .B1(n10541), .B2(n7274), .C1(n9007), .C2(n8855), .ZN(P1_U3345) );
  INV_X1 U8503 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U8504 ( .A1(P2_U3966), .A2(n8394), .ZN(n7275) );
  OAI21_X1 U8505 ( .B1(P2_U3966), .B2(n7292), .A(n7275), .ZN(P2_U3561) );
  NAND2_X1 U8506 ( .A1(P2_U3966), .A2(n8455), .ZN(n7276) );
  OAI21_X1 U8507 ( .B1(P2_U3966), .B2(n6665), .A(n7276), .ZN(P2_U3557) );
  INV_X1 U8508 ( .A(n7755), .ZN(n7277) );
  NAND2_X1 U8509 ( .A1(P2_U3966), .A2(n7277), .ZN(n7278) );
  OAI21_X1 U8510 ( .B1(P2_U3966), .B2(n5263), .A(n7278), .ZN(P2_U3552) );
  INV_X1 U8511 ( .A(n8541), .ZN(n7280) );
  OAI21_X1 U8512 ( .B1(n10552), .B2(n7280), .A(n7279), .ZN(n7283) );
  NAND2_X1 U8513 ( .A1(n10552), .A2(n7281), .ZN(n7282) );
  INV_X1 U8514 ( .A(n8373), .ZN(n10674) );
  NOR2_X1 U8515 ( .A1(n10674), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8516 ( .A(n7284), .ZN(n7291) );
  INV_X1 U8517 ( .A(n8831), .ZN(n7966) );
  AOI22_X1 U8518 ( .A1(n7596), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n7966), .ZN(n7285) );
  OAI21_X1 U8519 ( .B1(n7291), .B2(n8691), .A(n7285), .ZN(P2_U3349) );
  NAND2_X1 U8520 ( .A1(n9385), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7286) );
  OAI21_X1 U8521 ( .B1(n9385), .B2(n7287), .A(n7286), .ZN(P2_U3583) );
  INV_X1 U8522 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7289) );
  NAND2_X1 U8523 ( .A1(n7651), .A2(P1_U4006), .ZN(n7288) );
  OAI21_X1 U8524 ( .B1(P1_U4006), .B2(n7289), .A(n7288), .ZN(P1_U3555) );
  INV_X1 U8525 ( .A(n7290), .ZN(n7338) );
  OAI222_X1 U8526 ( .A1(n7338), .A2(P1_U3084), .B1(n8855), .B2(n7292), .C1(
        n7291), .C2(n10541), .ZN(P1_U3344) );
  INV_X1 U8527 ( .A(n7293), .ZN(n7296) );
  AOI22_X1 U8528 ( .A1(n7629), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n7966), .ZN(n7294) );
  OAI21_X1 U8529 ( .B1(n7296), .B2(n8691), .A(n7294), .ZN(P2_U3348) );
  AOI22_X1 U8530 ( .A1(n10228), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10539), .ZN(n7295) );
  OAI21_X1 U8531 ( .B1(n7296), .B2(n10541), .A(n7295), .ZN(P1_U3343) );
  NAND2_X1 U8532 ( .A1(n6655), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7299) );
  NAND2_X1 U8533 ( .A1(n7809), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7298) );
  NAND2_X1 U8534 ( .A1(n7810), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7297) );
  NAND2_X1 U8535 ( .A1(n10211), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7300) );
  OAI21_X1 U8536 ( .B1(n10012), .B2(n10211), .A(n7300), .ZN(P1_U3586) );
  NAND2_X1 U8537 ( .A1(n6655), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7303) );
  NAND2_X1 U8538 ( .A1(n7809), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7302) );
  NAND2_X1 U8539 ( .A1(n7810), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7301) );
  AND3_X1 U8540 ( .A1(n7303), .A2(n7302), .A3(n7301), .ZN(n10109) );
  NAND2_X1 U8541 ( .A1(n10211), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7304) );
  OAI21_X1 U8542 ( .B1(n10109), .B2(n10211), .A(n7304), .ZN(P1_U3585) );
  AOI211_X1 U8543 ( .C1(n7307), .C2(n7306), .A(n7305), .B(n10254), .ZN(n7315)
         );
  XNOR2_X1 U8544 ( .A(n7309), .B(n7308), .ZN(n7310) );
  OAI22_X1 U8545 ( .A1(n7311), .A2(n10249), .B1(n10651), .B2(n7310), .ZN(n7314) );
  INV_X1 U8546 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7312) );
  NAND2_X1 U8547 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7947) );
  OAI21_X1 U8548 ( .B1(n7784), .B2(n7312), .A(n7947), .ZN(n7313) );
  OR3_X1 U8549 ( .A1(n7315), .A2(n7314), .A3(n7313), .ZN(P1_U3246) );
  INV_X1 U8550 ( .A(n10254), .ZN(n10649) );
  OAI21_X1 U8551 ( .B1(n7318), .B2(n7317), .A(n7316), .ZN(n7323) );
  OAI21_X1 U8552 ( .B1(n7321), .B2(n7320), .A(n7319), .ZN(n7322) );
  AOI22_X1 U8553 ( .A1(n10649), .A2(n7323), .B1(n10216), .B2(n7322), .ZN(n7328) );
  INV_X1 U8554 ( .A(n10249), .ZN(n10657) );
  INV_X1 U8555 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U8556 ( .A1(n5013), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8127) );
  OAI21_X1 U8557 ( .B1(n7784), .B2(n7324), .A(n8127), .ZN(n7325) );
  AOI21_X1 U8558 ( .B1(n10657), .B2(n7326), .A(n7325), .ZN(n7327) );
  NAND2_X1 U8559 ( .A1(n7328), .A2(n7327), .ZN(P1_U3248) );
  INV_X1 U8560 ( .A(n7329), .ZN(n7332) );
  AOI22_X1 U8561 ( .A1(n7454), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10539), .ZN(n7330) );
  OAI21_X1 U8562 ( .B1(n7332), .B2(n10541), .A(n7330), .ZN(P1_U3342) );
  INV_X1 U8563 ( .A(n7630), .ZN(n7683) );
  INV_X1 U8564 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7331) );
  OAI222_X1 U8565 ( .A1(n8691), .A2(n7332), .B1(n7683), .B2(P2_U3152), .C1(
        n7331), .C2(n8831), .ZN(P2_U3347) );
  OAI21_X1 U8566 ( .B1(n7335), .B2(n7334), .A(n7333), .ZN(n7344) );
  NAND2_X1 U8567 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n7337) );
  NAND2_X1 U8568 ( .A1(n10648), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n7336) );
  OAI211_X1 U8569 ( .C1(n10249), .C2(n7338), .A(n7337), .B(n7336), .ZN(n7343)
         );
  AOI211_X1 U8570 ( .C1(n7341), .C2(n7340), .A(n7339), .B(n10651), .ZN(n7342)
         );
  AOI211_X1 U8571 ( .C1(n10649), .C2(n7344), .A(n7343), .B(n7342), .ZN(n7345)
         );
  INV_X1 U8572 ( .A(n7345), .ZN(P1_U3250) );
  NAND2_X1 U8573 ( .A1(n8335), .A2(P1_U4006), .ZN(n7346) );
  OAI21_X1 U8574 ( .B1(P1_U4006), .B2(n5628), .A(n7346), .ZN(P1_U3563) );
  OAI21_X1 U8575 ( .B1(n7349), .B2(n7348), .A(n7347), .ZN(n7359) );
  OAI21_X1 U8576 ( .B1(n7352), .B2(n7351), .A(n7350), .ZN(n7353) );
  NAND2_X1 U8577 ( .A1(n7353), .A2(n10216), .ZN(n7356) );
  INV_X1 U8578 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7354) );
  NOR2_X1 U8579 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7354), .ZN(n8228) );
  AOI21_X1 U8580 ( .B1(n10648), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n8228), .ZN(
        n7355) );
  OAI211_X1 U8581 ( .C1(n10249), .C2(n7357), .A(n7356), .B(n7355), .ZN(n7358)
         );
  AOI21_X1 U8582 ( .B1(n10649), .B2(n7359), .A(n7358), .ZN(n7360) );
  INV_X1 U8583 ( .A(n7360), .ZN(P1_U3249) );
  INV_X1 U8584 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7366) );
  OAI211_X1 U8585 ( .C1(n7363), .C2(n7362), .A(n10649), .B(n7361), .ZN(n7365)
         );
  INV_X1 U8586 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7848) );
  NOR2_X1 U8587 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7848), .ZN(n7702) );
  INV_X1 U8588 ( .A(n7702), .ZN(n7364) );
  OAI211_X1 U8589 ( .C1(n7366), .C2(n7784), .A(n7365), .B(n7364), .ZN(n7367)
         );
  INV_X1 U8590 ( .A(n7367), .ZN(n7372) );
  OAI211_X1 U8591 ( .C1(n7370), .C2(n7369), .A(n10216), .B(n7368), .ZN(n7371)
         );
  OAI211_X1 U8592 ( .C1(n10249), .C2(n7373), .A(n7372), .B(n7371), .ZN(
        P1_U3244) );
  INV_X1 U8593 ( .A(n7374), .ZN(n7376) );
  AOI22_X1 U8594 ( .A1(n7432), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10539), .ZN(n7375) );
  OAI21_X1 U8595 ( .B1(n7376), .B2(n10541), .A(n7375), .ZN(P1_U3341) );
  INV_X1 U8596 ( .A(n7625), .ZN(n7672) );
  OAI222_X1 U8597 ( .A1(n8831), .A2(n7377), .B1(n8691), .B2(n7376), .C1(
        P2_U3152), .C2(n7672), .ZN(P2_U3346) );
  AOI21_X1 U8598 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n7385) );
  INV_X1 U8599 ( .A(n9397), .ZN(n7763) );
  OAI22_X1 U8600 ( .A1(n7763), .A2(n9565), .B1(n7755), .B2(n9641), .ZN(n7862)
         );
  INV_X1 U8601 ( .A(n7381), .ZN(n8040) );
  NAND2_X1 U8602 ( .A1(n7382), .A2(n8040), .ZN(n7413) );
  AOI22_X1 U8603 ( .A1(n9373), .A2(n7862), .B1(n7413), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7384) );
  NAND2_X1 U8604 ( .A1(n9379), .A2(n8108), .ZN(n7383) );
  OAI211_X1 U8605 ( .C1(n7385), .C2(n9381), .A(n7384), .B(n7383), .ZN(P2_U3224) );
  NOR2_X1 U8606 ( .A1(n7651), .A2(n8799), .ZN(n7835) );
  AND2_X1 U8607 ( .A1(n7651), .A2(n8799), .ZN(n10046) );
  NOR2_X1 U8608 ( .A1(n7835), .A2(n10046), .ZN(n10153) );
  NAND2_X1 U8609 ( .A1(n7386), .A2(n7653), .ZN(n7389) );
  INV_X1 U8610 ( .A(n7836), .ZN(n7388) );
  INV_X1 U8611 ( .A(n10018), .ZN(n7387) );
  OAI22_X1 U8612 ( .A1(n10153), .A2(n7389), .B1(n7388), .B2(n10403), .ZN(
        n10698) );
  AOI21_X1 U8613 ( .B1(n7846), .B2(n10694), .A(n10698), .ZN(n7412) );
  OAI21_X1 U8614 ( .B1(n7393), .B2(P1_D_REG_1__SCAN_IN), .A(n7390), .ZN(n7396)
         );
  INV_X1 U8615 ( .A(n7391), .ZN(n7392) );
  OR2_X1 U8616 ( .A1(n7393), .A2(n7392), .ZN(n7394) );
  NAND3_X1 U8617 ( .A1(n7396), .A2(n7395), .A3(n7394), .ZN(n7400) );
  INV_X1 U8618 ( .A(n7397), .ZN(n7398) );
  NAND2_X1 U8619 ( .A1(n10975), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7401) );
  OAI21_X1 U8620 ( .B1(n7412), .B2(n10975), .A(n7401), .ZN(P1_U3523) );
  XNOR2_X1 U8621 ( .A(n7403), .B(n7402), .ZN(n7407) );
  AOI22_X1 U8622 ( .A1(n9379), .A2(n8061), .B1(n7413), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7406) );
  AOI22_X1 U8623 ( .A1(n9335), .A2(n7404), .B1(n9334), .B2(n9396), .ZN(n7405)
         );
  OAI211_X1 U8624 ( .C1(n7407), .C2(n9381), .A(n7406), .B(n7405), .ZN(P2_U3239) );
  INV_X1 U8625 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7410) );
  OR2_X1 U8626 ( .A1(n10981), .A2(n7410), .ZN(n7411) );
  OAI21_X1 U8627 ( .B1(n7412), .B2(n10978), .A(n7411), .ZN(P1_U3454) );
  AOI22_X1 U8628 ( .A1(n9379), .A2(n10701), .B1(n7413), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7417) );
  MUX2_X1 U8629 ( .A(n10701), .B(n7414), .S(n6274), .Z(n7415) );
  INV_X1 U8630 ( .A(n8034), .ZN(n7861) );
  OAI21_X1 U8631 ( .B1(n7415), .B2(n7861), .A(n9352), .ZN(n7416) );
  OAI211_X1 U8632 ( .C1(n9362), .C2(n6329), .A(n7417), .B(n7416), .ZN(P2_U3234) );
  XNOR2_X1 U8633 ( .A(n7419), .B(n7418), .ZN(n7421) );
  XNOR2_X1 U8634 ( .A(n7421), .B(n7420), .ZN(n7427) );
  AOI22_X1 U8635 ( .A1(n9906), .A2(n7830), .B1(n9923), .B2(n7651), .ZN(n7426)
         );
  INV_X1 U8636 ( .A(n7422), .ZN(n7744) );
  NAND3_X1 U8637 ( .A1(n7424), .A2(n7423), .A3(n7744), .ZN(n8796) );
  AOI22_X1 U8638 ( .A1(n9928), .A2(n7654), .B1(n8796), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7425) );
  OAI211_X1 U8639 ( .C1(n7427), .C2(n9931), .A(n7426), .B(n7425), .ZN(P1_U3220) );
  INV_X1 U8640 ( .A(n7428), .ZN(n7431) );
  AOI22_X1 U8641 ( .A1(n7780), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10539), .ZN(n7429) );
  OAI21_X1 U8642 ( .B1(n7431), .B2(n10541), .A(n7429), .ZN(P1_U3340) );
  AOI22_X1 U8643 ( .A1(n7723), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n7966), .ZN(n7430) );
  OAI21_X1 U8644 ( .B1(n7431), .B2(n8691), .A(n7430), .ZN(P2_U3345) );
  INV_X1 U8645 ( .A(n7432), .ZN(n7444) );
  OAI21_X1 U8646 ( .B1(n7435), .B2(n7434), .A(n7433), .ZN(n7439) );
  INV_X1 U8647 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7436) );
  NOR2_X1 U8648 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7436), .ZN(n8554) );
  INV_X1 U8649 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7437) );
  NOR2_X1 U8650 ( .A1(n7784), .A2(n7437), .ZN(n7438) );
  AOI211_X1 U8651 ( .C1(n10649), .C2(n7439), .A(n8554), .B(n7438), .ZN(n7443)
         );
  OAI211_X1 U8652 ( .C1(n7461), .C2(n7441), .A(n10216), .B(n7440), .ZN(n7442)
         );
  OAI211_X1 U8653 ( .C1(n10249), .C2(n7444), .A(n7443), .B(n7442), .ZN(
        P1_U3253) );
  XOR2_X1 U8654 ( .A(n7446), .B(n7445), .Z(n7449) );
  AOI22_X1 U8655 ( .A1(n9906), .A2(n10210), .B1(n9923), .B2(n7836), .ZN(n7448)
         );
  AOI22_X1 U8656 ( .A1(n9928), .A2(n10053), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n8796), .ZN(n7447) );
  OAI211_X1 U8657 ( .C1(n7449), .C2(n9931), .A(n7448), .B(n7447), .ZN(P1_U3235) );
  OAI21_X1 U8658 ( .B1(n7452), .B2(n7451), .A(n7450), .ZN(n7466) );
  INV_X1 U8659 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7458) );
  AND3_X1 U8660 ( .A1(n7453), .A2(n7460), .A3(P1_REG2_REG_11__SCAN_IN), .ZN(
        n7455) );
  OAI21_X1 U8661 ( .B1(n10657), .B2(n7455), .A(n7454), .ZN(n7457) );
  NAND2_X1 U8662 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(n5013), .ZN(n7456) );
  OAI211_X1 U8663 ( .C1(n7458), .C2(n7784), .A(n7457), .B(n7456), .ZN(n7465)
         );
  INV_X1 U8664 ( .A(n7459), .ZN(n7463) );
  INV_X1 U8665 ( .A(n7460), .ZN(n7462) );
  AOI211_X1 U8666 ( .C1(n7463), .C2(n7462), .A(n7461), .B(n10651), .ZN(n7464)
         );
  AOI211_X1 U8667 ( .C1(n10649), .C2(n7466), .A(n7465), .B(n7464), .ZN(n7467)
         );
  INV_X1 U8668 ( .A(n7467), .ZN(P1_U3252) );
  INV_X1 U8669 ( .A(n7468), .ZN(n7637) );
  AOI22_X1 U8670 ( .A1(n7972), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n7966), .ZN(n7469) );
  OAI21_X1 U8671 ( .B1(n7637), .B2(n8691), .A(n7469), .ZN(P2_U3344) );
  NAND2_X1 U8672 ( .A1(n10552), .A2(n7470), .ZN(n7473) );
  INV_X1 U8673 ( .A(n7471), .ZN(n7472) );
  NAND3_X1 U8674 ( .A1(n7473), .A2(n8541), .A3(n7472), .ZN(n7477) );
  NAND2_X1 U8675 ( .A1(n7477), .A2(n7475), .ZN(n7474) );
  NAND2_X1 U8676 ( .A1(n7474), .A2(n9385), .ZN(n7494) );
  INV_X1 U8677 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7487) );
  AND2_X1 U8678 ( .A1(n7475), .A2(n5941), .ZN(n7476) );
  NAND2_X1 U8679 ( .A1(n7477), .A2(n7476), .ZN(n9422) );
  XNOR2_X1 U8680 ( .A(n7696), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n7684) );
  NAND2_X1 U8681 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n7688) );
  INV_X1 U8682 ( .A(n7688), .ZN(n7478) );
  NAND2_X1 U8683 ( .A1(n7684), .A2(n7478), .ZN(n7685) );
  INV_X1 U8684 ( .A(n7696), .ZN(n7488) );
  NAND2_X1 U8685 ( .A1(n7488), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7479) );
  AND2_X1 U8686 ( .A1(n7685), .A2(n7479), .ZN(n10682) );
  NAND2_X1 U8687 ( .A1(n10679), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7480) );
  OAI21_X1 U8688 ( .B1(n10679), .B2(P2_REG1_REG_2__SCAN_IN), .A(n7480), .ZN(
        n10681) );
  OR2_X1 U8689 ( .A1(n10682), .A2(n10681), .ZN(n10683) );
  AND2_X1 U8690 ( .A1(n10683), .A2(n7480), .ZN(n7483) );
  OR2_X1 U8691 ( .A1(n7499), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7481) );
  NAND2_X1 U8692 ( .A1(n7499), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U8693 ( .A1(n7481), .A2(n7503), .ZN(n7482) );
  NOR2_X1 U8694 ( .A1(n7483), .A2(n7482), .ZN(n7501) );
  AOI21_X1 U8695 ( .B1(n7483), .B2(n7482), .A(n7501), .ZN(n7484) );
  NAND2_X1 U8696 ( .A1(n10684), .A2(n7484), .ZN(n7486) );
  NAND2_X1 U8697 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n7485) );
  OAI211_X1 U8698 ( .C1(n8373), .C2(n7487), .A(n7486), .B(n7485), .ZN(n7498)
         );
  XNOR2_X1 U8699 ( .A(n7696), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n7693) );
  AND2_X1 U8700 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7692) );
  NAND2_X1 U8701 ( .A1(n7693), .A2(n7692), .ZN(n7691) );
  NAND2_X1 U8702 ( .A1(n7488), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7489) );
  AND2_X1 U8703 ( .A1(n7691), .A2(n7489), .ZN(n10676) );
  NAND2_X1 U8704 ( .A1(n10679), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7490) );
  OAI21_X1 U8705 ( .B1(n10679), .B2(P2_REG2_REG_2__SCAN_IN), .A(n7490), .ZN(
        n10675) );
  OR2_X1 U8706 ( .A1(n10676), .A2(n10675), .ZN(n10678) );
  INV_X1 U8707 ( .A(n10678), .ZN(n7491) );
  AOI21_X1 U8708 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10679), .A(n7491), .ZN(
        n7496) );
  NAND2_X1 U8709 ( .A1(n7499), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7492) );
  OAI21_X1 U8710 ( .B1(n7499), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7492), .ZN(
        n7495) );
  NOR2_X1 U8711 ( .A1(n7496), .A2(n7495), .ZN(n7518) );
  NOR2_X1 U8712 ( .A1(n5940), .A2(n5941), .ZN(n7493) );
  AOI211_X1 U8713 ( .C1(n7496), .C2(n7495), .A(n7518), .B(n10689), .ZN(n7497)
         );
  AOI211_X1 U8714 ( .C1(n10680), .C2(n7499), .A(n7498), .B(n7497), .ZN(n7500)
         );
  INV_X1 U8715 ( .A(n7500), .ZN(P2_U3248) );
  INV_X1 U8716 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7517) );
  MUX2_X1 U8717 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6038), .S(n7608), .Z(n7604)
         );
  INV_X1 U8718 ( .A(n7501), .ZN(n7502) );
  NAND2_X1 U8719 ( .A1(n7503), .A2(n7502), .ZN(n7603) );
  NAND2_X1 U8720 ( .A1(n7604), .A2(n7603), .ZN(n7602) );
  NAND2_X1 U8721 ( .A1(n7608), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U8722 ( .A1(n7602), .A2(n7504), .ZN(n7539) );
  MUX2_X1 U8723 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6046), .S(n7545), .Z(n7540)
         );
  NAND2_X1 U8724 ( .A1(n7539), .A2(n7540), .ZN(n7538) );
  NAND2_X1 U8725 ( .A1(n7545), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7505) );
  NAND2_X1 U8726 ( .A1(n7538), .A2(n7505), .ZN(n7565) );
  MUX2_X1 U8727 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6057), .S(n7571), .Z(n7566)
         );
  NAND2_X1 U8728 ( .A1(n7565), .A2(n7566), .ZN(n7564) );
  NAND2_X1 U8729 ( .A1(n7571), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7506) );
  NAND2_X1 U8730 ( .A1(n7564), .A2(n7506), .ZN(n7578) );
  MUX2_X1 U8731 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6068), .S(n7583), .Z(n7579)
         );
  NAND2_X1 U8732 ( .A1(n7578), .A2(n7579), .ZN(n7577) );
  NAND2_X1 U8733 ( .A1(n7583), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U8734 ( .A1(n7577), .A2(n7507), .ZN(n7552) );
  MUX2_X1 U8735 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6078), .S(n7558), .Z(n7553)
         );
  NAND2_X1 U8736 ( .A1(n7552), .A2(n7553), .ZN(n7551) );
  NAND2_X1 U8737 ( .A1(n7558), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7508) );
  NAND2_X1 U8738 ( .A1(n7551), .A2(n7508), .ZN(n7590) );
  MUX2_X1 U8739 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6088), .S(n7596), .Z(n7591)
         );
  NAND2_X1 U8740 ( .A1(n7590), .A2(n7591), .ZN(n7589) );
  NAND2_X1 U8741 ( .A1(n7596), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7509) );
  AND2_X1 U8742 ( .A1(n7589), .A2(n7509), .ZN(n7512) );
  MUX2_X1 U8743 ( .A(n7510), .B(P2_REG1_REG_10__SCAN_IN), .S(n7629), .Z(n7511)
         );
  NOR2_X1 U8744 ( .A1(n7512), .A2(n7511), .ZN(n7616) );
  INV_X1 U8745 ( .A(n7616), .ZN(n7514) );
  NAND2_X1 U8746 ( .A1(n7512), .A2(n7511), .ZN(n7513) );
  NAND3_X1 U8747 ( .A1(n10684), .A2(n7514), .A3(n7513), .ZN(n7516) );
  NAND2_X1 U8748 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7515) );
  OAI211_X1 U8749 ( .C1(n8373), .C2(n7517), .A(n7516), .B(n7515), .ZN(n7536)
         );
  INV_X1 U8750 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8197) );
  INV_X1 U8751 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7522) );
  MUX2_X1 U8752 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7522), .S(n7608), .Z(n7611)
         );
  INV_X1 U8753 ( .A(n7518), .ZN(n7519) );
  OAI21_X1 U8754 ( .B1(n7521), .B2(n7520), .A(n7519), .ZN(n7610) );
  NAND2_X1 U8755 ( .A1(n7611), .A2(n7610), .ZN(n7609) );
  OAI21_X1 U8756 ( .B1(n7523), .B2(n7522), .A(n7609), .ZN(n7547) );
  MUX2_X1 U8757 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7525), .S(n7545), .Z(n7548)
         );
  NAND2_X1 U8758 ( .A1(n7547), .A2(n7548), .ZN(n7546) );
  OAI21_X1 U8759 ( .B1(n7525), .B2(n7524), .A(n7546), .ZN(n7573) );
  MUX2_X1 U8760 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7526), .S(n7571), .Z(n7574)
         );
  NAND2_X1 U8761 ( .A1(n7573), .A2(n7574), .ZN(n7572) );
  OAI21_X1 U8762 ( .B1(n7527), .B2(n7526), .A(n7572), .ZN(n7585) );
  MUX2_X1 U8763 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7529), .S(n7583), .Z(n7586)
         );
  NAND2_X1 U8764 ( .A1(n7585), .A2(n7586), .ZN(n7584) );
  OAI21_X1 U8765 ( .B1(n7529), .B2(n7528), .A(n7584), .ZN(n7560) );
  XNOR2_X1 U8766 ( .A(n7558), .B(n8197), .ZN(n7561) );
  NAND2_X1 U8767 ( .A1(n7560), .A2(n7561), .ZN(n7559) );
  OAI21_X1 U8768 ( .B1(n8197), .B2(n7530), .A(n7559), .ZN(n7598) );
  MUX2_X1 U8769 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8294), .S(n7596), .Z(n7599)
         );
  NAND2_X1 U8770 ( .A1(n7598), .A2(n7599), .ZN(n7597) );
  INV_X1 U8771 ( .A(n7597), .ZN(n7531) );
  AOI21_X1 U8772 ( .B1(n7596), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7531), .ZN(
        n7534) );
  NAND2_X1 U8773 ( .A1(n7629), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7532) );
  OAI21_X1 U8774 ( .B1(n7629), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7532), .ZN(
        n7533) );
  NOR2_X1 U8775 ( .A1(n7534), .A2(n7533), .ZN(n7628) );
  AOI211_X1 U8776 ( .C1(n7534), .C2(n7533), .A(n7628), .B(n10689), .ZN(n7535)
         );
  AOI211_X1 U8777 ( .C1(n10680), .C2(n7629), .A(n7536), .B(n7535), .ZN(n7537)
         );
  INV_X1 U8778 ( .A(n7537), .ZN(P2_U3255) );
  OAI21_X1 U8779 ( .B1(n7540), .B2(n7539), .A(n7538), .ZN(n7541) );
  NOR2_X1 U8780 ( .A1(n9422), .A2(n7541), .ZN(n7544) );
  INV_X1 U8781 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7542) );
  NAND2_X1 U8782 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7732) );
  OAI21_X1 U8783 ( .B1(n8373), .B2(n7542), .A(n7732), .ZN(n7543) );
  AOI211_X1 U8784 ( .C1(n10680), .C2(n7545), .A(n7544), .B(n7543), .ZN(n7550)
         );
  INV_X1 U8785 ( .A(n10689), .ZN(n10665) );
  OAI211_X1 U8786 ( .C1(n7548), .C2(n7547), .A(n10665), .B(n7546), .ZN(n7549)
         );
  NAND2_X1 U8787 ( .A1(n7550), .A2(n7549), .ZN(P2_U3250) );
  OAI21_X1 U8788 ( .B1(n7553), .B2(n7552), .A(n7551), .ZN(n7554) );
  NOR2_X1 U8789 ( .A1(n9422), .A2(n7554), .ZN(n7557) );
  INV_X1 U8790 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U8791 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7555) );
  OAI21_X1 U8792 ( .B1(n8373), .B2(n10586), .A(n7555), .ZN(n7556) );
  AOI211_X1 U8793 ( .C1(n10680), .C2(n7558), .A(n7557), .B(n7556), .ZN(n7563)
         );
  OAI211_X1 U8794 ( .C1(n7561), .C2(n7560), .A(n10665), .B(n7559), .ZN(n7562)
         );
  NAND2_X1 U8795 ( .A1(n7563), .A2(n7562), .ZN(P2_U3253) );
  OAI21_X1 U8796 ( .B1(n7566), .B2(n7565), .A(n7564), .ZN(n7567) );
  NOR2_X1 U8797 ( .A1(n9422), .A2(n7567), .ZN(n7570) );
  INV_X1 U8798 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7568) );
  NAND2_X1 U8799 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7819) );
  OAI21_X1 U8800 ( .B1(n8373), .B2(n7568), .A(n7819), .ZN(n7569) );
  AOI211_X1 U8801 ( .C1(n10680), .C2(n7571), .A(n7570), .B(n7569), .ZN(n7576)
         );
  OAI211_X1 U8802 ( .C1(n7574), .C2(n7573), .A(n10665), .B(n7572), .ZN(n7575)
         );
  NAND2_X1 U8803 ( .A1(n7576), .A2(n7575), .ZN(P2_U3251) );
  OAI21_X1 U8804 ( .B1(n7579), .B2(n7578), .A(n7577), .ZN(n7580) );
  NOR2_X1 U8805 ( .A1(n9422), .A2(n7580), .ZN(n7582) );
  INV_X1 U8806 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10581) );
  NAND2_X1 U8807 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7873) );
  OAI21_X1 U8808 ( .B1(n8373), .B2(n10581), .A(n7873), .ZN(n7581) );
  AOI211_X1 U8809 ( .C1(n10680), .C2(n7583), .A(n7582), .B(n7581), .ZN(n7588)
         );
  OAI211_X1 U8810 ( .C1(n7586), .C2(n7585), .A(n10665), .B(n7584), .ZN(n7587)
         );
  NAND2_X1 U8811 ( .A1(n7588), .A2(n7587), .ZN(P2_U3252) );
  OAI21_X1 U8812 ( .B1(n7591), .B2(n7590), .A(n7589), .ZN(n7592) );
  NOR2_X1 U8813 ( .A1(n9422), .A2(n7592), .ZN(n7595) );
  INV_X1 U8814 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U8815 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8097) );
  OAI21_X1 U8816 ( .B1(n8373), .B2(n7593), .A(n8097), .ZN(n7594) );
  AOI211_X1 U8817 ( .C1(n10680), .C2(n7596), .A(n7595), .B(n7594), .ZN(n7601)
         );
  OAI211_X1 U8818 ( .C1(n7599), .C2(n7598), .A(n10665), .B(n7597), .ZN(n7600)
         );
  NAND2_X1 U8819 ( .A1(n7601), .A2(n7600), .ZN(P2_U3254) );
  INV_X1 U8820 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7606) );
  OAI211_X1 U8821 ( .C1(n7604), .C2(n7603), .A(n10684), .B(n7602), .ZN(n7605)
         );
  NAND2_X1 U8822 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7708) );
  OAI211_X1 U8823 ( .C1(n8373), .C2(n7606), .A(n7605), .B(n7708), .ZN(n7607)
         );
  AOI21_X1 U8824 ( .B1(n7608), .B2(n10680), .A(n7607), .ZN(n7613) );
  OAI211_X1 U8825 ( .C1(n7611), .C2(n7610), .A(n10665), .B(n7609), .ZN(n7612)
         );
  NAND2_X1 U8826 ( .A1(n7613), .A2(n7612), .ZN(P2_U3249) );
  INV_X1 U8827 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7623) );
  MUX2_X1 U8828 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n7614), .S(n7723), .Z(n7620)
         );
  OR2_X1 U8829 ( .A1(n7625), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7618) );
  MUX2_X1 U8830 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7615), .S(n7625), .Z(n7665)
         );
  AOI21_X1 U8831 ( .B1(n7629), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7616), .ZN(
        n7679) );
  MUX2_X1 U8832 ( .A(n7617), .B(P2_REG1_REG_11__SCAN_IN), .S(n7630), .Z(n7678)
         );
  NOR2_X1 U8833 ( .A1(n7679), .A2(n7678), .ZN(n7677) );
  AOI21_X1 U8834 ( .B1(n7630), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7677), .ZN(
        n7666) );
  NAND2_X1 U8835 ( .A1(n7665), .A2(n7666), .ZN(n7664) );
  NAND2_X1 U8836 ( .A1(n7618), .A2(n7664), .ZN(n7619) );
  NAND2_X1 U8837 ( .A1(n7620), .A2(n7619), .ZN(n7715) );
  OAI21_X1 U8838 ( .B1(n7620), .B2(n7619), .A(n7715), .ZN(n7621) );
  NAND2_X1 U8839 ( .A1(n10684), .A2(n7621), .ZN(n7622) );
  NAND2_X1 U8840 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8529) );
  OAI211_X1 U8841 ( .C1(n8373), .C2(n7623), .A(n7622), .B(n8529), .ZN(n7624)
         );
  AOI21_X1 U8842 ( .B1(n7723), .B2(n10680), .A(n7624), .ZN(n7636) );
  MUX2_X1 U8843 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n8570), .S(n7723), .Z(n7633)
         );
  OR2_X1 U8844 ( .A1(n7625), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7631) );
  MUX2_X1 U8845 ( .A(n8509), .B(P2_REG2_REG_12__SCAN_IN), .S(n7625), .Z(n7626)
         );
  INV_X1 U8846 ( .A(n7626), .ZN(n7661) );
  NOR2_X1 U8847 ( .A1(n7630), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7627) );
  AOI21_X1 U8848 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n7630), .A(n7627), .ZN(
        n7675) );
  AOI21_X1 U8849 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7629), .A(n7628), .ZN(
        n7674) );
  NAND2_X1 U8850 ( .A1(n7675), .A2(n7674), .ZN(n7673) );
  OAI21_X1 U8851 ( .B1(n7630), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7673), .ZN(
        n7662) );
  NAND2_X1 U8852 ( .A1(n7661), .A2(n7662), .ZN(n7660) );
  NAND2_X1 U8853 ( .A1(n7631), .A2(n7660), .ZN(n7632) );
  NAND2_X1 U8854 ( .A1(n7633), .A2(n7632), .ZN(n7724) );
  OAI21_X1 U8855 ( .B1(n7633), .B2(n7632), .A(n7724), .ZN(n7634) );
  NAND2_X1 U8856 ( .A1(n10665), .A2(n7634), .ZN(n7635) );
  NAND2_X1 U8857 ( .A1(n7636), .A2(n7635), .ZN(P2_U3258) );
  INV_X1 U8858 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7638) );
  OAI222_X1 U8859 ( .A1(n8855), .A2(n7638), .B1(n10541), .B2(n7637), .C1(
        P1_U3084), .C2(n7804), .ZN(P1_U3339) );
  AOI21_X1 U8860 ( .B1(n7641), .B2(n7640), .A(n7639), .ZN(n7642) );
  OAI22_X1 U8861 ( .A1(n7643), .A2(n10249), .B1(n10651), .B2(n7642), .ZN(n7649) );
  XOR2_X1 U8862 ( .A(n7645), .B(n7644), .Z(n7647) );
  AND2_X1 U8863 ( .A1(n5013), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7892) );
  AOI21_X1 U8864 ( .B1(n10648), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n7892), .ZN(
        n7646) );
  OAI21_X1 U8865 ( .B1(n10254), .B2(n7647), .A(n7646), .ZN(n7648) );
  OR3_X1 U8866 ( .A1(n7650), .A2(n7649), .A3(n7648), .ZN(P1_U3245) );
  NAND2_X1 U8867 ( .A1(n7836), .A2(n7654), .ZN(n7825) );
  NAND2_X1 U8868 ( .A1(n7828), .A2(n7825), .ZN(n10152) );
  AND2_X1 U8869 ( .A1(n7651), .A2(n10694), .ZN(n7827) );
  XNOR2_X1 U8870 ( .A(n10152), .B(n7827), .ZN(n7748) );
  NAND2_X1 U8871 ( .A1(n10737), .A2(n10740), .ZN(n8848) );
  NAND2_X1 U8872 ( .A1(n10047), .A2(n8799), .ZN(n7930) );
  OAI211_X1 U8873 ( .C1(n10047), .C2(n8799), .A(n10973), .B(n7930), .ZN(n7738)
         );
  NAND2_X1 U8874 ( .A1(n7830), .A2(n10942), .ZN(n7739) );
  OAI211_X1 U8875 ( .C1(n10047), .C2(n10970), .A(n7738), .B(n7739), .ZN(n7658)
         );
  XOR2_X1 U8876 ( .A(n10152), .B(n7835), .Z(n7657) );
  OR2_X1 U8877 ( .A1(n8538), .A2(n10740), .ZN(n7655) );
  NAND2_X1 U8878 ( .A1(n10049), .A2(n10115), .ZN(n10016) );
  INV_X1 U8879 ( .A(n7651), .ZN(n7656) );
  OAI22_X1 U8880 ( .A1(n7657), .A2(n10873), .B1(n7656), .B2(n10401), .ZN(n7741) );
  AOI211_X1 U8881 ( .C1(n7748), .C2(n10952), .A(n7658), .B(n7741), .ZN(n7751)
         );
  NAND2_X1 U8882 ( .A1(n10975), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7659) );
  OAI21_X1 U8883 ( .B1(n7751), .B2(n10975), .A(n7659), .ZN(P1_U3524) );
  OAI21_X1 U8884 ( .B1(n7662), .B2(n7661), .A(n7660), .ZN(n7663) );
  NAND2_X1 U8885 ( .A1(n7663), .A2(n10665), .ZN(n7671) );
  OAI21_X1 U8886 ( .B1(n7666), .B2(n7665), .A(n7664), .ZN(n7669) );
  INV_X1 U8887 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U8888 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8439) );
  OAI21_X1 U8889 ( .B1(n8373), .B2(n7667), .A(n8439), .ZN(n7668) );
  AOI21_X1 U8890 ( .B1(n10684), .B2(n7669), .A(n7668), .ZN(n7670) );
  OAI211_X1 U8891 ( .C1(n10668), .C2(n7672), .A(n7671), .B(n7670), .ZN(
        P2_U3257) );
  OAI21_X1 U8892 ( .B1(n7675), .B2(n7674), .A(n7673), .ZN(n7676) );
  NAND2_X1 U8893 ( .A1(n7676), .A2(n10665), .ZN(n7682) );
  NOR2_X1 U8894 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8959), .ZN(n8264) );
  AOI211_X1 U8895 ( .C1(n7679), .C2(n7678), .A(n7677), .B(n9422), .ZN(n7680)
         );
  AOI211_X1 U8896 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n10674), .A(n8264), .B(
        n7680), .ZN(n7681) );
  OAI211_X1 U8897 ( .C1(n10668), .C2(n7683), .A(n7682), .B(n7681), .ZN(
        P2_U3256) );
  INV_X1 U8898 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8103) );
  NOR2_X1 U8899 ( .A1(n8103), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7690) );
  INV_X1 U8900 ( .A(n7684), .ZN(n7687) );
  INV_X1 U8901 ( .A(n7685), .ZN(n7686) );
  AOI211_X1 U8902 ( .C1(n7688), .C2(n7687), .A(n7686), .B(n9422), .ZN(n7689)
         );
  AOI211_X1 U8903 ( .C1(P2_ADDR_REG_1__SCAN_IN), .C2(n10674), .A(n7690), .B(
        n7689), .ZN(n7695) );
  OAI211_X1 U8904 ( .C1(n7693), .C2(n7692), .A(n10665), .B(n7691), .ZN(n7694)
         );
  OAI211_X1 U8905 ( .C1(n10668), .C2(n7696), .A(n7695), .B(n7694), .ZN(
        P2_U3246) );
  XNOR2_X1 U8906 ( .A(n7697), .B(n7698), .ZN(n7699) );
  NAND2_X1 U8907 ( .A1(n7699), .A2(n9893), .ZN(n7704) );
  INV_X1 U8908 ( .A(n7830), .ZN(n10054) );
  INV_X1 U8909 ( .A(n9923), .ZN(n7700) );
  OAI22_X1 U8910 ( .A1(n10054), .A2(n7700), .B1(n9903), .B2(n7832), .ZN(n7701)
         );
  AOI211_X1 U8911 ( .C1(n9906), .C2(n10209), .A(n7702), .B(n7701), .ZN(n7703)
         );
  OAI211_X1 U8912 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9926), .A(n7704), .B(
        n7703), .ZN(P1_U3216) );
  AOI21_X1 U8913 ( .B1(n7707), .B2(n7706), .A(n7705), .ZN(n7713) );
  INV_X1 U8914 ( .A(n8455), .ZN(n7820) );
  OAI21_X1 U8915 ( .B1(n9362), .B2(n7820), .A(n7708), .ZN(n7711) );
  INV_X1 U8916 ( .A(n9396), .ZN(n7709) );
  OAI22_X1 U8917 ( .A1(n9365), .A2(n7709), .B1(n9363), .B2(n8216), .ZN(n7710)
         );
  AOI211_X1 U8918 ( .C1(n9379), .C2(n8218), .A(n7711), .B(n7710), .ZN(n7712)
         );
  OAI21_X1 U8919 ( .B1(n7713), .B2(n9381), .A(n7712), .ZN(P2_U3232) );
  INV_X1 U8920 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7721) );
  MUX2_X1 U8921 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7714), .S(n7972), .Z(n7718)
         );
  OR2_X1 U8922 ( .A1(n7723), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U8923 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  NAND2_X1 U8924 ( .A1(n7718), .A2(n7717), .ZN(n7971) );
  OAI21_X1 U8925 ( .B1(n7718), .B2(n7717), .A(n7971), .ZN(n7719) );
  NAND2_X1 U8926 ( .A1(n10684), .A2(n7719), .ZN(n7720) );
  NAND2_X1 U8927 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8588) );
  OAI211_X1 U8928 ( .C1(n8373), .C2(n7721), .A(n7720), .B(n8588), .ZN(n7722)
         );
  AOI21_X1 U8929 ( .B1(n7972), .B2(n10680), .A(n7722), .ZN(n7730) );
  MUX2_X1 U8930 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n8612), .S(n7972), .Z(n7727)
         );
  OR2_X1 U8931 ( .A1(n7723), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U8932 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  NAND2_X1 U8933 ( .A1(n7727), .A2(n7726), .ZN(n7968) );
  OAI21_X1 U8934 ( .B1(n7727), .B2(n7726), .A(n7968), .ZN(n7728) );
  NAND2_X1 U8935 ( .A1(n10665), .A2(n7728), .ZN(n7729) );
  NAND2_X1 U8936 ( .A1(n7730), .A2(n7729), .ZN(P2_U3259) );
  XNOR2_X1 U8937 ( .A(n5093), .B(n7731), .ZN(n7737) );
  INV_X1 U8938 ( .A(n7732), .ZN(n7734) );
  OAI22_X1 U8939 ( .A1(n9365), .A2(n7791), .B1(n9363), .B2(n10752), .ZN(n7733)
         );
  AOI211_X1 U8940 ( .C1(n9334), .C2(n9394), .A(n7734), .B(n7733), .ZN(n7736)
         );
  NAND2_X1 U8941 ( .A1(n9379), .A2(n10753), .ZN(n7735) );
  OAI211_X1 U8942 ( .C1(n7737), .C2(n9381), .A(n7736), .B(n7735), .ZN(P2_U3229) );
  INV_X1 U8943 ( .A(n7738), .ZN(n7743) );
  INV_X1 U8944 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7740) );
  OAI21_X1 U8945 ( .B1(n10819), .B2(n7740), .A(n7739), .ZN(n7742) );
  AOI211_X1 U8946 ( .C1(n7743), .C2(n10740), .A(n7742), .B(n7741), .ZN(n7750)
         );
  NAND3_X1 U8947 ( .A1(n7746), .A2(n7745), .A3(n7744), .ZN(n8252) );
  INV_X1 U8948 ( .A(n10406), .ZN(n10964) );
  OAI22_X1 U8949 ( .A1(n10792), .A2(n10047), .B1(n6550), .B2(n10822), .ZN(
        n7747) );
  AOI21_X1 U8950 ( .B1(n7748), .B2(n10964), .A(n7747), .ZN(n7749) );
  OAI21_X1 U8951 ( .B1(n7750), .B2(n10969), .A(n7749), .ZN(P1_U3290) );
  INV_X1 U8952 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7753) );
  OR2_X1 U8953 ( .A1(n7751), .A2(n10978), .ZN(n7752) );
  OAI21_X1 U8954 ( .B1(n10981), .B2(n7753), .A(n7752), .ZN(P1_U3457) );
  NAND2_X1 U8955 ( .A1(n7866), .A2(n7867), .ZN(n7865) );
  OR2_X1 U8956 ( .A1(n7404), .A2(n8108), .ZN(n7757) );
  NAND2_X1 U8957 ( .A1(n7865), .A2(n7757), .ZN(n8053) );
  NAND2_X1 U8958 ( .A1(n8053), .A2(n8052), .ZN(n8055) );
  OR2_X1 U8959 ( .A1(n9397), .A2(n8061), .ZN(n7758) );
  NAND2_X1 U8960 ( .A1(n8055), .A2(n7758), .ZN(n7759) );
  NAND2_X1 U8961 ( .A1(n7759), .A2(n7765), .ZN(n7914) );
  OAI21_X1 U8962 ( .B1(n7759), .B2(n7765), .A(n7914), .ZN(n7771) );
  INV_X1 U8963 ( .A(n7771), .ZN(n8357) );
  INV_X1 U8964 ( .A(n10836), .ZN(n8316) );
  NAND2_X1 U8965 ( .A1(n6004), .A2(n7760), .ZN(n8042) );
  XNOR2_X1 U8966 ( .A(n8042), .B(n7761), .ZN(n7762) );
  NAND2_X1 U8967 ( .A1(n7762), .A2(n9407), .ZN(n8393) );
  INV_X1 U8968 ( .A(n8393), .ZN(n8293) );
  OAI22_X1 U8969 ( .A1(n7763), .A2(n9641), .B1(n7791), .B2(n9565), .ZN(n7770)
         );
  XOR2_X1 U8970 ( .A(n7765), .B(n7764), .Z(n7768) );
  NOR2_X1 U8971 ( .A1(n7768), .A2(n9561), .ZN(n7769) );
  AOI211_X1 U8972 ( .C1(n8293), .C2(n7771), .A(n7770), .B(n7769), .ZN(n8362)
         );
  AOI21_X1 U8973 ( .B1(n7912), .B2(n8064), .A(n8209), .ZN(n8360) );
  AOI22_X1 U8974 ( .A1(n8360), .A2(n9746), .B1(n9745), .B2(n7912), .ZN(n7772)
         );
  OAI211_X1 U8975 ( .C1(n8357), .C2(n8316), .A(n8362), .B(n7772), .ZN(n8074)
         );
  NAND2_X1 U8976 ( .A1(n8074), .A2(n10923), .ZN(n7773) );
  OAI21_X1 U8977 ( .B1(n10923), .B2(n6026), .A(n7773), .ZN(P2_U3523) );
  OAI211_X1 U8978 ( .C1(n7776), .C2(n7775), .A(n10216), .B(n7774), .ZN(n7788)
         );
  INV_X1 U8979 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7785) );
  OAI21_X1 U8980 ( .B1(n7779), .B2(n7778), .A(n7777), .ZN(n7781) );
  AOI22_X1 U8981 ( .A1(n10649), .A2(n7781), .B1(n10657), .B2(n7780), .ZN(n7783) );
  AND2_X1 U8982 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8669) );
  INV_X1 U8983 ( .A(n8669), .ZN(n7782) );
  OAI211_X1 U8984 ( .C1(n7785), .C2(n7784), .A(n7783), .B(n7782), .ZN(n7786)
         );
  INV_X1 U8985 ( .A(n7786), .ZN(n7787) );
  NAND2_X1 U8986 ( .A1(n7788), .A2(n7787), .ZN(P1_U3254) );
  XNOR2_X1 U8987 ( .A(n7790), .B(n7789), .ZN(n7795) );
  MUX2_X1 U8988 ( .A(n9374), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n7793) );
  OAI22_X1 U8989 ( .A1(n9362), .A2(n7791), .B1(n8356), .B2(n9358), .ZN(n7792)
         );
  AOI211_X1 U8990 ( .C1(n9335), .C2(n9397), .A(n7793), .B(n7792), .ZN(n7794)
         );
  OAI21_X1 U8991 ( .B1(n7795), .B2(n9381), .A(n7794), .ZN(P2_U3220) );
  AOI21_X1 U8992 ( .B1(n7804), .B2(n8677), .A(n7796), .ZN(n7798) );
  XNOR2_X1 U8993 ( .A(n7798), .B(n7797), .ZN(n7808) );
  OAI21_X1 U8994 ( .B1(n7801), .B2(n7800), .A(n7799), .ZN(n7806) );
  NOR2_X1 U8995 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7802), .ZN(n9805) );
  AOI21_X1 U8996 ( .B1(n10648), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n9805), .ZN(
        n7803) );
  OAI21_X1 U8997 ( .B1(n7804), .B2(n10249), .A(n7803), .ZN(n7805) );
  AOI21_X1 U8998 ( .B1(n7806), .B2(n10649), .A(n7805), .ZN(n7807) );
  OAI21_X1 U8999 ( .B1(n7808), .B2(n10651), .A(n7807), .ZN(P1_U3255) );
  NAND2_X1 U9000 ( .A1(n7809), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U9001 ( .A1(n6655), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7813) );
  OR2_X1 U9002 ( .A1(n7117), .A2(n8786), .ZN(n7812) );
  NAND2_X1 U9003 ( .A1(n7810), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7811) );
  NAND4_X1 U9004 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n8769)
         );
  NAND2_X1 U9005 ( .A1(n8769), .A2(P1_U4006), .ZN(n7815) );
  OAI21_X1 U9006 ( .B1(n5754), .B2(P1_U4006), .A(n7815), .ZN(P1_U3584) );
  INV_X1 U9007 ( .A(n8450), .ZN(n10768) );
  NAND2_X1 U9008 ( .A1(n7818), .A2(n9352), .ZN(n7824) );
  INV_X1 U9009 ( .A(n7819), .ZN(n7822) );
  OAI22_X1 U9010 ( .A1(n9365), .A2(n7820), .B1(n9363), .B2(n8448), .ZN(n7821)
         );
  AOI211_X1 U9011 ( .C1(n9334), .C2(n9393), .A(n7822), .B(n7821), .ZN(n7823)
         );
  OAI211_X1 U9012 ( .C1(n10768), .C2(n9358), .A(n7824), .B(n7823), .ZN(
        P2_U3241) );
  INV_X1 U9013 ( .A(n7825), .ZN(n7826) );
  AOI21_X1 U9014 ( .B1(n7828), .B2(n7827), .A(n7826), .ZN(n7926) );
  XNOR2_X1 U9015 ( .A(n7830), .B(n10708), .ZN(n10154) );
  NAND2_X1 U9016 ( .A1(n7926), .A2(n10154), .ZN(n7925) );
  NAND2_X1 U9017 ( .A1(n10054), .A2(n10708), .ZN(n7831) );
  INV_X1 U9018 ( .A(n10210), .ZN(n7982) );
  NAND2_X1 U9019 ( .A1(n10119), .A2(n8021), .ZN(n7833) );
  OAI21_X1 U9020 ( .B1(n7834), .B2(n7833), .A(n7984), .ZN(n7902) );
  OAI22_X1 U9021 ( .A1(n10054), .A2(n10401), .B1(n7985), .B2(n10403), .ZN(
        n7842) );
  NAND2_X1 U9022 ( .A1(n10152), .A2(n7835), .ZN(n7838) );
  OR2_X1 U9023 ( .A1(n7836), .A2(n10047), .ZN(n7837) );
  NAND2_X1 U9024 ( .A1(n7838), .A2(n7837), .ZN(n7924) );
  INV_X1 U9025 ( .A(n10154), .ZN(n7839) );
  NAND2_X1 U9026 ( .A1(n10054), .A2(n10053), .ZN(n10052) );
  XNOR2_X1 U9027 ( .A(n7833), .B(n10124), .ZN(n7840) );
  NOR2_X1 U9028 ( .A1(n7840), .A2(n10873), .ZN(n7841) );
  AOI211_X1 U9029 ( .C1(n10876), .C2(n7902), .A(n7842), .B(n7841), .ZN(n7906)
         );
  AND2_X1 U9030 ( .A1(n7843), .A2(n10366), .ZN(n7844) );
  NAND2_X1 U9031 ( .A1(n10822), .A2(n7844), .ZN(n10385) );
  INV_X1 U9032 ( .A(n10385), .ZN(n10887) );
  OR2_X1 U9033 ( .A1(n7930), .A2(n10053), .ZN(n7932) );
  AOI21_X1 U9034 ( .B1(n7903), .B2(n7932), .A(n7988), .ZN(n7904) );
  AND2_X1 U9035 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  NAND2_X1 U9036 ( .A1(n7904), .A2(n10786), .ZN(n7850) );
  INV_X1 U9037 ( .A(n10819), .ZN(n10957) );
  AOI22_X1 U9038 ( .A1(n10969), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10957), .B2(
        n7848), .ZN(n7849) );
  OAI211_X1 U9039 ( .C1(n7832), .C2(n10792), .A(n7850), .B(n7849), .ZN(n7851)
         );
  AOI21_X1 U9040 ( .B1(n10887), .B2(n7902), .A(n7851), .ZN(n7852) );
  OAI21_X1 U9041 ( .B1(n7906), .B2(n10969), .A(n7852), .ZN(P1_U3288) );
  INV_X1 U9042 ( .A(n7853), .ZN(n7855) );
  OAI222_X1 U9043 ( .A1(n8831), .A2(n7854), .B1(n8691), .B2(n7855), .C1(
        P2_U3152), .C2(n8185), .ZN(P2_U3343) );
  OAI222_X1 U9044 ( .A1(n8118), .A2(n5013), .B1(n10541), .B2(n7855), .C1(n9210), .C2(n8855), .ZN(P1_U3338) );
  INV_X1 U9045 ( .A(n7856), .ZN(n7859) );
  OAI222_X1 U9046 ( .A1(n8691), .A2(n7859), .B1(n8364), .B2(P2_U3152), .C1(
        n7857), .C2(n8831), .ZN(P2_U3342) );
  INV_X1 U9047 ( .A(n7858), .ZN(n8277) );
  OAI222_X1 U9048 ( .A1(n5013), .A2(n8277), .B1(n10541), .B2(n7859), .C1(n9209), .C2(n8855), .ZN(P1_U3337) );
  NAND2_X1 U9049 ( .A1(n10701), .A2(n8108), .ZN(n7860) );
  NAND2_X1 U9050 ( .A1(n8062), .A2(n7860), .ZN(n8104) );
  AOI21_X1 U9051 ( .B1(n7861), .B2(n7867), .A(n9561), .ZN(n7864) );
  AOI21_X1 U9052 ( .B1(n7864), .B2(n7863), .A(n7862), .ZN(n8111) );
  OAI21_X1 U9053 ( .B1(n7867), .B2(n7866), .A(n7865), .ZN(n8107) );
  NAND2_X1 U9054 ( .A1(n8107), .A2(n10921), .ZN(n7868) );
  OAI211_X1 U9055 ( .C1(n10916), .C2(n8104), .A(n8111), .B(n7868), .ZN(n8238)
         );
  NOR2_X1 U9056 ( .A1(n10923), .A2(n6007), .ZN(n7869) );
  AOI21_X1 U9057 ( .B1(n10923), .B2(n8238), .A(n7869), .ZN(n7870) );
  OAI21_X1 U9058 ( .B1(n8240), .B2(n9742), .A(n7870), .ZN(P2_U3521) );
  XNOR2_X1 U9059 ( .A(n7872), .B(n7871), .ZN(n7879) );
  INV_X1 U9060 ( .A(n7873), .ZN(n7876) );
  OAI22_X1 U9061 ( .A1(n9365), .A2(n7874), .B1(n9363), .B2(n8461), .ZN(n7875)
         );
  AOI211_X1 U9062 ( .C1(n9334), .C2(n9392), .A(n7876), .B(n7875), .ZN(n7878)
         );
  NAND2_X1 U9063 ( .A1(n9379), .A2(n8463), .ZN(n7877) );
  OAI211_X1 U9064 ( .C1(n7879), .C2(n9381), .A(n7878), .B(n7877), .ZN(P2_U3215) );
  INV_X1 U9065 ( .A(n7880), .ZN(n7883) );
  AOI22_X1 U9066 ( .A1(n10245), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10539), .ZN(n7881) );
  OAI21_X1 U9067 ( .B1(n7883), .B2(n10541), .A(n7881), .ZN(P1_U3336) );
  AOI22_X1 U9068 ( .A1(n9400), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n7966), .ZN(n7882) );
  OAI21_X1 U9069 ( .B1(n7883), .B2(n8691), .A(n7882), .ZN(P2_U3341) );
  XNOR2_X1 U9070 ( .A(n7885), .B(n7884), .ZN(n7890) );
  OAI22_X1 U9071 ( .A1(n7886), .A2(n9641), .B1(n8172), .B2(n9565), .ZN(n8088)
         );
  AOI22_X1 U9072 ( .A1(n9373), .A2(n8088), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n7887) );
  OAI21_X1 U9073 ( .B1(n9363), .B2(n8196), .A(n7887), .ZN(n7888) );
  AOI21_X1 U9074 ( .B1(n9379), .B2(n8281), .A(n7888), .ZN(n7889) );
  OAI21_X1 U9075 ( .B1(n7890), .B2(n9381), .A(n7889), .ZN(P2_U3223) );
  INV_X1 U9076 ( .A(n7891), .ZN(n7990) );
  INV_X1 U9077 ( .A(n7991), .ZN(n10724) );
  AOI21_X1 U9078 ( .B1(n9906), .B2(n10208), .A(n7892), .ZN(n7894) );
  NAND2_X1 U9079 ( .A1(n9923), .A2(n10210), .ZN(n7893) );
  OAI211_X1 U9080 ( .C1(n10724), .C2(n9903), .A(n7894), .B(n7893), .ZN(n7900)
         );
  INV_X1 U9081 ( .A(n7895), .ZN(n7896) );
  AOI211_X1 U9082 ( .C1(n7898), .C2(n7897), .A(n9931), .B(n7896), .ZN(n7899)
         );
  AOI211_X1 U9083 ( .C1(n7990), .C2(n9900), .A(n7900), .B(n7899), .ZN(n7901)
         );
  INV_X1 U9084 ( .A(n7901), .ZN(P1_U3228) );
  INV_X1 U9085 ( .A(n7902), .ZN(n7907) );
  AOI22_X1 U9086 ( .A1(n7904), .A2(n10973), .B1(n10802), .B2(n7903), .ZN(n7905) );
  OAI211_X1 U9087 ( .C1(n7907), .C2(n10520), .A(n7906), .B(n7905), .ZN(n7909)
         );
  NAND2_X1 U9088 ( .A1(n7909), .A2(n10977), .ZN(n7908) );
  OAI21_X1 U9089 ( .B1(n10977), .B2(n7145), .A(n7908), .ZN(P1_U3526) );
  INV_X1 U9090 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U9091 ( .A1(n7909), .A2(n10981), .ZN(n7910) );
  OAI21_X1 U9092 ( .B1(n10981), .B2(n7911), .A(n7910), .ZN(P1_U3463) );
  OR2_X1 U9093 ( .A1(n9396), .A2(n7912), .ZN(n7913) );
  XNOR2_X1 U9094 ( .A(n7953), .B(n7954), .ZN(n10760) );
  INV_X1 U9095 ( .A(n7916), .ZN(n8447) );
  AOI211_X1 U9096 ( .C1(n10753), .C2(n8211), .A(n10916), .B(n8447), .ZN(n10751) );
  NAND2_X1 U9097 ( .A1(n7917), .A2(n7918), .ZN(n7919) );
  NAND3_X1 U9098 ( .A1(n7920), .A2(n9644), .A3(n7919), .ZN(n7922) );
  AOI22_X1 U9099 ( .A1(n9619), .A2(n9395), .B1(n9394), .B2(n9638), .ZN(n7921)
         );
  NAND2_X1 U9100 ( .A1(n7922), .A2(n7921), .ZN(n10759) );
  AOI211_X1 U9101 ( .C1(n10921), .C2(n10760), .A(n10751), .B(n10759), .ZN(
        n8342) );
  INV_X1 U9102 ( .A(n9742), .ZN(n8432) );
  AOI22_X1 U9103 ( .A1(n8432), .A2(n10753), .B1(n10922), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7923) );
  OAI21_X1 U9104 ( .B1(n8342), .B2(n10922), .A(n7923), .ZN(P2_U3525) );
  XNOR2_X1 U9105 ( .A(n10154), .B(n7924), .ZN(n7929) );
  AOI22_X1 U9106 ( .A1(n10942), .A2(n10210), .B1(n7836), .B2(n10944), .ZN(
        n7928) );
  OAI21_X1 U9107 ( .B1(n7926), .B2(n10154), .A(n7925), .ZN(n10712) );
  NAND2_X1 U9108 ( .A1(n10712), .A2(n10876), .ZN(n7927) );
  OAI211_X1 U9109 ( .C1(n7929), .C2(n10873), .A(n7928), .B(n7927), .ZN(n10710)
         );
  INV_X1 U9110 ( .A(n10710), .ZN(n7939) );
  NAND2_X1 U9111 ( .A1(n7930), .A2(n10053), .ZN(n7931) );
  NAND2_X1 U9112 ( .A1(n7932), .A2(n7931), .ZN(n10709) );
  NOR2_X1 U9113 ( .A1(n10819), .A2(n7933), .ZN(n7935) );
  NOR2_X1 U9114 ( .A1(n10792), .A2(n10708), .ZN(n7934) );
  AOI211_X1 U9115 ( .C1(n10969), .C2(P1_REG2_REG_2__SCAN_IN), .A(n7935), .B(
        n7934), .ZN(n7936) );
  OAI21_X1 U9116 ( .B1(n10429), .B2(n10709), .A(n7936), .ZN(n7937) );
  AOI21_X1 U9117 ( .B1(n10887), .B2(n10712), .A(n7937), .ZN(n7938) );
  OAI21_X1 U9118 ( .B1(n7939), .B2(n10969), .A(n7938), .ZN(P1_U3289) );
  NAND2_X1 U9119 ( .A1(n7945), .A2(n7942), .ZN(n7943) );
  AOI22_X1 U9120 ( .A1(n7941), .A2(n7945), .B1(n7944), .B2(n7943), .ZN(n7951)
         );
  NOR2_X1 U9121 ( .A1(n9903), .A2(n8014), .ZN(n7949) );
  NAND2_X1 U9122 ( .A1(n9923), .A2(n10209), .ZN(n7946) );
  OAI211_X1 U9123 ( .C1(n8243), .C2(n9919), .A(n7947), .B(n7946), .ZN(n7948)
         );
  AOI211_X1 U9124 ( .C1(n10742), .C2(n9900), .A(n7949), .B(n7948), .ZN(n7950)
         );
  OAI21_X1 U9125 ( .B1(n7951), .B2(n9931), .A(n7950), .ZN(P1_U3225) );
  OR2_X1 U9126 ( .A1(n10753), .A2(n8455), .ZN(n7952) );
  NAND2_X1 U9127 ( .A1(n7953), .A2(n7952), .ZN(n7956) );
  NAND2_X1 U9128 ( .A1(n7954), .A2(n10753), .ZN(n7955) );
  NAND2_X1 U9129 ( .A1(n7956), .A2(n7955), .ZN(n8444) );
  NAND2_X1 U9130 ( .A1(n8450), .A2(n9394), .ZN(n7958) );
  XNOR2_X1 U9131 ( .A(n8079), .B(n8078), .ZN(n8469) );
  INV_X1 U9132 ( .A(n8090), .ZN(n7959) );
  OAI21_X1 U9133 ( .B1(n8344), .B2(n8445), .A(n7959), .ZN(n8465) );
  NOR2_X1 U9134 ( .A1(n8465), .A2(n10916), .ZN(n7963) );
  OAI211_X1 U9135 ( .C1(n8078), .C2(n7960), .A(n8082), .B(n9644), .ZN(n7962)
         );
  AOI22_X1 U9136 ( .A1(n9619), .A2(n9394), .B1(n9392), .B2(n9638), .ZN(n7961)
         );
  NAND2_X1 U9137 ( .A1(n7962), .A2(n7961), .ZN(n8466) );
  AOI211_X1 U9138 ( .C1(n8469), .C2(n10921), .A(n7963), .B(n8466), .ZN(n8347)
         );
  AOI22_X1 U9139 ( .A1(n8432), .A2(n8463), .B1(n10922), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7964) );
  OAI21_X1 U9140 ( .B1(n8347), .B2(n10922), .A(n7964), .ZN(P2_U3527) );
  INV_X1 U9141 ( .A(n7965), .ZN(n8033) );
  AOI22_X1 U9142 ( .A1(n9414), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7966), .ZN(n7967) );
  OAI21_X1 U9143 ( .B1(n8033), .B2(n8691), .A(n7967), .ZN(P2_U3340) );
  OAI21_X1 U9144 ( .B1(n7972), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7968), .ZN(
        n8184) );
  INV_X1 U9145 ( .A(n8184), .ZN(n7969) );
  XNOR2_X1 U9146 ( .A(n8185), .B(n7969), .ZN(n7970) );
  NAND2_X1 U9147 ( .A1(n7970), .A2(n8653), .ZN(n8186) );
  OAI21_X1 U9148 ( .B1(n7970), .B2(n8653), .A(n8186), .ZN(n7980) );
  INV_X1 U9149 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7977) );
  OAI21_X1 U9150 ( .B1(n7972), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7971), .ZN(
        n8177) );
  XNOR2_X1 U9151 ( .A(n8185), .B(n8177), .ZN(n7974) );
  NOR2_X1 U9152 ( .A1(n7973), .A2(n7974), .ZN(n8178) );
  AOI21_X1 U9153 ( .B1(n7974), .B2(n7973), .A(n8178), .ZN(n7975) );
  NAND2_X1 U9154 ( .A1(n10684), .A2(n7975), .ZN(n7976) );
  NAND2_X1 U9155 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8642) );
  OAI211_X1 U9156 ( .C1(n8373), .C2(n7977), .A(n7976), .B(n8642), .ZN(n7979)
         );
  NOR2_X1 U9157 ( .A1(n10668), .A2(n8185), .ZN(n7978) );
  AOI211_X1 U9158 ( .C1(n10665), .C2(n7980), .A(n7979), .B(n7978), .ZN(n7981)
         );
  INV_X1 U9159 ( .A(n7981), .ZN(P2_U3260) );
  NAND2_X1 U9160 ( .A1(n7982), .A2(n7832), .ZN(n7983) );
  NAND2_X1 U9161 ( .A1(n7984), .A2(n7983), .ZN(n7986) );
  NAND2_X1 U9162 ( .A1(n10209), .A2(n10724), .ZN(n10122) );
  OR2_X1 U9163 ( .A1(n7986), .A2(n10155), .ZN(n7987) );
  NAND2_X1 U9164 ( .A1(n8013), .A2(n7987), .ZN(n10728) );
  NAND2_X1 U9165 ( .A1(n7988), .A2(n10724), .ZN(n8152) );
  OR2_X1 U9166 ( .A1(n7988), .A2(n10724), .ZN(n7989) );
  NAND2_X1 U9167 ( .A1(n8152), .A2(n7989), .ZN(n10725) );
  AOI22_X1 U9168 ( .A1(n10959), .A2(n7991), .B1(n7990), .B2(n10957), .ZN(n7992) );
  OAI21_X1 U9169 ( .B1(n10725), .B2(n10429), .A(n7992), .ZN(n8000) );
  NAND2_X1 U9170 ( .A1(n10728), .A2(n10876), .ZN(n7998) );
  INV_X1 U9171 ( .A(n10119), .ZN(n7993) );
  NAND2_X1 U9172 ( .A1(n8022), .A2(n8021), .ZN(n7994) );
  XNOR2_X1 U9173 ( .A(n7994), .B(n10155), .ZN(n7995) );
  NAND2_X1 U9174 ( .A1(n7995), .A2(n10947), .ZN(n7997) );
  AOI22_X1 U9175 ( .A1(n10944), .A2(n10210), .B1(n10208), .B2(n10942), .ZN(
        n7996) );
  NAND3_X1 U9176 ( .A1(n7998), .A2(n7997), .A3(n7996), .ZN(n10726) );
  MUX2_X1 U9177 ( .A(n10726), .B(P1_REG2_REG_4__SCAN_IN), .S(n10969), .Z(n7999) );
  AOI211_X1 U9178 ( .C1(n10887), .C2(n10728), .A(n8000), .B(n7999), .ZN(n8001)
         );
  INV_X1 U9179 ( .A(n8001), .ZN(P1_U3287) );
  NAND2_X1 U9180 ( .A1(n7941), .A2(n8002), .ZN(n8123) );
  OAI21_X1 U9181 ( .B1(n8002), .B2(n7941), .A(n8123), .ZN(n8010) );
  AOI21_X1 U9182 ( .B1(n9906), .B2(n10206), .A(n8003), .ZN(n8008) );
  OR2_X1 U9183 ( .A1(n9903), .A2(n5305), .ZN(n8007) );
  INV_X1 U9184 ( .A(n8141), .ZN(n8004) );
  NAND2_X1 U9185 ( .A1(n9900), .A2(n8004), .ZN(n8006) );
  NAND2_X1 U9186 ( .A1(n9923), .A2(n10208), .ZN(n8005) );
  NAND4_X1 U9187 ( .A1(n8008), .A2(n8007), .A3(n8006), .A4(n8005), .ZN(n8009)
         );
  AOI21_X1 U9188 ( .B1(n8010), .B2(n9893), .A(n8009), .ZN(n8011) );
  INV_X1 U9189 ( .A(n8011), .ZN(P1_U3237) );
  NAND2_X1 U9190 ( .A1(n7985), .A2(n10724), .ZN(n8012) );
  INV_X1 U9191 ( .A(n10208), .ZN(n8136) );
  NAND2_X1 U9192 ( .A1(n8136), .A2(n10744), .ZN(n10125) );
  NAND2_X1 U9193 ( .A1(n10208), .A2(n8014), .ZN(n8023) );
  NAND2_X1 U9194 ( .A1(n10208), .A2(n10744), .ZN(n8016) );
  INV_X1 U9195 ( .A(n8134), .ZN(n8018) );
  NAND2_X1 U9196 ( .A1(n10207), .A2(n5305), .ZN(n9935) );
  NAND2_X1 U9197 ( .A1(n8243), .A2(n5305), .ZN(n8019) );
  NAND2_X1 U9198 ( .A1(n8132), .A2(n8019), .ZN(n8246) );
  INV_X1 U9199 ( .A(n10206), .ZN(n8137) );
  NAND2_X1 U9200 ( .A1(n8137), .A2(n8408), .ZN(n10043) );
  INV_X1 U9201 ( .A(n8408), .ZN(n8256) );
  NAND2_X1 U9202 ( .A1(n10206), .A2(n8256), .ZN(n9939) );
  NAND2_X1 U9203 ( .A1(n10043), .A2(n9939), .ZN(n10161) );
  NAND2_X1 U9204 ( .A1(n8137), .A2(n8256), .ZN(n8020) );
  NAND2_X1 U9205 ( .A1(n10776), .A2(n8335), .ZN(n10065) );
  INV_X1 U9206 ( .A(n8335), .ZN(n8244) );
  NAND2_X1 U9207 ( .A1(n8244), .A2(n8301), .ZN(n10042) );
  NAND2_X1 U9208 ( .A1(n10065), .A2(n10042), .ZN(n9942) );
  OAI21_X1 U9209 ( .B1(n5094), .B2(n9942), .A(n8303), .ZN(n10775) );
  AND2_X1 U9210 ( .A1(n8021), .A2(n10122), .ZN(n10123) );
  AND3_X1 U9211 ( .A1(n10126), .A2(n10125), .A3(n10120), .ZN(n10060) );
  INV_X1 U9212 ( .A(n8023), .ZN(n10127) );
  NAND2_X1 U9213 ( .A1(n10126), .A2(n10127), .ZN(n10058) );
  NAND2_X1 U9214 ( .A1(n10058), .A2(n9935), .ZN(n8024) );
  INV_X1 U9215 ( .A(n10161), .ZN(n8242) );
  NAND2_X1 U9216 ( .A1(n8306), .A2(n10043), .ZN(n8025) );
  XNOR2_X1 U9217 ( .A(n8025), .B(n9942), .ZN(n8026) );
  OAI222_X1 U9218 ( .A1(n10403), .A2(n8304), .B1(n10401), .B2(n8137), .C1(
        n8026), .C2(n10873), .ZN(n10778) );
  OAI21_X1 U9219 ( .B1(n8250), .B2(n10776), .A(n8310), .ZN(n10777) );
  OAI22_X1 U9220 ( .A1(n10822), .A2(n8027), .B1(n8227), .B2(n10819), .ZN(n8028) );
  AOI21_X1 U9221 ( .B1(n10959), .B2(n8301), .A(n8028), .ZN(n8029) );
  OAI21_X1 U9222 ( .B1(n10777), .B2(n10429), .A(n8029), .ZN(n8030) );
  AOI21_X1 U9223 ( .B1(n10778), .B2(n10822), .A(n8030), .ZN(n8031) );
  OAI21_X1 U9224 ( .B1(n10775), .B2(n10406), .A(n8031), .ZN(P1_U3283) );
  INV_X1 U9225 ( .A(n10658), .ZN(n10239) );
  INV_X1 U9226 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8032) );
  OAI222_X1 U9227 ( .A1(n10239), .A2(P1_U3084), .B1(n10541), .B2(n8033), .C1(
        n8032), .C2(n8855), .ZN(P1_U3335) );
  NAND2_X1 U9228 ( .A1(n8035), .A2(n8034), .ZN(n10703) );
  INV_X1 U9229 ( .A(n10703), .ZN(n8049) );
  INV_X1 U9230 ( .A(n8036), .ZN(n8037) );
  OR2_X1 U9231 ( .A1(n8042), .A2(n9407), .ZN(n8059) );
  NAND2_X1 U9232 ( .A1(n8393), .A2(n8059), .ZN(n10848) );
  AOI22_X1 U9233 ( .A1(n10703), .A2(n9644), .B1(n9638), .B2(n7404), .ZN(n10705) );
  OAI22_X1 U9234 ( .A1(n10705), .A2(n10851), .B1(n8043), .B2(n10860), .ZN(
        n8044) );
  AOI21_X1 U9235 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n10851), .A(n8044), .ZN(
        n8048) );
  INV_X1 U9236 ( .A(n10702), .ZN(n8045) );
  OAI21_X1 U9237 ( .B1(n9655), .B2(n9610), .A(n10701), .ZN(n8047) );
  OAI211_X1 U9238 ( .C1(n8049), .C2(n9602), .A(n8048), .B(n8047), .ZN(P2_U3296) );
  XNOR2_X1 U9239 ( .A(n8051), .B(n8050), .ZN(n8058) );
  OR2_X1 U9240 ( .A1(n8053), .A2(n8052), .ZN(n8054) );
  NAND2_X1 U9241 ( .A1(n8055), .A2(n8054), .ZN(n10720) );
  NAND2_X1 U9242 ( .A1(n10720), .A2(n8293), .ZN(n8057) );
  AOI22_X1 U9243 ( .A1(n9619), .A2(n7404), .B1(n9396), .B2(n9638), .ZN(n8056)
         );
  OAI211_X1 U9244 ( .C1(n8058), .C2(n9561), .A(n8057), .B(n8056), .ZN(n10718)
         );
  INV_X1 U9245 ( .A(n10718), .ZN(n8073) );
  INV_X1 U9246 ( .A(n8059), .ZN(n8060) );
  NAND2_X1 U9247 ( .A1(n10856), .A2(n8060), .ZN(n8404) );
  INV_X1 U9248 ( .A(n8404), .ZN(n8071) );
  NAND2_X1 U9249 ( .A1(n8062), .A2(n8061), .ZN(n8063) );
  NAND2_X1 U9250 ( .A1(n8064), .A2(n8063), .ZN(n10717) );
  INV_X1 U9251 ( .A(n10717), .ZN(n8066) );
  INV_X1 U9252 ( .A(n10860), .ZN(n10755) );
  AND2_X1 U9253 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(n10755), .ZN(n8065) );
  AOI21_X1 U9254 ( .B1(n9610), .B2(n8066), .A(n8065), .ZN(n8069) );
  OR2_X1 U9255 ( .A1(n10856), .A2(n8067), .ZN(n8068) );
  OAI211_X1 U9256 ( .C1(n10716), .C2(n9628), .A(n8069), .B(n8068), .ZN(n8070)
         );
  AOI21_X1 U9257 ( .B1(n8071), .B2(n10720), .A(n8070), .ZN(n8072) );
  OAI21_X1 U9258 ( .B1(n10851), .B2(n8073), .A(n8072), .ZN(P2_U3294) );
  INV_X1 U9259 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U9260 ( .A1(n8074), .A2(n5011), .ZN(n8075) );
  OAI21_X1 U9261 ( .B1(n5011), .B2(n8076), .A(n8075), .ZN(P2_U3460) );
  OR2_X1 U9262 ( .A1(n8463), .A2(n9393), .ZN(n8077) );
  NAND2_X1 U9263 ( .A1(n8081), .A2(n8083), .ZN(n8283) );
  OAI21_X1 U9264 ( .B1(n8081), .B2(n8083), .A(n8283), .ZN(n8195) );
  INV_X1 U9265 ( .A(n8082), .ZN(n8085) );
  OAI21_X1 U9266 ( .B1(n8085), .B2(n8084), .A(n8083), .ZN(n8087) );
  AOI21_X1 U9267 ( .B1(n8087), .B2(n8086), .A(n9561), .ZN(n8089) );
  NOR2_X1 U9268 ( .A1(n8089), .A2(n8088), .ZN(n8204) );
  OAI211_X1 U9269 ( .C1(n8090), .C2(n8351), .A(n9746), .B(n8295), .ZN(n8200)
         );
  OAI211_X1 U9270 ( .C1(n9750), .C2(n8195), .A(n8204), .B(n8200), .ZN(n8353)
         );
  OAI22_X1 U9271 ( .A1(n9742), .A2(n8351), .B1(n10923), .B2(n6078), .ZN(n8091)
         );
  AOI21_X1 U9272 ( .B1(n8353), .B2(n10923), .A(n8091), .ZN(n8092) );
  INV_X1 U9273 ( .A(n8092), .ZN(P2_U3528) );
  INV_X1 U9274 ( .A(n8385), .ZN(n8297) );
  OAI21_X1 U9275 ( .B1(n8095), .B2(n8094), .A(n8093), .ZN(n8096) );
  NAND2_X1 U9276 ( .A1(n8096), .A2(n9352), .ZN(n8101) );
  INV_X1 U9277 ( .A(n8097), .ZN(n8099) );
  OAI22_X1 U9278 ( .A1(n9365), .A2(n8285), .B1(n9363), .B2(n8296), .ZN(n8098)
         );
  AOI211_X1 U9279 ( .C1(n9334), .C2(n9391), .A(n8099), .B(n8098), .ZN(n8100)
         );
  OAI211_X1 U9280 ( .C1(n8297), .C2(n9358), .A(n8101), .B(n8100), .ZN(P2_U3233) );
  NOR2_X1 U9281 ( .A1(n10856), .A2(n8102), .ZN(n8106) );
  OAI22_X1 U9282 ( .A1(n8615), .A2(n8104), .B1(n8103), .B2(n10860), .ZN(n8105)
         );
  AOI211_X1 U9283 ( .C1(n9660), .C2(n8107), .A(n8106), .B(n8105), .ZN(n8110)
         );
  NAND2_X1 U9284 ( .A1(n9655), .A2(n8108), .ZN(n8109) );
  OAI211_X1 U9285 ( .C1(n10851), .C2(n8111), .A(n8110), .B(n8109), .ZN(
        P2_U3295) );
  AOI211_X1 U9286 ( .C1(n8113), .C2(n10932), .A(n8112), .B(n10254), .ZN(n8121)
         );
  AOI211_X1 U9287 ( .C1(n8116), .C2(n8115), .A(n8114), .B(n10651), .ZN(n8120)
         );
  NAND2_X1 U9288 ( .A1(n5013), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9918) );
  NAND2_X1 U9289 ( .A1(n10648), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n8117) );
  OAI211_X1 U9290 ( .C1(n10249), .C2(n8118), .A(n9918), .B(n8117), .ZN(n8119)
         );
  OR3_X1 U9291 ( .A1(n8121), .A2(n8120), .A3(n8119), .ZN(P1_U3256) );
  NAND2_X1 U9292 ( .A1(n8123), .A2(n8122), .ZN(n8124) );
  INV_X1 U9293 ( .A(n8125), .ZN(n8253) );
  NOR2_X1 U9294 ( .A1(n9903), .A2(n8256), .ZN(n8129) );
  NAND2_X1 U9295 ( .A1(n9923), .A2(n10207), .ZN(n8126) );
  OAI211_X1 U9296 ( .C1(n8244), .C2(n9919), .A(n8127), .B(n8126), .ZN(n8128)
         );
  AOI211_X1 U9297 ( .C1(n8253), .C2(n9900), .A(n8129), .B(n8128), .ZN(n8130)
         );
  OAI21_X1 U9298 ( .B1(n8131), .B2(n9931), .A(n8130), .ZN(P1_U3211) );
  INV_X1 U9299 ( .A(n8132), .ZN(n8133) );
  AOI21_X1 U9300 ( .B1(n10159), .B2(n8134), .A(n8133), .ZN(n10762) );
  AND2_X1 U9301 ( .A1(n8135), .A2(n10120), .ZN(n8155) );
  XNOR2_X1 U9302 ( .A(n9934), .B(n10159), .ZN(n8139) );
  OAI22_X1 U9303 ( .A1(n8137), .A2(n10403), .B1(n8136), .B2(n10401), .ZN(n8138) );
  AOI21_X1 U9304 ( .B1(n8139), .B2(n10947), .A(n8138), .ZN(n8140) );
  OAI21_X1 U9305 ( .B1(n10762), .B2(n8848), .A(n8140), .ZN(n10764) );
  NAND2_X1 U9306 ( .A1(n10764), .A2(n10822), .ZN(n8148) );
  OAI22_X1 U9307 ( .A1(n10822), .A2(n8142), .B1(n8141), .B2(n10819), .ZN(n8145) );
  NAND2_X1 U9308 ( .A1(n8153), .A2(n8146), .ZN(n8143) );
  NAND2_X1 U9309 ( .A1(n8251), .A2(n8143), .ZN(n10763) );
  NOR2_X1 U9310 ( .A1(n10763), .A2(n10429), .ZN(n8144) );
  AOI211_X1 U9311 ( .C1(n10959), .C2(n8146), .A(n8145), .B(n8144), .ZN(n8147)
         );
  OAI211_X1 U9312 ( .C1(n10762), .C2(n10385), .A(n8148), .B(n8147), .ZN(
        P1_U3285) );
  NAND2_X1 U9313 ( .A1(n8150), .A2(n10157), .ZN(n8151) );
  NAND2_X1 U9314 ( .A1(n8149), .A2(n8151), .ZN(n10739) );
  AOI21_X1 U9315 ( .B1(n8152), .B2(n10744), .A(n10927), .ZN(n8154) );
  AND2_X1 U9316 ( .A1(n8154), .A2(n8153), .ZN(n10741) );
  INV_X1 U9317 ( .A(n8155), .ZN(n8157) );
  NAND2_X1 U9318 ( .A1(n8157), .A2(n10157), .ZN(n8156) );
  OAI21_X1 U9319 ( .B1(n10157), .B2(n8157), .A(n8156), .ZN(n8158) );
  NAND2_X1 U9320 ( .A1(n8158), .A2(n10947), .ZN(n8160) );
  AOI22_X1 U9321 ( .A1(n10944), .A2(n10209), .B1(n10207), .B2(n10942), .ZN(
        n8159) );
  NAND2_X1 U9322 ( .A1(n8160), .A2(n8159), .ZN(n10749) );
  AOI211_X1 U9323 ( .C1(n10802), .C2(n10744), .A(n10741), .B(n10749), .ZN(
        n8161) );
  OAI21_X1 U9324 ( .B1(n10800), .B2(n10739), .A(n8161), .ZN(n8166) );
  NAND2_X1 U9325 ( .A1(n8166), .A2(n10977), .ZN(n8162) );
  OAI21_X1 U9326 ( .B1(n10977), .B2(n7150), .A(n8162), .ZN(P1_U3528) );
  INV_X1 U9327 ( .A(n8163), .ZN(n8164) );
  OAI222_X1 U9328 ( .A1(n10740), .A2(n5013), .B1(n10541), .B2(n8164), .C1(
        n8987), .C2(n8855), .ZN(P1_U3334) );
  OAI222_X1 U9329 ( .A1(n8831), .A2(n8165), .B1(n8691), .B2(n8164), .C1(n9407), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U9330 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U9331 ( .A1(n8166), .A2(n10981), .ZN(n8167) );
  OAI21_X1 U9332 ( .B1(n10981), .B2(n8168), .A(n8167), .ZN(P1_U3469) );
  XNOR2_X1 U9333 ( .A(n8170), .B(n8169), .ZN(n8176) );
  INV_X1 U9334 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8171) );
  OAI22_X1 U9335 ( .A1(n9362), .A2(n8506), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8171), .ZN(n8174) );
  OAI22_X1 U9336 ( .A1(n9365), .A2(n8172), .B1(n9363), .B2(n8398), .ZN(n8173)
         );
  AOI211_X1 U9337 ( .C1(n9379), .C2(n8416), .A(n8174), .B(n8173), .ZN(n8175)
         );
  OAI21_X1 U9338 ( .B1(n8176), .B2(n9381), .A(n8175), .ZN(P2_U3219) );
  NOR2_X1 U9339 ( .A1(n8185), .A2(n8177), .ZN(n8179) );
  NOR2_X1 U9340 ( .A1(n8179), .A2(n8178), .ZN(n8181) );
  XNOR2_X1 U9341 ( .A(n8364), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U9342 ( .A1(n8181), .A2(n8180), .ZN(n8365) );
  OAI21_X1 U9343 ( .B1(n8181), .B2(n8180), .A(n8365), .ZN(n8182) );
  INV_X1 U9344 ( .A(n8182), .ZN(n8194) );
  INV_X1 U9345 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U9346 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8697) );
  OAI21_X1 U9347 ( .B1(n8373), .B2(n8183), .A(n8697), .ZN(n8192) );
  NAND2_X1 U9348 ( .A1(n8185), .A2(n8184), .ZN(n8187) );
  NAND2_X1 U9349 ( .A1(n8187), .A2(n8186), .ZN(n8190) );
  NAND2_X1 U9350 ( .A1(n8377), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8188) );
  OAI21_X1 U9351 ( .B1(n8377), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8188), .ZN(
        n8189) );
  NOR2_X1 U9352 ( .A1(n8190), .A2(n8189), .ZN(n8376) );
  AOI211_X1 U9353 ( .C1(n8190), .C2(n8189), .A(n8376), .B(n10689), .ZN(n8191)
         );
  AOI211_X1 U9354 ( .C1(n8377), .C2(n10680), .A(n8192), .B(n8191), .ZN(n8193)
         );
  OAI21_X1 U9355 ( .B1(n8194), .B2(n9422), .A(n8193), .ZN(P2_U3261) );
  INV_X1 U9356 ( .A(n8195), .ZN(n8202) );
  AND2_X1 U9357 ( .A1(n10856), .A2(n9407), .ZN(n9633) );
  INV_X1 U9358 ( .A(n9633), .ZN(n9658) );
  OAI22_X1 U9359 ( .A1(n10856), .A2(n8197), .B1(n8196), .B2(n10860), .ZN(n8198) );
  AOI21_X1 U9360 ( .B1(n9655), .B2(n8281), .A(n8198), .ZN(n8199) );
  OAI21_X1 U9361 ( .B1(n8200), .B2(n9658), .A(n8199), .ZN(n8201) );
  AOI21_X1 U9362 ( .B1(n8202), .B2(n9660), .A(n8201), .ZN(n8203) );
  OAI21_X1 U9363 ( .B1(n8204), .B2(n10851), .A(n8203), .ZN(P2_U3288) );
  XNOR2_X1 U9364 ( .A(n8205), .B(n8215), .ZN(n8206) );
  NAND2_X1 U9365 ( .A1(n8206), .A2(n9644), .ZN(n8208) );
  AOI22_X1 U9366 ( .A1(n9619), .A2(n9396), .B1(n8455), .B2(n9638), .ZN(n8207)
         );
  NAND2_X1 U9367 ( .A1(n8208), .A2(n8207), .ZN(n10733) );
  OR2_X1 U9368 ( .A1(n8209), .A2(n10731), .ZN(n8210) );
  NAND2_X1 U9369 ( .A1(n8211), .A2(n8210), .ZN(n10732) );
  INV_X1 U9370 ( .A(n8212), .ZN(n8213) );
  AOI21_X1 U9371 ( .B1(n8215), .B2(n8214), .A(n8213), .ZN(n10735) );
  NAND2_X1 U9372 ( .A1(n10735), .A2(n9660), .ZN(n8220) );
  OAI22_X1 U9373 ( .A1(n10856), .A2(n7522), .B1(n8216), .B2(n10860), .ZN(n8217) );
  AOI21_X1 U9374 ( .B1(n9655), .B2(n8218), .A(n8217), .ZN(n8219) );
  OAI211_X1 U9375 ( .C1(n8615), .C2(n10732), .A(n8220), .B(n8219), .ZN(n8221)
         );
  AOI21_X1 U9376 ( .B1(n10856), .B2(n10733), .A(n8221), .ZN(n8222) );
  INV_X1 U9377 ( .A(n8222), .ZN(P2_U3292) );
  NAND2_X1 U9378 ( .A1(n8224), .A2(n8223), .ZN(n8225) );
  XOR2_X1 U9379 ( .A(n8226), .B(n8225), .Z(n8235) );
  INV_X1 U9380 ( .A(n8227), .ZN(n8233) );
  INV_X1 U9381 ( .A(n8228), .ZN(n8230) );
  NAND2_X1 U9382 ( .A1(n9923), .A2(n10206), .ZN(n8229) );
  OAI211_X1 U9383 ( .C1(n8304), .C2(n9919), .A(n8230), .B(n8229), .ZN(n8232)
         );
  NOR2_X1 U9384 ( .A1(n10776), .A2(n9903), .ZN(n8231) );
  AOI211_X1 U9385 ( .C1(n8233), .C2(n9900), .A(n8232), .B(n8231), .ZN(n8234)
         );
  OAI21_X1 U9386 ( .B1(n8235), .B2(n9931), .A(n8234), .ZN(P1_U3219) );
  INV_X1 U9387 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8236) );
  NOR2_X1 U9388 ( .A1(n5011), .A2(n8236), .ZN(n8237) );
  AOI21_X1 U9389 ( .B1(n5011), .B2(n8238), .A(n8237), .ZN(n8239) );
  OAI21_X1 U9390 ( .B1(n8240), .B2(n9786), .A(n8239), .ZN(P2_U3454) );
  OAI21_X1 U9391 ( .B1(n8242), .B2(n8241), .A(n8306), .ZN(n8249) );
  OAI22_X1 U9392 ( .A1(n8244), .A2(n10403), .B1(n8243), .B2(n10401), .ZN(n8248) );
  OAI21_X1 U9393 ( .B1(n8246), .B2(n10161), .A(n8245), .ZN(n8258) );
  INV_X1 U9394 ( .A(n8258), .ZN(n8411) );
  NOR2_X1 U9395 ( .A1(n8411), .A2(n8848), .ZN(n8247) );
  AOI211_X1 U9396 ( .C1(n10947), .C2(n8249), .A(n8248), .B(n8247), .ZN(n8410)
         );
  AOI211_X1 U9397 ( .C1(n8408), .C2(n8251), .A(n10927), .B(n8250), .ZN(n8407)
         );
  NOR2_X1 U9398 ( .A1(n8252), .A2(n10366), .ZN(n10962) );
  NAND2_X1 U9399 ( .A1(n8407), .A2(n10962), .ZN(n8255) );
  AOI22_X1 U9400 ( .A1(n10969), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n8253), .B2(
        n10957), .ZN(n8254) );
  OAI211_X1 U9401 ( .C1(n8256), .C2(n10792), .A(n8255), .B(n8254), .ZN(n8257)
         );
  AOI21_X1 U9402 ( .B1(n8258), .B2(n10887), .A(n8257), .ZN(n8259) );
  OAI21_X1 U9403 ( .B1(n8410), .B2(n10969), .A(n8259), .ZN(P1_U3284) );
  XNOR2_X1 U9404 ( .A(n8261), .B(n8260), .ZN(n8268) );
  NAND2_X1 U9405 ( .A1(n9389), .A2(n9638), .ZN(n8263) );
  NAND2_X1 U9406 ( .A1(n9391), .A2(n9619), .ZN(n8262) );
  AND2_X1 U9407 ( .A1(n8263), .A2(n8262), .ZN(n8426) );
  INV_X1 U9408 ( .A(n8426), .ZN(n10850) );
  AOI21_X1 U9409 ( .B1(n9373), .B2(n10850), .A(n8264), .ZN(n8265) );
  OAI21_X1 U9410 ( .B1(n9363), .B2(n10861), .A(n8265), .ZN(n8266) );
  AOI21_X1 U9411 ( .B1(n10852), .B2(n9379), .A(n8266), .ZN(n8267) );
  OAI21_X1 U9412 ( .B1(n8268), .B2(n9381), .A(n8267), .ZN(P2_U3238) );
  AOI211_X1 U9413 ( .C1(n8271), .C2(n8270), .A(n8269), .B(n10651), .ZN(n8280)
         );
  AOI211_X1 U9414 ( .C1(n8274), .C2(n8273), .A(n8272), .B(n10254), .ZN(n8279)
         );
  NAND2_X1 U9415 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(n5013), .ZN(n8276) );
  NAND2_X1 U9416 ( .A1(n10648), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8275) );
  OAI211_X1 U9417 ( .C1(n10249), .C2(n8277), .A(n8276), .B(n8275), .ZN(n8278)
         );
  OR3_X1 U9418 ( .A1(n8280), .A2(n8279), .A3(n8278), .ZN(P1_U3257) );
  NAND2_X1 U9419 ( .A1(n8281), .A2(n9392), .ZN(n8282) );
  OAI21_X1 U9420 ( .B1(n5095), .B2(n8289), .A(n8387), .ZN(n8292) );
  INV_X1 U9421 ( .A(n8292), .ZN(n8317) );
  OAI22_X1 U9422 ( .A1(n8285), .A2(n9641), .B1(n8284), .B2(n9565), .ZN(n8291)
         );
  INV_X1 U9423 ( .A(n8286), .ZN(n8287) );
  AOI211_X1 U9424 ( .C1(n8289), .C2(n8288), .A(n9561), .B(n8287), .ZN(n8290)
         );
  AOI211_X1 U9425 ( .C1(n8293), .C2(n8292), .A(n8291), .B(n8290), .ZN(n8315)
         );
  MUX2_X1 U9426 ( .A(n8294), .B(n8315), .S(n10856), .Z(n8300) );
  AOI21_X1 U9427 ( .B1(n8385), .B2(n8295), .A(n5090), .ZN(n8313) );
  OAI22_X1 U9428 ( .A1(n8297), .A2(n9628), .B1(n8296), .B2(n10860), .ZN(n8298)
         );
  AOI21_X1 U9429 ( .B1(n8313), .B2(n9610), .A(n8298), .ZN(n8299) );
  OAI211_X1 U9430 ( .C1(n8317), .C2(n8404), .A(n8300), .B(n8299), .ZN(P2_U3287) );
  NAND2_X1 U9431 ( .A1(n8301), .A2(n8335), .ZN(n8302) );
  OR2_X1 U9432 ( .A1(n8471), .A2(n8304), .ZN(n10064) );
  NAND2_X1 U9433 ( .A1(n8471), .A2(n8304), .ZN(n10037) );
  XNOR2_X1 U9434 ( .A(n8474), .B(n10162), .ZN(n10783) );
  INV_X1 U9435 ( .A(n10043), .ZN(n9941) );
  INV_X1 U9436 ( .A(n10162), .ZN(n8307) );
  OAI21_X1 U9437 ( .B1(n5091), .B2(n8307), .A(n8478), .ZN(n8308) );
  AOI222_X1 U9438 ( .A1(n10947), .A2(n8308), .B1(n10205), .B2(n10942), .C1(
        n8335), .C2(n10944), .ZN(n10784) );
  INV_X1 U9439 ( .A(n10803), .ZN(n8309) );
  AOI21_X1 U9440 ( .B1(n8471), .B2(n8310), .A(n8309), .ZN(n10787) );
  AOI22_X1 U9441 ( .A1(n10787), .A2(n10973), .B1(n10802), .B2(n8471), .ZN(
        n8311) );
  OAI211_X1 U9442 ( .C1(n10783), .C2(n10800), .A(n10784), .B(n8311), .ZN(n8320) );
  NAND2_X1 U9443 ( .A1(n8320), .A2(n10977), .ZN(n8312) );
  OAI21_X1 U9444 ( .B1(n10977), .B2(n7209), .A(n8312), .ZN(P1_U3532) );
  INV_X1 U9445 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8319) );
  AOI22_X1 U9446 ( .A1(n8313), .A2(n9746), .B1(n9745), .B2(n8385), .ZN(n8314)
         );
  OAI211_X1 U9447 ( .C1(n8317), .C2(n8316), .A(n8315), .B(n8314), .ZN(n8323)
         );
  NAND2_X1 U9448 ( .A1(n8323), .A2(n5011), .ZN(n8318) );
  OAI21_X1 U9449 ( .B1(n5011), .B2(n8319), .A(n8318), .ZN(P2_U3478) );
  INV_X1 U9450 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U9451 ( .A1(n8320), .A2(n10981), .ZN(n8321) );
  OAI21_X1 U9452 ( .B1(n10981), .B2(n8322), .A(n8321), .ZN(P1_U3481) );
  NAND2_X1 U9453 ( .A1(n8323), .A2(n10923), .ZN(n8324) );
  OAI21_X1 U9454 ( .B1(n10923), .B2(n6088), .A(n8324), .ZN(P2_U3529) );
  INV_X1 U9455 ( .A(n8325), .ZN(n8406) );
  OAI222_X1 U9456 ( .A1(P1_U3084), .A2(n8327), .B1(n10541), .B2(n8406), .C1(
        n8326), .C2(n8855), .ZN(P1_U3333) );
  INV_X1 U9457 ( .A(n8471), .ZN(n10793) );
  OAI21_X1 U9458 ( .B1(n8330), .B2(n8329), .A(n8328), .ZN(n8331) );
  NAND2_X1 U9459 ( .A1(n8331), .A2(n9893), .ZN(n8337) );
  INV_X1 U9460 ( .A(n10205), .ZN(n8475) );
  OAI22_X1 U9461 ( .A1(n8475), .A2(n9919), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8332), .ZN(n8334) );
  NOR2_X1 U9462 ( .A1(n9926), .A2(n10788), .ZN(n8333) );
  AOI211_X1 U9463 ( .C1(n9923), .C2(n8335), .A(n8334), .B(n8333), .ZN(n8336)
         );
  OAI211_X1 U9464 ( .C1(n10793), .C2(n9903), .A(n8337), .B(n8336), .ZN(
        P1_U3229) );
  INV_X1 U9465 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8338) );
  OAI22_X1 U9466 ( .A1(n9786), .A2(n8339), .B1(n5011), .B2(n8338), .ZN(n8340)
         );
  INV_X1 U9467 ( .A(n8340), .ZN(n8341) );
  OAI21_X1 U9468 ( .B1(n8342), .B2(n10985), .A(n8341), .ZN(P2_U3466) );
  INV_X1 U9469 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8343) );
  OAI22_X1 U9470 ( .A1(n9786), .A2(n8344), .B1(n5011), .B2(n8343), .ZN(n8345)
         );
  INV_X1 U9471 ( .A(n8345), .ZN(n8346) );
  OAI21_X1 U9472 ( .B1(n8347), .B2(n10985), .A(n8346), .ZN(P2_U3472) );
  INV_X1 U9473 ( .A(n8348), .ZN(n8384) );
  OAI222_X1 U9474 ( .A1(n8691), .A2(n8384), .B1(P2_U3152), .B2(n8350), .C1(
        n8349), .C2(n8831), .ZN(P2_U3337) );
  OAI22_X1 U9475 ( .A1(n9786), .A2(n8351), .B1(n5011), .B2(n6075), .ZN(n8352)
         );
  AOI21_X1 U9476 ( .B1(n8353), .B2(n5011), .A(n8352), .ZN(n8354) );
  INV_X1 U9477 ( .A(n8354), .ZN(P2_U3475) );
  AOI22_X1 U9478 ( .A1(n10851), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n10755), .B2(
        n9139), .ZN(n8355) );
  OAI21_X1 U9479 ( .B1(n8356), .B2(n9628), .A(n8355), .ZN(n8359) );
  NOR2_X1 U9480 ( .A1(n8357), .A2(n8404), .ZN(n8358) );
  AOI211_X1 U9481 ( .C1(n8360), .C2(n9610), .A(n8359), .B(n8358), .ZN(n8361)
         );
  OAI21_X1 U9482 ( .B1(n8362), .B2(n10851), .A(n8361), .ZN(P2_U3293) );
  INV_X1 U9483 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8372) );
  XNOR2_X1 U9484 ( .A(n9400), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U9485 ( .A1(n8364), .A2(n8363), .ZN(n8366) );
  NAND2_X1 U9486 ( .A1(n8366), .A2(n8365), .ZN(n8367) );
  NOR2_X1 U9487 ( .A1(n8368), .A2(n8367), .ZN(n9399) );
  AOI21_X1 U9488 ( .B1(n8368), .B2(n8367), .A(n9399), .ZN(n8369) );
  NAND2_X1 U9489 ( .A1(n10684), .A2(n8369), .ZN(n8371) );
  NAND2_X1 U9490 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n8370) );
  OAI211_X1 U9491 ( .C1(n8373), .C2(n8372), .A(n8371), .B(n8370), .ZN(n8381)
         );
  INV_X1 U9492 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9630) );
  OR2_X1 U9493 ( .A1(n9400), .A2(n9630), .ZN(n8375) );
  NAND2_X1 U9494 ( .A1(n9400), .A2(n9630), .ZN(n8374) );
  AND2_X1 U9495 ( .A1(n8375), .A2(n8374), .ZN(n8379) );
  AOI21_X1 U9496 ( .B1(n8377), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8376), .ZN(
        n8378) );
  NOR2_X1 U9497 ( .A1(n8378), .A2(n8379), .ZN(n9398) );
  AOI211_X1 U9498 ( .C1(n8379), .C2(n8378), .A(n9398), .B(n10689), .ZN(n8380)
         );
  AOI211_X1 U9499 ( .C1(n10680), .C2(n9400), .A(n8381), .B(n8380), .ZN(n8382)
         );
  INV_X1 U9500 ( .A(n8382), .ZN(P2_U3262) );
  OAI222_X1 U9501 ( .A1(n5013), .A2(n10183), .B1(n10541), .B2(n8384), .C1(
        n8383), .C2(n8855), .ZN(P1_U3332) );
  OR2_X1 U9502 ( .A1(n8385), .A2(n8394), .ZN(n8386) );
  OAI21_X1 U9503 ( .B1(n8388), .B2(n8390), .A(n8418), .ZN(n10831) );
  NAND2_X1 U9504 ( .A1(n8391), .A2(n8390), .ZN(n8392) );
  AND2_X1 U9505 ( .A1(n5487), .A2(n8392), .ZN(n8397) );
  OR2_X1 U9506 ( .A1(n10831), .A2(n8393), .ZN(n8396) );
  AOI22_X1 U9507 ( .A1(n9619), .A2(n8394), .B1(n9390), .B2(n9638), .ZN(n8395)
         );
  OAI211_X1 U9508 ( .C1(n9561), .C2(n8397), .A(n8396), .B(n8395), .ZN(n10833)
         );
  NAND2_X1 U9509 ( .A1(n10833), .A2(n10856), .ZN(n8403) );
  OAI22_X1 U9510 ( .A1(n10856), .A2(n8399), .B1(n8398), .B2(n10860), .ZN(n8401) );
  OAI21_X1 U9511 ( .B1(n5090), .B2(n5352), .A(n8423), .ZN(n10832) );
  NOR2_X1 U9512 ( .A1(n10832), .A2(n8615), .ZN(n8400) );
  AOI211_X1 U9513 ( .C1(n9655), .C2(n8416), .A(n8401), .B(n8400), .ZN(n8402)
         );
  OAI211_X1 U9514 ( .C1(n10831), .C2(n8404), .A(n8403), .B(n8402), .ZN(
        P2_U3286) );
  OAI222_X1 U9515 ( .A1(n8691), .A2(n8406), .B1(P2_U3152), .B2(n6004), .C1(
        n8405), .C2(n8831), .ZN(P2_U3338) );
  AOI21_X1 U9516 ( .B1(n10802), .B2(n8408), .A(n8407), .ZN(n8409) );
  OAI211_X1 U9517 ( .C1(n8411), .C2(n10520), .A(n8410), .B(n8409), .ZN(n8413)
         );
  NAND2_X1 U9518 ( .A1(n8413), .A2(n10977), .ZN(n8412) );
  OAI21_X1 U9519 ( .B1(n10977), .B2(n6698), .A(n8412), .ZN(P1_U3530) );
  INV_X1 U9520 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U9521 ( .A1(n8413), .A2(n10981), .ZN(n8414) );
  OAI21_X1 U9522 ( .B1(n10981), .B2(n8415), .A(n8414), .ZN(P1_U3475) );
  NAND2_X1 U9523 ( .A1(n8416), .A2(n9391), .ZN(n8417) );
  XNOR2_X1 U9524 ( .A(n8500), .B(n8419), .ZN(n10849) );
  NAND2_X1 U9525 ( .A1(n5092), .A2(n8499), .ZN(n8421) );
  OAI211_X1 U9526 ( .C1(n8420), .C2(n8422), .A(n8421), .B(n9644), .ZN(n10854)
         );
  INV_X1 U9527 ( .A(n8507), .ZN(n8425) );
  AOI21_X1 U9528 ( .B1(n8423), .B2(n10852), .A(n10916), .ZN(n8424) );
  NAND2_X1 U9529 ( .A1(n8425), .A2(n8424), .ZN(n10855) );
  NAND3_X1 U9530 ( .A1(n10854), .A2(n8426), .A3(n10855), .ZN(n8427) );
  AOI21_X1 U9531 ( .B1(n10849), .B2(n10921), .A(n8427), .ZN(n8434) );
  INV_X1 U9532 ( .A(n9786), .ZN(n8430) );
  INV_X1 U9533 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8428) );
  NOR2_X1 U9534 ( .A1(n5011), .A2(n8428), .ZN(n8429) );
  AOI21_X1 U9535 ( .B1(n8430), .B2(n10852), .A(n8429), .ZN(n8431) );
  OAI21_X1 U9536 ( .B1(n8434), .B2(n10985), .A(n8431), .ZN(P2_U3484) );
  AOI22_X1 U9537 ( .A1(n8432), .A2(n10852), .B1(n10922), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n8433) );
  OAI21_X1 U9538 ( .B1(n8434), .B2(n10922), .A(n8433), .ZN(P2_U3531) );
  OAI21_X1 U9539 ( .B1(n8437), .B2(n8436), .A(n8435), .ZN(n8438) );
  NAND2_X1 U9540 ( .A1(n8438), .A2(n9352), .ZN(n8443) );
  INV_X1 U9541 ( .A(n8439), .ZN(n8441) );
  OAI22_X1 U9542 ( .A1(n9365), .A2(n8506), .B1(n9363), .B2(n8508), .ZN(n8440)
         );
  AOI211_X1 U9543 ( .C1(n9334), .C2(n9388), .A(n8441), .B(n8440), .ZN(n8442)
         );
  OAI211_X1 U9544 ( .C1(n10892), .C2(n9358), .A(n8443), .B(n8442), .ZN(
        P2_U3226) );
  XNOR2_X1 U9545 ( .A(n8444), .B(n8453), .ZN(n10772) );
  INV_X1 U9546 ( .A(n8445), .ZN(n8446) );
  OAI21_X1 U9547 ( .B1(n10768), .B2(n8447), .A(n8446), .ZN(n10769) );
  INV_X1 U9548 ( .A(n8448), .ZN(n8449) );
  AOI22_X1 U9549 ( .A1(n9655), .A2(n8450), .B1(n8449), .B2(n10755), .ZN(n8451)
         );
  OAI21_X1 U9550 ( .B1(n10769), .B2(n8615), .A(n8451), .ZN(n8459) );
  OAI211_X1 U9551 ( .C1(n8454), .C2(n8453), .A(n8452), .B(n9644), .ZN(n8457)
         );
  AOI22_X1 U9552 ( .A1(n9619), .A2(n8455), .B1(n9393), .B2(n9638), .ZN(n8456)
         );
  NAND2_X1 U9553 ( .A1(n8457), .A2(n8456), .ZN(n10770) );
  MUX2_X1 U9554 ( .A(n10770), .B(P2_REG2_REG_6__SCAN_IN), .S(n10851), .Z(n8458) );
  AOI211_X1 U9555 ( .C1(n9660), .C2(n10772), .A(n8459), .B(n8458), .ZN(n8460)
         );
  INV_X1 U9556 ( .A(n8460), .ZN(P2_U3290) );
  INV_X1 U9557 ( .A(n8461), .ZN(n8462) );
  AOI22_X1 U9558 ( .A1(n9655), .A2(n8463), .B1(n10755), .B2(n8462), .ZN(n8464)
         );
  OAI21_X1 U9559 ( .B1(n8465), .B2(n8615), .A(n8464), .ZN(n8468) );
  MUX2_X1 U9560 ( .A(n8466), .B(P2_REG2_REG_7__SCAN_IN), .S(n10851), .Z(n8467)
         );
  AOI211_X1 U9561 ( .C1(n9660), .C2(n8469), .A(n8468), .B(n8467), .ZN(n8470)
         );
  INV_X1 U9562 ( .A(n8470), .ZN(P2_U3289) );
  AND2_X1 U9563 ( .A1(n8471), .A2(n10811), .ZN(n8473) );
  OR2_X1 U9564 ( .A1(n10828), .A2(n8475), .ZN(n10066) );
  NAND2_X1 U9565 ( .A1(n10828), .A2(n8475), .ZN(n10038) );
  NAND2_X1 U9566 ( .A1(n10066), .A2(n10038), .ZN(n10798) );
  NAND2_X1 U9567 ( .A1(n10799), .A2(n10798), .ZN(n8477) );
  OR2_X1 U9568 ( .A1(n10828), .A2(n10205), .ZN(n8476) );
  NAND2_X1 U9569 ( .A1(n8477), .A2(n8476), .ZN(n8625) );
  INV_X1 U9570 ( .A(n10871), .ZN(n8493) );
  OR2_X1 U9571 ( .A1(n8626), .A2(n8493), .ZN(n10068) );
  NAND2_X1 U9572 ( .A1(n8626), .A2(n8493), .ZN(n10041) );
  XNOR2_X1 U9573 ( .A(n8625), .B(n9948), .ZN(n10843) );
  INV_X1 U9574 ( .A(n10798), .ZN(n10809) );
  NAND2_X1 U9575 ( .A1(n10807), .A2(n10809), .ZN(n10808) );
  XNOR2_X1 U9576 ( .A(n8620), .B(n9948), .ZN(n8480) );
  AOI22_X1 U9577 ( .A1(n10944), .A2(n10205), .B1(n10204), .B2(n10942), .ZN(
        n8479) );
  OAI21_X1 U9578 ( .B1(n8480), .B2(n10873), .A(n8479), .ZN(n8481) );
  AOI21_X1 U9579 ( .B1(n10843), .B2(n10876), .A(n8481), .ZN(n10845) );
  INV_X1 U9580 ( .A(n8626), .ZN(n10840) );
  NOR2_X1 U9581 ( .A1(n10806), .A2(n10840), .ZN(n8482) );
  OR2_X1 U9582 ( .A1(n10866), .A2(n8482), .ZN(n10841) );
  OAI22_X1 U9583 ( .A1(n10822), .A2(n8483), .B1(n8521), .B2(n10819), .ZN(n8484) );
  AOI21_X1 U9584 ( .B1(n8626), .B2(n10959), .A(n8484), .ZN(n8485) );
  OAI21_X1 U9585 ( .B1(n10841), .B2(n10429), .A(n8485), .ZN(n8486) );
  AOI21_X1 U9586 ( .B1(n10843), .B2(n10887), .A(n8486), .ZN(n8487) );
  OAI21_X1 U9587 ( .B1(n10845), .B2(n10969), .A(n8487), .ZN(P1_U3280) );
  NAND2_X1 U9588 ( .A1(n8488), .A2(n8489), .ZN(n8491) );
  XNOR2_X1 U9589 ( .A(n8491), .B(n8490), .ZN(n8498) );
  NOR2_X1 U9590 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8492), .ZN(n10229) );
  NOR2_X1 U9591 ( .A1(n8493), .A2(n9919), .ZN(n8494) );
  AOI211_X1 U9592 ( .C1(n9923), .C2(n10811), .A(n10229), .B(n8494), .ZN(n8495)
         );
  OAI21_X1 U9593 ( .B1(n9926), .B2(n10820), .A(n8495), .ZN(n8496) );
  AOI21_X1 U9594 ( .B1(n10828), .B2(n9928), .A(n8496), .ZN(n8497) );
  OAI21_X1 U9595 ( .B1(n8498), .B2(n9931), .A(n8497), .ZN(P1_U3215) );
  XNOR2_X1 U9596 ( .A(n8562), .B(n8563), .ZN(n10896) );
  INV_X1 U9597 ( .A(n10896), .ZN(n8514) );
  INV_X1 U9598 ( .A(n8501), .ZN(n8504) );
  AOI21_X1 U9599 ( .B1(n8420), .B2(n8502), .A(n8563), .ZN(n8503) );
  NOR2_X1 U9600 ( .A1(n8504), .A2(n8503), .ZN(n8505) );
  OAI222_X1 U9601 ( .A1(n9565), .A2(n8604), .B1(n9641), .B2(n8506), .C1(n9561), 
        .C2(n8505), .ZN(n10894) );
  OAI21_X1 U9602 ( .B1(n8507), .B2(n10892), .A(n8572), .ZN(n10893) );
  OAI22_X1 U9603 ( .A1(n10856), .A2(n8509), .B1(n8508), .B2(n10860), .ZN(n8510) );
  AOI21_X1 U9604 ( .B1(n8564), .B2(n9655), .A(n8510), .ZN(n8511) );
  OAI21_X1 U9605 ( .B1(n10893), .B2(n8615), .A(n8511), .ZN(n8512) );
  AOI21_X1 U9606 ( .B1(n10894), .B2(n10856), .A(n8512), .ZN(n8513) );
  OAI21_X1 U9607 ( .B1(n9602), .B2(n8514), .A(n8513), .ZN(P2_U3284) );
  XOR2_X1 U9608 ( .A(n8516), .B(n8517), .Z(n8524) );
  INV_X1 U9609 ( .A(n10204), .ZN(n8621) );
  OAI22_X1 U9610 ( .A1(n8621), .A2(n9919), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8518), .ZN(n8519) );
  AOI21_X1 U9611 ( .B1(n9923), .B2(n10205), .A(n8519), .ZN(n8520) );
  OAI21_X1 U9612 ( .B1(n9926), .B2(n8521), .A(n8520), .ZN(n8522) );
  AOI21_X1 U9613 ( .B1(n8626), .B2(n9928), .A(n8522), .ZN(n8523) );
  OAI21_X1 U9614 ( .B1(n8524), .B2(n9931), .A(n8523), .ZN(P1_U3234) );
  INV_X1 U9615 ( .A(n8605), .ZN(n8535) );
  OAI21_X1 U9616 ( .B1(n8527), .B2(n8526), .A(n8525), .ZN(n8528) );
  NAND2_X1 U9617 ( .A1(n8528), .A2(n9352), .ZN(n8534) );
  INV_X1 U9618 ( .A(n8529), .ZN(n8532) );
  OAI22_X1 U9619 ( .A1(n9365), .A2(n8530), .B1(n9363), .B2(n8569), .ZN(n8531)
         );
  AOI211_X1 U9620 ( .C1(n9334), .C2(n9387), .A(n8532), .B(n8531), .ZN(n8533)
         );
  OAI211_X1 U9621 ( .C1(n8535), .C2(n9358), .A(n8534), .B(n8533), .ZN(P2_U3236) );
  INV_X1 U9622 ( .A(n8536), .ZN(n8539) );
  OAI222_X1 U9623 ( .A1(n8538), .A2(n5013), .B1(n10541), .B2(n8539), .C1(n8537), .C2(n8855), .ZN(P1_U3331) );
  OAI222_X1 U9624 ( .A1(n8831), .A2(n8540), .B1(n8691), .B2(n8539), .C1(n5939), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U9625 ( .A1(n8545), .A2(n9794), .ZN(n8542) );
  OAI211_X1 U9626 ( .C1(n8543), .C2(n8831), .A(n8542), .B(n8541), .ZN(P2_U3335) );
  NAND2_X1 U9627 ( .A1(n8545), .A2(n8544), .ZN(n8547) );
  OR2_X1 U9628 ( .A1(n8546), .A2(P1_U3084), .ZN(n10196) );
  OAI211_X1 U9629 ( .C1(n8548), .C2(n8855), .A(n8547), .B(n10196), .ZN(
        P1_U3330) );
  XNOR2_X1 U9630 ( .A(n8551), .B(n8550), .ZN(n8552) );
  XNOR2_X1 U9631 ( .A(n8549), .B(n8552), .ZN(n8558) );
  INV_X1 U9632 ( .A(n10870), .ZN(n8619) );
  NOR2_X1 U9633 ( .A1(n8619), .A2(n9919), .ZN(n8553) );
  AOI211_X1 U9634 ( .C1(n9923), .C2(n10871), .A(n8554), .B(n8553), .ZN(n8555)
         );
  OAI21_X1 U9635 ( .B1(n9926), .B2(n10882), .A(n8555), .ZN(n8556) );
  AOI21_X1 U9636 ( .B1(n10884), .B2(n9928), .A(n8556), .ZN(n8557) );
  OAI21_X1 U9637 ( .B1(n8558), .B2(n9931), .A(n8557), .ZN(P1_U3222) );
  OAI21_X1 U9638 ( .B1(n8567), .B2(n8560), .A(n8559), .ZN(n8561) );
  AOI222_X1 U9639 ( .A1(n9644), .A2(n8561), .B1(n9387), .B2(n9638), .C1(n9389), 
        .C2(n9619), .ZN(n8595) );
  INV_X1 U9640 ( .A(n8562), .ZN(n8566) );
  NOR2_X1 U9641 ( .A1(n8564), .A2(n9389), .ZN(n8565) );
  AOI21_X1 U9642 ( .B1(n8566), .B2(n6338), .A(n8565), .ZN(n8568) );
  NAND2_X1 U9643 ( .A1(n8568), .A2(n5291), .ZN(n8607) );
  OAI21_X1 U9644 ( .B1(n8568), .B2(n5291), .A(n8607), .ZN(n8596) );
  OAI22_X1 U9645 ( .A1(n10856), .A2(n8570), .B1(n8569), .B2(n10860), .ZN(n8571) );
  AOI21_X1 U9646 ( .B1(n8605), .B2(n9655), .A(n8571), .ZN(n8575) );
  NAND2_X1 U9647 ( .A1(n8572), .A2(n8605), .ZN(n8573) );
  AND2_X1 U9648 ( .A1(n8608), .A2(n8573), .ZN(n8593) );
  NAND2_X1 U9649 ( .A1(n8593), .A2(n9610), .ZN(n8574) );
  OAI211_X1 U9650 ( .C1(n8596), .C2(n9602), .A(n8575), .B(n8574), .ZN(n8576)
         );
  INV_X1 U9651 ( .A(n8576), .ZN(n8577) );
  OAI21_X1 U9652 ( .B1(n10851), .B2(n8595), .A(n8577), .ZN(P2_U3283) );
  INV_X1 U9653 ( .A(n8578), .ZN(n8582) );
  OAI222_X1 U9654 ( .A1(n8691), .A2(n8582), .B1(P2_U3152), .B2(n8580), .C1(
        n8579), .C2(n8831), .ZN(P2_U3334) );
  OAI222_X1 U9655 ( .A1(n8583), .A2(P1_U3084), .B1(n10541), .B2(n8582), .C1(
        n8581), .C2(n8855), .ZN(P1_U3329) );
  INV_X1 U9656 ( .A(n8656), .ZN(n10915) );
  OAI21_X1 U9657 ( .B1(n8586), .B2(n8585), .A(n8584), .ZN(n8587) );
  NAND2_X1 U9658 ( .A1(n8587), .A2(n9352), .ZN(n8592) );
  INV_X1 U9659 ( .A(n8588), .ZN(n8590) );
  OAI22_X1 U9660 ( .A1(n9365), .A2(n8604), .B1(n9363), .B2(n8611), .ZN(n8589)
         );
  AOI211_X1 U9661 ( .C1(n9334), .C2(n9386), .A(n8590), .B(n8589), .ZN(n8591)
         );
  OAI211_X1 U9662 ( .C1(n10915), .C2(n9358), .A(n8592), .B(n8591), .ZN(
        P2_U3217) );
  INV_X1 U9663 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8598) );
  AOI22_X1 U9664 ( .A1(n8593), .A2(n9746), .B1(n9745), .B2(n8605), .ZN(n8594)
         );
  OAI211_X1 U9665 ( .C1(n8596), .C2(n9750), .A(n8595), .B(n8594), .ZN(n8599)
         );
  NAND2_X1 U9666 ( .A1(n8599), .A2(n5011), .ZN(n8597) );
  OAI21_X1 U9667 ( .B1(n5011), .B2(n8598), .A(n8597), .ZN(P2_U3490) );
  NAND2_X1 U9668 ( .A1(n8599), .A2(n10923), .ZN(n8600) );
  OAI21_X1 U9669 ( .B1(n10923), .B2(n7614), .A(n8600), .ZN(P2_U3533) );
  XNOR2_X1 U9670 ( .A(n8602), .B(n8601), .ZN(n8603) );
  OAI222_X1 U9671 ( .A1(n9565), .A2(n9642), .B1(n9641), .B2(n8604), .C1(n9561), 
        .C2(n8603), .ZN(n10918) );
  INV_X1 U9672 ( .A(n10918), .ZN(n8618) );
  NAND2_X1 U9673 ( .A1(n8605), .A2(n9388), .ZN(n8606) );
  NAND2_X1 U9674 ( .A1(n8607), .A2(n8606), .ZN(n8659) );
  XNOR2_X1 U9675 ( .A(n8659), .B(n8658), .ZN(n10920) );
  INV_X1 U9676 ( .A(n8608), .ZN(n8610) );
  INV_X1 U9677 ( .A(n8609), .ZN(n8650) );
  OAI21_X1 U9678 ( .B1(n10915), .B2(n8610), .A(n8650), .ZN(n10917) );
  OAI22_X1 U9679 ( .A1(n10856), .A2(n8612), .B1(n8611), .B2(n10860), .ZN(n8613) );
  AOI21_X1 U9680 ( .B1(n8656), .B2(n9655), .A(n8613), .ZN(n8614) );
  OAI21_X1 U9681 ( .B1(n10917), .B2(n8615), .A(n8614), .ZN(n8616) );
  AOI21_X1 U9682 ( .B1(n10920), .B2(n9660), .A(n8616), .ZN(n8617) );
  OAI21_X1 U9683 ( .B1(n8618), .B2(n10851), .A(n8617), .ZN(P2_U3282) );
  OR2_X1 U9684 ( .A1(n8683), .A2(n8619), .ZN(n10076) );
  NAND2_X1 U9685 ( .A1(n8683), .A2(n8619), .ZN(n10074) );
  OR2_X1 U9686 ( .A1(n10884), .A2(n8621), .ZN(n10069) );
  INV_X1 U9687 ( .A(n10069), .ZN(n8622) );
  NAND2_X1 U9688 ( .A1(n10884), .A2(n8621), .ZN(n10073) );
  OAI21_X1 U9689 ( .B1(n10166), .B2(n8623), .A(n8675), .ZN(n8624) );
  AOI222_X1 U9690 ( .A1(n10947), .A2(n8624), .B1(n10203), .B2(n10942), .C1(
        n10204), .C2(n10944), .ZN(n10901) );
  NAND2_X1 U9691 ( .A1(n8625), .A2(n9948), .ZN(n8628) );
  OR2_X1 U9692 ( .A1(n8626), .A2(n10871), .ZN(n8627) );
  INV_X1 U9693 ( .A(n10862), .ZN(n8630) );
  NAND2_X1 U9694 ( .A1(n10884), .A2(n10204), .ZN(n8631) );
  OAI21_X1 U9695 ( .B1(n5083), .B2(n5385), .A(n8684), .ZN(n10904) );
  NAND2_X1 U9696 ( .A1(n10904), .A2(n10964), .ZN(n8637) );
  OAI22_X1 U9697 ( .A1(n10822), .A2(n8632), .B1(n8671), .B2(n10819), .ZN(n8635) );
  INV_X1 U9698 ( .A(n10884), .ZN(n10867) );
  INV_X1 U9699 ( .A(n10865), .ZN(n8633) );
  INV_X1 U9700 ( .A(n8683), .ZN(n10899) );
  OAI21_X1 U9701 ( .B1(n8633), .B2(n10899), .A(n8678), .ZN(n10900) );
  NOR2_X1 U9702 ( .A1(n10900), .A2(n10429), .ZN(n8634) );
  AOI211_X1 U9703 ( .C1(n10959), .C2(n8683), .A(n8635), .B(n8634), .ZN(n8636)
         );
  OAI211_X1 U9704 ( .C1(n10969), .C2(n10901), .A(n8637), .B(n8636), .ZN(
        P1_U3278) );
  OAI21_X1 U9705 ( .B1(n8640), .B2(n8639), .A(n8638), .ZN(n8641) );
  NAND2_X1 U9706 ( .A1(n8641), .A2(n9352), .ZN(n8647) );
  INV_X1 U9707 ( .A(n8642), .ZN(n8645) );
  OAI22_X1 U9708 ( .A1(n9365), .A2(n8643), .B1(n9363), .B2(n8652), .ZN(n8644)
         );
  AOI211_X1 U9709 ( .C1(n9334), .C2(n9618), .A(n8645), .B(n8644), .ZN(n8646)
         );
  OAI211_X1 U9710 ( .C1(n8651), .C2(n9358), .A(n8647), .B(n8646), .ZN(P2_U3243) );
  XNOR2_X1 U9711 ( .A(n8648), .B(n8660), .ZN(n8649) );
  AOI222_X1 U9712 ( .A1(n9644), .A2(n8649), .B1(n9618), .B2(n9638), .C1(n9387), 
        .C2(n9619), .ZN(n9749) );
  AOI21_X1 U9713 ( .B1(n9744), .B2(n8650), .A(n9651), .ZN(n9747) );
  NOR2_X1 U9714 ( .A1(n8651), .A2(n9628), .ZN(n8655) );
  OAI22_X1 U9715 ( .A1(n10856), .A2(n8653), .B1(n8652), .B2(n10860), .ZN(n8654) );
  AOI211_X1 U9716 ( .C1(n9747), .C2(n9610), .A(n8655), .B(n8654), .ZN(n8663)
         );
  OR2_X1 U9717 ( .A1(n8656), .A2(n9387), .ZN(n8657) );
  OAI21_X1 U9718 ( .B1(n8661), .B2(n8660), .A(n8801), .ZN(n9743) );
  NAND2_X1 U9719 ( .A1(n9743), .A2(n9660), .ZN(n8662) );
  OAI211_X1 U9720 ( .C1(n9749), .C2(n10851), .A(n8663), .B(n8662), .ZN(
        P2_U3281) );
  AOI21_X1 U9721 ( .B1(n8667), .B2(n8665), .A(n8664), .ZN(n8666) );
  AOI21_X1 U9722 ( .B1(n5085), .B2(n8667), .A(n8666), .ZN(n8674) );
  INV_X1 U9723 ( .A(n10203), .ZN(n8719) );
  NOR2_X1 U9724 ( .A1(n8719), .A2(n9919), .ZN(n8668) );
  AOI211_X1 U9725 ( .C1(n9923), .C2(n10204), .A(n8669), .B(n8668), .ZN(n8670)
         );
  OAI21_X1 U9726 ( .B1(n9926), .B2(n8671), .A(n8670), .ZN(n8672) );
  AOI21_X1 U9727 ( .B1(n8683), .B2(n9928), .A(n8672), .ZN(n8673) );
  OAI21_X1 U9728 ( .B1(n8674), .B2(n9931), .A(n8673), .ZN(P1_U3232) );
  NAND2_X1 U9729 ( .A1(n9809), .A2(n8719), .ZN(n10035) );
  XOR2_X1 U9730 ( .A(n8714), .B(n10168), .Z(n8676) );
  AOI222_X1 U9731 ( .A1(n10947), .A2(n8676), .B1(n10945), .B2(n10942), .C1(
        n10870), .C2(n10944), .ZN(n10908) );
  OAI22_X1 U9732 ( .A1(n10822), .A2(n8677), .B1(n9807), .B2(n10819), .ZN(n8682) );
  INV_X1 U9733 ( .A(n9809), .ZN(n10909) );
  INV_X1 U9734 ( .A(n8678), .ZN(n8679) );
  OAI211_X1 U9735 ( .C1(n10909), .C2(n8679), .A(n5325), .B(n10973), .ZN(n10907) );
  INV_X1 U9736 ( .A(n10962), .ZN(n8680) );
  NOR2_X1 U9737 ( .A1(n10907), .A2(n8680), .ZN(n8681) );
  AOI211_X1 U9738 ( .C1(n10959), .C2(n9809), .A(n8682), .B(n8681), .ZN(n8686)
         );
  XNOR2_X1 U9739 ( .A(n8709), .B(n10168), .ZN(n10911) );
  NAND2_X1 U9740 ( .A1(n10911), .A2(n10964), .ZN(n8685) );
  OAI211_X1 U9741 ( .C1(n10908), .C2(n10969), .A(n8686), .B(n8685), .ZN(
        P1_U3277) );
  INV_X1 U9742 ( .A(n8687), .ZN(n8690) );
  OAI222_X1 U9743 ( .A1(P1_U3084), .A2(n8688), .B1(n10541), .B2(n8690), .C1(
        n9195), .C2(n8855), .ZN(P1_U3328) );
  OAI222_X1 U9744 ( .A1(n8831), .A2(n8692), .B1(n8691), .B2(n8690), .C1(n8689), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI21_X1 U9745 ( .B1(n8695), .B2(n8694), .A(n8693), .ZN(n8696) );
  NAND2_X1 U9746 ( .A1(n8696), .A2(n9352), .ZN(n8701) );
  INV_X1 U9747 ( .A(n8697), .ZN(n8699) );
  OAI22_X1 U9748 ( .A1(n9365), .A2(n9642), .B1(n9363), .B2(n9652), .ZN(n8698)
         );
  AOI211_X1 U9749 ( .C1(n9334), .C2(n9639), .A(n8699), .B(n8698), .ZN(n8700)
         );
  OAI211_X1 U9750 ( .C1(n9787), .C2(n9358), .A(n8701), .B(n8700), .ZN(P2_U3228) );
  INV_X1 U9751 ( .A(n8702), .ZN(n8705) );
  OAI222_X1 U9752 ( .A1(n8691), .A2(n8705), .B1(P2_U3152), .B2(n8704), .C1(
        n8703), .C2(n8831), .ZN(P2_U3332) );
  OAI222_X1 U9753 ( .A1(n8706), .A2(n5013), .B1(n10541), .B2(n8705), .C1(n9191), .C2(n8855), .ZN(P1_U3327) );
  INV_X1 U9754 ( .A(n8707), .ZN(n8727) );
  OAI222_X1 U9755 ( .A1(n8691), .A2(n8727), .B1(n5941), .B2(P2_U3152), .C1(
        n8708), .C2(n8831), .ZN(P2_U3331) );
  INV_X1 U9756 ( .A(n10945), .ZN(n9803) );
  OR2_X1 U9757 ( .A1(n9929), .A2(n9803), .ZN(n10081) );
  NAND2_X1 U9758 ( .A1(n9929), .A2(n9803), .ZN(n10036) );
  NAND2_X1 U9759 ( .A1(n8709), .A2(n10168), .ZN(n8711) );
  OR2_X1 U9760 ( .A1(n9809), .A2(n10203), .ZN(n8710) );
  INV_X1 U9761 ( .A(n8752), .ZN(n8712) );
  AOI21_X1 U9762 ( .B1(n9964), .B2(n8713), .A(n8712), .ZN(n10931) );
  INV_X1 U9763 ( .A(n10931), .ZN(n8726) );
  INV_X1 U9764 ( .A(n10436), .ZN(n9920) );
  INV_X1 U9765 ( .A(n9964), .ZN(n10169) );
  NAND2_X1 U9766 ( .A1(n8715), .A2(n10077), .ZN(n8717) );
  OR2_X2 U9767 ( .A1(n8717), .A2(n10169), .ZN(n8771) );
  INV_X1 U9768 ( .A(n8771), .ZN(n8716) );
  AOI21_X1 U9769 ( .B1(n10169), .B2(n8717), .A(n8716), .ZN(n8718) );
  OAI222_X1 U9770 ( .A1(n10403), .A2(n9920), .B1(n10401), .B2(n8719), .C1(
        n10873), .C2(n8718), .ZN(n10929) );
  INV_X1 U9771 ( .A(n9929), .ZN(n10926) );
  INV_X1 U9772 ( .A(n10949), .ZN(n8720) );
  OAI21_X1 U9773 ( .B1(n10926), .B2(n8721), .A(n8720), .ZN(n10928) );
  OAI22_X1 U9774 ( .A1(n10822), .A2(n8115), .B1(n9925), .B2(n10819), .ZN(n8722) );
  AOI21_X1 U9775 ( .B1(n9929), .B2(n10959), .A(n8722), .ZN(n8723) );
  OAI21_X1 U9776 ( .B1(n10928), .B2(n10429), .A(n8723), .ZN(n8724) );
  AOI21_X1 U9777 ( .B1(n10929), .B2(n10822), .A(n8724), .ZN(n8725) );
  OAI21_X1 U9778 ( .B1(n8726), .B2(n10406), .A(n8725), .ZN(P1_U3276) );
  OAI222_X1 U9779 ( .A1(n5013), .A2(n7155), .B1(n10541), .B2(n8727), .C1(n9190), .C2(n8855), .ZN(P1_U3326) );
  NAND2_X1 U9780 ( .A1(n8834), .A2(n6723), .ZN(n8729) );
  INV_X1 U9781 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8856) );
  OR2_X1 U9782 ( .A1(n8823), .A2(n8856), .ZN(n8728) );
  NAND2_X1 U9783 ( .A1(n10457), .A2(n7058), .ZN(n8731) );
  INV_X1 U9784 ( .A(n10272), .ZN(n10200) );
  NAND2_X1 U9785 ( .A1(n10200), .A2(n6977), .ZN(n8730) );
  NAND2_X1 U9786 ( .A1(n8731), .A2(n8730), .ZN(n8733) );
  XNOR2_X1 U9787 ( .A(n8733), .B(n8732), .ZN(n8737) );
  NOR2_X1 U9788 ( .A1(n10272), .A2(n6764), .ZN(n8734) );
  AOI21_X1 U9789 ( .B1(n10457), .B2(n8735), .A(n8734), .ZN(n8736) );
  XNOR2_X1 U9790 ( .A(n8737), .B(n8736), .ZN(n8743) );
  INV_X1 U9791 ( .A(n8743), .ZN(n8738) );
  NAND2_X1 U9792 ( .A1(n8738), .A2(n9893), .ZN(n8749) );
  INV_X1 U9793 ( .A(n8739), .ZN(n8742) );
  NAND4_X1 U9794 ( .A1(n8748), .A2(n9893), .A3(n8742), .A4(n8743), .ZN(n8747)
         );
  AOI22_X1 U9795 ( .A1(n9906), .A2(n8769), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8741) );
  NAND2_X1 U9796 ( .A1(n9923), .A2(n10287), .ZN(n8740) );
  OAI211_X1 U9797 ( .C1(n9926), .C2(n8849), .A(n8741), .B(n8740), .ZN(n8745)
         );
  NOR3_X1 U9798 ( .A1(n8743), .A2(n8742), .A3(n9931), .ZN(n8744) );
  AOI211_X1 U9799 ( .C1(n9928), .C2(n10457), .A(n8745), .B(n8744), .ZN(n8746)
         );
  OAI211_X1 U9800 ( .C1(n8749), .C2(n8748), .A(n8747), .B(n8746), .ZN(P1_U3218) );
  INV_X1 U9801 ( .A(n8766), .ZN(n8793) );
  OAI222_X1 U9802 ( .A1(n8691), .A2(n8793), .B1(n8831), .B2(n5754), .C1(
        P2_U3152), .C2(n8750), .ZN(P2_U3329) );
  NAND2_X1 U9803 ( .A1(n9929), .A2(n10945), .ZN(n8751) );
  OR2_X1 U9804 ( .A1(n10960), .A2(n9920), .ZN(n10082) );
  NAND2_X1 U9805 ( .A1(n10960), .A2(n9920), .ZN(n10031) );
  NAND2_X1 U9806 ( .A1(n10082), .A2(n10031), .ZN(n10936) );
  NAND2_X1 U9807 ( .A1(n10960), .A2(n10436), .ZN(n8753) );
  INV_X1 U9808 ( .A(n10943), .ZN(n8754) );
  NAND2_X1 U9809 ( .A1(n10516), .A2(n8754), .ZN(n10032) );
  INV_X1 U9810 ( .A(n10435), .ZN(n10400) );
  OR2_X1 U9811 ( .A1(n10426), .A2(n10400), .ZN(n10025) );
  NAND2_X1 U9812 ( .A1(n10426), .A2(n10400), .ZN(n10034) );
  OR2_X1 U9813 ( .A1(n10516), .A2(n10943), .ZN(n10409) );
  AND2_X1 U9814 ( .A1(n10414), .A2(n10409), .ZN(n8755) );
  INV_X1 U9815 ( .A(n10506), .ZN(n10391) );
  XNOR2_X1 U9816 ( .A(n10500), .B(n10359), .ZN(n10372) );
  INV_X1 U9817 ( .A(n10359), .ZN(n10402) );
  INV_X1 U9818 ( .A(n10500), .ZN(n10383) );
  INV_X1 U9819 ( .A(n10374), .ZN(n10347) );
  OR2_X1 U9820 ( .A1(n10496), .A2(n10347), .ZN(n9978) );
  NAND2_X1 U9821 ( .A1(n10496), .A2(n10347), .ZN(n9977) );
  NAND2_X1 U9822 ( .A1(n9978), .A2(n9977), .ZN(n10357) );
  NAND2_X1 U9823 ( .A1(n10491), .A2(n10335), .ZN(n8761) );
  INV_X1 U9824 ( .A(n10491), .ZN(n8760) );
  INV_X1 U9825 ( .A(n10335), .ZN(n10362) );
  NAND2_X1 U9826 ( .A1(n10323), .A2(n8762), .ZN(n8763) );
  INV_X1 U9827 ( .A(n10481), .ZN(n8784) );
  INV_X1 U9828 ( .A(n10334), .ZN(n10302) );
  NOR2_X1 U9829 ( .A1(n8784), .A2(n10302), .ZN(n8764) );
  NAND2_X1 U9830 ( .A1(n10474), .A2(n10315), .ZN(n10105) );
  INV_X1 U9831 ( .A(n10474), .ZN(n10298) );
  INV_X1 U9832 ( .A(n10469), .ZN(n10283) );
  NAND2_X1 U9833 ( .A1(n10283), .A2(n10303), .ZN(n8765) );
  NAND2_X1 U9834 ( .A1(n10464), .A2(n8843), .ZN(n10101) );
  NAND2_X1 U9835 ( .A1(n8839), .A2(n5595), .ZN(n8770) );
  NAND2_X1 U9836 ( .A1(n8766), .A2(n6723), .ZN(n8768) );
  INV_X1 U9837 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8792) );
  OR2_X1 U9838 ( .A1(n8823), .A2(n8792), .ZN(n8767) );
  INV_X1 U9839 ( .A(n8769), .ZN(n8844) );
  NAND2_X1 U9840 ( .A1(n8785), .A2(n8844), .ZN(n10144) );
  NAND2_X1 U9841 ( .A1(n10005), .A2(n10144), .ZN(n10151) );
  NAND2_X1 U9842 ( .A1(n8771), .A2(n10036), .ZN(n10940) );
  INV_X1 U9843 ( .A(n10936), .ZN(n10941) );
  INV_X1 U9844 ( .A(n10034), .ZN(n8773) );
  OR2_X1 U9845 ( .A1(n10506), .A2(n9898), .ZN(n10027) );
  NAND2_X1 U9846 ( .A1(n10506), .A2(n9898), .ZN(n10132) );
  NAND2_X1 U9847 ( .A1(n10027), .A2(n10132), .ZN(n10397) );
  INV_X1 U9848 ( .A(n10132), .ZN(n8774) );
  OR2_X1 U9849 ( .A1(n10500), .A2(n10402), .ZN(n10355) );
  AND2_X1 U9850 ( .A1(n9978), .A2(n10355), .ZN(n10030) );
  INV_X1 U9851 ( .A(n9977), .ZN(n9975) );
  NAND2_X1 U9852 ( .A1(n10491), .A2(n10362), .ZN(n10090) );
  OR2_X1 U9853 ( .A1(n10484), .A2(n10348), .ZN(n9988) );
  OR2_X1 U9854 ( .A1(n10491), .A2(n10362), .ZN(n10330) );
  AND2_X1 U9855 ( .A1(n9988), .A2(n10330), .ZN(n10117) );
  NAND2_X1 U9856 ( .A1(n10481), .A2(n10302), .ZN(n9991) );
  NAND2_X1 U9857 ( .A1(n10484), .A2(n10348), .ZN(n10310) );
  AND2_X1 U9858 ( .A1(n9991), .A2(n10310), .ZN(n10138) );
  NOR2_X1 U9859 ( .A1(n10481), .A2(n10302), .ZN(n10023) );
  INV_X1 U9860 ( .A(n10020), .ZN(n8775) );
  OR2_X1 U9861 ( .A1(n10469), .A2(n10303), .ZN(n10021) );
  NAND2_X1 U9862 ( .A1(n10469), .A2(n10303), .ZN(n10098) );
  INV_X1 U9863 ( .A(n10100), .ZN(n10001) );
  NOR2_X1 U9864 ( .A1(n8842), .A2(n10178), .ZN(n8841) );
  INV_X1 U9865 ( .A(n10004), .ZN(n8776) );
  XNOR2_X1 U9866 ( .A(n8777), .B(n10151), .ZN(n8781) );
  INV_X1 U9867 ( .A(P1_B_REG_SCAN_IN), .ZN(n10199) );
  NOR2_X1 U9868 ( .A1(n7155), .A2(n10199), .ZN(n8778) );
  OR2_X1 U9869 ( .A1(n10403), .A2(n8778), .ZN(n8826) );
  OAI21_X1 U9870 ( .B1(n8781), .B2(n10873), .A(n8780), .ZN(n10454) );
  INV_X1 U9871 ( .A(n10960), .ZN(n10950) );
  NAND2_X1 U9872 ( .A1(n10949), .A2(n10950), .ZN(n10948) );
  INV_X1 U9873 ( .A(n8783), .ZN(n10354) );
  NOR2_X2 U9874 ( .A1(n10469), .A2(n10294), .ZN(n10279) );
  INV_X1 U9875 ( .A(n8785), .ZN(n10451) );
  OAI21_X1 U9876 ( .B1(n5031), .B2(n10451), .A(n10257), .ZN(n10452) );
  NOR2_X1 U9877 ( .A1(n10452), .A2(n10429), .ZN(n8790) );
  INV_X1 U9878 ( .A(n8786), .ZN(n8787) );
  AOI22_X1 U9879 ( .A1(n10969), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n10957), 
        .B2(n8787), .ZN(n8788) );
  OAI21_X1 U9880 ( .B1(n10451), .B2(n10792), .A(n8788), .ZN(n8789) );
  AOI211_X1 U9881 ( .C1(n10454), .C2(n10822), .A(n8790), .B(n8789), .ZN(n8791)
         );
  OAI21_X1 U9882 ( .B1(n10455), .B2(n10406), .A(n8791), .ZN(P1_U3355) );
  OAI222_X1 U9883 ( .A1(P1_U3084), .A2(n8794), .B1(n10541), .B2(n8793), .C1(
        n8792), .C2(n8855), .ZN(P1_U3324) );
  NAND2_X1 U9884 ( .A1(n8795), .A2(n9893), .ZN(n8798) );
  AOI22_X1 U9885 ( .A1(n9906), .A2(n7836), .B1(n8796), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n8797) );
  OAI211_X1 U9886 ( .C1(n9903), .C2(n8799), .A(n8798), .B(n8797), .ZN(P1_U3230) );
  INV_X1 U9887 ( .A(n9700), .ZN(n9527) );
  OR2_X1 U9888 ( .A1(n9744), .A2(n9386), .ZN(n8800) );
  OR2_X1 U9889 ( .A1(n9727), .A2(n9620), .ZN(n8803) );
  OAI21_X1 U9890 ( .B1(n9444), .B2(n9679), .A(n8808), .ZN(n9435) );
  INV_X1 U9891 ( .A(n9674), .ZN(n9440) );
  AOI22_X1 U9892 ( .A1(n9435), .A2(n8809), .B1(n8862), .B2(n9440), .ZN(n8810)
         );
  XNOR2_X1 U9893 ( .A(n8810), .B(n8815), .ZN(n9673) );
  AOI21_X1 U9894 ( .B1(n9668), .B2(n9436), .A(n9431), .ZN(n9669) );
  INV_X1 U9895 ( .A(n9668), .ZN(n8814) );
  INV_X1 U9896 ( .A(n8811), .ZN(n8812) );
  AOI22_X1 U9897 ( .A1(n8812), .A2(n10755), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10851), .ZN(n8813) );
  OAI21_X1 U9898 ( .B1(n8814), .B2(n9628), .A(n8813), .ZN(n8818) );
  INV_X1 U9899 ( .A(n8862), .ZN(n9468) );
  NOR2_X1 U9900 ( .A1(n9671), .A2(n10851), .ZN(n8817) );
  AOI211_X1 U9901 ( .C1(n9669), .C2(n9610), .A(n8818), .B(n8817), .ZN(n8819)
         );
  OAI21_X1 U9902 ( .B1(n9673), .B2(n9602), .A(n8819), .ZN(P2_U3267) );
  NAND2_X1 U9903 ( .A1(n8830), .A2(n6723), .ZN(n8821) );
  INV_X1 U9904 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8837) );
  OR2_X1 U9905 ( .A1(n8823), .A2(n8837), .ZN(n8820) );
  NAND2_X1 U9906 ( .A1(n10537), .A2(n6723), .ZN(n8825) );
  INV_X1 U9907 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8822) );
  OR2_X1 U9908 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  XNOR2_X1 U9909 ( .A(n10256), .B(n10011), .ZN(n10450) );
  NOR2_X1 U9910 ( .A1(n10012), .A2(n8826), .ZN(n10972) );
  INV_X1 U9911 ( .A(n10972), .ZN(n8827) );
  NOR2_X1 U9912 ( .A1(n8827), .A2(n10969), .ZN(n10259) );
  NOR2_X1 U9913 ( .A1(n10011), .A2(n10792), .ZN(n8828) );
  AOI211_X1 U9914 ( .C1(n10969), .C2(P1_REG2_REG_31__SCAN_IN), .A(n10259), .B(
        n8828), .ZN(n8829) );
  OAI21_X1 U9915 ( .B1(n10429), .B2(n10450), .A(n8829), .ZN(P1_U3261) );
  INV_X1 U9916 ( .A(n8830), .ZN(n8838) );
  OAI222_X1 U9917 ( .A1(n8691), .A2(n8838), .B1(n8833), .B2(P2_U3152), .C1(
        n8832), .C2(n8831), .ZN(P2_U3328) );
  INV_X1 U9918 ( .A(n8834), .ZN(n8857) );
  OAI222_X1 U9919 ( .A1(n8691), .A2(n8857), .B1(n5940), .B2(P2_U3152), .C1(
        n8835), .C2(n8831), .ZN(P2_U3330) );
  OAI222_X1 U9920 ( .A1(n5013), .A2(n8836), .B1(n10541), .B2(n8838), .C1(n8837), .C2(n8855), .ZN(P1_U3323) );
  AOI211_X1 U9921 ( .C1(n8842), .C2(n10178), .A(n10873), .B(n8841), .ZN(n8846)
         );
  OAI22_X1 U9922 ( .A1(n8844), .A2(n10403), .B1(n8843), .B2(n10401), .ZN(n8845) );
  NOR2_X1 U9923 ( .A1(n8846), .A2(n8845), .ZN(n8847) );
  OAI21_X1 U9924 ( .B1(n10460), .B2(n8848), .A(n8847), .ZN(n10456) );
  NAND2_X1 U9925 ( .A1(n10456), .A2(n10822), .ZN(n8854) );
  AOI21_X1 U9926 ( .B1(n10457), .B2(n10263), .A(n5031), .ZN(n10458) );
  INV_X1 U9927 ( .A(n8849), .ZN(n8850) );
  AOI22_X1 U9928 ( .A1(n10969), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n10957), 
        .B2(n8850), .ZN(n8851) );
  OAI21_X1 U9929 ( .B1(n5333), .B2(n10792), .A(n8851), .ZN(n8852) );
  AOI21_X1 U9930 ( .B1(n10458), .B2(n10786), .A(n8852), .ZN(n8853) );
  OAI211_X1 U9931 ( .C1(n10385), .C2(n10460), .A(n8854), .B(n8853), .ZN(
        P1_U3263) );
  OAI222_X1 U9932 ( .A1(P1_U3084), .A2(n7127), .B1(n10541), .B2(n8857), .C1(
        n8856), .C2(n8855), .ZN(P1_U3325) );
  XNOR2_X1 U9933 ( .A(n8859), .B(n8858), .ZN(n8865) );
  OAI22_X1 U9934 ( .A1(n9455), .A2(n9363), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8923), .ZN(n8860) );
  AOI21_X1 U9935 ( .B1(n9335), .B2(n9384), .A(n8860), .ZN(n8861) );
  OAI21_X1 U9936 ( .B1(n8862), .B2(n9362), .A(n8861), .ZN(n8863) );
  AOI21_X1 U9937 ( .B1(n9679), .B2(n9379), .A(n8863), .ZN(n8864) );
  OAI21_X1 U9938 ( .B1(n8865), .B2(n9381), .A(n8864), .ZN(n9290) );
  XNOR2_X1 U9939 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .ZN(n8868) );
  XNOR2_X1 U9940 ( .A(SI_31_), .B(keyinput_129), .ZN(n8867) );
  XNOR2_X1 U9941 ( .A(SI_30_), .B(keyinput_130), .ZN(n8866) );
  OAI21_X1 U9942 ( .B1(n8868), .B2(n8867), .A(n8866), .ZN(n8871) );
  XNOR2_X1 U9943 ( .A(n9075), .B(keyinput_131), .ZN(n8870) );
  XNOR2_X1 U9944 ( .A(SI_28_), .B(keyinput_132), .ZN(n8869) );
  AOI21_X1 U9945 ( .B1(n8871), .B2(n8870), .A(n8869), .ZN(n8880) );
  XNOR2_X1 U9946 ( .A(n8872), .B(keyinput_134), .ZN(n8879) );
  XNOR2_X1 U9947 ( .A(SI_27_), .B(keyinput_133), .ZN(n8876) );
  XNOR2_X1 U9948 ( .A(SI_23_), .B(keyinput_137), .ZN(n8875) );
  XNOR2_X1 U9949 ( .A(SI_25_), .B(keyinput_135), .ZN(n8874) );
  XNOR2_X1 U9950 ( .A(SI_22_), .B(keyinput_138), .ZN(n8873) );
  NAND4_X1 U9951 ( .A1(n8876), .A2(n8875), .A3(n8874), .A4(n8873), .ZN(n8878)
         );
  XNOR2_X1 U9952 ( .A(SI_24_), .B(keyinput_136), .ZN(n8877) );
  NOR4_X1 U9953 ( .A1(n8880), .A2(n8879), .A3(n8878), .A4(n8877), .ZN(n8889)
         );
  XNOR2_X1 U9954 ( .A(n8881), .B(keyinput_139), .ZN(n8888) );
  XNOR2_X1 U9955 ( .A(SI_18_), .B(keyinput_142), .ZN(n8887) );
  XNOR2_X1 U9956 ( .A(n8882), .B(keyinput_140), .ZN(n8885) );
  XNOR2_X1 U9957 ( .A(n8883), .B(keyinput_141), .ZN(n8884) );
  NAND2_X1 U9958 ( .A1(n8885), .A2(n8884), .ZN(n8886) );
  NOR4_X1 U9959 ( .A1(n8889), .A2(n8888), .A3(n8887), .A4(n8886), .ZN(n8897)
         );
  XNOR2_X1 U9960 ( .A(SI_17_), .B(keyinput_143), .ZN(n8896) );
  XNOR2_X1 U9961 ( .A(n9094), .B(keyinput_147), .ZN(n8894) );
  XNOR2_X1 U9962 ( .A(n8890), .B(keyinput_145), .ZN(n8893) );
  XNOR2_X1 U9963 ( .A(SI_16_), .B(keyinput_144), .ZN(n8892) );
  XNOR2_X1 U9964 ( .A(SI_14_), .B(keyinput_146), .ZN(n8891) );
  NOR4_X1 U9965 ( .A1(n8894), .A2(n8893), .A3(n8892), .A4(n8891), .ZN(n8895)
         );
  OAI21_X1 U9966 ( .B1(n8897), .B2(n8896), .A(n8895), .ZN(n8902) );
  XNOR2_X1 U9967 ( .A(n9102), .B(keyinput_149), .ZN(n8901) );
  XNOR2_X1 U9968 ( .A(n8898), .B(keyinput_150), .ZN(n8900) );
  XNOR2_X1 U9969 ( .A(n9101), .B(keyinput_148), .ZN(n8899) );
  NAND4_X1 U9970 ( .A1(n8902), .A2(n8901), .A3(n8900), .A4(n8899), .ZN(n8905)
         );
  XNOR2_X1 U9971 ( .A(SI_9_), .B(keyinput_151), .ZN(n8904) );
  XNOR2_X1 U9972 ( .A(SI_8_), .B(keyinput_152), .ZN(n8903) );
  AOI21_X1 U9973 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8919) );
  XOR2_X1 U9974 ( .A(SI_7_), .B(keyinput_153), .Z(n8918) );
  INV_X1 U9975 ( .A(keyinput_160), .ZN(n8912) );
  AOI22_X1 U9976 ( .A1(SI_4_), .A2(keyinput_156), .B1(n9119), .B2(keyinput_157), .ZN(n8908) );
  AOI22_X1 U9977 ( .A1(n8906), .A2(keyinput_160), .B1(n8909), .B2(keyinput_155), .ZN(n8907) );
  OAI211_X1 U9978 ( .C1(SI_4_), .C2(keyinput_156), .A(n8908), .B(n8907), .ZN(
        n8911) );
  OAI22_X1 U9979 ( .A1(keyinput_155), .A2(n8909), .B1(n9119), .B2(keyinput_157), .ZN(n8910) );
  AOI211_X1 U9980 ( .C1(SI_0_), .C2(n8912), .A(n8911), .B(n8910), .ZN(n8916)
         );
  XNOR2_X1 U9981 ( .A(SI_2_), .B(keyinput_158), .ZN(n8915) );
  XNOR2_X1 U9982 ( .A(SI_6_), .B(keyinput_154), .ZN(n8914) );
  XNOR2_X1 U9983 ( .A(SI_1_), .B(keyinput_159), .ZN(n8913) );
  AND4_X1 U9984 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), .ZN(n8917)
         );
  OAI21_X1 U9985 ( .B1(n8919), .B2(n8918), .A(n8917), .ZN(n8922) );
  XOR2_X1 U9986 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_161), .Z(n8921) );
  XNOR2_X1 U9987 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_162), .ZN(n8920) );
  AOI21_X1 U9988 ( .B1(n8922), .B2(n8921), .A(n8920), .ZN(n8930) );
  XNOR2_X1 U9989 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n8929) );
  XOR2_X1 U9990 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .Z(n8927) );
  XNOR2_X1 U9991 ( .A(n8923), .B(keyinput_164), .ZN(n8926) );
  XNOR2_X1 U9992 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n8925)
         );
  XNOR2_X1 U9993 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n8924)
         );
  NOR4_X1 U9994 ( .A1(n8927), .A2(n8926), .A3(n8925), .A4(n8924), .ZN(n8928)
         );
  OAI21_X1 U9995 ( .B1(n8930), .B2(n8929), .A(n8928), .ZN(n8933) );
  XNOR2_X1 U9996 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n8932) );
  XNOR2_X1 U9997 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n8931)
         );
  AOI21_X1 U9998 ( .B1(n8933), .B2(n8932), .A(n8931), .ZN(n8937) );
  XNOR2_X1 U9999 ( .A(n8934), .B(keyinput_170), .ZN(n8936) );
  XNOR2_X1 U10000 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n8935)
         );
  OAI21_X1 U10001 ( .B1(n8937), .B2(n8936), .A(n8935), .ZN(n8942) );
  XOR2_X1 U10002 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .Z(n8941) );
  XNOR2_X1 U10003 ( .A(n8938), .B(keyinput_174), .ZN(n8940) );
  XNOR2_X1 U10004 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n8939)
         );
  AOI211_X1 U10005 ( .C1(n8942), .C2(n8941), .A(n8940), .B(n8939), .ZN(n8945)
         );
  XNOR2_X1 U10006 ( .A(n9320), .B(keyinput_175), .ZN(n8944) );
  XNOR2_X1 U10007 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n8943)
         );
  NOR3_X1 U10008 ( .A1(n8945), .A2(n8944), .A3(n8943), .ZN(n8953) );
  XNOR2_X1 U10009 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_177), .ZN(n8952)
         );
  XNOR2_X1 U10010 ( .A(n8946), .B(keyinput_181), .ZN(n8950) );
  XNOR2_X1 U10011 ( .A(n9156), .B(keyinput_180), .ZN(n8949) );
  XNOR2_X1 U10012 ( .A(n9157), .B(keyinput_179), .ZN(n8948) );
  XNOR2_X1 U10013 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n8947)
         );
  NOR4_X1 U10014 ( .A1(n8950), .A2(n8949), .A3(n8948), .A4(n8947), .ZN(n8951)
         );
  OAI21_X1 U10015 ( .B1(n8953), .B2(n8952), .A(n8951), .ZN(n8963) );
  XNOR2_X1 U10016 ( .A(n8954), .B(keyinput_184), .ZN(n8958) );
  XNOR2_X1 U10017 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_185), .ZN(n8957)
         );
  XNOR2_X1 U10018 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_183), .ZN(n8956)
         );
  XNOR2_X1 U10019 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n8955)
         );
  NOR4_X1 U10020 ( .A1(n8958), .A2(n8957), .A3(n8956), .A4(n8955), .ZN(n8962)
         );
  XNOR2_X1 U10021 ( .A(n8959), .B(keyinput_186), .ZN(n8961) );
  XNOR2_X1 U10022 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .ZN(n8960)
         );
  AOI211_X1 U10023 ( .C1(n8963), .C2(n8962), .A(n8961), .B(n8960), .ZN(n8966)
         );
  XNOR2_X1 U10024 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n8965)
         );
  XNOR2_X1 U10025 ( .A(n9175), .B(keyinput_189), .ZN(n8964) );
  OAI21_X1 U10026 ( .B1(n8966), .B2(n8965), .A(n8964), .ZN(n8971) );
  XNOR2_X1 U10027 ( .A(n9179), .B(keyinput_191), .ZN(n8970) );
  XNOR2_X1 U10028 ( .A(n8967), .B(keyinput_190), .ZN(n8969) );
  XNOR2_X1 U10029 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .ZN(n8968) );
  NAND4_X1 U10030 ( .A1(n8971), .A2(n8970), .A3(n8969), .A4(n8968), .ZN(n8974)
         );
  XOR2_X1 U10031 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .Z(n8973)
         );
  XOR2_X1 U10032 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .Z(n8972)
         );
  NAND3_X1 U10033 ( .A1(n8974), .A2(n8973), .A3(n8972), .ZN(n8977) );
  XNOR2_X1 U10034 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .ZN(n8976)
         );
  XNOR2_X1 U10035 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n8975)
         );
  NAND3_X1 U10036 ( .A1(n8977), .A2(n8976), .A3(n8975), .ZN(n8980) );
  XNOR2_X1 U10037 ( .A(n9190), .B(keyinput_197), .ZN(n8979) );
  XNOR2_X1 U10038 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .ZN(n8978)
         );
  NAND3_X1 U10039 ( .A1(n8980), .A2(n8979), .A3(n8978), .ZN(n8983) );
  XNOR2_X1 U10040 ( .A(n9195), .B(keyinput_199), .ZN(n8982) );
  XOR2_X1 U10041 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .Z(n8981)
         );
  AOI21_X1 U10042 ( .B1(n8983), .B2(n8982), .A(n8981), .ZN(n8986) );
  XNOR2_X1 U10043 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n8985)
         );
  XNOR2_X1 U10044 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .ZN(n8984)
         );
  NOR3_X1 U10045 ( .A1(n8986), .A2(n8985), .A3(n8984), .ZN(n8994) );
  XOR2_X1 U10046 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .Z(n8991)
         );
  XNOR2_X1 U10047 ( .A(n8987), .B(keyinput_205), .ZN(n8990) );
  XNOR2_X1 U10048 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_204), .ZN(n8989)
         );
  XNOR2_X1 U10049 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .ZN(n8988)
         );
  NAND4_X1 U10050 ( .A1(n8991), .A2(n8990), .A3(n8989), .A4(n8988), .ZN(n8993)
         );
  XNOR2_X1 U10051 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n8992)
         );
  OAI21_X1 U10052 ( .B1(n8994), .B2(n8993), .A(n8992), .ZN(n8997) );
  XNOR2_X1 U10053 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .ZN(n8996)
         );
  XNOR2_X1 U10054 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n8995)
         );
  NAND3_X1 U10055 ( .A1(n8997), .A2(n8996), .A3(n8995), .ZN(n9002) );
  XOR2_X1 U10056 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .Z(n9001)
         );
  XNOR2_X1 U10057 ( .A(n8998), .B(keyinput_211), .ZN(n9000) );
  XNOR2_X1 U10058 ( .A(n9214), .B(keyinput_212), .ZN(n8999) );
  AOI211_X1 U10059 ( .C1(n9002), .C2(n9001), .A(n9000), .B(n8999), .ZN(n9005)
         );
  XOR2_X1 U10060 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .Z(n9004)
         );
  XNOR2_X1 U10061 ( .A(n9219), .B(keyinput_214), .ZN(n9003) );
  OAI21_X1 U10062 ( .B1(n9005), .B2(n9004), .A(n9003), .ZN(n9012) );
  OAI22_X1 U10063 ( .A1(n9007), .A2(keyinput_216), .B1(keyinput_215), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n9006) );
  AOI221_X1 U10064 ( .B1(n9007), .B2(keyinput_216), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput_215), .A(n9006), .ZN(n9011) );
  XNOR2_X1 U10065 ( .A(n10637), .B(keyinput_219), .ZN(n9010) );
  OAI22_X1 U10066 ( .A1(n5193), .A2(keyinput_218), .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_217), .ZN(n9008) );
  AOI221_X1 U10067 ( .B1(n5193), .B2(keyinput_218), .C1(keyinput_217), .C2(
        P2_DATAO_REG_7__SCAN_IN), .A(n9008), .ZN(n9009) );
  NAND4_X1 U10068 ( .A1(n9012), .A2(n9011), .A3(n9010), .A4(n9009), .ZN(n9022)
         );
  XNOR2_X1 U10069 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_220), .ZN(n9021) );
  INV_X1 U10070 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9014) );
  OAI22_X1 U10071 ( .A1(n9014), .A2(keyinput_223), .B1(P1_IR_REG_3__SCAN_IN), 
        .B2(keyinput_222), .ZN(n9013) );
  AOI221_X1 U10072 ( .B1(n9014), .B2(keyinput_223), .C1(keyinput_222), .C2(
        P1_IR_REG_3__SCAN_IN), .A(n9013), .ZN(n9019) );
  XNOR2_X1 U10073 ( .A(n9015), .B(keyinput_225), .ZN(n9018) );
  XNOR2_X1 U10074 ( .A(n6662), .B(keyinput_224), .ZN(n9017) );
  XNOR2_X1 U10075 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_221), .ZN(n9016) );
  NAND4_X1 U10076 ( .A1(n9019), .A2(n9018), .A3(n9017), .A4(n9016), .ZN(n9020)
         );
  AOI21_X1 U10077 ( .B1(n9022), .B2(n9021), .A(n9020), .ZN(n9025) );
  XNOR2_X1 U10078 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_226), .ZN(n9024) );
  XNOR2_X1 U10079 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_227), .ZN(n9023) );
  OAI21_X1 U10080 ( .B1(n9025), .B2(n9024), .A(n9023), .ZN(n9030) );
  XOR2_X1 U10081 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_228), .Z(n9029) );
  XNOR2_X1 U10082 ( .A(n9026), .B(keyinput_230), .ZN(n9028) );
  XNOR2_X1 U10083 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_229), .ZN(n9027) );
  AOI211_X1 U10084 ( .C1(n9030), .C2(n9029), .A(n9028), .B(n9027), .ZN(n9037)
         );
  XNOR2_X1 U10085 ( .A(n6841), .B(keyinput_232), .ZN(n9036) );
  XNOR2_X1 U10086 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_233), .ZN(n9035) );
  XNOR2_X1 U10087 ( .A(n9251), .B(keyinput_234), .ZN(n9033) );
  XNOR2_X1 U10088 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_231), .ZN(n9032) );
  XNOR2_X1 U10089 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_235), .ZN(n9031) );
  NAND3_X1 U10090 ( .A1(n9033), .A2(n9032), .A3(n9031), .ZN(n9034) );
  NOR4_X1 U10091 ( .A1(n9037), .A2(n9036), .A3(n9035), .A4(n9034), .ZN(n9040)
         );
  XNOR2_X1 U10092 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_236), .ZN(n9039) );
  XNOR2_X1 U10093 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_237), .ZN(n9038) );
  NOR3_X1 U10094 ( .A1(n9040), .A2(n9039), .A3(n9038), .ZN(n9043) );
  XNOR2_X1 U10095 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_238), .ZN(n9042) );
  XOR2_X1 U10096 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_239), .Z(n9041) );
  OAI21_X1 U10097 ( .B1(n9043), .B2(n9042), .A(n9041), .ZN(n9047) );
  XNOR2_X1 U10098 ( .A(n9262), .B(keyinput_240), .ZN(n9046) );
  XNOR2_X1 U10099 ( .A(n9044), .B(keyinput_241), .ZN(n9045) );
  NAND3_X1 U10100 ( .A1(n9047), .A2(n9046), .A3(n9045), .ZN(n9052) );
  XNOR2_X1 U10101 ( .A(n9048), .B(keyinput_242), .ZN(n9051) );
  XNOR2_X1 U10102 ( .A(n9266), .B(keyinput_244), .ZN(n9050) );
  XNOR2_X1 U10103 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_243), .ZN(n9049) );
  NAND4_X1 U10104 ( .A1(n9052), .A2(n9051), .A3(n9050), .A4(n9049), .ZN(n9064)
         );
  XNOR2_X1 U10105 ( .A(n9053), .B(keyinput_245), .ZN(n9057) );
  XNOR2_X1 U10106 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_247), .ZN(n9056) );
  XNOR2_X1 U10107 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_248), .ZN(n9055) );
  XNOR2_X1 U10108 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_246), .ZN(n9054) );
  NOR4_X1 U10109 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9054), .ZN(n9063)
         );
  XOR2_X1 U10110 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_249), .Z(n9061) );
  XOR2_X1 U10111 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_252), .Z(n9060) );
  XNOR2_X1 U10112 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_251), .ZN(n9059) );
  XNOR2_X1 U10113 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_250), .ZN(n9058) );
  NAND4_X1 U10114 ( .A1(n9061), .A2(n9060), .A3(n9059), .A4(n9058), .ZN(n9062)
         );
  AOI21_X1 U10115 ( .B1(n9064), .B2(n9063), .A(n9062), .ZN(n9067) );
  INV_X1 U10116 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10545) );
  XNOR2_X1 U10117 ( .A(n10545), .B(keyinput_253), .ZN(n9066) );
  INV_X1 U10118 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10546) );
  XNOR2_X1 U10119 ( .A(n10546), .B(keyinput_254), .ZN(n9065) );
  NOR3_X1 U10120 ( .A1(n9067), .A2(n9066), .A3(n9065), .ZN(n9070) );
  INV_X1 U10121 ( .A(n9070), .ZN(n9069) );
  INV_X1 U10122 ( .A(keyinput_127), .ZN(n9068) );
  AOI21_X1 U10123 ( .B1(n9069), .B2(keyinput_255), .A(n9068), .ZN(n9288) );
  INV_X1 U10124 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10547) );
  NOR2_X1 U10125 ( .A1(n9070), .A2(keyinput_255), .ZN(n9071) );
  OAI21_X1 U10126 ( .B1(n9071), .B2(keyinput_127), .A(n10547), .ZN(n9287) );
  XNOR2_X1 U10127 ( .A(SI_31_), .B(keyinput_1), .ZN(n9074) );
  XNOR2_X1 U10128 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n9073) );
  XOR2_X1 U10129 ( .A(SI_30_), .B(keyinput_2), .Z(n9072) );
  OAI21_X1 U10130 ( .B1(n9074), .B2(n9073), .A(n9072), .ZN(n9078) );
  XNOR2_X1 U10131 ( .A(n9075), .B(keyinput_3), .ZN(n9077) );
  XNOR2_X1 U10132 ( .A(SI_28_), .B(keyinput_4), .ZN(n9076) );
  AOI21_X1 U10133 ( .B1(n9078), .B2(n9077), .A(n9076), .ZN(n9086) );
  XNOR2_X1 U10134 ( .A(SI_27_), .B(keyinput_5), .ZN(n9085) );
  XNOR2_X1 U10135 ( .A(SI_23_), .B(keyinput_9), .ZN(n9084) );
  XNOR2_X1 U10136 ( .A(SI_26_), .B(keyinput_6), .ZN(n9082) );
  XNOR2_X1 U10137 ( .A(SI_24_), .B(keyinput_8), .ZN(n9081) );
  XNOR2_X1 U10138 ( .A(SI_25_), .B(keyinput_7), .ZN(n9080) );
  XNOR2_X1 U10139 ( .A(SI_22_), .B(keyinput_10), .ZN(n9079) );
  NAND4_X1 U10140 ( .A1(n9082), .A2(n9081), .A3(n9080), .A4(n9079), .ZN(n9083)
         );
  NOR4_X1 U10141 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(n9093)
         );
  XNOR2_X1 U10142 ( .A(SI_20_), .B(keyinput_12), .ZN(n9090) );
  XNOR2_X1 U10143 ( .A(SI_21_), .B(keyinput_11), .ZN(n9089) );
  XNOR2_X1 U10144 ( .A(SI_19_), .B(keyinput_13), .ZN(n9088) );
  XNOR2_X1 U10145 ( .A(SI_18_), .B(keyinput_14), .ZN(n9087) );
  NAND4_X1 U10146 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n9092)
         );
  XNOR2_X1 U10147 ( .A(SI_17_), .B(keyinput_15), .ZN(n9091) );
  OAI21_X1 U10148 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(n9108) );
  XNOR2_X1 U10149 ( .A(n9094), .B(keyinput_19), .ZN(n9100) );
  XNOR2_X1 U10150 ( .A(n9095), .B(keyinput_18), .ZN(n9099) );
  XNOR2_X1 U10151 ( .A(n9096), .B(keyinput_16), .ZN(n9098) );
  XNOR2_X1 U10152 ( .A(SI_15_), .B(keyinput_17), .ZN(n9097) );
  NOR4_X1 U10153 ( .A1(n9100), .A2(n9099), .A3(n9098), .A4(n9097), .ZN(n9107)
         );
  XNOR2_X1 U10154 ( .A(n9101), .B(keyinput_20), .ZN(n9105) );
  XNOR2_X1 U10155 ( .A(n9102), .B(keyinput_21), .ZN(n9104) );
  XNOR2_X1 U10156 ( .A(SI_10_), .B(keyinput_22), .ZN(n9103) );
  NAND3_X1 U10157 ( .A1(n9105), .A2(n9104), .A3(n9103), .ZN(n9106) );
  AOI21_X1 U10158 ( .B1(n9108), .B2(n9107), .A(n9106), .ZN(n9113) );
  XNOR2_X1 U10159 ( .A(n9109), .B(keyinput_23), .ZN(n9112) );
  XNOR2_X1 U10160 ( .A(n9110), .B(keyinput_24), .ZN(n9111) );
  OAI21_X1 U10161 ( .B1(n9113), .B2(n9112), .A(n9111), .ZN(n9127) );
  XOR2_X1 U10162 ( .A(SI_7_), .B(keyinput_25), .Z(n9126) );
  INV_X1 U10163 ( .A(keyinput_29), .ZN(n9118) );
  AOI22_X1 U10164 ( .A1(SI_4_), .A2(keyinput_28), .B1(SI_6_), .B2(keyinput_26), 
        .ZN(n9115) );
  AOI22_X1 U10165 ( .A1(SI_0_), .A2(keyinput_32), .B1(SI_3_), .B2(keyinput_29), 
        .ZN(n9114) );
  OAI211_X1 U10166 ( .C1(SI_4_), .C2(keyinput_28), .A(n9115), .B(n9114), .ZN(
        n9117) );
  OAI22_X1 U10167 ( .A1(SI_0_), .A2(keyinput_32), .B1(SI_6_), .B2(keyinput_26), 
        .ZN(n9116) );
  AOI211_X1 U10168 ( .C1(n9119), .C2(n9118), .A(n9117), .B(n9116), .ZN(n9124)
         );
  XNOR2_X1 U10169 ( .A(n9120), .B(keyinput_30), .ZN(n9123) );
  XNOR2_X1 U10170 ( .A(SI_1_), .B(keyinput_31), .ZN(n9122) );
  XNOR2_X1 U10171 ( .A(SI_5_), .B(keyinput_27), .ZN(n9121) );
  NAND4_X1 U10172 ( .A1(n9124), .A2(n9123), .A3(n9122), .A4(n9121), .ZN(n9125)
         );
  AOI21_X1 U10173 ( .B1(n9127), .B2(n9126), .A(n9125), .ZN(n9130) );
  XNOR2_X1 U10174 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n9129) );
  XNOR2_X1 U10175 ( .A(P2_U3152), .B(keyinput_34), .ZN(n9128) );
  OAI21_X1 U10176 ( .B1(n9130), .B2(n9129), .A(n9128), .ZN(n9138) );
  XOR2_X1 U10177 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .Z(n9137) );
  XOR2_X1 U10178 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .Z(n9135) );
  XNOR2_X1 U10179 ( .A(n9293), .B(keyinput_38), .ZN(n9134) );
  XNOR2_X1 U10180 ( .A(n9131), .B(keyinput_37), .ZN(n9133) );
  XNOR2_X1 U10181 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n9132)
         );
  NAND4_X1 U10182 ( .A1(n9135), .A2(n9134), .A3(n9133), .A4(n9132), .ZN(n9136)
         );
  AOI21_X1 U10183 ( .B1(n9138), .B2(n9137), .A(n9136), .ZN(n9143) );
  XNOR2_X1 U10184 ( .A(n9139), .B(keyinput_40), .ZN(n9142) );
  XNOR2_X1 U10185 ( .A(n9140), .B(keyinput_41), .ZN(n9141) );
  OAI21_X1 U10186 ( .B1(n9143), .B2(n9142), .A(n9141), .ZN(n9147) );
  XNOR2_X1 U10187 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n9146)
         );
  XNOR2_X1 U10188 ( .A(n9144), .B(keyinput_43), .ZN(n9145) );
  AOI21_X1 U10189 ( .B1(n9147), .B2(n9146), .A(n9145), .ZN(n9151) );
  XOR2_X1 U10190 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n9150) );
  XOR2_X1 U10191 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .Z(n9149) );
  XNOR2_X1 U10192 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n9148)
         );
  OAI211_X1 U10193 ( .C1(n9151), .C2(n9150), .A(n9149), .B(n9148), .ZN(n9154)
         );
  XNOR2_X1 U10194 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_48), .ZN(n9153)
         );
  XNOR2_X1 U10195 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n9152)
         );
  NAND3_X1 U10196 ( .A1(n9154), .A2(n9153), .A3(n9152), .ZN(n9164) );
  XNOR2_X1 U10197 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n9163) );
  XNOR2_X1 U10198 ( .A(n9155), .B(keyinput_50), .ZN(n9161) );
  XNOR2_X1 U10199 ( .A(n9156), .B(keyinput_52), .ZN(n9160) );
  XNOR2_X1 U10200 ( .A(n9157), .B(keyinput_51), .ZN(n9159) );
  XNOR2_X1 U10201 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n9158) );
  NAND4_X1 U10202 ( .A1(n9161), .A2(n9160), .A3(n9159), .A4(n9158), .ZN(n9162)
         );
  AOI21_X1 U10203 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(n9173) );
  XOR2_X1 U10204 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n9169) );
  XNOR2_X1 U10205 ( .A(n9165), .B(keyinput_57), .ZN(n9168) );
  XNOR2_X1 U10206 ( .A(n9343), .B(keyinput_55), .ZN(n9167) );
  XNOR2_X1 U10207 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_56), .ZN(n9166)
         );
  NAND4_X1 U10208 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .ZN(n9172)
         );
  XOR2_X1 U10209 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .Z(n9171) );
  XNOR2_X1 U10210 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n9170)
         );
  OAI211_X1 U10211 ( .C1(n9173), .C2(n9172), .A(n9171), .B(n9170), .ZN(n9178)
         );
  XNOR2_X1 U10212 ( .A(n9174), .B(keyinput_60), .ZN(n9177) );
  XNOR2_X1 U10213 ( .A(n9175), .B(keyinput_61), .ZN(n9176) );
  AOI21_X1 U10214 ( .B1(n9178), .B2(n9177), .A(n9176), .ZN(n9186) );
  XOR2_X1 U10215 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .Z(n9182) );
  XNOR2_X1 U10216 ( .A(n9179), .B(keyinput_63), .ZN(n9181) );
  XNOR2_X1 U10217 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n9180)
         );
  NAND3_X1 U10218 ( .A1(n9182), .A2(n9181), .A3(n9180), .ZN(n9185) );
  XOR2_X1 U10219 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .Z(n9184) );
  XNOR2_X1 U10220 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .ZN(n9183)
         );
  OAI211_X1 U10221 ( .C1(n9186), .C2(n9185), .A(n9184), .B(n9183), .ZN(n9189)
         );
  XOR2_X1 U10222 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .Z(n9188) );
  XNOR2_X1 U10223 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .ZN(n9187)
         );
  NAND3_X1 U10224 ( .A1(n9189), .A2(n9188), .A3(n9187), .ZN(n9194) );
  XNOR2_X1 U10225 ( .A(n9190), .B(keyinput_69), .ZN(n9193) );
  XNOR2_X1 U10226 ( .A(n9191), .B(keyinput_70), .ZN(n9192) );
  NAND3_X1 U10227 ( .A1(n9194), .A2(n9193), .A3(n9192), .ZN(n9198) );
  XNOR2_X1 U10228 ( .A(n9195), .B(keyinput_71), .ZN(n9197) );
  XNOR2_X1 U10229 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .ZN(n9196)
         );
  AOI21_X1 U10230 ( .B1(n9198), .B2(n9197), .A(n9196), .ZN(n9201) );
  XNOR2_X1 U10231 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n9200)
         );
  XNOR2_X1 U10232 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n9199)
         );
  NOR3_X1 U10233 ( .A1(n9201), .A2(n9200), .A3(n9199), .ZN(n9208) );
  XOR2_X1 U10234 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n9205) );
  XOR2_X1 U10235 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n9204) );
  XNOR2_X1 U10236 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n9203)
         );
  XNOR2_X1 U10237 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n9202)
         );
  NAND4_X1 U10238 ( .A1(n9205), .A2(n9204), .A3(n9203), .A4(n9202), .ZN(n9207)
         );
  XOR2_X1 U10239 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .Z(n9206) );
  OAI21_X1 U10240 ( .B1(n9208), .B2(n9207), .A(n9206), .ZN(n9213) );
  XNOR2_X1 U10241 ( .A(n9209), .B(keyinput_80), .ZN(n9212) );
  XNOR2_X1 U10242 ( .A(n9210), .B(keyinput_81), .ZN(n9211) );
  NAND3_X1 U10243 ( .A1(n9213), .A2(n9212), .A3(n9211), .ZN(n9218) );
  XNOR2_X1 U10244 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n9217)
         );
  XNOR2_X1 U10245 ( .A(n9214), .B(keyinput_84), .ZN(n9216) );
  XNOR2_X1 U10246 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n9215)
         );
  AOI211_X1 U10247 ( .C1(n9218), .C2(n9217), .A(n9216), .B(n9215), .ZN(n9222)
         );
  XOR2_X1 U10248 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .Z(n9221) );
  XNOR2_X1 U10249 ( .A(n9219), .B(keyinput_86), .ZN(n9220) );
  OAI21_X1 U10250 ( .B1(n9222), .B2(n9221), .A(n9220), .ZN(n9229) );
  XNOR2_X1 U10251 ( .A(n10637), .B(keyinput_91), .ZN(n9228) );
  XNOR2_X1 U10252 ( .A(n7292), .B(keyinput_87), .ZN(n9227) );
  XOR2_X1 U10253 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n9225) );
  XNOR2_X1 U10254 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n9224)
         );
  XNOR2_X1 U10255 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .ZN(n9223)
         );
  NOR3_X1 U10256 ( .A1(n9225), .A2(n9224), .A3(n9223), .ZN(n9226) );
  NAND4_X1 U10257 ( .A1(n9229), .A2(n9228), .A3(n9227), .A4(n9226), .ZN(n9238)
         );
  XNOR2_X1 U10258 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_92), .ZN(n9237) );
  XNOR2_X1 U10259 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_95), .ZN(n9231) );
  XNOR2_X1 U10260 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_96), .ZN(n9230) );
  NOR2_X1 U10261 ( .A1(n9231), .A2(n9230), .ZN(n9235) );
  XNOR2_X1 U10262 ( .A(n9015), .B(keyinput_97), .ZN(n9234) );
  XNOR2_X1 U10263 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_94), .ZN(n9233) );
  XNOR2_X1 U10264 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_93), .ZN(n9232) );
  NAND4_X1 U10265 ( .A1(n9235), .A2(n9234), .A3(n9233), .A4(n9232), .ZN(n9236)
         );
  AOI21_X1 U10266 ( .B1(n9238), .B2(n9237), .A(n9236), .ZN(n9241) );
  XNOR2_X1 U10267 ( .A(n6725), .B(keyinput_98), .ZN(n9240) );
  XOR2_X1 U10268 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_99), .Z(n9239) );
  OAI21_X1 U10269 ( .B1(n9241), .B2(n9240), .A(n9239), .ZN(n9245) );
  XNOR2_X1 U10270 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_100), .ZN(n9244) );
  XNOR2_X1 U10271 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_102), .ZN(n9243) );
  XNOR2_X1 U10272 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_101), .ZN(n9242) );
  AOI211_X1 U10273 ( .C1(n9245), .C2(n9244), .A(n9243), .B(n9242), .ZN(n9258)
         );
  XNOR2_X1 U10274 ( .A(n9246), .B(keyinput_103), .ZN(n9250) );
  XNOR2_X1 U10275 ( .A(n9247), .B(keyinput_105), .ZN(n9249) );
  XNOR2_X1 U10276 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_107), .ZN(n9248) );
  NOR3_X1 U10277 ( .A1(n9250), .A2(n9249), .A3(n9248), .ZN(n9254) );
  XNOR2_X1 U10278 ( .A(n6841), .B(keyinput_104), .ZN(n9253) );
  XNOR2_X1 U10279 ( .A(n9251), .B(keyinput_106), .ZN(n9252) );
  NAND3_X1 U10280 ( .A1(n9254), .A2(n9253), .A3(n9252), .ZN(n9257) );
  XNOR2_X1 U10281 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_109), .ZN(n9256) );
  XNOR2_X1 U10282 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_108), .ZN(n9255) );
  OAI211_X1 U10283 ( .C1(n9258), .C2(n9257), .A(n9256), .B(n9255), .ZN(n9261)
         );
  XNOR2_X1 U10284 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_110), .ZN(n9260) );
  XOR2_X1 U10285 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_111), .Z(n9259) );
  AOI21_X1 U10286 ( .B1(n9261), .B2(n9260), .A(n9259), .ZN(n9265) );
  XNOR2_X1 U10287 ( .A(n9262), .B(keyinput_112), .ZN(n9264) );
  XNOR2_X1 U10288 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_113), .ZN(n9263) );
  NOR3_X1 U10289 ( .A1(n9265), .A2(n9264), .A3(n9263), .ZN(n9270) );
  XNOR2_X1 U10290 ( .A(n9266), .B(keyinput_116), .ZN(n9269) );
  XNOR2_X1 U10291 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_114), .ZN(n9268) );
  XNOR2_X1 U10292 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_115), .ZN(n9267) );
  NOR4_X1 U10293 ( .A1(n9270), .A2(n9269), .A3(n9268), .A4(n9267), .ZN(n9282)
         );
  XNOR2_X1 U10294 ( .A(n9271), .B(keyinput_118), .ZN(n9275) );
  XNOR2_X1 U10295 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_120), .ZN(n9274) );
  XNOR2_X1 U10296 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_117), .ZN(n9273) );
  XNOR2_X1 U10297 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_119), .ZN(n9272) );
  NAND4_X1 U10298 ( .A1(n9275), .A2(n9274), .A3(n9273), .A4(n9272), .ZN(n9281)
         );
  XOR2_X1 U10299 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_122), .Z(n9279) );
  XOR2_X1 U10300 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_123), .Z(n9278) );
  XNOR2_X1 U10301 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_124), .ZN(n9277) );
  XNOR2_X1 U10302 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_121), .ZN(n9276) );
  NOR4_X1 U10303 ( .A1(n9279), .A2(n9278), .A3(n9277), .A4(n9276), .ZN(n9280)
         );
  OAI21_X1 U10304 ( .B1(n9282), .B2(n9281), .A(n9280), .ZN(n9285) );
  XNOR2_X1 U10305 ( .A(n10545), .B(keyinput_125), .ZN(n9284) );
  XNOR2_X1 U10306 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_126), .ZN(n9283) );
  NAND3_X1 U10307 ( .A1(n9285), .A2(n9284), .A3(n9283), .ZN(n9286) );
  OAI211_X1 U10308 ( .C1(n9288), .C2(n10547), .A(n9287), .B(n9286), .ZN(n9289)
         );
  XNOR2_X1 U10309 ( .A(n9290), .B(n9289), .ZN(P2_U3216) );
  XNOR2_X1 U10310 ( .A(n9292), .B(n9291), .ZN(n9298) );
  OAI22_X1 U10311 ( .A1(n9564), .A2(n9365), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9293), .ZN(n9296) );
  OAI22_X1 U10312 ( .A1(n9294), .A2(n9362), .B1(n9524), .B2(n9363), .ZN(n9295)
         );
  AOI211_X1 U10313 ( .C1(n9700), .C2(n9379), .A(n9296), .B(n9295), .ZN(n9297)
         );
  OAI21_X1 U10314 ( .B1(n9298), .B2(n9381), .A(n9297), .ZN(P2_U3218) );
  OAI21_X1 U10315 ( .B1(n9301), .B2(n9300), .A(n9299), .ZN(n9302) );
  NAND2_X1 U10316 ( .A1(n9302), .A2(n9352), .ZN(n9305) );
  AND2_X1 U10317 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9419) );
  OAI22_X1 U10318 ( .A1(n9365), .A2(n9593), .B1(n9363), .B2(n9597), .ZN(n9303)
         );
  AOI211_X1 U10319 ( .C1(n9334), .C2(n9591), .A(n9419), .B(n9303), .ZN(n9304)
         );
  OAI211_X1 U10320 ( .C1(n9777), .C2(n9358), .A(n9305), .B(n9304), .ZN(
        P2_U3221) );
  XNOR2_X1 U10321 ( .A(n9307), .B(n9306), .ZN(n9313) );
  OAI22_X1 U10322 ( .A1(n9564), .A2(n9362), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9308), .ZN(n9311) );
  INV_X1 U10323 ( .A(n9566), .ZN(n9309) );
  OAI22_X1 U10324 ( .A1(n9365), .A2(n9563), .B1(n9363), .B2(n9309), .ZN(n9310)
         );
  AOI211_X1 U10325 ( .C1(n9557), .C2(n9379), .A(n9311), .B(n9310), .ZN(n9312)
         );
  OAI21_X1 U10326 ( .B1(n9313), .B2(n9381), .A(n9312), .ZN(P2_U3225) );
  OAI21_X1 U10327 ( .B1(n9316), .B2(n9315), .A(n9314), .ZN(n9317) );
  NAND2_X1 U10328 ( .A1(n9317), .A2(n9352), .ZN(n9324) );
  NAND2_X1 U10329 ( .A1(n9384), .A2(n9638), .ZN(n9319) );
  NAND2_X1 U10330 ( .A1(n9530), .A2(n9619), .ZN(n9318) );
  NAND2_X1 U10331 ( .A1(n9319), .A2(n9318), .ZN(n9493) );
  INV_X1 U10332 ( .A(n9499), .ZN(n9321) );
  OAI22_X1 U10333 ( .A1(n9321), .A2(n9363), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9320), .ZN(n9322) );
  AOI21_X1 U10334 ( .B1(n9493), .B2(n9373), .A(n9322), .ZN(n9323) );
  OAI211_X1 U10335 ( .C1(n9765), .C2(n9358), .A(n9324), .B(n9323), .ZN(
        P2_U3227) );
  XNOR2_X1 U10336 ( .A(n9326), .B(n9325), .ZN(n9331) );
  OAI22_X1 U10337 ( .A1(n9362), .A2(n9593), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9155), .ZN(n9329) );
  OAI22_X1 U10338 ( .A1(n9365), .A2(n9327), .B1(n9363), .B2(n9629), .ZN(n9328)
         );
  AOI211_X1 U10339 ( .C1(n9627), .C2(n9379), .A(n9329), .B(n9328), .ZN(n9330)
         );
  OAI21_X1 U10340 ( .B1(n9331), .B2(n9381), .A(n9330), .ZN(P2_U3230) );
  XNOR2_X1 U10341 ( .A(n9332), .B(n9333), .ZN(n9340) );
  NAND2_X1 U10342 ( .A1(n9513), .A2(n9334), .ZN(n9337) );
  AOI22_X1 U10343 ( .A1(n9512), .A2(n9335), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n9336) );
  OAI211_X1 U10344 ( .C1(n9363), .C2(n9507), .A(n9337), .B(n9336), .ZN(n9338)
         );
  AOI21_X1 U10345 ( .B1(n9695), .B2(n9379), .A(n9338), .ZN(n9339) );
  OAI21_X1 U10346 ( .B1(n9340), .B2(n9381), .A(n9339), .ZN(P2_U3231) );
  XNOR2_X1 U10347 ( .A(n9342), .B(n9341), .ZN(n9348) );
  OAI22_X1 U10348 ( .A1(n9365), .A2(n9361), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9343), .ZN(n9346) );
  INV_X1 U10349 ( .A(n9574), .ZN(n9344) );
  OAI22_X1 U10350 ( .A1(n9547), .A2(n9362), .B1(n9363), .B2(n9344), .ZN(n9345)
         );
  AOI211_X1 U10351 ( .C1(n9716), .C2(n9379), .A(n9346), .B(n9345), .ZN(n9347)
         );
  OAI21_X1 U10352 ( .B1(n9348), .B2(n9381), .A(n9347), .ZN(P2_U3235) );
  OAI21_X1 U10353 ( .B1(n9351), .B2(n9350), .A(n9349), .ZN(n9353) );
  NAND2_X1 U10354 ( .A1(n9353), .A2(n9352), .ZN(n9357) );
  OAI22_X1 U10355 ( .A1(n9547), .A2(n9365), .B1(n9541), .B2(n9363), .ZN(n9355)
         );
  NOR2_X1 U10356 ( .A1(n9548), .A2(n9362), .ZN(n9354) );
  AOI211_X1 U10357 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n9355), 
        .B(n9354), .ZN(n9356) );
  OAI211_X1 U10358 ( .C1(n9544), .C2(n9358), .A(n9357), .B(n9356), .ZN(
        P2_U3237) );
  XNOR2_X1 U10359 ( .A(n9360), .B(n9359), .ZN(n9369) );
  NAND2_X1 U10360 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9401) );
  OAI21_X1 U10361 ( .B1(n9362), .B2(n9361), .A(n9401), .ZN(n9367) );
  OAI22_X1 U10362 ( .A1(n9365), .A2(n9364), .B1(n9363), .B2(n9606), .ZN(n9366)
         );
  AOI211_X1 U10363 ( .C1(n9727), .C2(n9379), .A(n9367), .B(n9366), .ZN(n9368)
         );
  OAI21_X1 U10364 ( .B1(n9369), .B2(n9381), .A(n9368), .ZN(P2_U3240) );
  XNOR2_X1 U10365 ( .A(n9371), .B(n9370), .ZN(n9382) );
  AND2_X1 U10366 ( .A1(n9513), .A2(n9619), .ZN(n9372) );
  AOI21_X1 U10367 ( .B1(n9444), .B2(n9638), .A(n9372), .ZN(n9478) );
  INV_X1 U10368 ( .A(n9373), .ZN(n9377) );
  INV_X1 U10369 ( .A(n9481), .ZN(n9375) );
  AOI22_X1 U10370 ( .A1(n9375), .A2(n9374), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n9376) );
  OAI21_X1 U10371 ( .B1(n9478), .B2(n9377), .A(n9376), .ZN(n9378) );
  AOI21_X1 U10372 ( .B1(n9684), .B2(n9379), .A(n9378), .ZN(n9380) );
  OAI21_X1 U10373 ( .B1(n9382), .B2(n9381), .A(n9380), .ZN(P2_U3242) );
  MUX2_X1 U10374 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9383), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10375 ( .A(n9445), .B(P2_DATAO_REG_29__SCAN_IN), .S(n9385), .Z(
        P2_U3581) );
  MUX2_X1 U10376 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9468), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U10377 ( .A(n9444), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9385), .Z(
        P2_U3579) );
  MUX2_X1 U10378 ( .A(n9384), .B(P2_DATAO_REG_26__SCAN_IN), .S(n9385), .Z(
        P2_U3578) );
  MUX2_X1 U10379 ( .A(n9513), .B(P2_DATAO_REG_25__SCAN_IN), .S(n9385), .Z(
        P2_U3577) );
  MUX2_X1 U10380 ( .A(n9530), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9385), .Z(
        P2_U3576) );
  MUX2_X1 U10381 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9512), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U10382 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9531), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10383 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9579), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10384 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9591), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10385 ( .A(n9604), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9385), .Z(
        P2_U3571) );
  MUX2_X1 U10386 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9620), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10387 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9639), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10388 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9618), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10389 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9386), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10390 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9387), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10391 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9388), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10392 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9389), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10393 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9390), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10394 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9391), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10395 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n9392), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10396 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n9393), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10397 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n9394), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10398 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n9395), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10399 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9396), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10400 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n9397), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10401 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n7404), .S(P2_U3966), .Z(
        P2_U3553) );
  XNOR2_X1 U10402 ( .A(n9414), .B(P2_REG2_REG_18__SCAN_IN), .ZN(n9410) );
  AOI21_X1 U10403 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n9400), .A(n9398), .ZN(
        n9408) );
  XNOR2_X1 U10404 ( .A(n9410), .B(n9408), .ZN(n9406) );
  XNOR2_X1 U10405 ( .A(n9414), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9416) );
  AOI21_X1 U10406 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9400), .A(n9399), .ZN(
        n9413) );
  XNOR2_X1 U10407 ( .A(n9416), .B(n9413), .ZN(n9403) );
  NAND2_X1 U10408 ( .A1(n10674), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n9402) );
  OAI211_X1 U10409 ( .C1(n9403), .C2(n9422), .A(n9402), .B(n9401), .ZN(n9404)
         );
  AOI21_X1 U10410 ( .B1(n9414), .B2(n10680), .A(n9404), .ZN(n9405) );
  OAI21_X1 U10411 ( .B1(n9406), .B2(n10689), .A(n9405), .ZN(P2_U3263) );
  MUX2_X1 U10412 ( .A(n6191), .B(P2_REG2_REG_19__SCAN_IN), .S(n9407), .Z(n9412) );
  INV_X1 U10413 ( .A(n9408), .ZN(n9409) );
  OAI22_X1 U10414 ( .A1(n9410), .A2(n9409), .B1(n9414), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n9411) );
  XOR2_X1 U10415 ( .A(n9412), .B(n9411), .Z(n9425) );
  XNOR2_X1 U10416 ( .A(n6002), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9418) );
  INV_X1 U10417 ( .A(n9413), .ZN(n9415) );
  OAI22_X1 U10418 ( .A1(n9416), .A2(n9415), .B1(n9414), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n9417) );
  XNOR2_X1 U10419 ( .A(n9418), .B(n9417), .ZN(n9421) );
  AOI21_X1 U10420 ( .B1(n10674), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n9419), .ZN(
        n9420) );
  OAI21_X1 U10421 ( .B1(n9422), .B2(n9421), .A(n9420), .ZN(n9423) );
  AOI21_X1 U10422 ( .B1(n6002), .B2(n10680), .A(n9423), .ZN(n9424) );
  OAI21_X1 U10423 ( .B1(n10689), .B2(n9425), .A(n9424), .ZN(P2_U3264) );
  NAND2_X1 U10424 ( .A1(n9426), .A2(n9610), .ZN(n9429) );
  INV_X1 U10425 ( .A(n9427), .ZN(n9665) );
  NOR2_X1 U10426 ( .A1(n10851), .A2(n9665), .ZN(n9432) );
  AOI21_X1 U10427 ( .B1(n10851), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9432), .ZN(
        n9428) );
  OAI211_X1 U10428 ( .C1(n9430), .C2(n9628), .A(n9429), .B(n9428), .ZN(
        P2_U3265) );
  OR2_X1 U10429 ( .A1(n9755), .A2(n9431), .ZN(n9664) );
  NAND3_X1 U10430 ( .A1(n9664), .A2(n9663), .A3(n9610), .ZN(n9434) );
  AOI21_X1 U10431 ( .B1(n10851), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9432), .ZN(
        n9433) );
  OAI211_X1 U10432 ( .C1(n9755), .C2(n9628), .A(n9434), .B(n9433), .ZN(
        P2_U3266) );
  XNOR2_X1 U10433 ( .A(n9435), .B(n9442), .ZN(n9678) );
  INV_X1 U10434 ( .A(n9436), .ZN(n9437) );
  AOI21_X1 U10435 ( .B1(n9674), .B2(n9452), .A(n9437), .ZN(n9675) );
  AOI22_X1 U10436 ( .A1(n9438), .A2(n10755), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n10851), .ZN(n9439) );
  OAI21_X1 U10437 ( .B1(n9440), .B2(n9628), .A(n9439), .ZN(n9449) );
  OAI211_X1 U10438 ( .C1(n9443), .C2(n9442), .A(n9441), .B(n9644), .ZN(n9447)
         );
  AOI22_X1 U10439 ( .A1(n9445), .A2(n9638), .B1(n9444), .B2(n9619), .ZN(n9446)
         );
  NOR2_X1 U10440 ( .A1(n9677), .A2(n10851), .ZN(n9448) );
  AOI211_X1 U10441 ( .C1(n9610), .C2(n9675), .A(n9449), .B(n9448), .ZN(n9450)
         );
  OAI21_X1 U10442 ( .B1(n9678), .B2(n9602), .A(n9450), .ZN(P2_U3268) );
  XOR2_X1 U10443 ( .A(n9465), .B(n9451), .Z(n9683) );
  INV_X1 U10444 ( .A(n9452), .ZN(n9453) );
  AOI21_X1 U10445 ( .B1(n9679), .B2(n9454), .A(n9453), .ZN(n9680) );
  INV_X1 U10446 ( .A(n9455), .ZN(n9456) );
  AOI22_X1 U10447 ( .A1(n9456), .A2(n10755), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n10851), .ZN(n9457) );
  OAI21_X1 U10448 ( .B1(n9458), .B2(n9628), .A(n9457), .ZN(n9470) );
  NOR2_X1 U10449 ( .A1(n9459), .A2(n9641), .ZN(n9467) );
  NAND2_X1 U10450 ( .A1(n9460), .A2(n9461), .ZN(n9464) );
  INV_X1 U10451 ( .A(n9462), .ZN(n9463) );
  AOI211_X1 U10452 ( .C1(n9465), .C2(n9464), .A(n9561), .B(n9463), .ZN(n9466)
         );
  AOI211_X1 U10453 ( .C1(n9638), .C2(n9468), .A(n9467), .B(n9466), .ZN(n9682)
         );
  NOR2_X1 U10454 ( .A1(n9682), .A2(n10851), .ZN(n9469) );
  AOI211_X1 U10455 ( .C1(n9610), .C2(n9680), .A(n9470), .B(n9469), .ZN(n9471)
         );
  OAI21_X1 U10456 ( .B1(n9683), .B2(n9602), .A(n9471), .ZN(P2_U3269) );
  OAI21_X1 U10457 ( .B1(n9473), .B2(n9477), .A(n9472), .ZN(n9687) );
  INV_X1 U10458 ( .A(n9687), .ZN(n9486) );
  AOI22_X1 U10459 ( .A1(n9684), .A2(n9655), .B1(n10851), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U10460 ( .A1(n9490), .A2(n9474), .ZN(n9476) );
  INV_X1 U10461 ( .A(n9460), .ZN(n9475) );
  AOI21_X1 U10462 ( .B1(n9477), .B2(n9476), .A(n9475), .ZN(n9479) );
  OAI21_X1 U10463 ( .B1(n9479), .B2(n9561), .A(n9478), .ZN(n9685) );
  AOI211_X1 U10464 ( .C1(n9684), .C2(n9496), .A(n10916), .B(n9480), .ZN(n9686)
         );
  INV_X1 U10465 ( .A(n9686), .ZN(n9482) );
  OAI22_X1 U10466 ( .A1(n9482), .A2(n6002), .B1(n10860), .B2(n9481), .ZN(n9483) );
  OAI21_X1 U10467 ( .B1(n9685), .B2(n9483), .A(n10856), .ZN(n9484) );
  OAI211_X1 U10468 ( .C1(n9486), .C2(n9602), .A(n9485), .B(n9484), .ZN(
        P2_U3270) );
  OAI21_X1 U10469 ( .B1(n9489), .B2(n9488), .A(n9487), .ZN(n9692) );
  INV_X1 U10470 ( .A(n9692), .ZN(n9504) );
  OAI211_X1 U10471 ( .C1(n9492), .C2(n9491), .A(n9490), .B(n9644), .ZN(n9495)
         );
  INV_X1 U10472 ( .A(n9493), .ZN(n9494) );
  NAND2_X1 U10473 ( .A1(n9495), .A2(n9494), .ZN(n9690) );
  INV_X1 U10474 ( .A(n9496), .ZN(n9497) );
  AOI211_X1 U10475 ( .C1(n9498), .C2(n5343), .A(n10916), .B(n9497), .ZN(n9691)
         );
  NAND2_X1 U10476 ( .A1(n9691), .A2(n9633), .ZN(n9501) );
  AOI22_X1 U10477 ( .A1(n9499), .A2(n10755), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10851), .ZN(n9500) );
  OAI211_X1 U10478 ( .C1(n9765), .C2(n9628), .A(n9501), .B(n9500), .ZN(n9502)
         );
  AOI21_X1 U10479 ( .B1(n9690), .B2(n10856), .A(n9502), .ZN(n9503) );
  OAI21_X1 U10480 ( .B1(n9504), .B2(n9602), .A(n9503), .ZN(P2_U3271) );
  XOR2_X1 U10481 ( .A(n9511), .B(n9505), .Z(n9699) );
  AOI21_X1 U10482 ( .B1(n9695), .B2(n9522), .A(n9506), .ZN(n9696) );
  INV_X1 U10483 ( .A(n9507), .ZN(n9508) );
  AOI22_X1 U10484 ( .A1(n9508), .A2(n10755), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10851), .ZN(n9509) );
  OAI21_X1 U10485 ( .B1(n5341), .B2(n9628), .A(n9509), .ZN(n9517) );
  OAI211_X1 U10486 ( .C1(n5075), .C2(n9511), .A(n9510), .B(n9644), .ZN(n9515)
         );
  AOI22_X1 U10487 ( .A1(n9513), .A2(n9638), .B1(n9619), .B2(n9512), .ZN(n9514)
         );
  AND2_X1 U10488 ( .A1(n9515), .A2(n9514), .ZN(n9698) );
  NOR2_X1 U10489 ( .A1(n9698), .A2(n10851), .ZN(n9516) );
  AOI211_X1 U10490 ( .C1(n9696), .C2(n9610), .A(n9517), .B(n9516), .ZN(n9518)
         );
  OAI21_X1 U10491 ( .B1(n9699), .B2(n9602), .A(n9518), .ZN(P2_U3272) );
  OAI21_X1 U10492 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(n9704) );
  INV_X1 U10493 ( .A(n9522), .ZN(n9523) );
  AOI21_X1 U10494 ( .B1(n9700), .B2(n9538), .A(n9523), .ZN(n9701) );
  INV_X1 U10495 ( .A(n9524), .ZN(n9525) );
  AOI22_X1 U10496 ( .A1(n9525), .A2(n10755), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n10851), .ZN(n9526) );
  OAI21_X1 U10497 ( .B1(n9527), .B2(n9628), .A(n9526), .ZN(n9534) );
  OAI21_X1 U10498 ( .B1(n9529), .B2(n5076), .A(n9528), .ZN(n9532) );
  AOI222_X1 U10499 ( .A1(n9644), .A2(n9532), .B1(n9531), .B2(n9619), .C1(n9530), .C2(n9638), .ZN(n9703) );
  NOR2_X1 U10500 ( .A1(n9703), .A2(n10851), .ZN(n9533) );
  AOI211_X1 U10501 ( .C1(n9701), .C2(n9610), .A(n9534), .B(n9533), .ZN(n9535)
         );
  OAI21_X1 U10502 ( .B1(n9602), .B2(n9704), .A(n9535), .ZN(P2_U3273) );
  AOI21_X1 U10503 ( .B1(n9537), .B2(n9536), .A(n5051), .ZN(n9709) );
  INV_X1 U10504 ( .A(n9556), .ZN(n9540) );
  INV_X1 U10505 ( .A(n9538), .ZN(n9539) );
  AOI21_X1 U10506 ( .B1(n9705), .B2(n9540), .A(n9539), .ZN(n9706) );
  INV_X1 U10507 ( .A(n9541), .ZN(n9542) );
  AOI22_X1 U10508 ( .A1(n9542), .A2(n10755), .B1(n10851), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n9543) );
  OAI21_X1 U10509 ( .B1(n9544), .B2(n9628), .A(n9543), .ZN(n9553) );
  AOI21_X1 U10510 ( .B1(n9546), .B2(n9545), .A(n9561), .ZN(n9551) );
  OAI22_X1 U10511 ( .A1(n9548), .A2(n9565), .B1(n9547), .B2(n9641), .ZN(n9549)
         );
  AOI21_X1 U10512 ( .B1(n9551), .B2(n9550), .A(n9549), .ZN(n9708) );
  NOR2_X1 U10513 ( .A1(n9708), .A2(n10851), .ZN(n9552) );
  AOI211_X1 U10514 ( .C1(n9706), .C2(n9610), .A(n9553), .B(n9552), .ZN(n9554)
         );
  OAI21_X1 U10515 ( .B1(n9709), .B2(n9602), .A(n9554), .ZN(P2_U3274) );
  XOR2_X1 U10516 ( .A(n9560), .B(n9555), .Z(n9710) );
  AOI21_X1 U10517 ( .B1(n9557), .B2(n9572), .A(n9556), .ZN(n9713) );
  INV_X1 U10518 ( .A(n9557), .ZN(n9772) );
  INV_X1 U10519 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9558) );
  OAI22_X1 U10520 ( .A1(n9772), .A2(n9628), .B1(n10856), .B2(n9558), .ZN(n9569) );
  XOR2_X1 U10521 ( .A(n9560), .B(n9559), .Z(n9562) );
  OAI222_X1 U10522 ( .A1(n9565), .A2(n9564), .B1(n9641), .B2(n9563), .C1(n9562), .C2(n9561), .ZN(n9712) );
  AOI21_X1 U10523 ( .B1(n9566), .B2(n10755), .A(n9712), .ZN(n9567) );
  NOR2_X1 U10524 ( .A1(n9567), .A2(n10851), .ZN(n9568) );
  AOI211_X1 U10525 ( .C1(n9713), .C2(n9610), .A(n9569), .B(n9568), .ZN(n9570)
         );
  OAI21_X1 U10526 ( .B1(n9710), .B2(n9602), .A(n9570), .ZN(P2_U3275) );
  XNOR2_X1 U10527 ( .A(n9571), .B(n9577), .ZN(n9720) );
  INV_X1 U10528 ( .A(n9572), .ZN(n9573) );
  AOI21_X1 U10529 ( .B1(n9716), .B2(n9596), .A(n9573), .ZN(n9717) );
  INV_X1 U10530 ( .A(n9716), .ZN(n9576) );
  AOI22_X1 U10531 ( .A1(n10851), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9574), 
        .B2(n10755), .ZN(n9575) );
  OAI21_X1 U10532 ( .B1(n9576), .B2(n9628), .A(n9575), .ZN(n9582) );
  XNOR2_X1 U10533 ( .A(n9578), .B(n9577), .ZN(n9580) );
  AOI222_X1 U10534 ( .A1(n9644), .A2(n9580), .B1(n9579), .B2(n9638), .C1(n9604), .C2(n9619), .ZN(n9719) );
  NOR2_X1 U10535 ( .A1(n9719), .A2(n10851), .ZN(n9581) );
  AOI211_X1 U10536 ( .C1(n9717), .C2(n9610), .A(n9582), .B(n9581), .ZN(n9583)
         );
  OAI21_X1 U10537 ( .B1(n9602), .B2(n9720), .A(n9583), .ZN(P2_U3276) );
  NAND2_X1 U10538 ( .A1(n9585), .A2(n9584), .ZN(n9586) );
  NAND2_X1 U10539 ( .A1(n9587), .A2(n9586), .ZN(n9723) );
  AOI22_X1 U10540 ( .A1(n9588), .A2(n9655), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n10851), .ZN(n9601) );
  XNOR2_X1 U10541 ( .A(n9590), .B(n9589), .ZN(n9595) );
  NAND2_X1 U10542 ( .A1(n9591), .A2(n9638), .ZN(n9592) );
  OAI21_X1 U10543 ( .B1(n9593), .B2(n9641), .A(n9592), .ZN(n9594) );
  AOI21_X1 U10544 ( .B1(n9595), .B2(n9644), .A(n9594), .ZN(n9722) );
  INV_X1 U10545 ( .A(n9722), .ZN(n9599) );
  OAI211_X1 U10546 ( .C1(n9777), .C2(n5080), .A(n9746), .B(n9596), .ZN(n9721)
         );
  OAI22_X1 U10547 ( .A1(n9721), .A2(n6002), .B1(n10860), .B2(n9597), .ZN(n9598) );
  OAI21_X1 U10548 ( .B1(n9599), .B2(n9598), .A(n10856), .ZN(n9600) );
  OAI211_X1 U10549 ( .C1(n9723), .C2(n9602), .A(n9601), .B(n9600), .ZN(
        P2_U3277) );
  XNOR2_X1 U10550 ( .A(n9603), .B(n9612), .ZN(n9605) );
  AOI222_X1 U10551 ( .A1(n9644), .A2(n9605), .B1(n9604), .B2(n9638), .C1(n9639), .C2(n9619), .ZN(n9730) );
  AOI21_X1 U10552 ( .B1(n9727), .B2(n9625), .A(n5080), .ZN(n9728) );
  NOR2_X1 U10553 ( .A1(n5347), .A2(n9628), .ZN(n9609) );
  INV_X1 U10554 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9607) );
  OAI22_X1 U10555 ( .A1(n10856), .A2(n9607), .B1(n9606), .B2(n10860), .ZN(
        n9608) );
  AOI211_X1 U10556 ( .C1(n9728), .C2(n9610), .A(n9609), .B(n9608), .ZN(n9615)
         );
  OAI21_X1 U10557 ( .B1(n9613), .B2(n9612), .A(n9611), .ZN(n9726) );
  NAND2_X1 U10558 ( .A1(n9726), .A2(n9660), .ZN(n9614) );
  OAI211_X1 U10559 ( .C1(n9730), .C2(n10851), .A(n9615), .B(n9614), .ZN(
        P2_U3278) );
  XNOR2_X1 U10560 ( .A(n9616), .B(n9623), .ZN(n9617) );
  NAND2_X1 U10561 ( .A1(n9617), .A2(n9644), .ZN(n9622) );
  AOI22_X1 U10562 ( .A1(n9620), .A2(n9638), .B1(n9619), .B2(n9618), .ZN(n9621)
         );
  NAND2_X1 U10563 ( .A1(n9622), .A2(n9621), .ZN(n9732) );
  INV_X1 U10564 ( .A(n9732), .ZN(n9636) );
  XNOR2_X1 U10565 ( .A(n9624), .B(n9623), .ZN(n9734) );
  NAND2_X1 U10566 ( .A1(n9734), .A2(n9660), .ZN(n9635) );
  INV_X1 U10567 ( .A(n9625), .ZN(n9626) );
  AOI211_X1 U10568 ( .C1(n9627), .C2(n9650), .A(n10916), .B(n9626), .ZN(n9733)
         );
  INV_X1 U10569 ( .A(n9627), .ZN(n9782) );
  NOR2_X1 U10570 ( .A1(n9782), .A2(n9628), .ZN(n9632) );
  OAI22_X1 U10571 ( .A1(n10856), .A2(n9630), .B1(n9629), .B2(n10860), .ZN(
        n9631) );
  AOI211_X1 U10572 ( .C1(n9733), .C2(n9633), .A(n9632), .B(n9631), .ZN(n9634)
         );
  OAI211_X1 U10573 ( .C1(n10851), .C2(n9636), .A(n9635), .B(n9634), .ZN(
        P2_U3279) );
  XNOR2_X1 U10574 ( .A(n5081), .B(n9637), .ZN(n9645) );
  NAND2_X1 U10575 ( .A1(n9639), .A2(n9638), .ZN(n9640) );
  OAI21_X1 U10576 ( .B1(n9642), .B2(n9641), .A(n9640), .ZN(n9643) );
  AOI21_X1 U10577 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(n9738) );
  NAND2_X1 U10578 ( .A1(n9647), .A2(n9646), .ZN(n9648) );
  NAND2_X1 U10579 ( .A1(n9649), .A2(n9648), .ZN(n9739) );
  INV_X1 U10580 ( .A(n9739), .ZN(n9661) );
  OAI211_X1 U10581 ( .C1(n9787), .C2(n9651), .A(n9746), .B(n9650), .ZN(n9737)
         );
  OAI22_X1 U10582 ( .A1(n10856), .A2(n9653), .B1(n9652), .B2(n10860), .ZN(
        n9654) );
  AOI21_X1 U10583 ( .B1(n9656), .B2(n9655), .A(n9654), .ZN(n9657) );
  OAI21_X1 U10584 ( .B1(n9737), .B2(n9658), .A(n9657), .ZN(n9659) );
  AOI21_X1 U10585 ( .B1(n9661), .B2(n9660), .A(n9659), .ZN(n9662) );
  OAI21_X1 U10586 ( .B1(n10851), .B2(n9738), .A(n9662), .ZN(P2_U3280) );
  NAND3_X1 U10587 ( .A1(n9664), .A2(n9663), .A3(n9746), .ZN(n9666) );
  AND2_X1 U10588 ( .A1(n9666), .A2(n9665), .ZN(n9753) );
  MUX2_X1 U10589 ( .A(n9753), .B(n6356), .S(n10922), .Z(n9667) );
  OAI21_X1 U10590 ( .B1(n9755), .B2(n9742), .A(n9667), .ZN(P2_U3550) );
  AOI22_X1 U10591 ( .A1(n9669), .A2(n9746), .B1(n9745), .B2(n9668), .ZN(n9670)
         );
  OAI21_X1 U10592 ( .B1(n9673), .B2(n9750), .A(n9672), .ZN(n9756) );
  MUX2_X1 U10593 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9756), .S(n10923), .Z(
        P2_U3549) );
  AOI22_X1 U10594 ( .A1(n9675), .A2(n9746), .B1(n9745), .B2(n9674), .ZN(n9676)
         );
  OAI211_X1 U10595 ( .C1(n9678), .C2(n9750), .A(n9677), .B(n9676), .ZN(n9757)
         );
  MUX2_X1 U10596 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9757), .S(n10923), .Z(
        P2_U3548) );
  AOI22_X1 U10597 ( .A1(n9680), .A2(n9746), .B1(n9745), .B2(n9679), .ZN(n9681)
         );
  OAI211_X1 U10598 ( .C1(n9683), .C2(n9750), .A(n9682), .B(n9681), .ZN(n9758)
         );
  MUX2_X1 U10599 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9758), .S(n10923), .Z(
        P2_U3547) );
  AOI211_X1 U10600 ( .C1(n9687), .C2(n10921), .A(n9686), .B(n9685), .ZN(n9759)
         );
  MUX2_X1 U10601 ( .A(n9688), .B(n9759), .S(n10923), .Z(n9689) );
  OAI21_X1 U10602 ( .B1(n8806), .B2(n9742), .A(n9689), .ZN(P2_U3546) );
  AOI211_X1 U10603 ( .C1(n9692), .C2(n10921), .A(n9691), .B(n9690), .ZN(n9762)
         );
  MUX2_X1 U10604 ( .A(n9693), .B(n9762), .S(n10923), .Z(n9694) );
  OAI21_X1 U10605 ( .B1(n9765), .B2(n9742), .A(n9694), .ZN(P2_U3545) );
  AOI22_X1 U10606 ( .A1(n9696), .A2(n9746), .B1(n9745), .B2(n9695), .ZN(n9697)
         );
  OAI211_X1 U10607 ( .C1(n9699), .C2(n9750), .A(n9698), .B(n9697), .ZN(n9766)
         );
  MUX2_X1 U10608 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9766), .S(n10923), .Z(
        P2_U3544) );
  AOI22_X1 U10609 ( .A1(n9701), .A2(n9746), .B1(n9745), .B2(n9700), .ZN(n9702)
         );
  OAI211_X1 U10610 ( .C1(n9704), .C2(n9750), .A(n9703), .B(n9702), .ZN(n9767)
         );
  MUX2_X1 U10611 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9767), .S(n10923), .Z(
        P2_U3543) );
  AOI22_X1 U10612 ( .A1(n9706), .A2(n9746), .B1(n9745), .B2(n9705), .ZN(n9707)
         );
  OAI211_X1 U10613 ( .C1(n9709), .C2(n9750), .A(n9708), .B(n9707), .ZN(n9768)
         );
  MUX2_X1 U10614 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9768), .S(n10923), .Z(
        P2_U3542) );
  NOR2_X1 U10615 ( .A1(n9710), .A2(n9750), .ZN(n9711) );
  AOI211_X1 U10616 ( .C1(n9746), .C2(n9713), .A(n9712), .B(n9711), .ZN(n9769)
         );
  MUX2_X1 U10617 ( .A(n9714), .B(n9769), .S(n10923), .Z(n9715) );
  OAI21_X1 U10618 ( .B1(n9772), .B2(n9742), .A(n9715), .ZN(P2_U3541) );
  AOI22_X1 U10619 ( .A1(n9717), .A2(n9746), .B1(n9745), .B2(n9716), .ZN(n9718)
         );
  OAI211_X1 U10620 ( .C1(n9720), .C2(n9750), .A(n9719), .B(n9718), .ZN(n9773)
         );
  MUX2_X1 U10621 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9773), .S(n10923), .Z(
        P2_U3540) );
  OAI211_X1 U10622 ( .C1(n9723), .C2(n9750), .A(n9722), .B(n9721), .ZN(n9774)
         );
  MUX2_X1 U10623 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9774), .S(n10923), .Z(
        n9724) );
  INV_X1 U10624 ( .A(n9724), .ZN(n9725) );
  OAI21_X1 U10625 ( .B1(n9777), .B2(n9742), .A(n9725), .ZN(P2_U3539) );
  INV_X1 U10626 ( .A(n9726), .ZN(n9731) );
  AOI22_X1 U10627 ( .A1(n9728), .A2(n9746), .B1(n9745), .B2(n9727), .ZN(n9729)
         );
  OAI211_X1 U10628 ( .C1(n9731), .C2(n9750), .A(n9730), .B(n9729), .ZN(n9778)
         );
  MUX2_X1 U10629 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9778), .S(n10923), .Z(
        P2_U3538) );
  AOI211_X1 U10630 ( .C1(n9734), .C2(n10921), .A(n9733), .B(n9732), .ZN(n9779)
         );
  MUX2_X1 U10631 ( .A(n9735), .B(n9779), .S(n10923), .Z(n9736) );
  OAI21_X1 U10632 ( .B1(n9782), .B2(n9742), .A(n9736), .ZN(P2_U3537) );
  OAI211_X1 U10633 ( .C1(n9739), .C2(n9750), .A(n9738), .B(n9737), .ZN(n9783)
         );
  MUX2_X1 U10634 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9783), .S(n10923), .Z(
        n9740) );
  INV_X1 U10635 ( .A(n9740), .ZN(n9741) );
  OAI21_X1 U10636 ( .B1(n9787), .B2(n9742), .A(n9741), .ZN(P2_U3536) );
  INV_X1 U10637 ( .A(n9743), .ZN(n9751) );
  AOI22_X1 U10638 ( .A1(n9747), .A2(n9746), .B1(n9745), .B2(n9744), .ZN(n9748)
         );
  OAI211_X1 U10639 ( .C1(n9751), .C2(n9750), .A(n9749), .B(n9748), .ZN(n9788)
         );
  MUX2_X1 U10640 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9788), .S(n10923), .Z(
        P2_U3535) );
  INV_X1 U10641 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9752) );
  MUX2_X1 U10642 ( .A(n9753), .B(n9752), .S(n10985), .Z(n9754) );
  OAI21_X1 U10643 ( .B1(n9755), .B2(n9786), .A(n9754), .ZN(P2_U3518) );
  MUX2_X1 U10644 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9756), .S(n5011), .Z(
        P2_U3517) );
  MUX2_X1 U10645 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9757), .S(n5011), .Z(
        P2_U3516) );
  MUX2_X1 U10646 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9758), .S(n5011), .Z(
        P2_U3515) );
  INV_X1 U10647 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9760) );
  MUX2_X1 U10648 ( .A(n9760), .B(n9759), .S(n5011), .Z(n9761) );
  OAI21_X1 U10649 ( .B1(n8806), .B2(n9786), .A(n9761), .ZN(P2_U3514) );
  INV_X1 U10650 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9763) );
  MUX2_X1 U10651 ( .A(n9763), .B(n9762), .S(n5011), .Z(n9764) );
  OAI21_X1 U10652 ( .B1(n9765), .B2(n9786), .A(n9764), .ZN(P2_U3513) );
  MUX2_X1 U10653 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9766), .S(n5011), .Z(
        P2_U3512) );
  MUX2_X1 U10654 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9767), .S(n5011), .Z(
        P2_U3511) );
  MUX2_X1 U10655 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9768), .S(n5011), .Z(
        P2_U3510) );
  INV_X1 U10656 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9770) );
  MUX2_X1 U10657 ( .A(n9770), .B(n9769), .S(n5011), .Z(n9771) );
  OAI21_X1 U10658 ( .B1(n9772), .B2(n9786), .A(n9771), .ZN(P2_U3509) );
  MUX2_X1 U10659 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9773), .S(n5011), .Z(
        P2_U3508) );
  MUX2_X1 U10660 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9774), .S(n5011), .Z(n9775) );
  INV_X1 U10661 ( .A(n9775), .ZN(n9776) );
  OAI21_X1 U10662 ( .B1(n9777), .B2(n9786), .A(n9776), .ZN(P2_U3507) );
  MUX2_X1 U10663 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9778), .S(n5011), .Z(
        P2_U3505) );
  INV_X1 U10664 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9780) );
  MUX2_X1 U10665 ( .A(n9780), .B(n9779), .S(n5011), .Z(n9781) );
  OAI21_X1 U10666 ( .B1(n9782), .B2(n9786), .A(n9781), .ZN(P2_U3502) );
  MUX2_X1 U10667 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9783), .S(n5011), .Z(n9784) );
  INV_X1 U10668 ( .A(n9784), .ZN(n9785) );
  OAI21_X1 U10669 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(P2_U3499) );
  MUX2_X1 U10670 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9788), .S(n5011), .Z(
        P2_U3496) );
  NAND3_X1 U10671 ( .A1(n9789), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9791) );
  OAI22_X1 U10672 ( .A1(n9792), .A2(n9791), .B1(n9790), .B2(n8831), .ZN(n9793)
         );
  AOI21_X1 U10673 ( .B1(n10537), .B2(n9794), .A(n9793), .ZN(n9795) );
  INV_X1 U10674 ( .A(n9795), .ZN(P2_U3327) );
  INV_X1 U10675 ( .A(n9796), .ZN(n9797) );
  MUX2_X1 U10676 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9797), .S(P2_U3152), .Z(
        P2_U3358) );
  NAND2_X1 U10677 ( .A1(n9800), .A2(n9799), .ZN(n9801) );
  XOR2_X1 U10678 ( .A(n9802), .B(n9801), .Z(n9811) );
  NOR2_X1 U10679 ( .A1(n9803), .A2(n9919), .ZN(n9804) );
  AOI211_X1 U10680 ( .C1(n9923), .C2(n10870), .A(n9805), .B(n9804), .ZN(n9806)
         );
  OAI21_X1 U10681 ( .B1(n9926), .B2(n9807), .A(n9806), .ZN(n9808) );
  AOI21_X1 U10682 ( .B1(n9809), .B2(n9928), .A(n9808), .ZN(n9810) );
  OAI21_X1 U10683 ( .B1(n9811), .B2(n9931), .A(n9810), .ZN(P1_U3213) );
  INV_X1 U10684 ( .A(n9812), .ZN(n9813) );
  NOR2_X1 U10685 ( .A1(n9814), .A2(n9813), .ZN(n9816) );
  XNOR2_X1 U10686 ( .A(n9816), .B(n9815), .ZN(n9821) );
  AOI22_X1 U10687 ( .A1(n9906), .A2(n10334), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(n5013), .ZN(n9818) );
  NAND2_X1 U10688 ( .A1(n9923), .A2(n10335), .ZN(n9817) );
  OAI211_X1 U10689 ( .C1(n9926), .C2(n10326), .A(n9818), .B(n9817), .ZN(n9819)
         );
  AOI21_X1 U10690 ( .B1(n10484), .B2(n9928), .A(n9819), .ZN(n9820) );
  OAI21_X1 U10691 ( .B1(n9821), .B2(n9931), .A(n9820), .ZN(P1_U3214) );
  XNOR2_X1 U10692 ( .A(n5079), .B(n9822), .ZN(n9823) );
  XNOR2_X1 U10693 ( .A(n9824), .B(n9823), .ZN(n9829) );
  NOR2_X1 U10694 ( .A1(n9926), .A2(n10392), .ZN(n9827) );
  NAND2_X1 U10695 ( .A1(n9923), .A2(n10435), .ZN(n9825) );
  NAND2_X1 U10696 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10243)
         );
  OAI211_X1 U10697 ( .C1(n10402), .C2(n9919), .A(n9825), .B(n10243), .ZN(n9826) );
  AOI211_X1 U10698 ( .C1(n10506), .C2(n9928), .A(n9827), .B(n9826), .ZN(n9828)
         );
  OAI21_X1 U10699 ( .B1(n9829), .B2(n9931), .A(n9828), .ZN(P1_U3217) );
  NAND2_X1 U10700 ( .A1(n5087), .A2(n9831), .ZN(n9832) );
  XNOR2_X1 U10701 ( .A(n9830), .B(n9832), .ZN(n9837) );
  AOI22_X1 U10702 ( .A1(n9906), .A2(n10335), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9834) );
  NAND2_X1 U10703 ( .A1(n10359), .A2(n9923), .ZN(n9833) );
  OAI211_X1 U10704 ( .C1(n9926), .C2(n10361), .A(n9834), .B(n9833), .ZN(n9835)
         );
  AOI21_X1 U10705 ( .B1(n10496), .B2(n9928), .A(n9835), .ZN(n9836) );
  OAI21_X1 U10706 ( .B1(n9837), .B2(n9931), .A(n9836), .ZN(P1_U3221) );
  XNOR2_X1 U10707 ( .A(n9840), .B(n9839), .ZN(n9841) );
  XNOR2_X1 U10708 ( .A(n9838), .B(n9841), .ZN(n9846) );
  AOI22_X1 U10709 ( .A1(n9906), .A2(n10201), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(n5013), .ZN(n9843) );
  NAND2_X1 U10710 ( .A1(n9923), .A2(n10334), .ZN(n9842) );
  OAI211_X1 U10711 ( .C1(n9926), .C2(n10295), .A(n9843), .B(n9842), .ZN(n9844)
         );
  AOI21_X1 U10712 ( .B1(n10474), .B2(n9928), .A(n9844), .ZN(n9845) );
  OAI21_X1 U10713 ( .B1(n9846), .B2(n9931), .A(n9845), .ZN(P1_U3223) );
  INV_X1 U10714 ( .A(n9848), .ZN(n9849) );
  AOI21_X1 U10715 ( .B1(n9850), .B2(n9847), .A(n9849), .ZN(n9855) );
  AOI22_X1 U10716 ( .A1(n9906), .A2(n10943), .B1(P1_REG3_REG_16__SCAN_IN), 
        .B2(n5013), .ZN(n9852) );
  NAND2_X1 U10717 ( .A1(n9923), .A2(n10945), .ZN(n9851) );
  OAI211_X1 U10718 ( .C1(n9926), .C2(n10956), .A(n9852), .B(n9851), .ZN(n9853)
         );
  AOI21_X1 U10719 ( .B1(n10960), .B2(n9928), .A(n9853), .ZN(n9854) );
  OAI21_X1 U10720 ( .B1(n9855), .B2(n9931), .A(n9854), .ZN(P1_U3224) );
  XOR2_X1 U10721 ( .A(n9857), .B(n9858), .Z(n9863) );
  AOI22_X1 U10722 ( .A1(n9923), .A2(n10436), .B1(P1_REG3_REG_17__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9860) );
  NAND2_X1 U10723 ( .A1(n9906), .A2(n10435), .ZN(n9859) );
  OAI211_X1 U10724 ( .C1(n9926), .C2(n10442), .A(n9860), .B(n9859), .ZN(n9861)
         );
  AOI21_X1 U10725 ( .B1(n10516), .B2(n9928), .A(n9861), .ZN(n9862) );
  OAI21_X1 U10726 ( .B1(n9863), .B2(n9931), .A(n9862), .ZN(P1_U3226) );
  XOR2_X1 U10727 ( .A(n9865), .B(n9864), .Z(n9870) );
  AOI22_X1 U10728 ( .A1(n9906), .A2(n10288), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(n5013), .ZN(n9867) );
  NAND2_X1 U10729 ( .A1(n9923), .A2(n10202), .ZN(n9866) );
  OAI211_X1 U10730 ( .C1(n9926), .C2(n10318), .A(n9867), .B(n9866), .ZN(n9868)
         );
  AOI21_X1 U10731 ( .B1(n10481), .B2(n9928), .A(n9868), .ZN(n9869) );
  OAI21_X1 U10732 ( .B1(n9870), .B2(n9931), .A(n9869), .ZN(P1_U3227) );
  NOR2_X1 U10733 ( .A1(n9872), .A2(n5082), .ZN(n9873) );
  XNOR2_X1 U10734 ( .A(n9871), .B(n9873), .ZN(n9878) );
  NAND2_X1 U10735 ( .A1(n10374), .A2(n9906), .ZN(n9875) );
  AOI22_X1 U10736 ( .A1(n10418), .A2(n9923), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(n5013), .ZN(n9874) );
  OAI211_X1 U10737 ( .C1(n9926), .C2(n10380), .A(n9875), .B(n9874), .ZN(n9876)
         );
  AOI21_X1 U10738 ( .B1(n10500), .B2(n9928), .A(n9876), .ZN(n9877) );
  OAI21_X1 U10739 ( .B1(n9878), .B2(n9931), .A(n9877), .ZN(P1_U3231) );
  INV_X1 U10740 ( .A(n9880), .ZN(n9881) );
  NOR2_X1 U10741 ( .A1(n9882), .A2(n9881), .ZN(n9883) );
  XNOR2_X1 U10742 ( .A(n9879), .B(n9883), .ZN(n9888) );
  NAND2_X1 U10743 ( .A1(n10374), .A2(n9923), .ZN(n9885) );
  AOI22_X1 U10744 ( .A1(n9906), .A2(n10202), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9884) );
  OAI211_X1 U10745 ( .C1(n9926), .C2(n10341), .A(n9885), .B(n9884), .ZN(n9886)
         );
  AOI21_X1 U10746 ( .B1(n10491), .B2(n9928), .A(n9886), .ZN(n9887) );
  OAI21_X1 U10747 ( .B1(n9888), .B2(n9931), .A(n9887), .ZN(P1_U3233) );
  INV_X1 U10748 ( .A(n9889), .ZN(n9895) );
  OAI21_X1 U10749 ( .B1(n9890), .B2(n9894), .A(n9891), .ZN(n9892) );
  OAI211_X1 U10750 ( .C1(n9895), .C2(n9894), .A(n9893), .B(n9892), .ZN(n9902)
         );
  NOR2_X1 U10751 ( .A1(n9896), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10656) );
  AOI21_X1 U10752 ( .B1(n9923), .B2(n10943), .A(n10656), .ZN(n9897) );
  OAI21_X1 U10753 ( .B1(n9898), .B2(n9919), .A(n9897), .ZN(n9899) );
  AOI21_X1 U10754 ( .B1(n10425), .B2(n9900), .A(n9899), .ZN(n9901) );
  OAI211_X1 U10755 ( .C1(n8782), .C2(n9903), .A(n9902), .B(n9901), .ZN(
        P1_U3236) );
  XNOR2_X1 U10756 ( .A(n9905), .B(n9904), .ZN(n9911) );
  AOI22_X1 U10757 ( .A1(n9906), .A2(n10287), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9908) );
  NAND2_X1 U10758 ( .A1(n9923), .A2(n10288), .ZN(n9907) );
  OAI211_X1 U10759 ( .C1(n9926), .C2(n10280), .A(n9908), .B(n9907), .ZN(n9909)
         );
  AOI21_X1 U10760 ( .B1(n10469), .B2(n9928), .A(n9909), .ZN(n9910) );
  OAI21_X1 U10761 ( .B1(n9911), .B2(n9931), .A(n9910), .ZN(P1_U3238) );
  INV_X1 U10762 ( .A(n9847), .ZN(n9917) );
  NAND2_X1 U10763 ( .A1(n9913), .A2(n9914), .ZN(n9915) );
  AOI22_X1 U10764 ( .A1(n9917), .A2(n9913), .B1(n9916), .B2(n9915), .ZN(n9932)
         );
  INV_X1 U10765 ( .A(n9918), .ZN(n9922) );
  NOR2_X1 U10766 ( .A1(n9920), .A2(n9919), .ZN(n9921) );
  AOI211_X1 U10767 ( .C1(n9923), .C2(n10203), .A(n9922), .B(n9921), .ZN(n9924)
         );
  OAI21_X1 U10768 ( .B1(n9926), .B2(n9925), .A(n9924), .ZN(n9927) );
  AOI21_X1 U10769 ( .B1(n9929), .B2(n9928), .A(n9927), .ZN(n9930) );
  OAI21_X1 U10770 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(P1_U3239) );
  NOR2_X1 U10771 ( .A1(n10017), .A2(n10196), .ZN(n10198) );
  NOR3_X1 U10772 ( .A1(n9933), .A2(n7127), .A3(n7155), .ZN(n10197) );
  INV_X1 U10773 ( .A(n10007), .ZN(n10014) );
  OR2_X1 U10774 ( .A1(n10258), .A2(n10109), .ZN(n10111) );
  XNOR2_X1 U10775 ( .A(n9934), .B(n10007), .ZN(n9938) );
  NAND2_X1 U10776 ( .A1(n9939), .A2(n9935), .ZN(n10118) );
  NAND2_X1 U10777 ( .A1(n10043), .A2(n10126), .ZN(n9936) );
  MUX2_X1 U10778 ( .A(n10118), .B(n9936), .S(n10007), .Z(n9937) );
  AOI21_X1 U10779 ( .B1(n9938), .B2(n10159), .A(n9937), .ZN(n9944) );
  INV_X1 U10780 ( .A(n9939), .ZN(n9940) );
  MUX2_X1 U10781 ( .A(n9941), .B(n9940), .S(n10007), .Z(n9943) );
  INV_X1 U10782 ( .A(n9942), .ZN(n10158) );
  OAI21_X1 U10783 ( .B1(n9944), .B2(n9943), .A(n10158), .ZN(n9946) );
  MUX2_X1 U10784 ( .A(n10042), .B(n10065), .S(n10007), .Z(n9945) );
  AOI21_X1 U10785 ( .B1(n9946), .B2(n9945), .A(n10162), .ZN(n9951) );
  MUX2_X1 U10786 ( .A(n10037), .B(n10064), .S(n10007), .Z(n9947) );
  NAND2_X1 U10787 ( .A1(n10809), .A2(n9947), .ZN(n9950) );
  INV_X1 U10788 ( .A(n9948), .ZN(n10165) );
  MUX2_X1 U10789 ( .A(n10066), .B(n10038), .S(n10007), .Z(n9949) );
  OAI211_X1 U10790 ( .C1(n9951), .C2(n9950), .A(n10165), .B(n9949), .ZN(n9952)
         );
  OAI211_X1 U10791 ( .C1(n10041), .C2(n10007), .A(n9952), .B(n10868), .ZN(
        n9954) );
  AOI21_X1 U10792 ( .B1(n9954), .B2(n10069), .A(n5406), .ZN(n9957) );
  INV_X1 U10793 ( .A(n10068), .ZN(n9953) );
  OAI21_X1 U10794 ( .B1(n9954), .B2(n9953), .A(n10073), .ZN(n9955) );
  AND2_X1 U10795 ( .A1(n9955), .A2(n10076), .ZN(n9956) );
  MUX2_X1 U10796 ( .A(n9957), .B(n9956), .S(n10007), .Z(n9959) );
  MUX2_X1 U10797 ( .A(n10035), .B(n10077), .S(n10007), .Z(n9958) );
  OAI21_X1 U10798 ( .B1(n9959), .B2(n10168), .A(n9958), .ZN(n9965) );
  INV_X1 U10799 ( .A(n10076), .ZN(n9960) );
  NAND2_X1 U10800 ( .A1(n10035), .A2(n9960), .ZN(n9962) );
  NAND2_X1 U10801 ( .A1(n10077), .A2(n5406), .ZN(n9961) );
  MUX2_X1 U10802 ( .A(n9962), .B(n9961), .S(n10007), .Z(n9963) );
  MUX2_X1 U10803 ( .A(n10036), .B(n10081), .S(n10007), .Z(n9966) );
  MUX2_X1 U10804 ( .A(n10082), .B(n10031), .S(n10007), .Z(n9967) );
  AOI21_X1 U10805 ( .B1(n9968), .B2(n9967), .A(n5380), .ZN(n9972) );
  MUX2_X1 U10806 ( .A(n10024), .B(n10032), .S(n10007), .Z(n9969) );
  NAND2_X1 U10807 ( .A1(n10410), .A2(n9969), .ZN(n9971) );
  INV_X1 U10808 ( .A(n10397), .ZN(n10389) );
  MUX2_X1 U10809 ( .A(n10034), .B(n10025), .S(n10007), .Z(n9970) );
  MUX2_X1 U10810 ( .A(n10027), .B(n10132), .S(n10007), .Z(n9973) );
  AOI21_X1 U10811 ( .B1(n9974), .B2(n9973), .A(n10357), .ZN(n9982) );
  NOR2_X1 U10812 ( .A1(n10030), .A2(n9975), .ZN(n9980) );
  NAND2_X1 U10813 ( .A1(n10500), .A2(n10402), .ZN(n9976) );
  NAND2_X1 U10814 ( .A1(n9977), .A2(n9976), .ZN(n9979) );
  AND2_X1 U10815 ( .A1(n9979), .A2(n9978), .ZN(n10088) );
  MUX2_X1 U10816 ( .A(n9980), .B(n10088), .S(n10007), .Z(n9981) );
  NAND2_X1 U10817 ( .A1(n10330), .A2(n10090), .ZN(n10344) );
  AOI211_X1 U10818 ( .C1(n9982), .C2(n10372), .A(n9981), .B(n10344), .ZN(n9986) );
  XNOR2_X1 U10819 ( .A(n10484), .B(n10348), .ZN(n10332) );
  INV_X1 U10820 ( .A(n10330), .ZN(n9984) );
  INV_X1 U10821 ( .A(n10090), .ZN(n9983) );
  MUX2_X1 U10822 ( .A(n9984), .B(n9983), .S(n10014), .Z(n9985) );
  NOR3_X1 U10823 ( .A1(n9986), .A2(n10332), .A3(n9985), .ZN(n9994) );
  INV_X1 U10824 ( .A(n9991), .ZN(n9987) );
  NOR2_X1 U10825 ( .A1(n10023), .A2(n9987), .ZN(n10313) );
  MUX2_X1 U10826 ( .A(n9988), .B(n10310), .S(n10007), .Z(n9989) );
  NAND2_X1 U10827 ( .A1(n10313), .A2(n9989), .ZN(n9993) );
  INV_X1 U10828 ( .A(n10300), .ZN(n10175) );
  INV_X1 U10829 ( .A(n10023), .ZN(n9990) );
  MUX2_X1 U10830 ( .A(n9991), .B(n9990), .S(n10007), .Z(n9992) );
  MUX2_X1 U10831 ( .A(n10020), .B(n10105), .S(n10007), .Z(n9995) );
  NAND3_X1 U10832 ( .A1(n9996), .A2(n10286), .A3(n9995), .ZN(n9999) );
  INV_X1 U10833 ( .A(n10271), .ZN(n9998) );
  MUX2_X1 U10834 ( .A(n10021), .B(n10098), .S(n10014), .Z(n9997) );
  INV_X1 U10835 ( .A(n10101), .ZN(n10000) );
  NAND2_X1 U10836 ( .A1(n10003), .A2(n10005), .ZN(n10009) );
  NAND2_X1 U10837 ( .A1(n10005), .A2(n10004), .ZN(n10145) );
  OAI21_X1 U10838 ( .B1(n10006), .B2(n10145), .A(n10144), .ZN(n10008) );
  OR2_X1 U10839 ( .A1(n10012), .A2(n10109), .ZN(n10010) );
  NAND2_X1 U10840 ( .A1(n10258), .A2(n10010), .ZN(n10143) );
  NAND2_X1 U10841 ( .A1(n10448), .A2(n10012), .ZN(n10112) );
  OR2_X1 U10842 ( .A1(n10111), .A2(n10012), .ZN(n10013) );
  NAND2_X1 U10843 ( .A1(n10112), .A2(n10013), .ZN(n10116) );
  AOI22_X1 U10844 ( .A1(n10015), .A2(n10112), .B1(n10014), .B2(n10116), .ZN(
        n10019) );
  INV_X1 U10845 ( .A(n10182), .ZN(n10147) );
  AND2_X1 U10846 ( .A1(n10021), .A2(n10020), .ZN(n10022) );
  NAND2_X1 U10847 ( .A1(n10100), .A2(n10022), .ZN(n10106) );
  NOR2_X1 U10848 ( .A1(n10106), .A2(n10023), .ZN(n10142) );
  INV_X1 U10849 ( .A(n10142), .ZN(n10097) );
  NAND2_X1 U10850 ( .A1(n10025), .A2(n10024), .ZN(n10026) );
  NAND3_X1 U10851 ( .A1(n10132), .A2(n10034), .A3(n10026), .ZN(n10028) );
  AND2_X1 U10852 ( .A1(n10028), .A2(n10027), .ZN(n10029) );
  AND2_X1 U10853 ( .A1(n10030), .A2(n10029), .ZN(n10137) );
  INV_X1 U10854 ( .A(n10137), .ZN(n10093) );
  AND2_X1 U10855 ( .A1(n10032), .A2(n10031), .ZN(n10033) );
  NAND2_X1 U10856 ( .A1(n10034), .A2(n10033), .ZN(n10062) );
  NAND2_X1 U10857 ( .A1(n10036), .A2(n10035), .ZN(n10063) );
  NAND2_X1 U10858 ( .A1(n10038), .A2(n10037), .ZN(n10039) );
  NAND2_X1 U10859 ( .A1(n10039), .A2(n10066), .ZN(n10040) );
  AND2_X1 U10860 ( .A1(n10041), .A2(n10040), .ZN(n10067) );
  AND4_X1 U10861 ( .A1(n10073), .A2(n10067), .A3(n10043), .A4(n10042), .ZN(
        n10044) );
  NAND2_X1 U10862 ( .A1(n10074), .A2(n10044), .ZN(n10045) );
  OR3_X1 U10863 ( .A1(n10062), .A2(n10063), .A3(n10045), .ZN(n10129) );
  INV_X1 U10864 ( .A(n10046), .ZN(n10050) );
  NAND2_X1 U10865 ( .A1(n7836), .A2(n10047), .ZN(n10048) );
  NAND3_X1 U10866 ( .A1(n10050), .A2(n10049), .A3(n10048), .ZN(n10051) );
  NAND2_X1 U10867 ( .A1(n10052), .A2(n10051), .ZN(n10055) );
  OAI22_X1 U10868 ( .A1(n7924), .A2(n10055), .B1(n10054), .B2(n10053), .ZN(
        n10056) );
  NAND2_X1 U10869 ( .A1(n10056), .A2(n10119), .ZN(n10057) );
  NAND2_X1 U10870 ( .A1(n10057), .A2(n10123), .ZN(n10061) );
  INV_X1 U10871 ( .A(n10058), .ZN(n10059) );
  AOI211_X1 U10872 ( .C1(n10061), .C2(n10060), .A(n10059), .B(n10118), .ZN(
        n10086) );
  INV_X1 U10873 ( .A(n10062), .ZN(n10084) );
  INV_X1 U10874 ( .A(n10063), .ZN(n10079) );
  AND3_X1 U10875 ( .A1(n10066), .A2(n10065), .A3(n10064), .ZN(n10071) );
  INV_X1 U10876 ( .A(n10067), .ZN(n10070) );
  OAI211_X1 U10877 ( .C1(n10071), .C2(n10070), .A(n10069), .B(n10068), .ZN(
        n10072) );
  NAND3_X1 U10878 ( .A1(n10074), .A2(n10073), .A3(n10072), .ZN(n10075) );
  NAND3_X1 U10879 ( .A1(n10077), .A2(n10076), .A3(n10075), .ZN(n10078) );
  NAND2_X1 U10880 ( .A1(n10079), .A2(n10078), .ZN(n10080) );
  NAND3_X1 U10881 ( .A1(n10082), .A2(n10081), .A3(n10080), .ZN(n10083) );
  AND2_X1 U10882 ( .A1(n10084), .A2(n10083), .ZN(n10133) );
  INV_X1 U10883 ( .A(n10133), .ZN(n10085) );
  OAI21_X1 U10884 ( .B1(n10129), .B2(n10086), .A(n10085), .ZN(n10087) );
  AND2_X1 U10885 ( .A1(n10087), .A2(n10132), .ZN(n10092) );
  INV_X1 U10886 ( .A(n10088), .ZN(n10089) );
  NAND2_X1 U10887 ( .A1(n10090), .A2(n10089), .ZN(n10135) );
  INV_X1 U10888 ( .A(n10135), .ZN(n10091) );
  OAI21_X1 U10889 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(n10094) );
  NAND2_X1 U10890 ( .A1(n10117), .A2(n10094), .ZN(n10095) );
  AND2_X1 U10891 ( .A1(n10138), .A2(n10095), .ZN(n10096) );
  NOR2_X1 U10892 ( .A1(n10097), .A2(n10096), .ZN(n10108) );
  INV_X1 U10893 ( .A(n10098), .ZN(n10099) );
  NAND2_X1 U10894 ( .A1(n10100), .A2(n10099), .ZN(n10102) );
  AND2_X1 U10895 ( .A1(n10102), .A2(n10101), .ZN(n10104) );
  OAI211_X1 U10896 ( .C1(n10106), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        n10140) );
  INV_X1 U10897 ( .A(n10145), .ZN(n10107) );
  OAI21_X1 U10898 ( .B1(n10108), .B2(n10140), .A(n10107), .ZN(n10110) );
  NAND2_X1 U10899 ( .A1(n10258), .A2(n10109), .ZN(n10179) );
  AND3_X1 U10900 ( .A1(n10110), .A2(n10144), .A3(n10179), .ZN(n10113) );
  NAND2_X1 U10901 ( .A1(n10112), .A2(n10111), .ZN(n10184) );
  OR2_X1 U10902 ( .A1(n10113), .A2(n10184), .ZN(n10114) );
  NAND2_X1 U10903 ( .A1(n10114), .A2(n10182), .ZN(n10193) );
  AOI21_X1 U10904 ( .B1(n10193), .B2(n10366), .A(n10115), .ZN(n10189) );
  INV_X1 U10905 ( .A(n10116), .ZN(n10149) );
  INV_X1 U10906 ( .A(n10118), .ZN(n10131) );
  NAND2_X1 U10907 ( .A1(n10120), .A2(n10119), .ZN(n10121) );
  AOI22_X1 U10908 ( .A1(n10124), .A2(n10123), .B1(n10122), .B2(n10121), .ZN(
        n10128) );
  OAI211_X1 U10909 ( .C1(n10128), .C2(n10127), .A(n10126), .B(n10125), .ZN(
        n10130) );
  AOI21_X1 U10910 ( .B1(n10131), .B2(n10130), .A(n10129), .ZN(n10134) );
  OAI21_X1 U10911 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(n10136) );
  AOI21_X1 U10912 ( .B1(n10137), .B2(n10136), .A(n10135), .ZN(n10139) );
  OAI21_X1 U10913 ( .B1(n5393), .B2(n10139), .A(n10138), .ZN(n10141) );
  AOI21_X1 U10914 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(n10146) );
  OAI211_X1 U10915 ( .C1(n10146), .C2(n10145), .A(n10144), .B(n10143), .ZN(
        n10148) );
  AOI211_X1 U10916 ( .C1(n10149), .C2(n10148), .A(n10183), .B(n10147), .ZN(
        n10150) );
  NOR2_X1 U10917 ( .A1(n10150), .A2(n10366), .ZN(n10187) );
  INV_X1 U10918 ( .A(n10151), .ZN(n10181) );
  INV_X1 U10919 ( .A(n10286), .ZN(n10177) );
  INV_X1 U10920 ( .A(n10372), .ZN(n10370) );
  NAND2_X1 U10921 ( .A1(n10153), .A2(n10152), .ZN(n10156) );
  NOR4_X1 U10922 ( .A1(n10156), .A2(n10155), .A3(n7833), .A4(n10154), .ZN(
        n10160) );
  NAND4_X1 U10923 ( .A1(n10160), .A2(n10159), .A3(n10158), .A4(n10157), .ZN(
        n10163) );
  NOR4_X1 U10924 ( .A1(n10163), .A2(n10162), .A3(n10798), .A4(n10161), .ZN(
        n10164) );
  NAND4_X1 U10925 ( .A1(n10166), .A2(n10165), .A3(n10868), .A4(n10164), .ZN(
        n10167) );
  NOR4_X1 U10926 ( .A1(n10936), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10170) );
  NAND4_X1 U10927 ( .A1(n10389), .A2(n10171), .A3(n10410), .A4(n10170), .ZN(
        n10172) );
  NOR4_X1 U10928 ( .A1(n10344), .A2(n10357), .A3(n10370), .A4(n10172), .ZN(
        n10174) );
  INV_X1 U10929 ( .A(n10332), .ZN(n10173) );
  NAND4_X1 U10930 ( .A1(n10175), .A2(n10313), .A3(n10174), .A4(n10173), .ZN(
        n10176) );
  NOR4_X1 U10931 ( .A1(n10178), .A2(n10271), .A3(n10177), .A4(n10176), .ZN(
        n10180) );
  NAND4_X1 U10932 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10185) );
  OAI21_X1 U10933 ( .B1(n10185), .B2(n10184), .A(n10183), .ZN(n10186) );
  MUX2_X1 U10934 ( .A(n5604), .B(n10187), .S(n10186), .Z(n10188) );
  NOR4_X1 U10935 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n10195) );
  NOR2_X1 U10936 ( .A1(n10193), .A2(n10192), .ZN(n10194) );
  OAI33_X1 U10937 ( .A1(n10199), .A2(n10198), .A3(n10197), .B1(n10196), .B2(
        n10195), .B3(n10194), .ZN(P1_U3240) );
  MUX2_X1 U10938 ( .A(n10200), .B(P1_DATAO_REG_28__SCAN_IN), .S(n10211), .Z(
        P1_U3583) );
  MUX2_X1 U10939 ( .A(n10287), .B(P1_DATAO_REG_27__SCAN_IN), .S(n10211), .Z(
        P1_U3582) );
  MUX2_X1 U10940 ( .A(n10201), .B(P1_DATAO_REG_26__SCAN_IN), .S(n10211), .Z(
        P1_U3581) );
  MUX2_X1 U10941 ( .A(n10288), .B(P1_DATAO_REG_25__SCAN_IN), .S(n10211), .Z(
        P1_U3580) );
  MUX2_X1 U10942 ( .A(n10334), .B(P1_DATAO_REG_24__SCAN_IN), .S(n10211), .Z(
        P1_U3579) );
  MUX2_X1 U10943 ( .A(n10202), .B(P1_DATAO_REG_23__SCAN_IN), .S(n10211), .Z(
        P1_U3578) );
  MUX2_X1 U10944 ( .A(n10335), .B(P1_DATAO_REG_22__SCAN_IN), .S(n10211), .Z(
        P1_U3577) );
  MUX2_X1 U10945 ( .A(n10374), .B(P1_DATAO_REG_21__SCAN_IN), .S(n10211), .Z(
        P1_U3576) );
  MUX2_X1 U10946 ( .A(n10359), .B(P1_DATAO_REG_20__SCAN_IN), .S(n10211), .Z(
        P1_U3575) );
  MUX2_X1 U10947 ( .A(n10418), .B(P1_DATAO_REG_19__SCAN_IN), .S(n10211), .Z(
        P1_U3574) );
  MUX2_X1 U10948 ( .A(n10435), .B(P1_DATAO_REG_18__SCAN_IN), .S(n10211), .Z(
        P1_U3573) );
  MUX2_X1 U10949 ( .A(n10943), .B(P1_DATAO_REG_17__SCAN_IN), .S(n10211), .Z(
        P1_U3572) );
  MUX2_X1 U10950 ( .A(n10436), .B(P1_DATAO_REG_16__SCAN_IN), .S(n10211), .Z(
        P1_U3571) );
  MUX2_X1 U10951 ( .A(n10945), .B(P1_DATAO_REG_15__SCAN_IN), .S(n10211), .Z(
        P1_U3570) );
  MUX2_X1 U10952 ( .A(n10203), .B(P1_DATAO_REG_14__SCAN_IN), .S(n10211), .Z(
        P1_U3569) );
  MUX2_X1 U10953 ( .A(n10870), .B(P1_DATAO_REG_13__SCAN_IN), .S(n10211), .Z(
        P1_U3568) );
  MUX2_X1 U10954 ( .A(n10204), .B(P1_DATAO_REG_12__SCAN_IN), .S(n10211), .Z(
        P1_U3567) );
  MUX2_X1 U10955 ( .A(n10871), .B(P1_DATAO_REG_11__SCAN_IN), .S(n10211), .Z(
        P1_U3566) );
  MUX2_X1 U10956 ( .A(n10205), .B(P1_DATAO_REG_10__SCAN_IN), .S(n10211), .Z(
        P1_U3565) );
  MUX2_X1 U10957 ( .A(n10811), .B(P1_DATAO_REG_9__SCAN_IN), .S(n10211), .Z(
        P1_U3564) );
  MUX2_X1 U10958 ( .A(n10206), .B(P1_DATAO_REG_7__SCAN_IN), .S(n10211), .Z(
        P1_U3562) );
  MUX2_X1 U10959 ( .A(n10207), .B(P1_DATAO_REG_6__SCAN_IN), .S(n10211), .Z(
        P1_U3561) );
  MUX2_X1 U10960 ( .A(n10208), .B(P1_DATAO_REG_5__SCAN_IN), .S(n10211), .Z(
        P1_U3560) );
  MUX2_X1 U10961 ( .A(n10209), .B(P1_DATAO_REG_4__SCAN_IN), .S(n10211), .Z(
        P1_U3559) );
  MUX2_X1 U10962 ( .A(n10210), .B(P1_DATAO_REG_3__SCAN_IN), .S(n10211), .Z(
        P1_U3558) );
  MUX2_X1 U10963 ( .A(n7830), .B(P1_DATAO_REG_2__SCAN_IN), .S(n10211), .Z(
        P1_U3557) );
  MUX2_X1 U10964 ( .A(n7836), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10211), .Z(
        P1_U3556) );
  OAI211_X1 U10965 ( .C1(n10214), .C2(n10213), .A(n10649), .B(n10212), .ZN(
        n10223) );
  OAI211_X1 U10966 ( .C1(n10218), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        n10222) );
  AOI22_X1 U10967 ( .A1(n10648), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n5013), .ZN(n10221) );
  NAND2_X1 U10968 ( .A1(n10657), .A2(n10219), .ZN(n10220) );
  NAND4_X1 U10969 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        P1_U3242) );
  AOI211_X1 U10970 ( .C1(n10226), .C2(n10225), .A(n10224), .B(n10651), .ZN(
        n10227) );
  AOI21_X1 U10971 ( .B1(n10657), .B2(n10228), .A(n10227), .ZN(n10237) );
  INV_X1 U10972 ( .A(n10229), .ZN(n10236) );
  NAND2_X1 U10973 ( .A1(n10648), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n10235) );
  OAI21_X1 U10974 ( .B1(n10232), .B2(n10231), .A(n10230), .ZN(n10233) );
  NAND2_X1 U10975 ( .A1(n10649), .A2(n10233), .ZN(n10234) );
  NAND4_X1 U10976 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        P1_U3251) );
  AOI21_X1 U10977 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n10245), .A(n10238), 
        .ZN(n10647) );
  AOI22_X1 U10978 ( .A1(n10658), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n10240), 
        .B2(n10239), .ZN(n10646) );
  NAND2_X1 U10979 ( .A1(n10647), .A2(n10646), .ZN(n10645) );
  OAI21_X1 U10980 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n10658), .A(n10645), 
        .ZN(n10242) );
  XNOR2_X1 U10981 ( .A(n10366), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n10241) );
  XNOR2_X1 U10982 ( .A(n10242), .B(n10241), .ZN(n10255) );
  INV_X1 U10983 ( .A(n10243), .ZN(n10252) );
  MUX2_X1 U10984 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n10393), .S(n10366), .Z(
        n10248) );
  AOI21_X1 U10985 ( .B1(n10245), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10244), 
        .ZN(n10654) );
  NAND2_X1 U10986 ( .A1(n10658), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10246) );
  OAI21_X1 U10987 ( .B1(n10658), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10246), 
        .ZN(n10653) );
  NOR2_X1 U10988 ( .A1(n10654), .A2(n10653), .ZN(n10652) );
  AOI21_X1 U10989 ( .B1(n10658), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10652), 
        .ZN(n10247) );
  XOR2_X1 U10990 ( .A(n10248), .B(n10247), .Z(n10250) );
  OAI22_X1 U10991 ( .A1(n10250), .A2(n10651), .B1(n10249), .B2(n10740), .ZN(
        n10251) );
  AOI211_X1 U10992 ( .C1(P1_ADDR_REG_19__SCAN_IN), .C2(n10648), .A(n10252), 
        .B(n10251), .ZN(n10253) );
  OAI21_X1 U10993 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(P1_U3260) );
  AOI21_X1 U10994 ( .B1(n10258), .B2(n10257), .A(n10256), .ZN(n10974) );
  NAND2_X1 U10995 ( .A1(n10974), .A2(n10786), .ZN(n10261) );
  AOI21_X1 U10996 ( .B1(n10969), .B2(P1_REG2_REG_30__SCAN_IN), .A(n10259), 
        .ZN(n10260) );
  OAI211_X1 U10997 ( .C1(n5329), .C2(n10792), .A(n10261), .B(n10260), .ZN(
        P1_U3262) );
  XOR2_X1 U10998 ( .A(n10271), .B(n10262), .Z(n10468) );
  INV_X1 U10999 ( .A(n10279), .ZN(n10265) );
  INV_X1 U11000 ( .A(n10263), .ZN(n10264) );
  AOI21_X1 U11001 ( .B1(n10464), .B2(n10265), .A(n10264), .ZN(n10465) );
  AOI22_X1 U11002 ( .A1(n10969), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10266), 
        .B2(n10957), .ZN(n10267) );
  OAI21_X1 U11003 ( .B1(n10268), .B2(n10792), .A(n10267), .ZN(n10276) );
  AOI211_X1 U11004 ( .C1(n10271), .C2(n10270), .A(n10873), .B(n10269), .ZN(
        n10274) );
  OAI22_X1 U11005 ( .A1(n10303), .A2(n10401), .B1(n10272), .B2(n10403), .ZN(
        n10273) );
  NOR2_X1 U11006 ( .A1(n10274), .A2(n10273), .ZN(n10467) );
  NOR2_X1 U11007 ( .A1(n10467), .A2(n10969), .ZN(n10275) );
  AOI211_X1 U11008 ( .C1(n10786), .C2(n10465), .A(n10276), .B(n10275), .ZN(
        n10277) );
  OAI21_X1 U11009 ( .B1(n10468), .B2(n10406), .A(n10277), .ZN(P1_U3264) );
  XOR2_X1 U11010 ( .A(n10278), .B(n10286), .Z(n10473) );
  AOI21_X1 U11011 ( .B1(n10469), .B2(n10294), .A(n10279), .ZN(n10470) );
  INV_X1 U11012 ( .A(n10280), .ZN(n10281) );
  AOI22_X1 U11013 ( .A1(n10969), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n10281), 
        .B2(n10957), .ZN(n10282) );
  OAI21_X1 U11014 ( .B1(n10283), .B2(n10792), .A(n10282), .ZN(n10291) );
  OAI21_X1 U11015 ( .B1(n10286), .B2(n10285), .A(n10284), .ZN(n10289) );
  AOI222_X1 U11016 ( .A1(n10947), .A2(n10289), .B1(n10288), .B2(n10944), .C1(
        n10287), .C2(n10942), .ZN(n10472) );
  NOR2_X1 U11017 ( .A1(n10472), .A2(n10969), .ZN(n10290) );
  AOI211_X1 U11018 ( .C1(n10470), .C2(n10786), .A(n10291), .B(n10290), .ZN(
        n10292) );
  OAI21_X1 U11019 ( .B1(n10473), .B2(n10406), .A(n10292), .ZN(P1_U3265) );
  XOR2_X1 U11020 ( .A(n10293), .B(n10300), .Z(n10478) );
  AOI21_X1 U11021 ( .B1(n10474), .B2(n10316), .A(n5315), .ZN(n10475) );
  INV_X1 U11022 ( .A(n10295), .ZN(n10296) );
  AOI22_X1 U11023 ( .A1(n10969), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10296), 
        .B2(n10957), .ZN(n10297) );
  OAI21_X1 U11024 ( .B1(n10298), .B2(n10792), .A(n10297), .ZN(n10307) );
  AOI211_X1 U11025 ( .C1(n10301), .C2(n10300), .A(n10873), .B(n10299), .ZN(
        n10305) );
  OAI22_X1 U11026 ( .A1(n10303), .A2(n10403), .B1(n10302), .B2(n10401), .ZN(
        n10304) );
  NOR2_X1 U11027 ( .A1(n10305), .A2(n10304), .ZN(n10477) );
  NOR2_X1 U11028 ( .A1(n10477), .A2(n10969), .ZN(n10306) );
  AOI211_X1 U11029 ( .C1(n10475), .C2(n10786), .A(n10307), .B(n10306), .ZN(
        n10308) );
  OAI21_X1 U11030 ( .B1(n10478), .B2(n10406), .A(n10308), .ZN(P1_U3266) );
  XOR2_X1 U11031 ( .A(n10309), .B(n10313), .Z(n10483) );
  AOI22_X1 U11032 ( .A1(n10481), .A2(n10959), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10969), .ZN(n10322) );
  NAND2_X1 U11033 ( .A1(n10311), .A2(n10310), .ZN(n10312) );
  XOR2_X1 U11034 ( .A(n10313), .B(n10312), .Z(n10314) );
  OAI222_X1 U11035 ( .A1(n10403), .A2(n10315), .B1(n10401), .B2(n10348), .C1(
        n10314), .C2(n10873), .ZN(n10479) );
  INV_X1 U11036 ( .A(n10324), .ZN(n10317) );
  AOI211_X1 U11037 ( .C1(n10481), .C2(n10317), .A(n10927), .B(n5316), .ZN(
        n10480) );
  INV_X1 U11038 ( .A(n10480), .ZN(n10319) );
  OAI22_X1 U11039 ( .A1(n10319), .A2(n10366), .B1(n10819), .B2(n10318), .ZN(
        n10320) );
  OAI21_X1 U11040 ( .B1(n10479), .B2(n10320), .A(n10822), .ZN(n10321) );
  OAI211_X1 U11041 ( .C1(n10483), .C2(n10406), .A(n10322), .B(n10321), .ZN(
        P1_U3267) );
  XNOR2_X1 U11042 ( .A(n10323), .B(n10332), .ZN(n10488) );
  INV_X1 U11043 ( .A(n10343), .ZN(n10325) );
  AOI21_X1 U11044 ( .B1(n10484), .B2(n10325), .A(n10324), .ZN(n10485) );
  INV_X1 U11045 ( .A(n10326), .ZN(n10327) );
  AOI22_X1 U11046 ( .A1(n10969), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10327), 
        .B2(n10957), .ZN(n10328) );
  OAI21_X1 U11047 ( .B1(n10329), .B2(n10792), .A(n10328), .ZN(n10338) );
  NAND2_X1 U11048 ( .A1(n10331), .A2(n10330), .ZN(n10333) );
  XNOR2_X1 U11049 ( .A(n10333), .B(n10332), .ZN(n10336) );
  AOI222_X1 U11050 ( .A1(n10947), .A2(n10336), .B1(n10335), .B2(n10944), .C1(
        n10334), .C2(n10942), .ZN(n10487) );
  NOR2_X1 U11051 ( .A1(n10487), .A2(n10969), .ZN(n10337) );
  AOI211_X1 U11052 ( .C1(n10485), .C2(n10786), .A(n10338), .B(n10337), .ZN(
        n10339) );
  OAI21_X1 U11053 ( .B1(n10488), .B2(n10406), .A(n10339), .ZN(P1_U3268) );
  XOR2_X1 U11054 ( .A(n10340), .B(n10344), .Z(n10493) );
  INV_X1 U11055 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10342) );
  OAI22_X1 U11056 ( .A1(n10822), .A2(n10342), .B1(n10341), .B2(n10819), .ZN(
        n10351) );
  AOI211_X1 U11057 ( .C1(n10491), .C2(n10354), .A(n10927), .B(n10343), .ZN(
        n10490) );
  XOR2_X1 U11058 ( .A(n10345), .B(n10344), .Z(n10346) );
  OAI222_X1 U11059 ( .A1(n10403), .A2(n10348), .B1(n10401), .B2(n10347), .C1(
        n10346), .C2(n10873), .ZN(n10489) );
  AOI21_X1 U11060 ( .B1(n10490), .B2(n10740), .A(n10489), .ZN(n10349) );
  NOR2_X1 U11061 ( .A1(n10349), .A2(n10969), .ZN(n10350) );
  AOI211_X1 U11062 ( .C1(n10959), .C2(n10491), .A(n10351), .B(n10350), .ZN(
        n10352) );
  OAI21_X1 U11063 ( .B1(n10406), .B2(n10493), .A(n10352), .ZN(P1_U3269) );
  XNOR2_X1 U11064 ( .A(n10353), .B(n10357), .ZN(n10499) );
  AOI22_X1 U11065 ( .A1(n10496), .A2(n10959), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10969), .ZN(n10369) );
  AOI211_X1 U11066 ( .C1(n10496), .C2(n10378), .A(n10927), .B(n8783), .ZN(
        n10494) );
  INV_X1 U11067 ( .A(n10494), .ZN(n10365) );
  NAND2_X1 U11068 ( .A1(n10356), .A2(n10355), .ZN(n10358) );
  XNOR2_X1 U11069 ( .A(n10358), .B(n10357), .ZN(n10360) );
  AOI22_X1 U11070 ( .A1(n10360), .A2(n10947), .B1(n10944), .B2(n10359), .ZN(
        n10498) );
  INV_X1 U11071 ( .A(n10361), .ZN(n10363) );
  NOR2_X1 U11072 ( .A1(n10362), .A2(n10403), .ZN(n10495) );
  AOI21_X1 U11073 ( .B1(n10957), .B2(n10363), .A(n10495), .ZN(n10364) );
  OAI211_X1 U11074 ( .C1(n10366), .C2(n10365), .A(n10498), .B(n10364), .ZN(
        n10367) );
  NAND2_X1 U11075 ( .A1(n10367), .A2(n10822), .ZN(n10368) );
  OAI211_X1 U11076 ( .C1(n10499), .C2(n10406), .A(n10369), .B(n10368), .ZN(
        P1_U3270) );
  XNOR2_X1 U11077 ( .A(n10371), .B(n10370), .ZN(n10384) );
  XNOR2_X1 U11078 ( .A(n10373), .B(n10372), .ZN(n10376) );
  AOI22_X1 U11079 ( .A1(n10374), .A2(n10942), .B1(n10944), .B2(n10418), .ZN(
        n10375) );
  OAI21_X1 U11080 ( .B1(n10376), .B2(n10873), .A(n10375), .ZN(n10377) );
  AOI21_X1 U11081 ( .B1(n10384), .B2(n10876), .A(n10377), .ZN(n10503) );
  INV_X1 U11082 ( .A(n10378), .ZN(n10379) );
  AOI21_X1 U11083 ( .B1(n10500), .B2(n5314), .A(n10379), .ZN(n10501) );
  INV_X1 U11084 ( .A(n10380), .ZN(n10381) );
  AOI22_X1 U11085 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n10969), .B1(n10381), 
        .B2(n10957), .ZN(n10382) );
  OAI21_X1 U11086 ( .B1(n10383), .B2(n10792), .A(n10382), .ZN(n10387) );
  INV_X1 U11087 ( .A(n10384), .ZN(n10504) );
  NOR2_X1 U11088 ( .A1(n10504), .A2(n10385), .ZN(n10386) );
  AOI211_X1 U11089 ( .C1(n10501), .C2(n10786), .A(n10387), .B(n10386), .ZN(
        n10388) );
  OAI21_X1 U11090 ( .B1(n10969), .B2(n10503), .A(n10388), .ZN(P1_U3271) );
  XNOR2_X1 U11091 ( .A(n5376), .B(n10389), .ZN(n10510) );
  AOI21_X1 U11092 ( .B1(n10506), .B2(n10424), .A(n10390), .ZN(n10507) );
  NOR2_X1 U11093 ( .A1(n10391), .A2(n10792), .ZN(n10395) );
  OAI22_X1 U11094 ( .A1(n10822), .A2(n10393), .B1(n10392), .B2(n10819), .ZN(
        n10394) );
  AOI211_X1 U11095 ( .C1(n10507), .C2(n10786), .A(n10395), .B(n10394), .ZN(
        n10405) );
  AOI21_X1 U11096 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(n10399) );
  OAI222_X1 U11097 ( .A1(n10403), .A2(n10402), .B1(n10401), .B2(n10400), .C1(
        n10873), .C2(n10399), .ZN(n10505) );
  NAND2_X1 U11098 ( .A1(n10505), .A2(n10822), .ZN(n10404) );
  OAI211_X1 U11099 ( .C1(n10510), .C2(n10406), .A(n10405), .B(n10404), .ZN(
        P1_U3272) );
  NAND2_X1 U11100 ( .A1(n10408), .A2(n10409), .ZN(n10411) );
  AND2_X1 U11101 ( .A1(n10411), .A2(n10410), .ZN(n10413) );
  AND2_X1 U11102 ( .A1(n10415), .A2(n10414), .ZN(n10416) );
  OAI21_X1 U11103 ( .B1(n10417), .B2(n10416), .A(n10947), .ZN(n10420) );
  AOI22_X1 U11104 ( .A1(n10418), .A2(n10942), .B1(n10943), .B2(n10944), .ZN(
        n10419) );
  NAND2_X1 U11105 ( .A1(n10420), .A2(n10419), .ZN(n10421) );
  AOI21_X1 U11106 ( .B1(n5029), .B2(n10876), .A(n10421), .ZN(n10514) );
  INV_X1 U11107 ( .A(n10422), .ZN(n10440) );
  NAND2_X1 U11108 ( .A1(n10440), .A2(n10426), .ZN(n10423) );
  NAND2_X1 U11109 ( .A1(n10424), .A2(n10423), .ZN(n10511) );
  AOI22_X1 U11110 ( .A1(n10969), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10425), 
        .B2(n10957), .ZN(n10428) );
  NAND2_X1 U11111 ( .A1(n10426), .A2(n10959), .ZN(n10427) );
  OAI211_X1 U11112 ( .C1(n10511), .C2(n10429), .A(n10428), .B(n10427), .ZN(
        n10430) );
  AOI21_X1 U11113 ( .B1(n5029), .B2(n10887), .A(n10430), .ZN(n10431) );
  OAI21_X1 U11114 ( .B1(n10514), .B2(n10969), .A(n10431), .ZN(P1_U3273) );
  INV_X1 U11115 ( .A(n10432), .ZN(n10433) );
  OAI21_X1 U11116 ( .B1(n10433), .B2(n5380), .A(n10408), .ZN(n10515) );
  XNOR2_X1 U11117 ( .A(n10434), .B(n5380), .ZN(n10438) );
  AOI22_X1 U11118 ( .A1(n10944), .A2(n10436), .B1(n10435), .B2(n10942), .ZN(
        n10437) );
  OAI21_X1 U11119 ( .B1(n10438), .B2(n10873), .A(n10437), .ZN(n10439) );
  AOI21_X1 U11120 ( .B1(n10515), .B2(n10876), .A(n10439), .ZN(n10519) );
  AOI21_X1 U11121 ( .B1(n10516), .B2(n10948), .A(n10422), .ZN(n10517) );
  INV_X1 U11122 ( .A(n10516), .ZN(n10441) );
  NOR2_X1 U11123 ( .A1(n10441), .A2(n10792), .ZN(n10445) );
  INV_X1 U11124 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10443) );
  OAI22_X1 U11125 ( .A1(n10822), .A2(n10443), .B1(n10442), .B2(n10819), .ZN(
        n10444) );
  AOI211_X1 U11126 ( .C1(n10517), .C2(n10786), .A(n10445), .B(n10444), .ZN(
        n10447) );
  NAND2_X1 U11127 ( .A1(n10515), .A2(n10887), .ZN(n10446) );
  OAI211_X1 U11128 ( .C1(n10519), .C2(n10969), .A(n10447), .B(n10446), .ZN(
        P1_U3274) );
  AOI21_X1 U11129 ( .B1(n10448), .B2(n10802), .A(n10972), .ZN(n10449) );
  OAI21_X1 U11130 ( .B1(n10450), .B2(n10927), .A(n10449), .ZN(n10522) );
  MUX2_X1 U11131 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10522), .S(n10977), .Z(
        P1_U3554) );
  OAI22_X1 U11132 ( .A1(n10452), .A2(n10927), .B1(n10451), .B2(n10970), .ZN(
        n10453) );
  MUX2_X1 U11133 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10523), .S(n10977), .Z(
        P1_U3552) );
  INV_X1 U11134 ( .A(n10456), .ZN(n10463) );
  AOI22_X1 U11135 ( .A1(n10458), .A2(n10973), .B1(n10802), .B2(n10457), .ZN(
        n10459) );
  OAI21_X1 U11136 ( .B1(n10460), .B2(n10520), .A(n10459), .ZN(n10461) );
  INV_X1 U11137 ( .A(n10461), .ZN(n10462) );
  NAND2_X1 U11138 ( .A1(n10463), .A2(n10462), .ZN(n10524) );
  MUX2_X1 U11139 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10524), .S(n10977), .Z(
        P1_U3551) );
  AOI22_X1 U11140 ( .A1(n10465), .A2(n10973), .B1(n10802), .B2(n10464), .ZN(
        n10466) );
  OAI211_X1 U11141 ( .C1(n10468), .C2(n10800), .A(n10467), .B(n10466), .ZN(
        n10525) );
  MUX2_X1 U11142 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10525), .S(n10977), .Z(
        P1_U3550) );
  AOI22_X1 U11143 ( .A1(n10470), .A2(n10973), .B1(n10802), .B2(n10469), .ZN(
        n10471) );
  OAI211_X1 U11144 ( .C1(n10473), .C2(n10800), .A(n10472), .B(n10471), .ZN(
        n10526) );
  MUX2_X1 U11145 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10526), .S(n10977), .Z(
        P1_U3549) );
  AOI22_X1 U11146 ( .A1(n10475), .A2(n10973), .B1(n10802), .B2(n10474), .ZN(
        n10476) );
  OAI211_X1 U11147 ( .C1(n10478), .C2(n10800), .A(n10477), .B(n10476), .ZN(
        n10527) );
  MUX2_X1 U11148 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10527), .S(n10977), .Z(
        P1_U3548) );
  AOI211_X1 U11149 ( .C1(n10802), .C2(n10481), .A(n10480), .B(n10479), .ZN(
        n10482) );
  OAI21_X1 U11150 ( .B1(n10483), .B2(n10800), .A(n10482), .ZN(n10528) );
  MUX2_X1 U11151 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10528), .S(n10977), .Z(
        P1_U3547) );
  AOI22_X1 U11152 ( .A1(n10485), .A2(n10973), .B1(n10802), .B2(n10484), .ZN(
        n10486) );
  OAI211_X1 U11153 ( .C1(n10488), .C2(n10800), .A(n10487), .B(n10486), .ZN(
        n10529) );
  MUX2_X1 U11154 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10529), .S(n10977), .Z(
        P1_U3546) );
  AOI211_X1 U11155 ( .C1(n10802), .C2(n10491), .A(n10490), .B(n10489), .ZN(
        n10492) );
  OAI21_X1 U11156 ( .B1(n10493), .B2(n10800), .A(n10492), .ZN(n10530) );
  MUX2_X1 U11157 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10530), .S(n10977), .Z(
        P1_U3545) );
  AOI211_X1 U11158 ( .C1(n10802), .C2(n10496), .A(n10495), .B(n10494), .ZN(
        n10497) );
  OAI211_X1 U11159 ( .C1(n10499), .C2(n10800), .A(n10498), .B(n10497), .ZN(
        n10531) );
  MUX2_X1 U11160 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10531), .S(n10977), .Z(
        P1_U3544) );
  AOI22_X1 U11161 ( .A1(n10501), .A2(n10973), .B1(n10802), .B2(n10500), .ZN(
        n10502) );
  OAI211_X1 U11162 ( .C1(n10504), .C2(n10520), .A(n10503), .B(n10502), .ZN(
        n10532) );
  MUX2_X1 U11163 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10532), .S(n10977), .Z(
        P1_U3543) );
  INV_X1 U11164 ( .A(n10505), .ZN(n10509) );
  AOI22_X1 U11165 ( .A1(n10507), .A2(n10973), .B1(n10802), .B2(n10506), .ZN(
        n10508) );
  OAI211_X1 U11166 ( .C1(n10510), .C2(n10800), .A(n10509), .B(n10508), .ZN(
        n10533) );
  MUX2_X1 U11167 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10533), .S(n10977), .Z(
        P1_U3542) );
  OAI22_X1 U11168 ( .A1(n10511), .A2(n10927), .B1(n8782), .B2(n10970), .ZN(
        n10512) );
  AOI21_X1 U11169 ( .B1(n5029), .B2(n10879), .A(n10512), .ZN(n10513) );
  NAND2_X1 U11170 ( .A1(n10514), .A2(n10513), .ZN(n10534) );
  MUX2_X1 U11171 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10534), .S(n10977), .Z(
        P1_U3541) );
  INV_X1 U11172 ( .A(n10515), .ZN(n10521) );
  AOI22_X1 U11173 ( .A1(n10517), .A2(n10973), .B1(n10802), .B2(n10516), .ZN(
        n10518) );
  OAI211_X1 U11174 ( .C1(n10521), .C2(n10520), .A(n10519), .B(n10518), .ZN(
        n10535) );
  MUX2_X1 U11175 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10535), .S(n10977), .Z(
        P1_U3540) );
  MUX2_X1 U11176 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10522), .S(n10981), .Z(
        P1_U3522) );
  MUX2_X1 U11177 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10523), .S(n10981), .Z(
        P1_U3520) );
  MUX2_X1 U11178 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10524), .S(n10981), .Z(
        P1_U3519) );
  MUX2_X1 U11179 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10525), .S(n10981), .Z(
        P1_U3518) );
  MUX2_X1 U11180 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10526), .S(n10981), .Z(
        P1_U3517) );
  MUX2_X1 U11181 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10527), .S(n10981), .Z(
        P1_U3516) );
  MUX2_X1 U11182 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10528), .S(n10981), .Z(
        P1_U3515) );
  MUX2_X1 U11183 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10529), .S(n10981), .Z(
        P1_U3514) );
  MUX2_X1 U11184 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10530), .S(n10981), .Z(
        P1_U3513) );
  MUX2_X1 U11185 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10531), .S(n10981), .Z(
        P1_U3512) );
  MUX2_X1 U11186 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10532), .S(n10981), .Z(
        P1_U3511) );
  MUX2_X1 U11187 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10533), .S(n10981), .Z(
        P1_U3510) );
  MUX2_X1 U11188 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10534), .S(n10981), .Z(
        P1_U3508) );
  MUX2_X1 U11189 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10535), .S(n10981), .Z(
        P1_U3505) );
  MUX2_X1 U11190 ( .A(n10536), .B(P1_D_REG_0__SCAN_IN), .S(n10549), .Z(
        P1_U3440) );
  INV_X1 U11191 ( .A(n10537), .ZN(n10542) );
  NOR4_X1 U11192 ( .A1(n5590), .A2(P1_IR_REG_30__SCAN_IN), .A3(n6806), .A4(
        P1_U3084), .ZN(n10538) );
  AOI21_X1 U11193 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10539), .A(n10538), 
        .ZN(n10540) );
  OAI21_X1 U11194 ( .B1(n10542), .B2(n10541), .A(n10540), .ZN(P1_U3322) );
  INV_X1 U11195 ( .A(n10543), .ZN(n10544) );
  MUX2_X1 U11196 ( .A(n10544), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11197 ( .A(n10549), .ZN(n10548) );
  NOR2_X1 U11198 ( .A1(n10548), .A2(n10545), .ZN(P1_U3321) );
  NOR2_X1 U11199 ( .A1(n10548), .A2(n10546), .ZN(P1_U3320) );
  NOR2_X1 U11200 ( .A1(n10548), .A2(n10547), .ZN(P1_U3319) );
  AND2_X1 U11201 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10549), .ZN(P1_U3318) );
  AND2_X1 U11202 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10549), .ZN(P1_U3317) );
  AND2_X1 U11203 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10549), .ZN(P1_U3316) );
  AND2_X1 U11204 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10549), .ZN(P1_U3315) );
  AND2_X1 U11205 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10549), .ZN(P1_U3314) );
  AND2_X1 U11206 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10549), .ZN(P1_U3313) );
  AND2_X1 U11207 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10549), .ZN(P1_U3312) );
  AND2_X1 U11208 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10549), .ZN(P1_U3311) );
  AND2_X1 U11209 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10549), .ZN(P1_U3310) );
  AND2_X1 U11210 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10549), .ZN(P1_U3309) );
  AND2_X1 U11211 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10549), .ZN(P1_U3308) );
  AND2_X1 U11212 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10549), .ZN(P1_U3307) );
  AND2_X1 U11213 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10549), .ZN(P1_U3306) );
  AND2_X1 U11214 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10549), .ZN(P1_U3305) );
  AND2_X1 U11215 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10549), .ZN(P1_U3304) );
  AND2_X1 U11216 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10549), .ZN(P1_U3303) );
  AND2_X1 U11217 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10549), .ZN(P1_U3302) );
  AND2_X1 U11218 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10549), .ZN(P1_U3301) );
  AND2_X1 U11219 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10549), .ZN(P1_U3300) );
  AND2_X1 U11220 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10549), .ZN(P1_U3299) );
  AND2_X1 U11221 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10549), .ZN(P1_U3298) );
  AND2_X1 U11222 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10549), .ZN(P1_U3297) );
  AND2_X1 U11223 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10549), .ZN(P1_U3296) );
  AND2_X1 U11224 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10549), .ZN(P1_U3295) );
  AND2_X1 U11225 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10549), .ZN(P1_U3294) );
  AND2_X1 U11226 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10549), .ZN(P1_U3293) );
  AND2_X1 U11227 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10549), .ZN(P1_U3292) );
  INV_X1 U11228 ( .A(n10550), .ZN(n10551) );
  AOI22_X1 U11229 ( .A1(n10554), .A2(n10663), .B1(n10553), .B2(n10661), .ZN(
        P2_U3438) );
  AND2_X1 U11230 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10661), .ZN(P2_U3326) );
  AND2_X1 U11231 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10661), .ZN(P2_U3325) );
  AND2_X1 U11232 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10661), .ZN(P2_U3324) );
  AND2_X1 U11233 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10661), .ZN(P2_U3323) );
  AND2_X1 U11234 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10661), .ZN(P2_U3322) );
  AND2_X1 U11235 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10661), .ZN(P2_U3321) );
  AND2_X1 U11236 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10661), .ZN(P2_U3320) );
  AND2_X1 U11237 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10661), .ZN(P2_U3319) );
  AND2_X1 U11238 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10661), .ZN(P2_U3318) );
  AND2_X1 U11239 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10661), .ZN(P2_U3317) );
  AND2_X1 U11240 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10661), .ZN(P2_U3316) );
  AND2_X1 U11241 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10661), .ZN(P2_U3315) );
  AND2_X1 U11242 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10661), .ZN(P2_U3314) );
  AND2_X1 U11243 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10661), .ZN(P2_U3313) );
  AND2_X1 U11244 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10661), .ZN(P2_U3312) );
  AND2_X1 U11245 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10661), .ZN(P2_U3311) );
  AND2_X1 U11246 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10661), .ZN(P2_U3310) );
  AND2_X1 U11247 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10661), .ZN(P2_U3309) );
  AND2_X1 U11248 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10661), .ZN(P2_U3308) );
  AND2_X1 U11249 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10661), .ZN(P2_U3307) );
  AND2_X1 U11250 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10661), .ZN(P2_U3306) );
  AND2_X1 U11251 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10661), .ZN(P2_U3305) );
  AND2_X1 U11252 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10661), .ZN(P2_U3304) );
  AND2_X1 U11253 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10661), .ZN(P2_U3303) );
  AND2_X1 U11254 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10661), .ZN(P2_U3302) );
  AND2_X1 U11255 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10661), .ZN(P2_U3301) );
  AND2_X1 U11256 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10661), .ZN(P2_U3300) );
  AND2_X1 U11257 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10661), .ZN(P2_U3299) );
  AND2_X1 U11258 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10661), .ZN(P2_U3298) );
  AND2_X1 U11259 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10661), .ZN(P2_U3297) );
  XOR2_X1 U11260 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  NAND3_X1 U11261 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10557) );
  AOI21_X1 U11262 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10559) );
  INV_X1 U11263 ( .A(n10559), .ZN(n10555) );
  NAND2_X1 U11264 ( .A1(n10557), .A2(n10555), .ZN(n10556) );
  XNOR2_X1 U11265 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10556), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11266 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10561) );
  INV_X1 U11267 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10558) );
  OAI21_X1 U11268 ( .B1(n10559), .B2(n10558), .A(n10557), .ZN(n10560) );
  XOR2_X1 U11269 ( .A(n10561), .B(n10560), .Z(ADD_1071_U54) );
  XOR2_X1 U11270 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10565) );
  NAND2_X1 U11271 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10563) );
  NAND2_X1 U11272 ( .A1(n10561), .A2(n10560), .ZN(n10562) );
  NAND2_X1 U11273 ( .A1(n10563), .A2(n10562), .ZN(n10564) );
  XOR2_X1 U11274 ( .A(n10565), .B(n10564), .Z(ADD_1071_U53) );
  XNOR2_X1 U11275 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10569) );
  NAND2_X1 U11276 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10567) );
  NAND2_X1 U11277 ( .A1(n10565), .A2(n10564), .ZN(n10566) );
  NAND2_X1 U11278 ( .A1(n10567), .A2(n10566), .ZN(n10568) );
  XNOR2_X1 U11279 ( .A(n10569), .B(n10568), .ZN(ADD_1071_U52) );
  NOR2_X1 U11280 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10571) );
  NOR2_X1 U11281 ( .A1(n10569), .A2(n10568), .ZN(n10570) );
  NOR2_X1 U11282 ( .A1(n10571), .A2(n10570), .ZN(n10572) );
  AND2_X1 U11283 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10572), .ZN(n10574) );
  NOR2_X1 U11284 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10572), .ZN(n10576) );
  NOR2_X1 U11285 ( .A1(n10574), .A2(n10576), .ZN(n10573) );
  XOR2_X1 U11286 ( .A(n10573), .B(P2_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  NOR2_X1 U11287 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10574), .ZN(n10575) );
  XOR2_X1 U11288 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10577), .Z(n10578) );
  XOR2_X1 U11289 ( .A(n10578), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NAND2_X1 U11290 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10577), .ZN(n10580) );
  NAND2_X1 U11291 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10578), .ZN(n10579) );
  NAND2_X1 U11292 ( .A1(n10580), .A2(n10579), .ZN(n10582) );
  XOR2_X1 U11293 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10582), .Z(n10583) );
  XNOR2_X1 U11294 ( .A(n10583), .B(n10581), .ZN(ADD_1071_U49) );
  NAND2_X1 U11295 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10582), .ZN(n10585) );
  NAND2_X1 U11296 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10583), .ZN(n10584) );
  NAND2_X1 U11297 ( .A1(n10585), .A2(n10584), .ZN(n10587) );
  XOR2_X1 U11298 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10587), .Z(n10588) );
  XNOR2_X1 U11299 ( .A(n10588), .B(n10586), .ZN(ADD_1071_U48) );
  NAND2_X1 U11300 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10587), .ZN(n10590) );
  NAND2_X1 U11301 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10588), .ZN(n10589) );
  NAND2_X1 U11302 ( .A1(n10590), .A2(n10589), .ZN(n10591) );
  XOR2_X1 U11303 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n10591), .Z(n10592) );
  XOR2_X1 U11304 ( .A(n10592), .B(P2_ADDR_REG_9__SCAN_IN), .Z(ADD_1071_U47) );
  XOR2_X1 U11305 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10596) );
  NAND2_X1 U11306 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n10591), .ZN(n10594) );
  NAND2_X1 U11307 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10592), .ZN(n10593) );
  NAND2_X1 U11308 ( .A1(n10594), .A2(n10593), .ZN(n10595) );
  XOR2_X1 U11309 ( .A(n10596), .B(n10595), .Z(ADD_1071_U63) );
  XOR2_X1 U11310 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10600) );
  NAND2_X1 U11311 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10598) );
  NAND2_X1 U11312 ( .A1(n10596), .A2(n10595), .ZN(n10597) );
  NAND2_X1 U11313 ( .A1(n10598), .A2(n10597), .ZN(n10599) );
  XOR2_X1 U11314 ( .A(n10600), .B(n10599), .Z(ADD_1071_U62) );
  NAND2_X1 U11315 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10602) );
  NAND2_X1 U11316 ( .A1(n10600), .A2(n10599), .ZN(n10601) );
  NAND2_X1 U11317 ( .A1(n10602), .A2(n10601), .ZN(n10604) );
  XNOR2_X1 U11318 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10603) );
  XNOR2_X1 U11319 ( .A(n10604), .B(n10603), .ZN(ADD_1071_U61) );
  NOR2_X1 U11320 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10606) );
  XNOR2_X1 U11321 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10607) );
  XNOR2_X1 U11322 ( .A(n10608), .B(n10607), .ZN(ADD_1071_U60) );
  NOR2_X1 U11323 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10610) );
  XNOR2_X1 U11324 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10611) );
  XNOR2_X1 U11325 ( .A(n10612), .B(n10611), .ZN(ADD_1071_U59) );
  NOR2_X1 U11326 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10614) );
  NOR2_X1 U11327 ( .A1(n10612), .A2(n10611), .ZN(n10613) );
  NOR2_X1 U11328 ( .A1(n10614), .A2(n10613), .ZN(n10616) );
  XNOR2_X1 U11329 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10615) );
  XNOR2_X1 U11330 ( .A(n10616), .B(n10615), .ZN(ADD_1071_U58) );
  NOR2_X1 U11331 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10618) );
  NOR2_X1 U11332 ( .A1(n10616), .A2(n10615), .ZN(n10617) );
  NOR2_X1 U11333 ( .A1(n10618), .A2(n10617), .ZN(n10620) );
  XNOR2_X1 U11334 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10619) );
  XNOR2_X1 U11335 ( .A(n10620), .B(n10619), .ZN(ADD_1071_U57) );
  NOR2_X1 U11336 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10622) );
  NOR2_X1 U11337 ( .A1(n10620), .A2(n10619), .ZN(n10621) );
  NOR2_X1 U11338 ( .A1(n10622), .A2(n10621), .ZN(n10624) );
  XNOR2_X1 U11339 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10623) );
  XNOR2_X1 U11340 ( .A(n10624), .B(n10623), .ZN(ADD_1071_U56) );
  NOR2_X1 U11341 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10626) );
  NOR2_X1 U11342 ( .A1(n10624), .A2(n10623), .ZN(n10625) );
  NOR2_X1 U11343 ( .A1(n10626), .A2(n10625), .ZN(n10627) );
  NOR2_X1 U11344 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10627), .ZN(n10630) );
  AND2_X1 U11345 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10627), .ZN(n10629) );
  NOR2_X1 U11346 ( .A1(n10630), .A2(n10629), .ZN(n10628) );
  XOR2_X1 U11347 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10628), .Z(ADD_1071_U55)
         );
  NOR2_X1 U11348 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10629), .ZN(n10631) );
  NOR2_X1 U11349 ( .A1(n10631), .A2(n10630), .ZN(n10633) );
  XNOR2_X1 U11350 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n10632) );
  XNOR2_X1 U11351 ( .A(n10633), .B(n10632), .ZN(ADD_1071_U4) );
  INV_X1 U11352 ( .A(n10634), .ZN(n10636) );
  INV_X1 U11353 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10635) );
  NAND2_X1 U11354 ( .A1(n7155), .A2(n10635), .ZN(n10638) );
  NAND2_X1 U11355 ( .A1(n10636), .A2(n10638), .ZN(n10639) );
  MUX2_X1 U11356 ( .A(n10639), .B(n10638), .S(n10637), .Z(n10641) );
  NAND2_X1 U11357 ( .A1(n10641), .A2(n10640), .ZN(n10643) );
  AOI22_X1 U11358 ( .A1(n10648), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10642) );
  OAI21_X1 U11359 ( .B1(n10644), .B2(n10643), .A(n10642), .ZN(P1_U3241) );
  OAI21_X1 U11360 ( .B1(n10647), .B2(n10646), .A(n10645), .ZN(n10650) );
  AOI22_X1 U11361 ( .A1(n10650), .A2(n10649), .B1(n10648), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n10660) );
  AOI211_X1 U11362 ( .C1(n10654), .C2(n10653), .A(n10652), .B(n10651), .ZN(
        n10655) );
  AOI211_X1 U11363 ( .C1(n10658), .C2(n10657), .A(n10656), .B(n10655), .ZN(
        n10659) );
  NAND2_X1 U11364 ( .A1(n10660), .A2(n10659), .ZN(P1_U3259) );
  AOI22_X1 U11365 ( .A1(n10664), .A2(n10663), .B1(n10662), .B2(n10661), .ZN(
        P2_U3437) );
  AOI22_X1 U11366 ( .A1(n10665), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10684), .ZN(n10672) );
  INV_X1 U11367 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10666) );
  NAND2_X1 U11368 ( .A1(n10684), .A2(n10666), .ZN(n10667) );
  OAI211_X1 U11369 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n10689), .A(n10668), .B(
        n10667), .ZN(n10669) );
  INV_X1 U11370 ( .A(n10669), .ZN(n10671) );
  AOI22_X1 U11371 ( .A1(n10674), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10670) );
  OAI221_X1 U11372 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10672), .C1(n5271), .C2(
        n10671), .A(n10670), .ZN(P2_U3245) );
  AOI22_X1 U11373 ( .A1(n10674), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10693) );
  NAND2_X1 U11374 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  NAND2_X1 U11375 ( .A1(n10678), .A2(n10677), .ZN(n10690) );
  NAND2_X1 U11376 ( .A1(n10680), .A2(n10679), .ZN(n10688) );
  INV_X1 U11377 ( .A(n10681), .ZN(n10686) );
  INV_X1 U11378 ( .A(n10682), .ZN(n10685) );
  OAI211_X1 U11379 ( .C1(n10686), .C2(n10685), .A(n10684), .B(n10683), .ZN(
        n10687) );
  OAI211_X1 U11380 ( .C1(n10690), .C2(n10689), .A(n10688), .B(n10687), .ZN(
        n10691) );
  INV_X1 U11381 ( .A(n10691), .ZN(n10692) );
  NAND2_X1 U11382 ( .A1(n10693), .A2(n10692), .ZN(P2_U3247) );
  XNOR2_X1 U11383 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11384 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10700) );
  OAI21_X1 U11385 ( .B1(n10959), .B2(n10786), .A(n10694), .ZN(n10695) );
  OAI21_X1 U11386 ( .B1(n10822), .B2(n10696), .A(n10695), .ZN(n10697) );
  AOI21_X1 U11387 ( .B1(n10698), .B2(n10822), .A(n10697), .ZN(n10699) );
  OAI21_X1 U11388 ( .B1(n10819), .B2(n10700), .A(n10699), .ZN(P1_U3291) );
  AOI22_X1 U11389 ( .A1(n10703), .A2(n10921), .B1(n10702), .B2(n10701), .ZN(
        n10704) );
  AND2_X1 U11390 ( .A1(n10705), .A2(n10704), .ZN(n10707) );
  AOI22_X1 U11391 ( .A1(n10923), .A2(n10707), .B1(n10666), .B2(n10922), .ZN(
        P2_U3520) );
  INV_X1 U11392 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U11393 ( .A1(n5011), .A2(n10707), .B1(n10706), .B2(n10985), .ZN(
        P2_U3451) );
  OAI22_X1 U11394 ( .A1(n10709), .A2(n10927), .B1(n10708), .B2(n10970), .ZN(
        n10711) );
  AOI211_X1 U11395 ( .C1(n10879), .C2(n10712), .A(n10711), .B(n10710), .ZN(
        n10715) );
  INV_X1 U11396 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U11397 ( .A1(n10977), .A2(n10715), .B1(n10713), .B2(n10975), .ZN(
        P1_U3525) );
  INV_X1 U11398 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U11399 ( .A1(n10981), .A2(n10715), .B1(n10714), .B2(n10978), .ZN(
        P1_U3460) );
  OAI22_X1 U11400 ( .A1(n10717), .A2(n10916), .B1(n10716), .B2(n10914), .ZN(
        n10719) );
  AOI211_X1 U11401 ( .C1(n10836), .C2(n10720), .A(n10719), .B(n10718), .ZN(
        n10723) );
  INV_X1 U11402 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U11403 ( .A1(n10923), .A2(n10723), .B1(n10721), .B2(n10922), .ZN(
        P2_U3522) );
  INV_X1 U11404 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U11405 ( .A1(n5011), .A2(n10723), .B1(n10722), .B2(n10985), .ZN(
        P2_U3457) );
  OAI22_X1 U11406 ( .A1(n10725), .A2(n10927), .B1(n10724), .B2(n10970), .ZN(
        n10727) );
  AOI211_X1 U11407 ( .C1(n10879), .C2(n10728), .A(n10727), .B(n10726), .ZN(
        n10730) );
  AOI22_X1 U11408 ( .A1(n10977), .A2(n10730), .B1(n7147), .B2(n10975), .ZN(
        P1_U3527) );
  INV_X1 U11409 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U11410 ( .A1(n10981), .A2(n10730), .B1(n10729), .B2(n10978), .ZN(
        P1_U3466) );
  OAI22_X1 U11411 ( .A1(n10732), .A2(n10916), .B1(n10731), .B2(n10914), .ZN(
        n10734) );
  AOI211_X1 U11412 ( .C1(n10735), .C2(n10921), .A(n10734), .B(n10733), .ZN(
        n10736) );
  AOI22_X1 U11413 ( .A1(n10923), .A2(n10736), .B1(n6038), .B2(n10922), .ZN(
        P2_U3524) );
  AOI22_X1 U11414 ( .A1(n5011), .A2(n10736), .B1(n6035), .B2(n10985), .ZN(
        P2_U3463) );
  INV_X1 U11415 ( .A(n10737), .ZN(n10738) );
  NOR2_X1 U11416 ( .A1(n10739), .A2(n10738), .ZN(n10748) );
  NAND2_X1 U11417 ( .A1(n10741), .A2(n10740), .ZN(n10746) );
  AOI22_X1 U11418 ( .A1(n10744), .A2(n10743), .B1(n10957), .B2(n10742), .ZN(
        n10745) );
  NAND2_X1 U11419 ( .A1(n10746), .A2(n10745), .ZN(n10747) );
  NOR3_X1 U11420 ( .A1(n10749), .A2(n10748), .A3(n10747), .ZN(n10750) );
  AOI22_X1 U11421 ( .A1(n10969), .A2(n7173), .B1(n10750), .B2(n10822), .ZN(
        P1_U3286) );
  INV_X1 U11422 ( .A(n10751), .ZN(n10757) );
  INV_X1 U11423 ( .A(n10752), .ZN(n10754) );
  AOI22_X1 U11424 ( .A1(n10755), .A2(n10754), .B1(n5600), .B2(n10753), .ZN(
        n10756) );
  OAI21_X1 U11425 ( .B1(n10757), .B2(n6002), .A(n10756), .ZN(n10758) );
  AOI211_X1 U11426 ( .C1(n10848), .C2(n10760), .A(n10759), .B(n10758), .ZN(
        n10761) );
  AOI22_X1 U11427 ( .A1(n10851), .A2(n7525), .B1(n10761), .B2(n10856), .ZN(
        P2_U3291) );
  INV_X1 U11428 ( .A(n10762), .ZN(n10766) );
  OAI22_X1 U11429 ( .A1(n10763), .A2(n10927), .B1(n5305), .B2(n10970), .ZN(
        n10765) );
  AOI211_X1 U11430 ( .C1(n10879), .C2(n10766), .A(n10765), .B(n10764), .ZN(
        n10767) );
  AOI22_X1 U11431 ( .A1(n10977), .A2(n10767), .B1(n6676), .B2(n10975), .ZN(
        P1_U3529) );
  AOI22_X1 U11432 ( .A1(n10981), .A2(n10767), .B1(n6679), .B2(n10978), .ZN(
        P1_U3472) );
  OAI22_X1 U11433 ( .A1(n10769), .A2(n10916), .B1(n10768), .B2(n10914), .ZN(
        n10771) );
  AOI211_X1 U11434 ( .C1(n10772), .C2(n10921), .A(n10771), .B(n10770), .ZN(
        n10774) );
  AOI22_X1 U11435 ( .A1(n10923), .A2(n10774), .B1(n6057), .B2(n10922), .ZN(
        P2_U3526) );
  INV_X1 U11436 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U11437 ( .A1(n5011), .A2(n10774), .B1(n10773), .B2(n10985), .ZN(
        P2_U3469) );
  INV_X1 U11438 ( .A(n10775), .ZN(n10780) );
  OAI22_X1 U11439 ( .A1(n10777), .A2(n10927), .B1(n10776), .B2(n10970), .ZN(
        n10779) );
  AOI211_X1 U11440 ( .C1(n10780), .C2(n10952), .A(n10779), .B(n10778), .ZN(
        n10782) );
  AOI22_X1 U11441 ( .A1(n10977), .A2(n10782), .B1(n6731), .B2(n10975), .ZN(
        P1_U3531) );
  INV_X1 U11442 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10781) );
  AOI22_X1 U11443 ( .A1(n10981), .A2(n10782), .B1(n10781), .B2(n10978), .ZN(
        P1_U3478) );
  INV_X1 U11444 ( .A(n10783), .ZN(n10795) );
  INV_X1 U11445 ( .A(n10784), .ZN(n10785) );
  AOI21_X1 U11446 ( .B1(n10876), .B2(n10795), .A(n10785), .ZN(n10797) );
  NAND2_X1 U11447 ( .A1(n10787), .A2(n10786), .ZN(n10791) );
  INV_X1 U11448 ( .A(n10788), .ZN(n10789) );
  AOI22_X1 U11449 ( .A1(n10969), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n10789), 
        .B2(n10957), .ZN(n10790) );
  OAI211_X1 U11450 ( .C1(n10793), .C2(n10792), .A(n10791), .B(n10790), .ZN(
        n10794) );
  AOI21_X1 U11451 ( .B1(n10795), .B2(n10887), .A(n10794), .ZN(n10796) );
  OAI21_X1 U11452 ( .B1(n10969), .B2(n10797), .A(n10796), .ZN(P1_U3282) );
  XNOR2_X1 U11453 ( .A(n10799), .B(n10798), .ZN(n10824) );
  INV_X1 U11454 ( .A(n10824), .ZN(n10801) );
  NOR2_X1 U11455 ( .A1(n10801), .A2(n10800), .ZN(n10815) );
  AND2_X1 U11456 ( .A1(n10828), .A2(n10802), .ZN(n10814) );
  NAND2_X1 U11457 ( .A1(n10803), .A2(n10828), .ZN(n10804) );
  NAND2_X1 U11458 ( .A1(n10804), .A2(n10973), .ZN(n10805) );
  NOR2_X1 U11459 ( .A1(n10806), .A2(n10805), .ZN(n10818) );
  OAI21_X1 U11460 ( .B1(n10809), .B2(n10807), .A(n10808), .ZN(n10810) );
  NAND2_X1 U11461 ( .A1(n10810), .A2(n10947), .ZN(n10813) );
  AOI22_X1 U11462 ( .A1(n10942), .A2(n10871), .B1(n10811), .B2(n10944), .ZN(
        n10812) );
  NAND2_X1 U11463 ( .A1(n10813), .A2(n10812), .ZN(n10823) );
  NOR4_X1 U11464 ( .A1(n10815), .A2(n10814), .A3(n10818), .A4(n10823), .ZN(
        n10817) );
  AOI22_X1 U11465 ( .A1(n10977), .A2(n10817), .B1(n7208), .B2(n10975), .ZN(
        P1_U3533) );
  INV_X1 U11466 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U11467 ( .A1(n10981), .A2(n10817), .B1(n10816), .B2(n10978), .ZN(
        P1_U3484) );
  AOI22_X1 U11468 ( .A1(n10824), .A2(n10887), .B1(n10962), .B2(n10818), .ZN(
        n10830) );
  INV_X1 U11469 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10821) );
  OAI22_X1 U11470 ( .A1(n10822), .A2(n10821), .B1(n10820), .B2(n10819), .ZN(
        n10827) );
  AOI21_X1 U11471 ( .B1(n10824), .B2(n10876), .A(n10823), .ZN(n10825) );
  NOR2_X1 U11472 ( .A1(n10825), .A2(n10969), .ZN(n10826) );
  AOI211_X1 U11473 ( .C1(n10959), .C2(n10828), .A(n10827), .B(n10826), .ZN(
        n10829) );
  NAND2_X1 U11474 ( .A1(n10830), .A2(n10829), .ZN(P1_U3281) );
  INV_X1 U11475 ( .A(n10831), .ZN(n10835) );
  OAI22_X1 U11476 ( .A1(n10832), .A2(n10916), .B1(n5352), .B2(n10914), .ZN(
        n10834) );
  AOI211_X1 U11477 ( .C1(n10836), .C2(n10835), .A(n10834), .B(n10833), .ZN(
        n10838) );
  AOI22_X1 U11478 ( .A1(n10923), .A2(n10838), .B1(n7510), .B2(n10922), .ZN(
        P2_U3530) );
  INV_X1 U11479 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U11480 ( .A1(n5011), .A2(n10838), .B1(n10837), .B2(n10985), .ZN(
        P2_U3481) );
  OAI22_X1 U11481 ( .A1(n10841), .A2(n10927), .B1(n10840), .B2(n10970), .ZN(
        n10842) );
  AOI21_X1 U11482 ( .B1(n10843), .B2(n10879), .A(n10842), .ZN(n10844) );
  AND2_X1 U11483 ( .A1(n10845), .A2(n10844), .ZN(n10847) );
  AOI22_X1 U11484 ( .A1(n10977), .A2(n10847), .B1(n7207), .B2(n10975), .ZN(
        P1_U3534) );
  INV_X1 U11485 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U11486 ( .A1(n10981), .A2(n10847), .B1(n10846), .B2(n10978), .ZN(
        P1_U3487) );
  AND2_X1 U11487 ( .A1(n10849), .A2(n10848), .ZN(n10858) );
  AOI211_X1 U11488 ( .C1(n10852), .C2(n5600), .A(n10851), .B(n10850), .ZN(
        n10853) );
  OAI211_X1 U11489 ( .C1(n6002), .C2(n10855), .A(n10854), .B(n10853), .ZN(
        n10857) );
  OAI22_X1 U11490 ( .A1(n10858), .A2(n10857), .B1(P2_REG2_REG_11__SCAN_IN), 
        .B2(n10856), .ZN(n10859) );
  OAI21_X1 U11491 ( .B1(n10861), .B2(n10860), .A(n10859), .ZN(P2_U3285) );
  INV_X1 U11492 ( .A(n10863), .ZN(n10864) );
  AOI21_X1 U11493 ( .B1(n10868), .B2(n10862), .A(n10864), .ZN(n10888) );
  OAI211_X1 U11494 ( .C1(n10866), .C2(n10867), .A(n10973), .B(n10865), .ZN(
        n10885) );
  OAI21_X1 U11495 ( .B1(n10867), .B2(n10970), .A(n10885), .ZN(n10878) );
  XNOR2_X1 U11496 ( .A(n10869), .B(n10868), .ZN(n10874) );
  AOI22_X1 U11497 ( .A1(n10944), .A2(n10871), .B1(n10870), .B2(n10942), .ZN(
        n10872) );
  OAI21_X1 U11498 ( .B1(n10874), .B2(n10873), .A(n10872), .ZN(n10875) );
  AOI21_X1 U11499 ( .B1(n10888), .B2(n10876), .A(n10875), .ZN(n10891) );
  INV_X1 U11500 ( .A(n10891), .ZN(n10877) );
  AOI211_X1 U11501 ( .C1(n10879), .C2(n10888), .A(n10878), .B(n10877), .ZN(
        n10881) );
  AOI22_X1 U11502 ( .A1(n10977), .A2(n10881), .B1(n7206), .B2(n10975), .ZN(
        P1_U3535) );
  INV_X1 U11503 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U11504 ( .A1(n10981), .A2(n10881), .B1(n10880), .B2(n10978), .ZN(
        P1_U3490) );
  INV_X1 U11505 ( .A(n10882), .ZN(n10883) );
  AOI222_X1 U11506 ( .A1(n10884), .A2(n10959), .B1(n10883), .B2(n10957), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(n10969), .ZN(n10890) );
  INV_X1 U11507 ( .A(n10885), .ZN(n10886) );
  AOI22_X1 U11508 ( .A1(n10888), .A2(n10887), .B1(n10962), .B2(n10886), .ZN(
        n10889) );
  OAI211_X1 U11509 ( .C1(n10969), .C2(n10891), .A(n10890), .B(n10889), .ZN(
        P1_U3279) );
  OAI22_X1 U11510 ( .A1(n10893), .A2(n10916), .B1(n10892), .B2(n10914), .ZN(
        n10895) );
  AOI211_X1 U11511 ( .C1(n10896), .C2(n10921), .A(n10895), .B(n10894), .ZN(
        n10898) );
  AOI22_X1 U11512 ( .A1(n10923), .A2(n10898), .B1(n7615), .B2(n10922), .ZN(
        P2_U3532) );
  INV_X1 U11513 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U11514 ( .A1(n5011), .A2(n10898), .B1(n10897), .B2(n10985), .ZN(
        P2_U3487) );
  OAI22_X1 U11515 ( .A1(n10900), .A2(n10927), .B1(n10899), .B2(n10970), .ZN(
        n10903) );
  INV_X1 U11516 ( .A(n10901), .ZN(n10902) );
  AOI211_X1 U11517 ( .C1(n10952), .C2(n10904), .A(n10903), .B(n10902), .ZN(
        n10906) );
  AOI22_X1 U11518 ( .A1(n10977), .A2(n10906), .B1(n7205), .B2(n10975), .ZN(
        P1_U3536) );
  INV_X1 U11519 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U11520 ( .A1(n10981), .A2(n10906), .B1(n10905), .B2(n10978), .ZN(
        P1_U3493) );
  OAI211_X1 U11521 ( .C1(n10909), .C2(n10970), .A(n10908), .B(n10907), .ZN(
        n10910) );
  AOI21_X1 U11522 ( .B1(n10952), .B2(n10911), .A(n10910), .ZN(n10913) );
  AOI22_X1 U11523 ( .A1(n10977), .A2(n10913), .B1(n6849), .B2(n10975), .ZN(
        P1_U3537) );
  INV_X1 U11524 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U11525 ( .A1(n10981), .A2(n10913), .B1(n10912), .B2(n10978), .ZN(
        P1_U3496) );
  OAI22_X1 U11526 ( .A1(n10917), .A2(n10916), .B1(n10915), .B2(n10914), .ZN(
        n10919) );
  AOI211_X1 U11527 ( .C1(n10921), .C2(n10920), .A(n10919), .B(n10918), .ZN(
        n10925) );
  AOI22_X1 U11528 ( .A1(n10923), .A2(n10925), .B1(n7714), .B2(n10922), .ZN(
        P2_U3534) );
  INV_X1 U11529 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U11530 ( .A1(n5011), .A2(n10925), .B1(n10924), .B2(n10985), .ZN(
        P2_U3493) );
  OAI22_X1 U11531 ( .A1(n10928), .A2(n10927), .B1(n10926), .B2(n10970), .ZN(
        n10930) );
  AOI211_X1 U11532 ( .C1(n10931), .C2(n10952), .A(n10930), .B(n10929), .ZN(
        n10934) );
  AOI22_X1 U11533 ( .A1(n10977), .A2(n10934), .B1(n10932), .B2(n10975), .ZN(
        P1_U3538) );
  INV_X1 U11534 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U11535 ( .A1(n10981), .A2(n10934), .B1(n10933), .B2(n10978), .ZN(
        P1_U3499) );
  OAI21_X1 U11536 ( .B1(n10937), .B2(n10936), .A(n10935), .ZN(n10938) );
  INV_X1 U11537 ( .A(n10938), .ZN(n10965) );
  OAI21_X1 U11538 ( .B1(n10941), .B2(n10940), .A(n10939), .ZN(n10946) );
  AOI222_X1 U11539 ( .A1(n10947), .A2(n10946), .B1(n10945), .B2(n10944), .C1(
        n10943), .C2(n10942), .ZN(n10968) );
  OAI211_X1 U11540 ( .C1(n10949), .C2(n10950), .A(n10973), .B(n10948), .ZN(
        n10961) );
  OAI211_X1 U11541 ( .C1(n10950), .C2(n10970), .A(n10968), .B(n10961), .ZN(
        n10951) );
  AOI21_X1 U11542 ( .B1(n10965), .B2(n10952), .A(n10951), .ZN(n10955) );
  AOI22_X1 U11543 ( .A1(n10977), .A2(n10955), .B1(n10953), .B2(n10975), .ZN(
        P1_U3539) );
  INV_X1 U11544 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U11545 ( .A1(n10981), .A2(n10955), .B1(n10954), .B2(n10978), .ZN(
        P1_U3502) );
  INV_X1 U11546 ( .A(n10956), .ZN(n10958) );
  AOI222_X1 U11547 ( .A1(n10960), .A2(n10959), .B1(n10958), .B2(n10957), .C1(
        P1_REG2_REG_16__SCAN_IN), .C2(n10969), .ZN(n10967) );
  INV_X1 U11548 ( .A(n10961), .ZN(n10963) );
  AOI22_X1 U11549 ( .A1(n10965), .A2(n10964), .B1(n10963), .B2(n10962), .ZN(
        n10966) );
  OAI211_X1 U11550 ( .C1(n10969), .C2(n10968), .A(n10967), .B(n10966), .ZN(
        P1_U3275) );
  NOR2_X1 U11551 ( .A1(n5329), .A2(n10970), .ZN(n10971) );
  AOI211_X1 U11552 ( .C1(n10974), .C2(n10973), .A(n10972), .B(n10971), .ZN(
        n10980) );
  INV_X1 U11553 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U11554 ( .A1(n10977), .A2(n10980), .B1(n10976), .B2(n10975), .ZN(
        P1_U3553) );
  INV_X1 U11555 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U11556 ( .A1(n10981), .A2(n10980), .B1(n10979), .B2(n10978), .ZN(
        P1_U3521) );
  XNOR2_X1 U11557 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X2 U5078 ( .A(n6754), .Z(n7809) );
  CLKBUF_X2 U5084 ( .A(n6708), .Z(n7030) );
  NAND2_X1 U5087 ( .A1(n10373), .A2(n10372), .ZN(n10356) );
  CLKBUF_X1 U5089 ( .A(n6708), .Z(n8735) );
  AND4_X1 U5099 ( .A1(n5802), .A2(n5804), .A3(n5952), .A4(n5954), .ZN(n10984)
         );
  OR2_X1 U6110 ( .A1(n5987), .A2(n5986), .ZN(n10985) );
endmodule

