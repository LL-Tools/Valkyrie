

module b17_C_SARLock_k_128_4 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9724, n9725, n9726, n9727,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356;

  AOI21_X1 U11151 ( .B1(n15410), .B2(n15408), .A(n15387), .ZN(n15402) );
  NAND2_X1 U11152 ( .A1(n17366), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n17347) );
  NAND2_X1 U11154 ( .A1(n15804), .A2(n15803), .ZN(n14262) );
  NAND2_X1 U11155 ( .A1(n10356), .A2(n13668), .ZN(n9864) );
  NOR3_X1 U11157 ( .A1(n13136), .A2(n13135), .A3(n13134), .ZN(n17559) );
  CLKBUF_X2 U11158 ( .A(n10292), .Z(n11271) );
  INV_X2 U11160 ( .A(n13090), .ZN(n17334) );
  CLKBUF_X2 U11161 ( .A(n11619), .Z(n11585) );
  CLKBUF_X2 U11162 ( .A(n11854), .Z(n12983) );
  CLKBUF_X2 U11163 ( .A(n11741), .Z(n12659) );
  BUF_X4 U11164 ( .A(n10114), .Z(n9720) );
  CLKBUF_X1 U11165 ( .A(n11820), .Z(n20257) );
  NAND4_X2 U11166 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n20243) );
  BUF_X1 U11167 ( .A(n11819), .Z(n12192) );
  BUF_X1 U11168 ( .A(n11765), .Z(n11837) );
  AND2_X1 U11169 ( .A1(n13753), .A2(n15044), .ZN(n11854) );
  AND2_X1 U11170 ( .A1(n15045), .A2(n11701), .ZN(n11741) );
  AND2_X1 U11171 ( .A1(n13755), .A2(n15045), .ZN(n11859) );
  AND2_X1 U11172 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11701) );
  INV_X1 U11174 ( .A(n21356), .ZN(n9707) );
  AND3_X1 U11175 ( .A1(n13745), .A2(n11821), .A3(n12314), .ZN(n11839) );
  CLKBUF_X2 U11178 ( .A(n11800), .Z(n12838) );
  AND2_X1 U11179 ( .A1(n11683), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11700) );
  OR2_X1 U11180 ( .A1(n12147), .A2(n12217), .ZN(n13745) );
  NAND2_X1 U11181 ( .A1(n11913), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9928) );
  AND2_X2 U11182 ( .A1(n11694), .A2(n15044), .ZN(n12610) );
  AND2_X1 U11183 ( .A1(n13753), .A2(n15045), .ZN(n11868) );
  AND2_X1 U11184 ( .A1(n10681), .A2(n10618), .ZN(n10714) );
  AND2_X1 U11185 ( .A1(n11428), .A2(n10367), .ZN(n11457) );
  INV_X1 U11186 ( .A(n10116), .ZN(n11461) );
  AND2_X1 U11187 ( .A1(n10801), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11463) );
  AND2_X1 U11188 ( .A1(n11618), .A2(n15872), .ZN(n11450) );
  AND2_X1 U11189 ( .A1(n10970), .A2(n10604), .ZN(n10262) );
  OR2_X1 U11190 ( .A1(n10334), .A2(n10335), .ZN(n10481) );
  NAND2_X1 U11192 ( .A1(n20266), .A2(n20243), .ZN(n12300) );
  AND4_X1 U11193 ( .A1(n11808), .A2(n11807), .A3(n11806), .A4(n11805), .ZN(
        n11809) );
  AND4_X2 U11194 ( .A1(n11709), .A2(n11708), .A3(n11707), .A4(n11706), .ZN(
        n13019) );
  AND3_X1 U11195 ( .A1(n11815), .A2(n13863), .A3(n11836), .ZN(n12309) );
  OR2_X1 U11196 ( .A1(n12011), .A2(n15038), .ZN(n12014) );
  BUF_X1 U11197 ( .A(n11822), .Z(n20275) );
  INV_X1 U11198 ( .A(n10257), .ZN(n10607) );
  NOR2_X1 U11199 ( .A1(n12920), .A2(n15396), .ZN(n12347) );
  AND2_X1 U11200 ( .A1(n10303), .A2(n10304), .ZN(n10318) );
  NAND2_X1 U11201 ( .A1(n9849), .A2(n9848), .ZN(n11004) );
  AND2_X1 U11203 ( .A1(n13739), .A2(n10329), .ZN(n13998) );
  INV_X1 U11205 ( .A(n12088), .ZN(n9721) );
  INV_X1 U11206 ( .A(n11819), .ZN(n20266) );
  NOR2_X1 U11207 ( .A1(n10732), .A2(n10749), .ZN(n10753) );
  AOI21_X2 U11208 ( .B1(n15464), .B2(n15462), .A(n15379), .ZN(n15456) );
  NOR3_X1 U11209 ( .A1(n18393), .A2(n13292), .A3(n15910), .ZN(n15911) );
  INV_X1 U11210 ( .A(n13089), .ZN(n13140) );
  AND3_X1 U11211 ( .A1(n13063), .A2(n18986), .A3(n17044), .ZN(n10114) );
  INV_X1 U11212 ( .A(n17914), .ZN(n17864) );
  BUF_X1 U11213 ( .A(n12211), .Z(n14026) );
  OR2_X1 U11214 ( .A1(n13446), .A2(n15091), .ZN(n15093) );
  INV_X1 U11215 ( .A(n11007), .ZN(n11284) );
  INV_X1 U11216 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16484) );
  INV_X1 U11217 ( .A(n17002), .ZN(n17025) );
  NAND2_X1 U11218 ( .A1(n17393), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17386) );
  INV_X1 U11219 ( .A(n14002), .ZN(n15276) );
  INV_X1 U11220 ( .A(n11288), .ZN(n15835) );
  AOI211_X1 U11221 ( .C1(n17332), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n13150), .B(n13149), .ZN(n17552) );
  INV_X1 U11222 ( .A(n17953), .ZN(n17971) );
  AND2_X1 U11223 ( .A1(n10252), .A2(n11013), .ZN(n9708) );
  AND3_X1 U11224 ( .A1(n10122), .A2(n10124), .A3(n10123), .ZN(n9709) );
  INV_X1 U11225 ( .A(n17229), .ZN(n9724) );
  AND2_X1 U11226 ( .A1(n10511), .A2(n10510), .ZN(n9710) );
  AND2_X1 U11227 ( .A1(n15500), .A2(n10671), .ZN(n9711) );
  AND2_X1 U11228 ( .A1(n13668), .A2(n10345), .ZN(n9712) );
  AND2_X1 U11229 ( .A1(n11886), .A2(n11884), .ZN(n11850) );
  AND2_X1 U11230 ( .A1(n15044), .A2(n11701), .ZN(n11747) );
  CLKBUF_X1 U11231 ( .A(n11747), .Z(n12986) );
  INV_X2 U11232 ( .A(n17579), .ZN(n18379) );
  AND2_X1 U11233 ( .A1(n13755), .A2(n11699), .ZN(n11800) );
  NAND2_X2 U11235 ( .A1(n10261), .A2(n10260), .ZN(n11233) );
  AND2_X1 U11236 ( .A1(n11699), .A2(n11694), .ZN(n11724) );
  CLKBUF_X1 U11237 ( .A(n11724), .Z(n12861) );
  AND2_X1 U11238 ( .A1(n11694), .A2(n15044), .ZN(n9713) );
  AND2_X1 U11239 ( .A1(n11694), .A2(n15044), .ZN(n9714) );
  INV_X1 U11240 ( .A(n10292), .ZN(n10808) );
  AOI211_X2 U11241 ( .C1(n16252), .C2(n14814), .A(n14813), .B(n14812), .ZN(
        n14815) );
  AND2_X4 U11242 ( .A1(n15870), .A2(n10362), .ZN(n10371) );
  OAI211_X2 U11243 ( .C1(n10635), .C2(n10634), .A(n10633), .B(n10632), .ZN(
        n10661) );
  CLKBUF_X1 U11244 ( .A(n11782), .Z(n9715) );
  AND2_X1 U11245 ( .A1(n11700), .A2(n11694), .ZN(n11782) );
  CLKBUF_X1 U11246 ( .A(n11782), .Z(n12985) );
  NAND2_X2 U11247 ( .A1(n10082), .A2(n10550), .ZN(n10569) );
  AOI21_X4 U11248 ( .B1(n10763), .B2(n10762), .A(n15353), .ZN(n15342) );
  INV_X1 U11249 ( .A(n17295), .ZN(n9716) );
  INV_X2 U11250 ( .A(n17295), .ZN(n9717) );
  OAI21_X2 U11251 ( .B1(n15456), .B2(n15453), .A(n15452), .ZN(n15700) );
  AND2_X1 U11252 ( .A1(n13969), .A2(n9819), .ZN(n14204) );
  NOR2_X2 U11253 ( .A1(n13976), .A2(n13975), .ZN(n13969) );
  INV_X4 U11254 ( .A(n15914), .ZN(n17199) );
  XNOR2_X2 U11255 ( .A(n10470), .B(n10471), .ZN(n15825) );
  NOR3_X2 U11257 ( .A1(n12348), .A2(n15371), .A3(n9906), .ZN(n12951) );
  INV_X1 U11258 ( .A(n13292), .ZN(n9719) );
  INV_X1 U11259 ( .A(n18410), .ZN(n17478) );
  AND2_X2 U11260 ( .A1(n11605), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10453) );
  NAND2_X2 U11261 ( .A1(n10200), .A2(n10199), .ZN(n19425) );
  INV_X1 U11262 ( .A(n11300), .ZN(n10328) );
  AOI21_X2 U11263 ( .B1(n15478), .B2(n10101), .A(n10095), .ZN(n11247) );
  INV_X4 U11264 ( .A(n13250), .ZN(n17332) );
  OR2_X1 U11265 ( .A1(n15528), .A2(n16436), .ZN(n9895) );
  XNOR2_X1 U11266 ( .A(n15300), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15528) );
  AOI21_X1 U11267 ( .B1(n13044), .B2(n13012), .A(n13043), .ZN(n14794) );
  NAND2_X1 U11268 ( .A1(n9852), .A2(n15627), .ZN(n15424) );
  NAND2_X1 U11269 ( .A1(n10913), .A2(n11240), .ZN(n15689) );
  NOR3_X1 U11270 ( .A1(n15098), .A2(n11658), .A3(n9971), .ZN(n9973) );
  INV_X2 U11271 ( .A(n10635), .ZN(n9868) );
  AND2_X1 U11272 ( .A1(n17468), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17466) );
  AND4_X1 U11273 ( .A1(n10344), .A2(n10342), .A3(n10343), .A4(n10341), .ZN(
        n10360) );
  XNOR2_X1 U11274 ( .A(n13737), .B(n13738), .ZN(n19503) );
  AOI22_X1 U11275 ( .A1(n18047), .A2(n9878), .B1(n17968), .B2(n18240), .ZN(
        n17956) );
  NAND2_X1 U11276 ( .A1(n10317), .A2(n10318), .ZN(n10316) );
  OAI211_X1 U11277 ( .C1(n9928), .C2(n9926), .A(n9925), .B(n9924), .ZN(n11852)
         );
  NAND2_X1 U11278 ( .A1(n11818), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11912) );
  INV_X2 U11279 ( .A(n11212), .ZN(n11009) );
  OR2_X1 U11280 ( .A1(n13342), .A2(n18821), .ZN(n15910) );
  NOR2_X1 U11281 ( .A1(n12183), .A2(n14025), .ZN(n12205) );
  INV_X1 U11282 ( .A(n16080), .ZN(n18053) );
  INV_X1 U11283 ( .A(n17572), .ZN(n13163) );
  INV_X4 U11284 ( .A(n10932), .ZN(n10263) );
  NOR2_X2 U11285 ( .A1(n12192), .A2(n20261), .ZN(n13863) );
  CLKBUF_X2 U11286 ( .A(n11026), .Z(n12889) );
  OR2_X1 U11287 ( .A1(n10437), .A2(n10436), .ZN(n11033) );
  NAND2_X1 U11288 ( .A1(n11739), .A2(n9788), .ZN(n11814) );
  NAND4_X2 U11289 ( .A1(n11812), .A2(n11811), .A3(n11810), .A4(n11809), .ZN(
        n12211) );
  INV_X4 U11290 ( .A(n17322), .ZN(n17367) );
  CLKBUF_X2 U11291 ( .A(n11997), .Z(n12994) );
  CLKBUF_X2 U11292 ( .A(n11868), .Z(n12715) );
  INV_X2 U11293 ( .A(n17298), .ZN(n17377) );
  INV_X2 U11294 ( .A(n9785), .ZN(n17274) );
  INV_X4 U11295 ( .A(n17373), .ZN(n17215) );
  INV_X4 U11296 ( .A(n17338), .ZN(n13113) );
  NAND2_X2 U11297 ( .A1(n19014), .A2(n9732), .ZN(n17056) );
  INV_X8 U11298 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13208) );
  INV_X1 U11299 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n9747) );
  INV_X1 U11300 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15872) );
  INV_X2 U11301 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10362) );
  INV_X1 U11302 ( .A(n15405), .ZN(n15378) );
  XNOR2_X1 U11303 ( .A(n15305), .B(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15536) );
  NAND2_X1 U11304 ( .A1(n14787), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12385) );
  AOI22_X1 U11305 ( .A1(n16260), .A2(n16360), .B1(n16367), .B2(n16259), .ZN(
        n16268) );
  AND2_X2 U11306 ( .A1(n15304), .A2(n9958), .ZN(n15300) );
  NAND2_X1 U11307 ( .A1(n12384), .A2(n12383), .ZN(n14787) );
  NOR2_X2 U11308 ( .A1(n15424), .A2(n21279), .ZN(n15417) );
  AND2_X2 U11309 ( .A1(n15320), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15304) );
  NAND2_X1 U11310 ( .A1(n12379), .A2(n10093), .ZN(n14788) );
  XNOR2_X1 U11311 ( .A(n14809), .B(n16264), .ZN(n16258) );
  AND2_X1 U11312 ( .A1(n12120), .A2(n12381), .ZN(n12379) );
  XNOR2_X1 U11313 ( .A(n10048), .B(n10047), .ZN(n14576) );
  NOR2_X2 U11314 ( .A1(n15690), .A2(n15687), .ZN(n15661) );
  NOR2_X2 U11315 ( .A1(n15347), .A2(n21297), .ZN(n15328) );
  AND2_X1 U11316 ( .A1(n15785), .A2(n9744), .ZN(n15761) );
  INV_X1 U11317 ( .A(n15689), .ZN(n9852) );
  OAI21_X1 U11318 ( .B1(n14807), .B2(n12119), .A(n9721), .ZN(n12120) );
  AND2_X1 U11319 ( .A1(n10076), .A2(n10074), .ZN(n15432) );
  CLKBUF_X1 U11320 ( .A(n10913), .Z(n15785) );
  AND2_X1 U11321 ( .A1(n10078), .A2(n10746), .ZN(n15410) );
  AND2_X1 U11322 ( .A1(n9756), .A2(n10575), .ZN(n9733) );
  NAND2_X2 U11324 ( .A1(n15342), .A2(n15332), .ZN(n15307) );
  OR2_X1 U11325 ( .A1(n9758), .A2(n10570), .ZN(n9757) );
  CLKBUF_X1 U11326 ( .A(n15499), .Z(n9729) );
  AND2_X1 U11327 ( .A1(n15186), .A2(n9985), .ZN(n15193) );
  NAND2_X1 U11328 ( .A1(n9948), .A2(n9721), .ZN(n16191) );
  INV_X1 U11329 ( .A(n14851), .ZN(n9950) );
  NOR2_X1 U11330 ( .A1(n14861), .A2(n12113), .ZN(n14951) );
  AOI211_X1 U11331 ( .C1(n15551), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15550), .B(n15549), .ZN(n15552) );
  NAND2_X1 U11332 ( .A1(n15198), .A2(n15197), .ZN(n15196) );
  AND2_X1 U11333 ( .A1(n11679), .A2(n11678), .ZN(n11680) );
  AOI211_X1 U11334 ( .C1(n17715), .C2(n16566), .A(n16577), .B(n18074), .ZN(
        n16573) );
  OR2_X1 U11335 ( .A1(n13388), .A2(n17958), .ZN(n13202) );
  AND2_X1 U11336 ( .A1(n11632), .A2(n11631), .ZN(n11633) );
  NAND2_X1 U11337 ( .A1(n12112), .A2(n12111), .ZN(n14861) );
  AND2_X1 U11338 ( .A1(n11276), .A2(n11269), .ZN(n9870) );
  INV_X1 U11339 ( .A(n13203), .ZN(n13389) );
  AND2_X1 U11340 ( .A1(n12893), .A2(n11659), .ZN(n15516) );
  OR2_X1 U11341 ( .A1(n17704), .A2(n17703), .ZN(n17705) );
  NAND4_X1 U11342 ( .A1(n9842), .A2(n9773), .A3(n9841), .A4(n9839), .ZN(n14449) );
  XNOR2_X1 U11343 ( .A(n11275), .B(n11274), .ZN(n14525) );
  AOI21_X1 U11344 ( .B1(n10902), .B2(n15080), .A(n11275), .ZN(n15515) );
  INV_X1 U11345 ( .A(n16560), .ZN(n17715) );
  AND2_X1 U11346 ( .A1(n10901), .A2(n10011), .ZN(n11275) );
  OAI21_X1 U11347 ( .B1(n14294), .B2(n9951), .A(n9952), .ZN(n14865) );
  NOR2_X1 U11348 ( .A1(n9745), .A2(n14450), .ZN(n9871) );
  NAND2_X1 U11349 ( .A1(n9996), .A2(n9995), .ZN(n9998) );
  AOI211_X1 U11350 ( .C1(n16398), .C2(n16457), .A(n15568), .B(n15567), .ZN(
        n15569) );
  INV_X1 U11351 ( .A(n15093), .ZN(n10901) );
  NAND2_X1 U11352 ( .A1(n12084), .A2(n12083), .ZN(n14294) );
  INV_X1 U11353 ( .A(n10572), .ZN(n10574) );
  NOR2_X1 U11354 ( .A1(n13448), .A2(n13449), .ZN(n11651) );
  AND2_X1 U11355 ( .A1(n13195), .A2(n17958), .ZN(n13196) );
  NAND2_X1 U11356 ( .A1(n10512), .A2(n10990), .ZN(n9762) );
  AND2_X1 U11357 ( .A1(n11471), .A2(n11495), .ZN(n11472) );
  NOR2_X1 U11358 ( .A1(n15221), .A2(n15220), .ZN(n15219) );
  INV_X1 U11359 ( .A(n17441), .ZN(n17437) );
  XNOR2_X1 U11360 ( .A(n13056), .B(n13055), .ZN(n14913) );
  XNOR2_X1 U11361 ( .A(n9994), .B(n9993), .ZN(n15221) );
  NAND2_X1 U11362 ( .A1(n9991), .A2(n9780), .ZN(n9994) );
  NAND2_X1 U11363 ( .A1(n9923), .A2(n13192), .ZN(n17825) );
  INV_X1 U11364 ( .A(n15233), .ZN(n9991) );
  NAND2_X1 U11365 ( .A1(n9823), .A2(n10115), .ZN(n15233) );
  NOR2_X2 U11366 ( .A1(n15164), .A2(n15149), .ZN(n15151) );
  NOR2_X1 U11367 ( .A1(n17832), .A2(n13193), .ZN(n17794) );
  AND2_X1 U11368 ( .A1(n15120), .A2(n11262), .ZN(n10786) );
  OR2_X1 U11369 ( .A1(n15161), .A2(n15162), .ZN(n15164) );
  AND2_X1 U11370 ( .A1(n10778), .A2(n10777), .ZN(n15120) );
  NAND2_X1 U11371 ( .A1(n15651), .A2(n15650), .ZN(n14331) );
  NAND2_X1 U11372 ( .A1(n9917), .A2(n17847), .ZN(n13188) );
  NAND4_X1 U11373 ( .A1(n10496), .A2(n10494), .A3(n10495), .A4(n10493), .ZN(
        n10511) );
  NAND2_X1 U11374 ( .A1(n12408), .A2(n12407), .ZN(n13837) );
  OAI21_X1 U11375 ( .B1(n12448), .B2(n12558), .A(n12447), .ZN(n13936) );
  AND4_X1 U11376 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10494) );
  AND2_X1 U11377 ( .A1(n10755), .A2(n15216), .ZN(n10776) );
  AND4_X1 U11378 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10529) );
  CLKBUF_X1 U11379 ( .A(n12076), .Z(n12087) );
  AND4_X1 U11380 ( .A1(n10414), .A2(n10413), .A3(n10412), .A4(n10411), .ZN(
        n10423) );
  NAND2_X1 U11381 ( .A1(n12035), .A2(n9809), .ZN(n12076) );
  OAI21_X1 U11382 ( .B1(n13948), .B2(n13947), .A(n11968), .ZN(n11994) );
  OAI22_X1 U11383 ( .A1(n19478), .A2(n10476), .B1(n11160), .B2(n9847), .ZN(
        n10477) );
  NAND2_X1 U11384 ( .A1(n12014), .A2(n11990), .ZN(n20241) );
  NAND2_X1 U11385 ( .A1(n15724), .A2(n15725), .ZN(n15711) );
  AND2_X1 U11386 ( .A1(n11309), .A2(n13785), .ZN(n13738) );
  NAND2_X1 U11388 ( .A1(n17257), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n17240) );
  AND2_X1 U11389 ( .A1(n10737), .A2(n10863), .ZN(n15420) );
  NOR2_X2 U11390 ( .A1(n18887), .A2(n18049), .ZN(n17914) );
  NOR2_X2 U11391 ( .A1(n17243), .A2(n17242), .ZN(n17257) );
  NOR2_X2 U11392 ( .A1(n17548), .A2(n18057), .ZN(n17968) );
  NOR2_X2 U11393 ( .A1(n13347), .A2(n18057), .ZN(n17953) );
  NOR2_X1 U11394 ( .A1(n18163), .A2(n17927), .ZN(n16563) );
  INV_X1 U11395 ( .A(n10355), .ZN(n10356) );
  OR2_X2 U11396 ( .A1(n10334), .A2(n10331), .ZN(n10480) );
  NAND2_X1 U11397 ( .A1(n18054), .A2(n17895), .ZN(n17837) );
  NAND2_X1 U11398 ( .A1(n18054), .A2(n18017), .ZN(n18049) );
  NAND2_X1 U11399 ( .A1(n13348), .A2(n17642), .ZN(n18057) );
  NOR2_X1 U11400 ( .A1(n13809), .A2(n13810), .ZN(n13808) );
  NAND2_X1 U11401 ( .A1(n11283), .A2(n11282), .ZN(n11297) );
  AND2_X1 U11402 ( .A1(n13598), .A2(n11294), .ZN(n13665) );
  NAND2_X1 U11403 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n13185), .ZN(
        n17927) );
  NAND2_X1 U11404 ( .A1(n11989), .A2(n11988), .ZN(n15035) );
  INV_X1 U11405 ( .A(n16680), .ZN(n13348) );
  NOR2_X2 U11406 ( .A1(n17642), .A2(n16680), .ZN(n18047) );
  CLKBUF_X1 U11407 ( .A(n13743), .Z(n20563) );
  NOR2_X2 U11408 ( .A1(n13037), .A2(n20239), .ZN(n13035) );
  NAND2_X1 U11409 ( .A1(n13815), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13814) );
  NAND2_X1 U11410 ( .A1(n9856), .A2(n9854), .ZN(n16680) );
  XNOR2_X1 U11411 ( .A(n11969), .B(n20406), .ZN(n13743) );
  NOR2_X1 U11412 ( .A1(n14436), .A2(n14435), .ZN(n14475) );
  NAND2_X1 U11413 ( .A1(n11052), .A2(n11051), .ZN(n15804) );
  OR2_X1 U11414 ( .A1(n18808), .A2(n9857), .ZN(n9856) );
  NAND2_X1 U11415 ( .A1(n10320), .A2(n10319), .ZN(n10321) );
  NAND2_X1 U11416 ( .A1(n11291), .A2(n11290), .ZN(n15849) );
  NOR2_X1 U11417 ( .A1(n17429), .A2(n17428), .ZN(n17554) );
  NAND2_X2 U11418 ( .A1(n20153), .A2(n20286), .ZN(n14728) );
  NOR2_X2 U11419 ( .A1(n17642), .A2(n18270), .ZN(n18808) );
  AND2_X2 U11420 ( .A1(n13047), .A2(n14575), .ZN(n20153) );
  NAND2_X1 U11421 ( .A1(n10714), .A2(n9808), .ZN(n10710) );
  AND2_X1 U11422 ( .A1(n10337), .A2(n10327), .ZN(n11289) );
  AND2_X1 U11423 ( .A1(n10811), .A2(n10315), .ZN(n10813) );
  NAND2_X1 U11424 ( .A1(n18002), .A2(n13177), .ZN(n17985) );
  NOR2_X2 U11425 ( .A1(n18828), .A2(n18818), .ZN(n9863) );
  NOR2_X1 U11426 ( .A1(n14399), .A2(n14131), .ZN(n14446) );
  INV_X1 U11427 ( .A(n11852), .ZN(n20371) );
  NAND2_X1 U11428 ( .A1(n18003), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18002) );
  INV_X2 U11429 ( .A(n15229), .ZN(n13900) );
  OAI21_X1 U11430 ( .B1(n13367), .B2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n17998), .ZN(n13370) );
  AND2_X1 U11431 ( .A1(n10308), .A2(n10307), .ZN(n10311) );
  AND2_X1 U11432 ( .A1(n16003), .A2(n16002), .ZN(n16697) );
  AOI21_X1 U11433 ( .B1(n11914), .B2(n21244), .A(n11915), .ZN(n11920) );
  XNOR2_X1 U11434 ( .A(n11029), .B(n11030), .ZN(n13630) );
  AND2_X1 U11435 ( .A1(n13316), .A2(n13315), .ZN(n16003) );
  NAND2_X1 U11436 ( .A1(n10617), .A2(n10616), .ZN(n10686) );
  INV_X1 U11437 ( .A(n9927), .ZN(n9926) );
  CLKBUF_X1 U11438 ( .A(n16428), .Z(n19409) );
  AOI21_X1 U11439 ( .B1(n14322), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10254), 
        .ZN(n10255) );
  INV_X1 U11440 ( .A(n10663), .ZN(n10617) );
  NAND2_X1 U11441 ( .A1(n10253), .A2(n9787), .ZN(n14322) );
  NOR2_X1 U11442 ( .A1(n18022), .A2(n13361), .ZN(n13363) );
  XNOR2_X1 U11443 ( .A(n13607), .B(n11020), .ZN(n13828) );
  AND2_X1 U11444 ( .A1(n10266), .A2(n10265), .ZN(n10267) );
  AND2_X1 U11445 ( .A1(n10283), .A2(n9787), .ZN(n10260) );
  INV_X2 U11446 ( .A(n11270), .ZN(n10896) );
  AND3_X1 U11447 ( .A1(n11041), .A2(n11040), .A3(n11039), .ZN(n14116) );
  OR2_X1 U11448 ( .A1(n10998), .A2(n13571), .ZN(n10270) );
  AND2_X1 U11449 ( .A1(n10975), .A2(n10229), .ZN(n10274) );
  CLKBUF_X1 U11450 ( .A(n10283), .Z(n14315) );
  OR2_X1 U11451 ( .A1(n17556), .A2(n13173), .ZN(n13178) );
  AOI21_X1 U11452 ( .B1(n12205), .B2(n11816), .A(n12309), .ZN(n11817) );
  AND3_X1 U11453 ( .A1(n11845), .A2(n11844), .A3(n11843), .ZN(n11849) );
  NAND2_X1 U11454 ( .A1(n13324), .A2(n13404), .ZN(n13327) );
  NOR4_X1 U11455 ( .A1(n18393), .A2(n18389), .A3(n13317), .A4(n13319), .ZN(
        n13329) );
  AND2_X2 U11456 ( .A1(n11629), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10292) );
  AND2_X1 U11457 ( .A1(n10250), .A2(n9708), .ZN(n9748) );
  CLKBUF_X1 U11458 ( .A(n11634), .Z(n9750) );
  INV_X1 U11459 ( .A(n10662), .ZN(n10616) );
  NAND2_X1 U11460 ( .A1(n17432), .A2(n17435), .ZN(n13342) );
  AND3_X2 U11461 ( .A1(n10264), .A2(n10263), .A3(n10262), .ZN(n11629) );
  NOR2_X1 U11462 ( .A1(n17562), .A2(n13166), .ZN(n13170) );
  INV_X1 U11463 ( .A(n10262), .ZN(n10981) );
  INV_X1 U11464 ( .A(n18404), .ZN(n17432) );
  AND2_X1 U11465 ( .A1(n10604), .A2(n11013), .ZN(n10805) );
  OR2_X1 U11466 ( .A1(n9898), .A2(n9897), .ZN(n12925) );
  NAND3_X1 U11467 ( .A1(n9793), .A2(n13111), .A3(n13110), .ZN(n17572) );
  AND2_X1 U11468 ( .A1(n13269), .A2(n13268), .ZN(n18404) );
  NAND2_X1 U11469 ( .A1(n10215), .A2(n10080), .ZN(n10972) );
  OAI211_X1 U11470 ( .C1(n17322), .C2(n17405), .A(n13243), .B(n13242), .ZN(
        n18398) );
  INV_X1 U11471 ( .A(n17567), .ZN(n13125) );
  INV_X1 U11472 ( .A(n18389), .ZN(n13326) );
  CLKBUF_X1 U11473 ( .A(n11836), .Z(n14023) );
  AND2_X1 U11474 ( .A1(n13099), .A2(n9919), .ZN(n17562) );
  OR2_X1 U11475 ( .A1(n10406), .A2(n10405), .ZN(n10583) );
  AOI211_X1 U11476 ( .C1(n13113), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n13277), .B(n13276), .ZN(n13278) );
  INV_X1 U11478 ( .A(n20243), .ZN(n14025) );
  AND2_X2 U11479 ( .A1(n11004), .A2(n11002), .ZN(n11032) );
  INV_X1 U11480 ( .A(n11814), .ZN(n12193) );
  INV_X1 U11481 ( .A(n11765), .ZN(n12398) );
  INV_X2 U11482 ( .A(n14076), .ZN(n9722) );
  INV_X1 U11483 ( .A(n10202), .ZN(n10230) );
  OR2_X1 U11484 ( .A1(n12929), .A2(n10907), .ZN(n12944) );
  NAND2_X2 U11485 ( .A1(n10147), .A2(n10146), .ZN(n10257) );
  OR2_X2 U11486 ( .A1(n11753), .A2(n11752), .ZN(n11822) );
  OR2_X1 U11487 ( .A1(n11897), .A2(n11896), .ZN(n12090) );
  AND2_X2 U11488 ( .A1(n10172), .A2(n10171), .ZN(n10202) );
  OR2_X2 U11489 ( .A1(n11719), .A2(n11718), .ZN(n20286) );
  OR2_X1 U11490 ( .A1(n11730), .A2(n11729), .ZN(n11765) );
  NAND2_X2 U11491 ( .A1(n10185), .A2(n10184), .ZN(n11013) );
  AND4_X1 U11492 ( .A1(n11734), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(
        n11739) );
  AND4_X1 U11493 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11812) );
  AND4_X1 U11494 ( .A1(n11804), .A2(n11803), .A3(n11802), .A4(n11801), .ZN(
        n11810) );
  AND4_X1 U11495 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n11790) );
  AND4_X1 U11496 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11789) );
  AND4_X1 U11497 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n11788) );
  AND4_X1 U11498 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n11709) );
  AND4_X1 U11499 ( .A1(n11693), .A2(n11692), .A3(n11691), .A4(n11690), .ZN(
        n11708) );
  AND4_X1 U11500 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11707) );
  AND4_X1 U11501 ( .A1(n11705), .A2(n11704), .A3(n11703), .A4(n11702), .ZN(
        n11706) );
  NOR2_X2 U11502 ( .A1(n20239), .A2(n20238), .ZN(n20240) );
  AND2_X2 U11503 ( .A1(n10193), .A2(n15872), .ZN(n11456) );
  NAND2_X2 U11504 ( .A1(n20052), .A2(n19950), .ZN(n19995) );
  NAND2_X2 U11505 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20052), .ZN(n19993) );
  AND2_X1 U11506 ( .A1(n10195), .A2(n10196), .ZN(n9743) );
  AOI22_X1 U11507 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11724), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11750) );
  AND4_X1 U11508 ( .A1(n11786), .A2(n11785), .A3(n11784), .A4(n11783), .ZN(
        n11787) );
  AND2_X2 U11509 ( .A1(n11585), .A2(n15872), .ZN(n11448) );
  NOR2_X2 U11510 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18593), .ZN(
        n18608) );
  INV_X2 U11511 ( .A(n16664), .ZN(U215) );
  INV_X4 U11512 ( .A(n17371), .ZN(n17086) );
  INV_X4 U11513 ( .A(n10111), .ZN(n17368) );
  NAND2_X2 U11514 ( .A1(n19041), .A2(n18913), .ZN(n18964) );
  NOR2_X1 U11515 ( .A1(n18887), .A2(n18891), .ZN(n19030) );
  BUF_X2 U11516 ( .A(n12589), .Z(n12993) );
  BUF_X2 U11517 ( .A(n11859), .Z(n12987) );
  INV_X1 U11518 ( .A(n10193), .ZN(n9725) );
  BUF_X2 U11520 ( .A(n12589), .Z(n12839) );
  NAND3_X1 U11521 ( .A1(n13063), .A2(n18986), .A3(n13064), .ZN(n17371) );
  OR2_X2 U11522 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13066), .ZN(
        n13090) );
  NAND2_X1 U11523 ( .A1(n13064), .A2(n13067), .ZN(n17295) );
  INV_X2 U11524 ( .A(n20053), .ZN(n20052) );
  OAI221_X1 U11525 ( .B1(n21088), .B2(keyinput35), .C1(n21087), .C2(keyinput28), .A(n21086), .ZN(n21101) );
  INV_X2 U11526 ( .A(n16668), .ZN(n16670) );
  BUF_X2 U11527 ( .A(n10371), .Z(n11618) );
  AND2_X1 U11528 ( .A1(n10908), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10254) );
  AND2_X2 U11529 ( .A1(n11682), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13753) );
  AND2_X1 U11530 ( .A1(n18986), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13065) );
  INV_X2 U11531 ( .A(n10178), .ZN(n9726) );
  AND2_X1 U11532 ( .A1(n9982), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14323) );
  NAND2_X2 U11533 ( .A1(n20004), .A2(n10908), .ZN(n19214) );
  NAND2_X1 U11534 ( .A1(n12935), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12932) );
  INV_X1 U11535 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9732) );
  NAND3_X1 U11536 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16008) );
  NOR2_X2 U11537 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15852) );
  AND2_X1 U11538 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15870) );
  INV_X2 U11539 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13063) );
  INV_X1 U11540 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19408) );
  AND2_X1 U11541 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17044) );
  NOR2_X2 U11542 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20689) );
  CLKBUF_X1 U11543 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n21244) );
  AND2_X1 U11544 ( .A1(n10201), .A2(n9801), .ZN(n9727) );
  AOI22_X1 U11545 ( .A1(n10484), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n19725), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10342) );
  XNOR2_X1 U11546 ( .A(n10569), .B(n10567), .ZN(n15499) );
  NAND2_X1 U11547 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U11548 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n9731) );
  AND2_X1 U11549 ( .A1(n9730), .A2(n9731), .ZN(n13153) );
  INV_X2 U11550 ( .A(n14149), .ZN(n19242) );
  OR2_X1 U11551 ( .A1(n19759), .A2(n11339), .ZN(n10341) );
  NOR2_X1 U11552 ( .A1(n16014), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13388) );
  NAND2_X1 U11553 ( .A1(n10328), .A2(n9712), .ZN(n19451) );
  NAND2_X1 U11554 ( .A1(n10232), .A2(n10951), .ZN(n9734) );
  NAND2_X1 U11555 ( .A1(n10232), .A2(n10951), .ZN(n9956) );
  NAND2_X1 U11556 ( .A1(n10953), .A2(n10249), .ZN(n9735) );
  NAND2_X1 U11557 ( .A1(n10953), .A2(n10249), .ZN(n10996) );
  INV_X1 U11558 ( .A(n9722), .ZN(n9736) );
  NAND2_X2 U11559 ( .A1(n9851), .A2(n9850), .ZN(n14076) );
  NAND2_X1 U11561 ( .A1(n15500), .A2(n9741), .ZN(n9738) );
  AND2_X2 U11562 ( .A1(n9738), .A2(n9739), .ZN(n15478) );
  OR2_X1 U11563 ( .A1(n9740), .A2(n10691), .ZN(n9739) );
  INV_X1 U11564 ( .A(n10069), .ZN(n9740) );
  AND2_X1 U11565 ( .A1(n10671), .A2(n10069), .ZN(n9741) );
  INV_X1 U11566 ( .A(n10248), .ZN(n9742) );
  NAND3_X1 U11567 ( .A1(n10197), .A2(n9743), .A3(n10194), .ZN(n10198) );
  INV_X1 U11568 ( .A(n10248), .ZN(n16515) );
  NAND2_X1 U11569 ( .A1(n15500), .A2(n10671), .ZN(n15484) );
  NOR2_X2 U11570 ( .A1(n11022), .A2(n11021), .ZN(n11029) );
  NOR2_X2 U11571 ( .A1(n15275), .A2(n15113), .ZN(n15112) );
  XNOR2_X2 U11572 ( .A(n12893), .B(n12892), .ZN(n14528) );
  NOR2_X1 U11573 ( .A1(n18986), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13067) );
  BUF_X4 U11574 ( .A(n13140), .Z(n17314) );
  NAND2_X1 U11575 ( .A1(n10125), .A2(n9709), .ZN(n10126) );
  AND2_X1 U11576 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9744) );
  NAND2_X2 U11577 ( .A1(n15378), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15377) );
  NAND2_X1 U11578 ( .A1(n15417), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15405) );
  AND2_X2 U11579 ( .A1(n10639), .A2(n9866), .ZN(n9745) );
  INV_X1 U11580 ( .A(n9745), .ZN(n14452) );
  AOI21_X1 U11581 ( .B1(n10297), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10310), .ZN(n10312) );
  AOI21_X1 U11582 ( .B1(n10297), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10298), .ZN(n10301) );
  XNOR2_X1 U11583 ( .A(n11994), .B(n14187), .ZN(n13940) );
  XNOR2_X2 U11584 ( .A(n11902), .B(n11937), .ZN(n12423) );
  NAND2_X1 U11585 ( .A1(n10230), .A2(n11013), .ZN(n9746) );
  OR2_X2 U11586 ( .A1(n10305), .A2(n9747), .ZN(n10296) );
  NAND2_X1 U11587 ( .A1(n10262), .A2(n9748), .ZN(n9787) );
  INV_X1 U11588 ( .A(n15844), .ZN(n9749) );
  NAND2_X1 U11589 ( .A1(n10231), .A2(n19425), .ZN(n9751) );
  NAND2_X1 U11590 ( .A1(n9752), .A2(n9751), .ZN(n10246) );
  AND2_X1 U11591 ( .A1(n10109), .A2(n10201), .ZN(n9752) );
  NAND2_X1 U11592 ( .A1(n10660), .A2(n14301), .ZN(n9753) );
  NAND2_X1 U11593 ( .A1(n10511), .A2(n10510), .ZN(n9754) );
  NAND2_X1 U11594 ( .A1(n10511), .A2(n10510), .ZN(n9755) );
  NAND2_X1 U11596 ( .A1(n10660), .A2(n14301), .ZN(n14451) );
  OR2_X1 U11597 ( .A1(n10551), .A2(n10626), .ZN(n10572) );
  NAND2_X1 U11598 ( .A1(n15499), .A2(n9759), .ZN(n9756) );
  INV_X1 U11599 ( .A(n16444), .ZN(n9758) );
  AND2_X1 U11600 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n16444), .ZN(
        n9759) );
  OAI21_X2 U11601 ( .B1(n15307), .B2(n10780), .A(n9837), .ZN(n9865) );
  NAND2_X1 U11602 ( .A1(n10571), .A2(n10570), .ZN(n16443) );
  NAND2_X1 U11603 ( .A1(n10324), .A2(n10323), .ZN(n10337) );
  NOR2_X2 U11604 ( .A1(n14369), .A2(n14433), .ZN(n14432) );
  NAND2_X2 U11605 ( .A1(n12011), .A2(n11958), .ZN(n12414) );
  OAI22_X2 U11606 ( .A1(n13860), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11961), 
        .B2(n11977), .ZN(n11936) );
  NOR2_X2 U11607 ( .A1(n14593), .A2(n14594), .ZN(n12875) );
  NOR2_X2 U11608 ( .A1(n14641), .A2(n10038), .ZN(n14606) );
  INV_X1 U11609 ( .A(n9764), .ZN(n9760) );
  INV_X1 U11610 ( .A(n9760), .ZN(n9761) );
  INV_X1 U11611 ( .A(n9762), .ZN(n14304) );
  CLKBUF_X1 U11612 ( .A(n14300), .Z(n9763) );
  INV_X1 U11613 ( .A(n9761), .ZN(n14303) );
  NOR2_X2 U11614 ( .A1(n17956), .A2(n18163), .ZN(n17833) );
  INV_X2 U11615 ( .A(n11277), .ZN(n13668) );
  AND2_X2 U11616 ( .A1(n15478), .A2(n10718), .ZN(n15464) );
  AND2_X2 U11617 ( .A1(n10474), .A2(n10473), .ZN(n9764) );
  NAND2_X2 U11618 ( .A1(n10159), .A2(n10158), .ZN(n10242) );
  INV_X1 U11619 ( .A(n9735), .ZN(n10253) );
  AND2_X1 U11620 ( .A1(n10222), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11077) );
  OAI21_X1 U11621 ( .B1(n9775), .B2(n21220), .A(n13194), .ZN(n17732) );
  NOR2_X2 U11622 ( .A1(n17944), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17931) );
  OR2_X2 U11623 ( .A1(n17838), .A2(n17958), .ZN(n13192) );
  NOR2_X2 U11624 ( .A1(n13198), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16561) );
  INV_X2 U11625 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15855) );
  INV_X4 U11626 ( .A(n17229), .ZN(n9765) );
  NAND2_X1 U11627 ( .A1(n13068), .A2(n13065), .ZN(n17229) );
  INV_X2 U11628 ( .A(n10178), .ZN(n9766) );
  NOR3_X2 U11629 ( .A1(n13124), .A2(n13123), .A3(n13122), .ZN(n17567) );
  NOR2_X1 U11630 ( .A1(n10932), .A2(n12955), .ZN(n10280) );
  OAI21_X2 U11631 ( .B1(n10305), .B2(n15833), .A(n10267), .ZN(n10287) );
  INV_X2 U11632 ( .A(n10305), .ZN(n10886) );
  INV_X4 U11633 ( .A(n17205), .ZN(n9767) );
  XNOR2_X2 U11634 ( .A(n10288), .B(n10287), .ZN(n10322) );
  NOR2_X4 U11635 ( .A1(n14331), .A2(n14332), .ZN(n14330) );
  INV_X2 U11636 ( .A(n10328), .ZN(n13739) );
  AND2_X1 U11637 ( .A1(n10361), .A2(n15872), .ZN(n11451) );
  AND2_X1 U11638 ( .A1(n10361), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10424) );
  AND2_X2 U11639 ( .A1(n15328), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15320) );
  AND2_X1 U11640 ( .A1(n14321), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9768) );
  AOI21_X1 U11641 ( .B1(n10361), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n10209), .ZN(n10213) );
  BUF_X4 U11642 ( .A(n10221), .Z(n10361) );
  NAND2_X2 U11643 ( .A1(n10913), .A2(n9957), .ZN(n15347) );
  NAND2_X2 U11644 ( .A1(n9733), .A2(n9757), .ZN(n10913) );
  INV_X4 U11645 ( .A(n10611), .ZN(n19435) );
  BUF_X4 U11646 ( .A(n10607), .Z(n10611) );
  NAND3_X2 U11647 ( .A1(n9853), .A2(n10468), .A3(n10450), .ZN(n14169) );
  NOR2_X4 U11648 ( .A1(n15377), .A2(n10915), .ZN(n15368) );
  NAND2_X1 U11649 ( .A1(n9722), .A2(n11007), .ZN(n10926) );
  INV_X2 U11650 ( .A(n10242), .ZN(n10187) );
  NAND2_X2 U11651 ( .A1(n14169), .A2(n10452), .ZN(n10470) );
  NAND2_X2 U11652 ( .A1(n11233), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10305) );
  INV_X2 U11653 ( .A(n10134), .ZN(n9769) );
  INV_X1 U11654 ( .A(n10134), .ZN(n9770) );
  INV_X1 U11656 ( .A(n10134), .ZN(n10193) );
  NAND2_X2 U11657 ( .A1(n10370), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10134) );
  NAND2_X2 U11658 ( .A1(n14076), .A2(n11004), .ZN(n10932) );
  INV_X2 U11659 ( .A(n10240), .ZN(n10604) );
  NAND2_X1 U11660 ( .A1(n13345), .A2(n13327), .ZN(n13332) );
  AOI21_X1 U11661 ( .B1(n13215), .B2(n13214), .A(n13213), .ZN(n13337) );
  INV_X2 U11662 ( .A(n10615), .ZN(n11262) );
  CLKBUF_X1 U11663 ( .A(n11927), .Z(n12984) );
  OR2_X1 U11665 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20236), .ZN(
        n12130) );
  NAND2_X1 U11666 ( .A1(n10589), .A2(n10588), .ZN(n10595) );
  NAND2_X1 U11667 ( .A1(n14606), .A2(n14608), .ZN(n14593) );
  AOI21_X1 U11668 ( .B1(n14865), .B2(n12109), .A(n12088), .ZN(n12110) );
  AOI21_X1 U11669 ( .B1(n9938), .B2(n9939), .A(n9791), .ZN(n9934) );
  XNOR2_X1 U11670 ( .A(n12076), .B(n12075), .ZN(n12465) );
  NAND2_X1 U11671 ( .A1(n13048), .A2(n13683), .ZN(n12306) );
  NAND2_X1 U11672 ( .A1(n13019), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11977) );
  OR2_X1 U11673 ( .A1(n20243), .A2(n11887), .ZN(n11976) );
  OR2_X1 U11674 ( .A1(n11941), .A2(n11940), .ZN(n11942) );
  NOR2_X1 U11675 ( .A1(n10005), .A2(n14044), .ZN(n10004) );
  INV_X1 U11676 ( .A(n13970), .ZN(n10005) );
  AOI211_X1 U11677 ( .C1(n11561), .C2(n11559), .A(n13783), .B(n15184), .ZN(
        n11560) );
  NAND2_X1 U11678 ( .A1(n11539), .A2(n9987), .ZN(n9986) );
  NOR2_X2 U11679 ( .A1(n9887), .A2(n9790), .ZN(n10615) );
  NAND2_X1 U11680 ( .A1(n10566), .A2(n9888), .ZN(n9887) );
  NAND2_X1 U11681 ( .A1(n11277), .A2(n15835), .ZN(n10353) );
  NAND2_X1 U11682 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17978), .ZN(
        n13377) );
  NAND3_X2 U11683 ( .A1(n13063), .A2(n18986), .A3(n13068), .ZN(n17322) );
  INV_X1 U11684 ( .A(n14569), .ZN(n14565) );
  AND2_X1 U11685 ( .A1(n21011), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13013) );
  OAI22_X1 U11686 ( .A1(n12916), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12955), 
        .B2(n11254), .ZN(n14149) );
  NAND2_X1 U11687 ( .A1(n11285), .A2(n10187), .ZN(n13783) );
  AND2_X1 U11688 ( .A1(n11284), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11285) );
  NAND3_X1 U11689 ( .A1(n9892), .A2(n15306), .A3(n9890), .ZN(n15294) );
  NAND3_X1 U11690 ( .A1(n9891), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n10779), .ZN(n9890) );
  NAND2_X1 U11691 ( .A1(n9970), .A2(n15693), .ZN(n9969) );
  INV_X1 U11692 ( .A(n15712), .ZN(n9970) );
  NAND2_X1 U11693 ( .A1(n10969), .A2(n19927), .ZN(n11249) );
  OR2_X1 U11694 ( .A1(n19503), .A2(n20035), .ZN(n19730) );
  AOI21_X1 U11695 ( .B1(n16000), .B2(n18809), .A(n15911), .ZN(n16077) );
  OR2_X1 U11696 ( .A1(n20045), .A2(n10807), .ZN(n16435) );
  NAND2_X1 U11697 ( .A1(n10231), .A2(n10230), .ZN(n10955) );
  INV_X1 U11698 ( .A(n12013), .ZN(n12010) );
  AOI21_X1 U11699 ( .B1(n12088), .B2(n12114), .A(n12284), .ZN(n9947) );
  INV_X1 U11700 ( .A(n12095), .ZN(n9954) );
  NOR2_X1 U11701 ( .A1(n9941), .A2(n20257), .ZN(n9940) );
  INV_X1 U11702 ( .A(n11951), .ZN(n9941) );
  NAND2_X1 U11703 ( .A1(n12193), .A2(n11822), .ZN(n11880) );
  NAND2_X1 U11704 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11803) );
  OR2_X1 U11705 ( .A1(n11865), .A2(n11864), .ZN(n11960) );
  INV_X1 U11706 ( .A(n12167), .ZN(n12173) );
  INV_X1 U11707 ( .A(n15209), .ZN(n9997) );
  AND2_X1 U11708 ( .A1(n10630), .A2(n10615), .ZN(n10631) );
  NAND2_X1 U11709 ( .A1(n10230), .A2(n11013), .ZN(n10949) );
  AND2_X1 U11710 ( .A1(n11426), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10209) );
  NOR2_X1 U11711 ( .A1(n19033), .A2(n17579), .ZN(n13318) );
  NAND2_X1 U11712 ( .A1(n17572), .A2(n13125), .ZN(n13166) );
  INV_X1 U11713 ( .A(n17562), .ZN(n13353) );
  NOR2_X1 U11714 ( .A1(n13340), .A2(n13318), .ZN(n13346) );
  OAI22_X1 U11715 ( .A1(n13063), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18855), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U11716 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17332), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13251) );
  NAND2_X1 U11717 ( .A1(n12784), .A2(n10041), .ZN(n10040) );
  INV_X1 U11718 ( .A(n14643), .ZN(n10041) );
  NOR2_X1 U11719 ( .A1(n14657), .A2(n10044), .ZN(n10043) );
  INV_X1 U11720 ( .A(n14717), .ZN(n10044) );
  INV_X1 U11721 ( .A(n13009), .ZN(n12869) );
  NAND2_X1 U11722 ( .A1(n15048), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13009) );
  AND2_X1 U11723 ( .A1(n14432), .A2(n12609), .ZN(n14470) );
  INV_X1 U11724 ( .A(n14089), .ZN(n12457) );
  NAND2_X1 U11725 ( .A1(n9950), .A2(n9947), .ZN(n9945) );
  NAND2_X1 U11726 ( .A1(n9947), .A2(n9721), .ZN(n9944) );
  INV_X1 U11727 ( .A(n14407), .ZN(n10061) );
  INV_X1 U11728 ( .A(n14408), .ZN(n10062) );
  AND2_X1 U11729 ( .A1(n14216), .A2(n16349), .ZN(n10059) );
  NAND2_X1 U11730 ( .A1(n13683), .A2(n12293), .ZN(n12298) );
  OR2_X1 U11731 ( .A1(n11987), .A2(n11986), .ZN(n12016) );
  NAND2_X1 U11732 ( .A1(n12216), .A2(n12215), .ZN(n12220) );
  OR2_X1 U11733 ( .A1(n11878), .A2(n11877), .ZN(n11959) );
  NOR2_X1 U11734 ( .A1(n11933), .A2(n11932), .ZN(n11961) );
  XNOR2_X1 U11735 ( .A(n11953), .B(n11949), .ZN(n12415) );
  INV_X1 U11736 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13752) );
  OAI21_X1 U11737 ( .B1(n16059), .B2(n16379), .A(n15064), .ZN(n20242) );
  AOI21_X1 U11738 ( .B1(n10595), .B2(n10594), .A(n10593), .ZN(n10598) );
  NAND2_X1 U11739 ( .A1(n10776), .A2(n9894), .ZN(n10764) );
  AND2_X1 U11740 ( .A1(n15207), .A2(n16391), .ZN(n9894) );
  NAND2_X1 U11741 ( .A1(n10592), .A2(n10591), .ZN(n10610) );
  NAND2_X1 U11742 ( .A1(n11033), .A2(n10263), .ZN(n10592) );
  AND2_X1 U11743 ( .A1(n11429), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10801) );
  INV_X1 U11744 ( .A(n13783), .ZN(n11536) );
  INV_X1 U11745 ( .A(n14485), .ZN(n9976) );
  AOI22_X1 U11746 ( .A1(n11426), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10138) );
  NOR2_X1 U11747 ( .A1(n10257), .A2(n11013), .ZN(n10215) );
  INV_X1 U11748 ( .A(n10186), .ZN(n10080) );
  INV_X1 U11749 ( .A(n14239), .ZN(n10001) );
  OR2_X1 U11750 ( .A1(n19237), .A2(n19408), .ZN(n10905) );
  INV_X1 U11751 ( .A(n12932), .ZN(n9901) );
  AND2_X1 U11752 ( .A1(n15136), .A2(n11262), .ZN(n15356) );
  NAND2_X1 U11753 ( .A1(n9980), .A2(n15795), .ZN(n9979) );
  INV_X1 U11754 ( .A(n14264), .ZN(n9980) );
  NAND2_X1 U11755 ( .A1(n9844), .A2(n9843), .ZN(n9842) );
  NAND2_X1 U11756 ( .A1(n10636), .A2(n10615), .ZN(n10639) );
  INV_X1 U11757 ( .A(n14116), .ZN(n9964) );
  INV_X1 U11758 ( .A(n19425), .ZN(n10970) );
  NAND2_X1 U11759 ( .A1(n10237), .A2(n9727), .ZN(n9981) );
  NAND2_X1 U11760 ( .A1(n10328), .A2(n10348), .ZN(n10352) );
  AOI22_X1 U11761 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10221), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U11762 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10197) );
  AND4_X1 U11763 ( .A1(n10607), .A2(n10202), .A3(n10187), .A4(n19425), .ZN(
        n10243) );
  NAND2_X1 U11764 ( .A1(n18834), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13334) );
  INV_X1 U11765 ( .A(n17056), .ZN(n13068) );
  NAND2_X1 U11766 ( .A1(n17878), .A2(n18195), .ZN(n9917) );
  NOR2_X1 U11767 ( .A1(n17989), .A2(n13371), .ZN(n13374) );
  AND2_X1 U11768 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13360), .ZN(
        n13361) );
  XNOR2_X1 U11769 ( .A(n13166), .B(n13353), .ZN(n13168) );
  NAND2_X1 U11770 ( .A1(n16080), .A2(n17572), .ZN(n13355) );
  OAI22_X1 U11771 ( .A1(n13208), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18833), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13333) );
  CLKBUF_X1 U11772 ( .A(n12195), .Z(n12196) );
  OR2_X1 U11773 ( .A1(n21016), .A2(n14017), .ZN(n20116) );
  AND2_X1 U11774 ( .A1(n12224), .A2(n12223), .ZN(n13953) );
  NAND2_X1 U11775 ( .A1(n13825), .A2(n12433), .ZN(n13838) );
  NOR2_X1 U11776 ( .A1(n10046), .A2(n13044), .ZN(n10045) );
  INV_X1 U11777 ( .A(n12876), .ZN(n10046) );
  NOR2_X1 U11778 ( .A1(n12761), .A2(n16092), .ZN(n12762) );
  NAND2_X1 U11779 ( .A1(n12762), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12802) );
  NOR2_X1 U11780 ( .A1(n12710), .A2(n12709), .ZN(n12711) );
  NAND2_X1 U11781 ( .A1(n12711), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12761) );
  NAND2_X1 U11782 ( .A1(n14951), .A2(n9949), .ZN(n9948) );
  AND2_X1 U11783 ( .A1(n16069), .A2(n16063), .ZN(n9949) );
  CLKBUF_X1 U11784 ( .A(n14087), .Z(n14088) );
  AND2_X1 U11785 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12438), .ZN(
        n12444) );
  AOI21_X1 U11786 ( .B1(n12413), .B2(n12558), .A(n10037), .ZN(n10036) );
  INV_X1 U11787 ( .A(n12433), .ZN(n10037) );
  INV_X1 U11788 ( .A(n20057), .ZN(n14575) );
  NAND2_X1 U11789 ( .A1(n14597), .A2(n12307), .ZN(n13049) );
  NAND2_X1 U11790 ( .A1(n14649), .A2(n12367), .ZN(n14628) );
  AND3_X1 U11791 ( .A1(n12263), .A2(n12278), .A3(n12262), .ZN(n14374) );
  NAND2_X1 U11792 ( .A1(n14969), .A2(n14974), .ZN(n16338) );
  NAND2_X1 U11793 ( .A1(n9935), .A2(n9934), .ZN(n12084) );
  NAND2_X1 U11794 ( .A1(n10066), .A2(n10064), .ZN(n14090) );
  AND3_X1 U11795 ( .A1(n10063), .A2(n12234), .A3(n13962), .ZN(n10064) );
  INV_X1 U11796 ( .A(n13988), .ZN(n10066) );
  OR2_X1 U11797 ( .A1(n13988), .A2(n10065), .ZN(n13964) );
  NAND2_X1 U11798 ( .A1(n10063), .A2(n13962), .ZN(n10065) );
  XNOR2_X1 U11799 ( .A(n11906), .B(n13814), .ZN(n13912) );
  BUF_X1 U11800 ( .A(n12205), .Z(n14567) );
  NOR2_X1 U11801 ( .A1(n20566), .A2(n20412), .ZN(n20808) );
  NAND2_X1 U11802 ( .A1(n11887), .A2(n20242), .ZN(n20412) );
  AOI21_X1 U11803 ( .B1(n20759), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20412), 
        .ZN(n20859) );
  AND2_X1 U11804 ( .A1(n12182), .A2(n12181), .ZN(n14569) );
  NAND2_X1 U11805 ( .A1(n10926), .A2(n10932), .ZN(n11634) );
  AND2_X1 U11806 ( .A1(n10753), .A2(n10752), .ZN(n10755) );
  NAND2_X1 U11807 ( .A1(n10623), .A2(n10622), .ZN(n10728) );
  NOR2_X1 U11808 ( .A1(n10640), .A2(n10637), .ZN(n9881) );
  INV_X1 U11809 ( .A(n10641), .ZN(n9880) );
  NAND2_X1 U11810 ( .A1(n15151), .A2(n10008), .ZN(n15213) );
  AND2_X1 U11811 ( .A1(n10010), .A2(n10009), .ZN(n10008) );
  INV_X1 U11812 ( .A(n15215), .ZN(n10009) );
  NAND2_X1 U11813 ( .A1(n11311), .A2(n9988), .ZN(n13787) );
  NOR2_X1 U11814 ( .A1(n11313), .A2(n9989), .ZN(n9988) );
  INV_X1 U11815 ( .A(n11310), .ZN(n9989) );
  NAND2_X1 U11816 ( .A1(n9983), .A2(n11560), .ZN(n15186) );
  NAND2_X1 U11817 ( .A1(n15124), .A2(n11644), .ZN(n15275) );
  INV_X1 U11818 ( .A(n11495), .ZN(n9993) );
  AND2_X1 U11819 ( .A1(n11365), .A2(n9803), .ZN(n9999) );
  AND2_X1 U11820 ( .A1(n11364), .A2(n13967), .ZN(n11365) );
  INV_X1 U11821 ( .A(n20020), .ZN(n14275) );
  NAND2_X1 U11822 ( .A1(n11003), .A2(n9974), .ZN(n13604) );
  AOI21_X1 U11823 ( .B1(n11284), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n9975), .ZN(n9974) );
  OAI21_X1 U11824 ( .B1(n11013), .B2(n13499), .A(n20033), .ZN(n9975) );
  NAND2_X1 U11825 ( .A1(n12917), .A2(n9784), .ZN(n9909) );
  NAND2_X1 U11826 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9906) );
  NAND2_X1 U11827 ( .A1(n15409), .A2(n15386), .ZN(n15387) );
  INV_X1 U11828 ( .A(n15420), .ZN(n15386) );
  NOR2_X1 U11829 ( .A1(n12944), .A2(n19184), .ZN(n12943) );
  AND2_X1 U11830 ( .A1(n10900), .A2(n10012), .ZN(n10011) );
  INV_X1 U11831 ( .A(n10902), .ZN(n10012) );
  NOR2_X1 U11832 ( .A1(n15301), .A2(n10781), .ZN(n9958) );
  NAND2_X1 U11833 ( .A1(n15304), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15305) );
  NOR2_X1 U11834 ( .A1(n10788), .A2(n10768), .ZN(n15332) );
  NOR2_X1 U11835 ( .A1(n15434), .A2(n10075), .ZN(n10074) );
  INV_X1 U11836 ( .A(n15381), .ZN(n10075) );
  NAND2_X1 U11837 ( .A1(n10077), .A2(n10079), .ZN(n10076) );
  INV_X1 U11838 ( .A(n15444), .ZN(n10077) );
  NOR2_X1 U11839 ( .A1(n9969), .A2(n9967), .ZN(n9966) );
  INV_X1 U11840 ( .A(n15711), .ZN(n9968) );
  INV_X1 U11841 ( .A(n15679), .ZN(n9967) );
  NOR2_X1 U11842 ( .A1(n15475), .A2(n10070), .ZN(n10069) );
  INV_X1 U11843 ( .A(n10108), .ZN(n10070) );
  XNOR2_X1 U11844 ( .A(n15849), .B(n11292), .ZN(n13600) );
  XNOR2_X1 U11845 ( .A(n11297), .B(n11295), .ZN(n13666) );
  NAND2_X1 U11846 ( .A1(n14069), .A2(n11002), .ZN(n9838) );
  NAND2_X1 U11847 ( .A1(n14275), .A2(n14061), .ZN(n19550) );
  INV_X1 U11848 ( .A(n19851), .ZN(n19765) );
  OR2_X1 U11849 ( .A1(n19503), .A2(n19277), .ZN(n19690) );
  NAND2_X1 U11850 ( .A1(n10031), .A2(n10029), .ZN(n10033) );
  NOR2_X1 U11851 ( .A1(n17025), .A2(n10030), .ZN(n10029) );
  NAND2_X1 U11852 ( .A1(n16754), .A2(n10032), .ZN(n10031) );
  NOR2_X1 U11853 ( .A1(n17698), .A2(n17002), .ZN(n10030) );
  AND2_X1 U11854 ( .A1(n10033), .A2(n16542), .ZN(n16734) );
  OR2_X1 U11855 ( .A1(n17002), .A2(n17730), .ZN(n10027) );
  OR2_X1 U11856 ( .A1(n16773), .A2(n9829), .ZN(n10026) );
  OR2_X1 U11857 ( .A1(n16773), .A2(n16774), .ZN(n10028) );
  OR2_X1 U11858 ( .A1(n17002), .A2(n17761), .ZN(n10023) );
  OR2_X1 U11859 ( .A1(n16809), .A2(n10024), .ZN(n10022) );
  OR2_X1 U11860 ( .A1(n17778), .A2(n17761), .ZN(n10024) );
  OR2_X1 U11861 ( .A1(n16809), .A2(n17778), .ZN(n10025) );
  NAND2_X1 U11862 ( .A1(n19044), .A2(n17579), .ZN(n16702) );
  INV_X1 U11863 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17372) );
  INV_X1 U11864 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17313) );
  BUF_X1 U11865 ( .A(n13250), .Z(n17327) );
  NAND2_X1 U11866 ( .A1(n13286), .A2(n10099), .ZN(n13287) );
  NAND2_X1 U11867 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13286) );
  INV_X1 U11868 ( .A(n13100), .ZN(n9920) );
  AOI21_X1 U11869 ( .B1(n9765), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(n13117), .ZN(n13118) );
  NOR2_X1 U11870 ( .A1(n17373), .A2(n17416), .ZN(n13117) );
  AND2_X1 U11871 ( .A1(n16079), .A2(n18867), .ZN(n17427) );
  NAND2_X1 U11872 ( .A1(n9862), .A2(n9861), .ZN(n17641) );
  INV_X1 U11873 ( .A(n13332), .ZN(n9862) );
  NOR2_X1 U11874 ( .A1(n17779), .A2(n16709), .ZN(n17762) );
  AND2_X1 U11875 ( .A1(n17744), .A2(n10120), .ZN(n13194) );
  NAND2_X1 U11876 ( .A1(n17749), .A2(n17847), .ZN(n17744) );
  NAND2_X1 U11877 ( .A1(n13188), .A2(n13187), .ZN(n17839) );
  INV_X1 U11878 ( .A(n13186), .ZN(n13187) );
  OAI22_X1 U11879 ( .A1(n16563), .A2(n18182), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17847), .ZN(n13186) );
  XNOR2_X1 U11880 ( .A(n17572), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18045) );
  NAND2_X1 U11881 ( .A1(n13563), .A2(n13593), .ZN(n21016) );
  AND2_X1 U11882 ( .A1(n14038), .A2(n14031), .ZN(n20133) );
  AND2_X1 U11883 ( .A1(n14038), .A2(n14027), .ZN(n20127) );
  NAND2_X1 U11884 ( .A1(n20153), .A2(n13057), .ZN(n14727) );
  XNOR2_X1 U11885 ( .A(n12365), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14831) );
  NAND2_X1 U11886 ( .A1(n14788), .A2(n9933), .ZN(n9929) );
  AND2_X1 U11887 ( .A1(n15052), .A2(n12380), .ZN(n9933) );
  INV_X1 U11888 ( .A(n16341), .ZN(n16367) );
  INV_X1 U11889 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20998) );
  CLKBUF_X1 U11890 ( .A(n14100), .Z(n14101) );
  CLKBUF_X1 U11891 ( .A(n13860), .Z(n13861) );
  NOR2_X1 U11892 ( .A1(n9913), .A2(n19242), .ZN(n16386) );
  INV_X1 U11893 ( .A(n10337), .ZN(n10338) );
  AND2_X1 U11894 ( .A1(n19057), .A2(n12960), .ZN(n19273) );
  XNOR2_X1 U11895 ( .A(n10796), .B(n10795), .ZN(n15513) );
  INV_X1 U11896 ( .A(n15636), .ZN(n10084) );
  OAI211_X1 U11897 ( .C1(P2_STATE2_REG_0__SCAN_IN), .C2(n20034), .A(n16435), 
        .B(n16436), .ZN(n16428) );
  NAND2_X1 U11898 ( .A1(n19409), .A2(n13621), .ZN(n16455) );
  INV_X1 U11899 ( .A(n16435), .ZN(n19400) );
  INV_X1 U11900 ( .A(n16455), .ZN(n19398) );
  INV_X1 U11901 ( .A(n15509), .ZN(n19403) );
  XNOR2_X1 U11902 ( .A(n11265), .B(n11264), .ZN(n12912) );
  OR2_X1 U11903 ( .A1(n15575), .A2(n12903), .ZN(n15543) );
  NAND2_X1 U11904 ( .A1(n15406), .A2(n15405), .ZN(n15636) );
  OR2_X1 U11905 ( .A1(n15417), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15406) );
  OR2_X1 U11906 ( .A1(n11249), .A2(n11234), .ZN(n15834) );
  AND2_X1 U11907 ( .A1(n11250), .A2(n20044), .ZN(n16471) );
  OR2_X1 U11908 ( .A1(n15849), .A2(n13589), .ZN(n20035) );
  CLKBUF_X1 U11909 ( .A(n11002), .Z(n20033) );
  INV_X1 U11910 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20024) );
  INV_X1 U11911 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20017) );
  INV_X1 U11912 ( .A(n20004), .ZN(n20013) );
  OR2_X1 U11913 ( .A1(n16501), .A2(n20033), .ZN(n15882) );
  AND2_X1 U11914 ( .A1(n10804), .A2(n10803), .ZN(n20045) );
  NOR2_X1 U11915 ( .A1(n18811), .A2(n17640), .ZN(n19044) );
  AOI21_X1 U11916 ( .B1(n9858), .B2(n9855), .A(n18883), .ZN(n9854) );
  INV_X1 U11917 ( .A(n18809), .ZN(n9855) );
  INV_X1 U11918 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n21122) );
  NOR2_X1 U11919 ( .A1(n17520), .A2(n17694), .ZN(n17516) );
  NAND2_X1 U11920 ( .A1(n17554), .A2(P3_EAX_REG_7__SCAN_IN), .ZN(n17549) );
  AOI21_X1 U11921 ( .B1(n17914), .B2(n17002), .A(n16553), .ZN(n9860) );
  INV_X1 U11922 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18866) );
  OR2_X1 U11923 ( .A1(n11842), .A2(n13019), .ZN(n11821) );
  NAND2_X1 U11924 ( .A1(n11825), .A2(n11824), .ZN(n12199) );
  AND2_X1 U11925 ( .A1(n12189), .A2(n13019), .ZN(n11824) );
  NAND2_X1 U11926 ( .A1(n9868), .A2(n9710), .ZN(n10551) );
  OR2_X1 U11927 ( .A1(n13214), .A2(n13215), .ZN(n13210) );
  CLKBUF_X1 U11928 ( .A(n11724), .Z(n12714) );
  OR2_X1 U11929 ( .A1(n12059), .A2(n12058), .ZN(n12077) );
  NAND2_X1 U11930 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U11931 ( .A1(n12199), .A2(n12313), .ZN(n11846) );
  NOR2_X1 U11932 ( .A1(n12131), .A2(n12130), .ZN(n12172) );
  OR3_X1 U11933 ( .A1(n12164), .A2(n12163), .A3(n12162), .ZN(n12165) );
  NOR2_X1 U11934 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11428) );
  INV_X1 U11935 ( .A(n14501), .ZN(n9992) );
  AND4_X1 U11936 ( .A1(n10555), .A2(n10554), .A3(n10553), .A4(n10552), .ZN(
        n10566) );
  NOR2_X1 U11937 ( .A1(n9797), .A2(n9889), .ZN(n9888) );
  INV_X1 U11938 ( .A(n10565), .ZN(n9889) );
  NAND2_X1 U11939 ( .A1(n10546), .A2(n10547), .ZN(n10549) );
  OAI22_X1 U11940 ( .A1(n19478), .A2(n10513), .B1(n11420), .B2(n9847), .ZN(
        n10514) );
  NAND2_X1 U11941 ( .A1(n14069), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10346) );
  OR2_X1 U11942 ( .A1(n10305), .A2(n14164), .ZN(n10308) );
  AOI22_X1 U11943 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10219) );
  AND2_X1 U11944 ( .A1(n11791), .A2(n10121), .ZN(n12195) );
  NAND2_X1 U11945 ( .A1(n9806), .A2(n10050), .ZN(n10049) );
  OR2_X1 U11946 ( .A1(n12529), .A2(n14356), .ZN(n10050) );
  OR2_X1 U11947 ( .A1(n12088), .A2(n15017), .ZN(n14892) );
  NAND2_X1 U11948 ( .A1(n14357), .A2(n14356), .ZN(n14358) );
  NAND2_X1 U11949 ( .A1(n12490), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12494) );
  OAI21_X1 U11950 ( .B1(n9950), .B2(n9721), .A(n9947), .ZN(n12117) );
  NAND2_X1 U11951 ( .A1(n14710), .A2(n10051), .ZN(n10055) );
  AND2_X1 U11952 ( .A1(n10052), .A2(n9832), .ZN(n10051) );
  NOR2_X1 U11953 ( .A1(n14705), .A2(n10053), .ZN(n10052) );
  INV_X1 U11954 ( .A(n14709), .ZN(n10053) );
  NOR2_X1 U11955 ( .A1(n14965), .A2(n14866), .ZN(n12106) );
  INV_X1 U11956 ( .A(n9953), .ZN(n9952) );
  OR2_X1 U11957 ( .A1(n12094), .A2(n9954), .ZN(n9951) );
  OAI21_X1 U11958 ( .B1(n12093), .B2(n9954), .A(n12096), .ZN(n9953) );
  OR2_X1 U11959 ( .A1(n12088), .A2(n15030), .ZN(n12095) );
  OR2_X1 U11960 ( .A1(n14292), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12093) );
  INV_X1 U11961 ( .A(n11938), .ZN(n12085) );
  INV_X1 U11962 ( .A(n13989), .ZN(n10063) );
  NAND2_X1 U11963 ( .A1(n11950), .A2(n9940), .ZN(n11883) );
  NAND2_X1 U11964 ( .A1(n12195), .A2(n20257), .ZN(n12203) );
  NAND2_X1 U11965 ( .A1(n11835), .A2(n11834), .ZN(n11886) );
  INV_X1 U11966 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13867) );
  INV_X1 U11967 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11684) );
  INV_X1 U11968 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U11969 ( .A1(n13743), .A2(n11887), .ZN(n11989) );
  AND2_X1 U11970 ( .A1(n11972), .A2(n20910), .ZN(n20565) );
  NAND2_X1 U11971 ( .A1(n9927), .A2(n11832), .ZN(n9925) );
  NAND2_X1 U11972 ( .A1(n11741), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11778) );
  INV_X1 U11973 ( .A(n12211), .ZN(n11820) );
  INV_X1 U11974 ( .A(n13019), .ZN(n12206) );
  INV_X1 U11975 ( .A(n15035), .ZN(n15038) );
  NOR2_X1 U11976 ( .A1(n12167), .A2(n12141), .ZN(n12170) );
  NAND2_X1 U11977 ( .A1(n11977), .A2(n11976), .ZN(n12145) );
  AND2_X1 U11978 ( .A1(n12129), .A2(n12130), .ZN(n12142) );
  OR2_X1 U11979 ( .A1(n12131), .A2(n12128), .ZN(n12129) );
  NOR2_X1 U11980 ( .A1(n10730), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10748) );
  OR2_X2 U11981 ( .A1(n10710), .A2(n9807), .ZN(n10724) );
  NAND2_X1 U11982 ( .A1(n10688), .A2(n9896), .ZN(n10694) );
  AND2_X1 U11983 ( .A1(n13974), .A2(n19192), .ZN(n9896) );
  NAND2_X1 U11984 ( .A1(n9886), .A2(n9885), .ZN(n10666) );
  NAND2_X1 U11985 ( .A1(n10611), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U11986 ( .A1(n10615), .A2(n19435), .ZN(n9886) );
  AND2_X1 U11987 ( .A1(n11231), .A2(n15123), .ZN(n10010) );
  AND2_X1 U11988 ( .A1(n10004), .A2(n10003), .ZN(n10002) );
  INV_X1 U11989 ( .A(n14243), .ZN(n10003) );
  NAND2_X1 U11990 ( .A1(n9972), .A2(n15081), .ZN(n9971) );
  INV_X1 U11991 ( .A(n15097), .ZN(n9972) );
  CLKBUF_X1 U11992 ( .A(n10361), .Z(n11604) );
  AOI21_X1 U11993 ( .B1(n11472), .B2(n9997), .A(n9824), .ZN(n9996) );
  NAND2_X1 U11994 ( .A1(n15219), .A2(n9997), .ZN(n9995) );
  INV_X1 U11995 ( .A(n10926), .ZN(n10250) );
  BUF_X1 U11996 ( .A(n10248), .Z(n10941) );
  NOR2_X1 U11997 ( .A1(n15296), .A2(n9908), .ZN(n9907) );
  NOR2_X1 U11998 ( .A1(n15413), .A2(n9903), .ZN(n9902) );
  NAND2_X1 U11999 ( .A1(n12927), .A2(n9815), .ZN(n9898) );
  INV_X1 U12000 ( .A(n10583), .ZN(n11025) );
  INV_X1 U12001 ( .A(n14441), .ZN(n10862) );
  AND2_X1 U12002 ( .A1(n11217), .A2(n11216), .ZN(n14223) );
  AND2_X1 U12003 ( .A1(n10845), .A2(n10844), .ZN(n14044) );
  AND2_X1 U12004 ( .A1(n10838), .A2(n10837), .ZN(n13975) );
  NOR2_X1 U12005 ( .A1(n10543), .A2(n10542), .ZN(n11046) );
  NAND2_X1 U12006 ( .A1(n10631), .A2(n10635), .ZN(n10632) );
  AND2_X1 U12007 ( .A1(n10629), .A2(n19223), .ZN(n10633) );
  OR2_X1 U12008 ( .A1(n10390), .A2(n10389), .ZN(n11017) );
  NAND2_X1 U12009 ( .A1(n10316), .A2(n10304), .ZN(n10814) );
  NAND3_X1 U12010 ( .A1(n20004), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19851), 
        .ZN(n14001) );
  INV_X1 U12011 ( .A(n17698), .ZN(n10032) );
  NOR2_X2 U12012 ( .A1(n13208), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13064) );
  NAND2_X1 U12013 ( .A1(n13318), .A2(n16672), .ZN(n15998) );
  NAND2_X1 U12014 ( .A1(n17725), .A2(n9783), .ZN(n13350) );
  NAND2_X1 U12015 ( .A1(n17762), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17739) );
  INV_X1 U12016 ( .A(n16003), .ZN(n18844) );
  NAND2_X1 U12017 ( .A1(n18393), .A2(n18404), .ZN(n18822) );
  INV_X1 U12018 ( .A(n16001), .ZN(n16002) );
  OAI211_X1 U12019 ( .C1(n17322), .C2(n17416), .A(n13279), .B(n13278), .ZN(
        n13340) );
  NOR2_X1 U12020 ( .A1(n13254), .A2(n13253), .ZN(n13255) );
  NAND2_X1 U12021 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  NAND2_X1 U12022 ( .A1(n13265), .A2(n13264), .ZN(n13266) );
  AOI21_X1 U12023 ( .B1(n9765), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(n13263), .ZN(n13264) );
  NOR2_X1 U12024 ( .A1(n17327), .A2(n17259), .ZN(n13263) );
  INV_X1 U12025 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16159) );
  INV_X1 U12026 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20083) );
  AND2_X1 U12027 ( .A1(n14720), .A2(n14658), .ZN(n14710) );
  AND2_X1 U12028 ( .A1(n12257), .A2(n12256), .ZN(n14445) );
  AOI21_X1 U12029 ( .B1(n12443), .B2(n12582), .A(n12442), .ZN(n13961) );
  CLKBUF_X1 U12030 ( .A(n13933), .Z(n13934) );
  NAND2_X1 U12031 ( .A1(n12399), .A2(n12582), .ZN(n12408) );
  INV_X1 U12032 ( .A(n20239), .ZN(n20237) );
  AND3_X1 U12033 ( .A1(n13650), .A2(n13649), .A3(n14565), .ZN(n20154) );
  AND2_X1 U12034 ( .A1(n12982), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14018) );
  AND2_X1 U12035 ( .A1(n14814), .A2(n12872), .ZN(n12829) );
  AND2_X1 U12036 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n12803), .ZN(
        n12804) );
  NAND2_X1 U12037 ( .A1(n10039), .A2(n14620), .ZN(n10038) );
  INV_X1 U12038 ( .A(n10040), .ZN(n10039) );
  INV_X1 U12039 ( .A(n14832), .ZN(n12362) );
  OR2_X1 U12040 ( .A1(n12764), .A2(n12763), .ZN(n14643) );
  CLKBUF_X1 U12041 ( .A(n14641), .Z(n14693) );
  AND2_X1 U12042 ( .A1(n12713), .A2(n12712), .ZN(n14756) );
  AND2_X1 U12043 ( .A1(n12694), .A2(n12693), .ZN(n14699) );
  NOR2_X1 U12044 ( .A1(n12674), .A2(n14855), .ZN(n12675) );
  AND2_X1 U12045 ( .A1(n10043), .A2(n12678), .ZN(n10042) );
  NAND2_X1 U12046 ( .A1(n12641), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12674) );
  NOR2_X1 U12047 ( .A1(n21087), .A2(n12622), .ZN(n12641) );
  NOR2_X1 U12048 ( .A1(n12605), .A2(n12604), .ZN(n12606) );
  NAND2_X1 U12049 ( .A1(n12606), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12622) );
  CLKBUF_X1 U12050 ( .A(n14470), .Z(n14471) );
  NAND2_X1 U12051 ( .A1(n12573), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12605) );
  INV_X1 U12052 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12604) );
  NOR2_X1 U12053 ( .A1(n12559), .A2(n14413), .ZN(n12573) );
  OR2_X1 U12054 ( .A1(n12553), .A2(n16159), .ZN(n12559) );
  CLKBUF_X1 U12055 ( .A(n14367), .Z(n14368) );
  AND2_X1 U12056 ( .A1(n12513), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12514) );
  NOR2_X1 U12057 ( .A1(n12494), .A2(n20083), .ZN(n12513) );
  AND4_X1 U12058 ( .A1(n12479), .A2(n12478), .A3(n12477), .A4(n12476), .ZN(
        n14213) );
  AND2_X1 U12059 ( .A1(n12459), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12490) );
  AOI21_X1 U12060 ( .B1(n12456), .B2(n12582), .A(n12455), .ZN(n14089) );
  AND2_X1 U12061 ( .A1(n12444), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12449) );
  INV_X1 U12062 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12400) );
  INV_X1 U12063 ( .A(n13822), .ZN(n10035) );
  INV_X1 U12064 ( .A(n13683), .ZN(n14572) );
  INV_X1 U12065 ( .A(n9932), .ZN(n9931) );
  OAI21_X1 U12066 ( .B1(n10093), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n9932) );
  NOR2_X1 U12067 ( .A1(n9721), .A2(n12382), .ZN(n12383) );
  NOR2_X1 U12068 ( .A1(n14609), .A2(n14595), .ZN(n14597) );
  NAND2_X1 U12069 ( .A1(n10068), .A2(n10067), .ZN(n14609) );
  INV_X1 U12070 ( .A(n14611), .ZN(n10067) );
  AND2_X1 U12071 ( .A1(n9944), .A2(n9943), .ZN(n9942) );
  INV_X1 U12072 ( .A(n14797), .ZN(n9943) );
  NOR2_X1 U12073 ( .A1(n10055), .A2(n10054), .ZN(n14649) );
  INV_X1 U12074 ( .A(n14651), .ZN(n10054) );
  NAND2_X1 U12075 ( .A1(n14710), .A2(n10052), .ZN(n16096) );
  NOR2_X1 U12076 ( .A1(n9786), .A2(n14719), .ZN(n14720) );
  NAND2_X1 U12077 ( .A1(n14475), .A2(n14474), .ZN(n14725) );
  XNOR2_X1 U12078 ( .A(n12088), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14967) );
  INV_X1 U12079 ( .A(n12104), .ZN(n14965) );
  OR2_X1 U12080 ( .A1(n12088), .A2(n12102), .ZN(n14881) );
  AND2_X1 U12081 ( .A1(n16212), .A2(n12101), .ZN(n14879) );
  NAND2_X1 U12082 ( .A1(n10062), .A2(n9816), .ZN(n14436) );
  INV_X1 U12083 ( .A(n14374), .ZN(n10060) );
  NAND2_X1 U12084 ( .A1(n10062), .A2(n10061), .ZN(n14410) );
  OR2_X1 U12085 ( .A1(n12088), .A2(n15002), .ZN(n16212) );
  NOR2_X1 U12086 ( .A1(n12337), .A2(n13913), .ZN(n15016) );
  INV_X1 U12087 ( .A(n16338), .ZN(n12337) );
  NAND2_X1 U12088 ( .A1(n14361), .A2(n14362), .ZN(n14408) );
  CLKBUF_X1 U12089 ( .A(n14865), .Z(n14903) );
  NAND2_X1 U12090 ( .A1(n16350), .A2(n9813), .ZN(n14399) );
  INV_X1 U12091 ( .A(n14396), .ZN(n10056) );
  NAND2_X1 U12092 ( .A1(n16350), .A2(n10059), .ZN(n14397) );
  NAND2_X1 U12093 ( .A1(n9955), .A2(n12093), .ZN(n14378) );
  OR2_X1 U12094 ( .A1(n14294), .A2(n12094), .ZN(n9955) );
  NAND2_X1 U12095 ( .A1(n9937), .A2(n16242), .ZN(n9936) );
  INV_X1 U12096 ( .A(n12048), .ZN(n9937) );
  INV_X1 U12097 ( .A(n16242), .ZN(n9939) );
  AND2_X1 U12098 ( .A1(n12243), .A2(n12242), .ZN(n16349) );
  NOR2_X1 U12099 ( .A1(n10058), .A2(n10057), .ZN(n16352) );
  INV_X1 U12100 ( .A(n16349), .ZN(n10057) );
  INV_X1 U12101 ( .A(n16350), .ZN(n10058) );
  AND2_X1 U12102 ( .A1(n12238), .A2(n12237), .ZN(n14091) );
  NOR2_X1 U12103 ( .A1(n14090), .A2(n14091), .ZN(n16350) );
  NAND2_X1 U12104 ( .A1(n12226), .A2(n12225), .ZN(n13988) );
  INV_X1 U12105 ( .A(n13954), .ZN(n12226) );
  NOR2_X1 U12106 ( .A1(n13988), .A2(n13989), .ZN(n13987) );
  AOI21_X1 U12107 ( .B1(n15036), .B2(n12081), .A(n11966), .ZN(n13947) );
  AND2_X2 U12108 ( .A1(n12211), .A2(n20243), .ZN(n13683) );
  NOR2_X1 U12109 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13818), .ZN(
        n13913) );
  OR2_X1 U12110 ( .A1(n12331), .A2(n13751), .ZN(n16333) );
  OR2_X1 U12111 ( .A1(n12331), .A2(n12327), .ZN(n14974) );
  OR2_X1 U12112 ( .A1(n12331), .A2(n13868), .ZN(n14969) );
  NAND2_X1 U12113 ( .A1(n11905), .A2(n11904), .ZN(n13815) );
  OR2_X1 U12114 ( .A1(n12423), .A2(n12141), .ZN(n11905) );
  CLKBUF_X1 U12115 ( .A(n12203), .Z(n12204) );
  NAND2_X1 U12116 ( .A1(n12300), .A2(n12293), .ZN(n13804) );
  OR2_X1 U12117 ( .A1(n11953), .A2(n11952), .ZN(n11954) );
  NAND2_X1 U12118 ( .A1(n11950), .A2(n11951), .ZN(n12417) );
  CLKBUF_X1 U12119 ( .A(n12986), .Z(n12813) );
  AND2_X1 U12120 ( .A1(n13774), .A2(n13773), .ZN(n13879) );
  NOR2_X1 U12121 ( .A1(n20370), .A2(n13889), .ZN(n20306) );
  OR2_X1 U12122 ( .A1(n12414), .A2(n15035), .ZN(n20532) );
  INV_X1 U12123 ( .A(n20637), .ZN(n20691) );
  AND2_X1 U12124 ( .A1(n20857), .A2(n20721), .ZN(n20758) );
  CLKBUF_X1 U12125 ( .A(n12206), .Z(n20270) );
  AND2_X1 U12126 ( .A1(n13889), .A2(n20757), .ZN(n20690) );
  NAND3_X1 U12128 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n11887), .A3(n20242), 
        .ZN(n20281) );
  AND2_X1 U12129 ( .A1(n14021), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16054) );
  NAND2_X1 U12130 ( .A1(n10600), .A2(n10599), .ZN(n10937) );
  NOR2_X1 U12131 ( .A1(n10783), .A2(n10782), .ZN(n10791) );
  INV_X1 U12132 ( .A(n10764), .ZN(n10770) );
  OR2_X1 U12133 ( .A1(n10663), .A2(n10611), .ZN(n10774) );
  NOR2_X1 U12134 ( .A1(n16402), .A2(n16403), .ZN(n16401) );
  NAND2_X1 U12135 ( .A1(n14330), .A2(n10102), .ZN(n15166) );
  AND2_X1 U12136 ( .A1(n14330), .A2(n9825), .ZN(n14486) );
  NAND2_X1 U12137 ( .A1(n10623), .A2(n9893), .ZN(n10730) );
  NOR2_X1 U12138 ( .A1(n10720), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n9893) );
  AND2_X1 U12139 ( .A1(n10704), .A2(n10709), .ZN(n19143) );
  AND2_X1 U12140 ( .A1(n10714), .A2(n10713), .ZN(n10716) );
  NAND2_X1 U12141 ( .A1(n10627), .A2(n9884), .ZN(n10663) );
  NOR2_X1 U12142 ( .A1(n10628), .A2(n10666), .ZN(n9884) );
  OR2_X1 U12143 ( .A1(n9883), .A2(n9882), .ZN(n10651) );
  INV_X1 U12144 ( .A(n10652), .ZN(n9883) );
  MUX2_X1 U12145 ( .A(n10608), .B(n14154), .S(n10611), .Z(n10649) );
  AND2_X1 U12146 ( .A1(n10858), .A2(n10857), .ZN(n14258) );
  NAND2_X1 U12147 ( .A1(n13969), .A2(n10002), .ZN(n14245) );
  AND3_X1 U12148 ( .A1(n11174), .A2(n11173), .A3(n11172), .ZN(n14249) );
  INV_X1 U12149 ( .A(n13979), .ZN(n10000) );
  NOR2_X1 U12150 ( .A1(n15098), .A2(n15097), .ZN(n15099) );
  INV_X1 U12151 ( .A(n11560), .ZN(n9984) );
  XNOR2_X1 U12152 ( .A(n11539), .B(n11540), .ZN(n15198) );
  XNOR2_X1 U12153 ( .A(n9998), .B(n11517), .ZN(n15206) );
  NAND2_X1 U12154 ( .A1(n15206), .A2(n15205), .ZN(n15204) );
  NAND2_X1 U12155 ( .A1(n14330), .A2(n9827), .ZN(n15127) );
  NAND2_X1 U12156 ( .A1(n10145), .A2(n10144), .ZN(n10146) );
  AND3_X1 U12157 ( .A1(n11195), .A2(n11194), .A3(n11193), .ZN(n15712) );
  INV_X1 U12158 ( .A(n10231), .ZN(n11639) );
  NAND2_X1 U12159 ( .A1(n12951), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12952) );
  AND2_X1 U12160 ( .A1(n10874), .A2(n10873), .ZN(n15149) );
  AND2_X1 U12161 ( .A1(n12927), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12948) );
  NAND2_X1 U12162 ( .A1(n12927), .A2(n9777), .ZN(n12949) );
  OR2_X1 U12163 ( .A1(n10906), .A2(n19209), .ZN(n10907) );
  NAND2_X1 U12164 ( .A1(n13894), .A2(n9799), .ZN(n13976) );
  INV_X1 U12165 ( .A(n9834), .ZN(n10007) );
  NAND2_X1 U12166 ( .A1(n13894), .A2(n9789), .ZN(n13920) );
  NOR2_X1 U12167 ( .A1(n10905), .A2(n19235), .ZN(n9900) );
  AND2_X1 U12168 ( .A1(n13894), .A2(n13930), .ZN(n13928) );
  NAND2_X1 U12169 ( .A1(n9901), .A2(n9899), .ZN(n12936) );
  INV_X1 U12170 ( .A(n10905), .ZN(n9899) );
  AND2_X1 U12171 ( .A1(n10820), .A2(n10819), .ZN(n13810) );
  OR3_X1 U12172 ( .A1(n12975), .A2(n10615), .A3(n15519), .ZN(n11256) );
  AND2_X1 U12173 ( .A1(n12901), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9957) );
  NAND2_X1 U12174 ( .A1(n15785), .A2(n12901), .ZN(n15350) );
  AND2_X1 U12175 ( .A1(n15177), .A2(n10736), .ZN(n15389) );
  NAND2_X1 U12176 ( .A1(n10073), .A2(n10072), .ZN(n10078) );
  AOI21_X1 U12177 ( .B1(n15445), .B2(n10074), .A(n15384), .ZN(n10072) );
  NAND2_X1 U12178 ( .A1(n15444), .A2(n10074), .ZN(n10073) );
  NAND2_X1 U12179 ( .A1(n9978), .A2(n15763), .ZN(n9977) );
  INV_X1 U12180 ( .A(n9979), .ZN(n9978) );
  NAND2_X1 U12181 ( .A1(n15785), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15784) );
  OR2_X1 U12182 ( .A1(n9711), .A2(n15485), .ZN(n15790) );
  NOR2_X1 U12183 ( .A1(n9867), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9866) );
  INV_X1 U12184 ( .A(n19238), .ZN(n9867) );
  NAND2_X1 U12185 ( .A1(n10547), .A2(n9840), .ZN(n9839) );
  NAND2_X1 U12186 ( .A1(n9965), .A2(n9963), .ZN(n9962) );
  AND2_X1 U12187 ( .A1(n14110), .A2(n9964), .ZN(n9963) );
  CLKBUF_X1 U12188 ( .A(n9735), .Z(n10997) );
  NOR2_X1 U12189 ( .A1(n11031), .A2(n9961), .ZN(n9960) );
  INV_X1 U12190 ( .A(n14110), .ZN(n9961) );
  NAND2_X1 U12191 ( .A1(n9853), .A2(n10468), .ZN(n14171) );
  OR2_X1 U12192 ( .A1(n11249), .A2(n10983), .ZN(n15667) );
  NOR2_X1 U12193 ( .A1(n10275), .A2(n12955), .ZN(n10276) );
  AOI21_X1 U12194 ( .B1(n11288), .B2(n11299), .A(n11287), .ZN(n13599) );
  NOR2_X1 U12195 ( .A1(n10961), .A2(n10938), .ZN(n16501) );
  NOR2_X1 U12196 ( .A1(n10937), .A2(n13571), .ZN(n10938) );
  CLKBUF_X1 U12197 ( .A(n10953), .Z(n10954) );
  NAND2_X1 U12198 ( .A1(n19503), .A2(n20035), .ZN(n19574) );
  NAND2_X1 U12199 ( .A1(n10208), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9850) );
  NAND2_X1 U12200 ( .A1(n10214), .A2(n15872), .ZN(n9851) );
  NAND2_X1 U12201 ( .A1(n10131), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10132) );
  NAND2_X1 U12202 ( .A1(n10192), .A2(n15872), .ZN(n10200) );
  NAND2_X1 U12203 ( .A1(n10177), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10185) );
  INV_X1 U12204 ( .A(n14010), .ZN(n19434) );
  NOR2_X2 U12205 ( .A1(n14002), .A2(n14001), .ZN(n19433) );
  NOR2_X2 U12206 ( .A1(n15276), .A2(n14001), .ZN(n19432) );
  NAND2_X1 U12207 ( .A1(n14275), .A2(n20026), .ZN(n19846) );
  AOI21_X1 U12208 ( .B1(n13337), .B2(n13336), .A(n13335), .ZN(n18812) );
  NOR2_X1 U12209 ( .A1(n16697), .A2(n16696), .ZN(n18811) );
  INV_X1 U12210 ( .A(n9858), .ZN(n9857) );
  NAND2_X1 U12211 ( .A1(n13425), .A2(n18813), .ZN(n9858) );
  NOR2_X1 U12212 ( .A1(n13350), .A2(n21104), .ZN(n13391) );
  NAND2_X1 U12213 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17197), .ZN(n17183) );
  NOR2_X1 U12214 ( .A1(n17432), .A2(n17435), .ZN(n18829) );
  OAI211_X1 U12215 ( .C1(n17327), .C2(n17372), .A(n13312), .B(n13311), .ZN(
        n17579) );
  AOI22_X1 U12216 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13312) );
  AOI211_X1 U12217 ( .C1(n17377), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n13310), .B(n13309), .ZN(n13311) );
  INV_X1 U12218 ( .A(n17636), .ZN(n17580) );
  AOI21_X1 U12219 ( .B1(n15998), .B2(n18869), .A(n19031), .ZN(n17578) );
  INV_X1 U12220 ( .A(n17641), .ZN(n17639) );
  INV_X1 U12221 ( .A(n17640), .ZN(n17638) );
  NOR2_X1 U12222 ( .A1(n17710), .A2(n10020), .ZN(n10019) );
  NAND2_X1 U12223 ( .A1(n17725), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17709) );
  NOR2_X1 U12224 ( .A1(n17739), .A2(n17740), .ZN(n17725) );
  NOR2_X1 U12225 ( .A1(n13397), .A2(n17862), .ZN(n17724) );
  NAND2_X1 U12226 ( .A1(n17836), .A2(n9778), .ZN(n17779) );
  NOR2_X1 U12227 ( .A1(n17814), .A2(n10017), .ZN(n10016) );
  NAND2_X1 U12228 ( .A1(n17836), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17812) );
  NOR2_X1 U12229 ( .A1(n17974), .A2(n16888), .ZN(n17892) );
  NAND2_X1 U12230 ( .A1(n17972), .A2(n13184), .ZN(n13185) );
  NOR2_X1 U12231 ( .A1(n10015), .A2(n17995), .ZN(n10014) );
  NOR2_X1 U12232 ( .A1(n17029), .A2(n18039), .ZN(n18018) );
  NAND2_X1 U12233 ( .A1(n17715), .A2(n9782), .ZN(n13203) );
  NOR2_X1 U12234 ( .A1(n16551), .A2(n18063), .ZN(n16534) );
  NOR2_X1 U12235 ( .A1(n13178), .A2(n17552), .ZN(n16566) );
  NAND2_X1 U12236 ( .A1(n9775), .A2(n9922), .ZN(n13195) );
  NAND2_X1 U12237 ( .A1(n17743), .A2(n9922), .ZN(n18064) );
  NOR2_X1 U12238 ( .A1(n9863), .A2(n9922), .ZN(n9875) );
  INV_X1 U12239 ( .A(n18065), .ZN(n9874) );
  NOR2_X1 U12240 ( .A1(n18097), .A2(n18082), .ZN(n17743) );
  NAND2_X1 U12241 ( .A1(n17869), .A2(n13381), .ZN(n18097) );
  NOR2_X1 U12242 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17795), .ZN(
        n17783) );
  OAI21_X1 U12243 ( .B1(n18821), .B2(n18844), .A(n18820), .ZN(n18828) );
  AND2_X1 U12244 ( .A1(n9878), .A2(n9877), .ZN(n17869) );
  INV_X1 U12245 ( .A(n18163), .ZN(n9877) );
  INV_X1 U12246 ( .A(n18828), .ZN(n18843) );
  NOR2_X1 U12247 ( .A1(n13376), .A2(n9879), .ZN(n17967) );
  AND2_X1 U12248 ( .A1(n13377), .A2(n13378), .ZN(n9879) );
  NOR2_X1 U12249 ( .A1(n17967), .A2(n9918), .ZN(n17966) );
  NAND2_X1 U12250 ( .A1(n13374), .A2(n13375), .ZN(n17978) );
  XNOR2_X1 U12251 ( .A(n13370), .B(n13369), .ZN(n17990) );
  NOR2_X1 U12252 ( .A1(n17990), .A2(n18297), .ZN(n17989) );
  NOR2_X1 U12253 ( .A1(n18012), .A2(n13364), .ZN(n17999) );
  XNOR2_X1 U12254 ( .A(n13363), .B(n18313), .ZN(n18013) );
  NOR2_X1 U12255 ( .A1(n18013), .A2(n18014), .ZN(n18012) );
  XNOR2_X1 U12256 ( .A(n13168), .B(n13167), .ZN(n18027) );
  NOR2_X1 U12257 ( .A1(n13359), .A2(n18333), .ZN(n18024) );
  NOR2_X1 U12258 ( .A1(n13413), .A2(n13408), .ZN(n13425) );
  XNOR2_X1 U12259 ( .A(n13355), .B(n13125), .ZN(n13358) );
  AOI211_X2 U12260 ( .C1(n13221), .C2(n13220), .A(n13337), .B(n13335), .ZN(
        n18809) );
  OAI211_X1 U12261 ( .C1(n17229), .C2(n17313), .A(n13302), .B(n13301), .ZN(
        n18389) );
  AOI211_X1 U12262 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n13300), .B(n13299), .ZN(n13301) );
  INV_X1 U12263 ( .A(n13341), .ZN(n18393) );
  AOI211_X1 U12264 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n13241), .B(n13240), .ZN(n13242) );
  NAND2_X1 U12265 ( .A1(n18871), .A2(n18377), .ZN(n18620) );
  AOI21_X1 U12266 ( .B1(n18808), .B2(n18809), .A(n9857), .ZN(n18817) );
  OR2_X1 U12267 ( .A1(n13560), .A2(n14569), .ZN(n13593) );
  AND2_X1 U12268 ( .A1(n14573), .A2(n12217), .ZN(n13566) );
  INV_X1 U12269 ( .A(n20099), .ZN(n16182) );
  AND2_X1 U12270 ( .A1(n20116), .A2(n14032), .ZN(n20131) );
  INV_X1 U12271 ( .A(n20131), .ZN(n16178) );
  NAND2_X1 U12272 ( .A1(n14038), .A2(n14037), .ZN(n20118) );
  INV_X1 U12273 ( .A(n20133), .ZN(n20095) );
  INV_X1 U12274 ( .A(n14727), .ZN(n20148) );
  INV_X1 U12275 ( .A(n14771), .ZN(n14782) );
  OR2_X1 U12276 ( .A1(n14767), .A2(n13821), .ZN(n14439) );
  NOR2_X1 U12277 ( .A1(n20154), .A2(n21019), .ZN(n20163) );
  BUF_X1 U12278 ( .A(n20163), .Z(n20177) );
  CLKBUF_X1 U12279 ( .A(n13850), .Z(n21019) );
  NAND2_X1 U12280 ( .A1(n9946), .A2(n12088), .ZN(n16190) );
  NAND2_X1 U12281 ( .A1(n9950), .A2(n12339), .ZN(n9946) );
  INV_X1 U12282 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n21087) );
  NOR2_X1 U12283 ( .A1(n14231), .A2(n14230), .ZN(n20145) );
  AND2_X1 U12284 ( .A1(n14212), .A2(n14122), .ZN(n20150) );
  OR2_X1 U12285 ( .A1(n20230), .A2(n12882), .ZN(n16256) );
  INV_X1 U12286 ( .A(n16256), .ZN(n20228) );
  NAND2_X1 U12287 ( .A1(n12049), .A2(n12048), .ZN(n16244) );
  INV_X1 U12288 ( .A(n16333), .ZN(n13958) );
  INV_X1 U12289 ( .A(n14969), .ZN(n13818) );
  INV_X1 U12290 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20759) );
  INV_X1 U12292 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20562) );
  OR2_X1 U12293 ( .A1(n13888), .A2(n13887), .ZN(n20996) );
  NOR2_X1 U12294 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15060) );
  INV_X1 U12295 ( .A(n20513), .ZN(n20510) );
  OAI22_X1 U12296 ( .A1(n20490), .A2(n20489), .B1(n20488), .B2(n20729), .ZN(
        n20517) );
  OAI22_X1 U12297 ( .A1(n20649), .A2(n20648), .B1(n20647), .B2(n20795), .ZN(
        n20672) );
  INV_X1 U12298 ( .A(n20645), .ZN(n20673) );
  INV_X1 U12299 ( .A(n20767), .ZN(n20791) );
  NOR2_X1 U12300 ( .A1(n20250), .A2(n20412), .ZN(n20800) );
  NOR2_X1 U12301 ( .A1(n20263), .A2(n20412), .ZN(n20819) );
  NOR2_X1 U12302 ( .A1(n20277), .A2(n20412), .ZN(n20833) );
  OAI211_X1 U12303 ( .C1(n20841), .C2(n20809), .A(n20808), .B(n20807), .ZN(
        n20845) );
  INV_X1 U12304 ( .A(n20810), .ZN(n20844) );
  INV_X1 U12305 ( .A(n20800), .ZN(n20854) );
  INV_X1 U12306 ( .A(n20827), .ZN(n20884) );
  INV_X1 U12307 ( .A(n20833), .ZN(n20891) );
  INV_X1 U12308 ( .A(n20906), .ZN(n20914) );
  NOR2_X1 U12309 ( .A1(n20726), .A2(n14569), .ZN(n16058) );
  INV_X1 U12310 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21011) );
  NAND2_X1 U12311 ( .A1(n11261), .A2(n10766), .ZN(n16395) );
  NAND2_X1 U12312 ( .A1(n10776), .A2(n15207), .ZN(n10765) );
  NOR2_X1 U12313 ( .A1(n19242), .A2(n15365), .ZN(n9914) );
  NOR2_X1 U12314 ( .A1(n16401), .A2(n19242), .ZN(n15117) );
  NOR2_X1 U12315 ( .A1(n15144), .A2(n19242), .ZN(n15133) );
  OAI21_X1 U12316 ( .B1(n15156), .B2(n9911), .A(n9910), .ZN(n15144) );
  NAND2_X1 U12317 ( .A1(n12349), .A2(n9912), .ZN(n9911) );
  NAND2_X1 U12318 ( .A1(n19242), .A2(n12349), .ZN(n9910) );
  INV_X1 U12319 ( .A(n15394), .ZN(n9912) );
  NOR2_X1 U12320 ( .A1(n19242), .A2(n15170), .ZN(n15156) );
  NOR2_X1 U12321 ( .A1(n15156), .A2(n15394), .ZN(n15155) );
  CLKBUF_X1 U12322 ( .A(n14149), .Z(n19226) );
  AND2_X1 U12323 ( .A1(n19057), .A2(n16517), .ZN(n19266) );
  OR2_X1 U12324 ( .A1(n19057), .A2(n12964), .ZN(n19222) );
  OR3_X1 U12325 ( .A1(n13463), .A2(n12970), .A3(n12969), .ZN(n19252) );
  INV_X1 U12326 ( .A(n19222), .ZN(n19265) );
  OR2_X1 U12327 ( .A1(n14046), .A2(n14045), .ZN(n14248) );
  OR2_X1 U12328 ( .A1(n11130), .A2(n11129), .ZN(n13967) );
  NAND2_X1 U12329 ( .A1(n11318), .A2(n11317), .ZN(n13978) );
  INV_X1 U12330 ( .A(n20026), .ZN(n14061) );
  INV_X1 U12331 ( .A(n11289), .ZN(n10348) );
  OR2_X1 U12332 ( .A1(n13900), .A2(n11676), .ZN(n15242) );
  NOR2_X1 U12333 ( .A1(n15219), .A2(n11472), .ZN(n15210) );
  INV_X1 U12334 ( .A(n19290), .ZN(n19284) );
  INV_X1 U12335 ( .A(n15284), .ZN(n19289) );
  AND2_X1 U12336 ( .A1(n13603), .A2(n14002), .ZN(n19291) );
  AND2_X1 U12337 ( .A1(n11638), .A2(n19927), .ZN(n19322) );
  OR2_X1 U12338 ( .A1(n13547), .A2(n11637), .ZN(n11638) );
  AND2_X1 U12339 ( .A1(n19297), .A2(n19324), .ZN(n19330) );
  NAND2_X1 U12340 ( .A1(n19322), .A2(n11639), .ZN(n19324) );
  NAND2_X1 U12341 ( .A1(n11311), .A2(n11310), .ZN(n13789) );
  OR2_X1 U12342 ( .A1(n13603), .A2(n19289), .ZN(n19314) );
  INV_X1 U12343 ( .A(n20035), .ZN(n19277) );
  AND2_X1 U12344 ( .A1(n19322), .A2(n11676), .ZN(n19339) );
  INV_X1 U12345 ( .A(n19322), .ZN(n19338) );
  INV_X1 U12346 ( .A(n19314), .ZN(n19347) );
  INV_X2 U12347 ( .A(n19357), .ZN(n19382) );
  AND2_X1 U12348 ( .A1(n13568), .A2(n13540), .ZN(n19394) );
  INV_X1 U12349 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19235) );
  OR2_X1 U12350 ( .A1(n15691), .A2(n11241), .ZN(n15639) );
  NAND2_X1 U12351 ( .A1(n10076), .A2(n15381), .ZN(n15433) );
  NOR2_X1 U12352 ( .A1(n15711), .A2(n9969), .ZN(n15678) );
  NAND2_X1 U12353 ( .A1(n10071), .A2(n10108), .ZN(n15474) );
  NAND2_X1 U12354 ( .A1(n11238), .A2(n15823), .ZN(n16463) );
  INV_X1 U12355 ( .A(n16476), .ZN(n16461) );
  OR2_X1 U12356 ( .A1(n11249), .A2(n16505), .ZN(n13627) );
  INV_X1 U12357 ( .A(n16482), .ZN(n15832) );
  AND2_X1 U12358 ( .A1(n13627), .A2(n15667), .ZN(n16482) );
  INV_X1 U12359 ( .A(n15834), .ZN(n16479) );
  INV_X1 U12360 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16493) );
  NAND2_X1 U12361 ( .A1(n11289), .A2(n11299), .ZN(n11291) );
  NAND2_X1 U12362 ( .A1(n13598), .A2(n13601), .ZN(n20026) );
  OR2_X1 U12363 ( .A1(n13600), .A2(n13599), .ZN(n13601) );
  NAND2_X1 U12364 ( .A1(n13664), .A2(n13667), .ZN(n20020) );
  INV_X1 U12365 ( .A(n19524), .ZN(n19533) );
  OAI21_X1 U12366 ( .B1(n15889), .B2(n15893), .A(n15888), .ZN(n19546) );
  OR2_X1 U12367 ( .A1(n19574), .A2(n19550), .ZN(n19563) );
  NOR2_X1 U12368 ( .A1(n19609), .A2(n19550), .ZN(n19599) );
  NAND2_X1 U12369 ( .A1(n19648), .A2(n19647), .ZN(n19666) );
  INV_X1 U12370 ( .A(n19663), .ZN(n19665) );
  NAND2_X1 U12371 ( .A1(n9838), .A2(n14064), .ZN(n14065) );
  INV_X1 U12372 ( .A(n19723), .ZN(n19714) );
  OAI21_X1 U12373 ( .B1(n19701), .B2(n19700), .A(n19699), .ZN(n19719) );
  INV_X1 U12374 ( .A(n9846), .ZN(n19696) );
  OAI21_X1 U12375 ( .B1(n19698), .B2(n19763), .A(n11002), .ZN(n9846) );
  OAI21_X1 U12376 ( .B1(n19785), .B2(n20033), .A(n19769), .ZN(n19788) );
  NOR2_X1 U12377 ( .A1(n19690), .A2(n19550), .ZN(n19807) );
  INV_X1 U12378 ( .A(n19866), .ZN(n19811) );
  AND2_X1 U12379 ( .A1(n11284), .A2(n19434), .ZN(n19859) );
  INV_X1 U12380 ( .A(n21353), .ZN(n19815) );
  AND2_X1 U12381 ( .A1(n19434), .A2(n10230), .ZN(n19882) );
  AND2_X1 U12382 ( .A1(n19435), .A2(n19434), .ZN(n19891) );
  OAI21_X1 U12383 ( .B1(n14278), .B2(n14281), .A(n14277), .ZN(n19833) );
  AND2_X1 U12384 ( .A1(n11013), .A2(n19434), .ZN(n19908) );
  INV_X1 U12385 ( .A(n19733), .ZN(n19854) );
  INV_X1 U12386 ( .A(n19736), .ZN(n19863) );
  INV_X1 U12387 ( .A(n19802), .ZN(n19877) );
  INV_X1 U12388 ( .A(n19744), .ZN(n19886) );
  INV_X1 U12389 ( .A(n19747), .ZN(n19895) );
  INV_X1 U12390 ( .A(n19751), .ZN(n19903) );
  NOR2_X2 U12391 ( .A1(n19690), .A2(n19846), .ZN(n19915) );
  NAND2_X1 U12392 ( .A1(n18867), .A2(n18812), .ZN(n17640) );
  INV_X1 U12393 ( .A(n10033), .ZN(n16735) );
  NOR2_X1 U12394 ( .A1(n16747), .A2(n17698), .ZN(n16746) );
  NOR2_X1 U12395 ( .A1(n16754), .A2(n17025), .ZN(n16747) );
  NAND2_X1 U12396 ( .A1(n10026), .A2(n10027), .ZN(n16766) );
  NAND2_X1 U12397 ( .A1(n10022), .A2(n10023), .ZN(n16792) );
  AND2_X1 U12398 ( .A1(n10025), .A2(n17002), .ZN(n16793) );
  NOR2_X1 U12399 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16935), .ZN(n16915) );
  NOR2_X1 U12400 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16942), .ZN(n16941) );
  NOR2_X2 U12401 ( .A1(n18983), .A2(n17058), .ZN(n17038) );
  INV_X1 U12402 ( .A(n17038), .ZN(n17059) );
  NOR2_X2 U12403 ( .A1(n18868), .A2(n16702), .ZN(n17051) );
  INV_X1 U12404 ( .A(n17051), .ZN(n17070) );
  OAI211_X1 U12405 ( .C1(n18871), .C2(n18872), .A(n16698), .B(n19046), .ZN(
        n17073) );
  NAND2_X1 U12406 ( .A1(n17258), .A2(P3_EBX_REG_14__SCAN_IN), .ZN(n17242) );
  NOR2_X1 U12407 ( .A1(n16912), .A2(n17289), .ZN(n17258) );
  NAND2_X1 U12408 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17310), .ZN(n17289) );
  INV_X1 U12409 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17390) );
  INV_X1 U12410 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17405) );
  NAND2_X1 U12411 ( .A1(n17424), .A2(n10107), .ZN(n17401) );
  INV_X1 U12412 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17407) );
  NOR2_X1 U12413 ( .A1(n17585), .A2(n17453), .ZN(n17446) );
  NAND2_X1 U12414 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17457), .ZN(n17453) );
  NAND2_X1 U12415 ( .A1(n17466), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17462) );
  NOR2_X1 U12416 ( .A1(n17603), .A2(n17505), .ZN(n17500) );
  OR3_X1 U12417 ( .A1(n17478), .A2(n17512), .A3(n17645), .ZN(n17505) );
  NAND2_X1 U12418 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17516), .ZN(n17512) );
  INV_X1 U12419 ( .A(n17480), .ZN(n17510) );
  INV_X1 U12420 ( .A(n17504), .ZN(n17511) );
  NAND2_X1 U12421 ( .A1(n17543), .A2(n17430), .ZN(n17520) );
  NOR2_X1 U12422 ( .A1(n13288), .A2(n13287), .ZN(n13289) );
  NAND4_X1 U12423 ( .A1(n13078), .A2(n13077), .A3(n13076), .A4(n13075), .ZN(
        n17548) );
  NAND2_X1 U12424 ( .A1(n17427), .A2(n10092), .ZN(n17429) );
  NOR2_X1 U12425 ( .A1(n9921), .A2(n9920), .ZN(n9919) );
  NOR2_X1 U12426 ( .A1(n13089), .A2(n21200), .ZN(n9921) );
  AND2_X1 U12427 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n13122) );
  NAND2_X1 U12428 ( .A1(n18829), .A2(n17427), .ZN(n17568) );
  NAND2_X1 U12429 ( .A1(n17427), .A2(n17478), .ZN(n17565) );
  INV_X1 U12430 ( .A(n17574), .ZN(n17571) );
  NAND2_X1 U12431 ( .A1(n17367), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13110) );
  INV_X1 U12432 ( .A(n17568), .ZN(n17573) );
  NOR2_X1 U12433 ( .A1(n17565), .A2(n18829), .ZN(n17574) );
  NOR2_X1 U12434 ( .A1(n19030), .A2(n17580), .ZN(n17628) );
  OAI211_X1 U12436 ( .C1(n19034), .C2(n19033), .A(n17639), .B(n17638), .ZN(
        n17659) );
  NOR3_X1 U12437 ( .A1(n17642), .A2(n17641), .A3(n17640), .ZN(n17673) );
  CLKBUF_X1 U12438 ( .A(n17673), .Z(n17684) );
  NOR2_X1 U12440 ( .A1(n17690), .A2(n19033), .ZN(n17691) );
  NOR2_X1 U12441 ( .A1(n17850), .A2(n17856), .ZN(n17836) );
  INV_X1 U12442 ( .A(n18693), .ZN(n18753) );
  INV_X1 U12443 ( .A(n17833), .ZN(n17862) );
  INV_X1 U12444 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17896) );
  NAND2_X1 U12445 ( .A1(n9772), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17974) );
  NAND2_X1 U12446 ( .A1(n10013), .A2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17996) );
  NOR2_X1 U12447 ( .A1(n18039), .A2(n10015), .ZN(n10013) );
  NAND2_X1 U12448 ( .A1(n18721), .A2(n15997), .ZN(n18693) );
  NAND2_X1 U12449 ( .A1(n16680), .A2(n9833), .ZN(n18054) );
  INV_X1 U12450 ( .A(n18270), .ZN(n16011) );
  NAND2_X1 U12451 ( .A1(n17715), .A2(n13199), .ZN(n16015) );
  INV_X1 U12452 ( .A(n17705), .ZN(n16577) );
  AOI21_X1 U12453 ( .B1(n18064), .B2(n18808), .A(n9872), .ZN(n18076) );
  NAND2_X1 U12454 ( .A1(n9876), .A2(n9873), .ZN(n9872) );
  NOR3_X1 U12455 ( .A1(n18084), .A2(n9875), .A3(n9874), .ZN(n9873) );
  NAND2_X1 U12456 ( .A1(n18063), .A2(n18191), .ZN(n9876) );
  NAND2_X1 U12457 ( .A1(n9863), .A2(n18267), .ZN(n18270) );
  INV_X1 U12458 ( .A(n18252), .ZN(n18237) );
  INV_X1 U12459 ( .A(n18263), .ZN(n18279) );
  XNOR2_X1 U12460 ( .A(n13358), .B(n18341), .ZN(n18334) );
  NOR2_X1 U12461 ( .A1(n18335), .A2(n18334), .ZN(n18333) );
  INV_X1 U12462 ( .A(n18357), .ZN(n18351) );
  INV_X1 U12463 ( .A(n18317), .ZN(n18355) );
  INV_X1 U12464 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18833) );
  INV_X1 U12465 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18855) );
  INV_X1 U12466 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18859) );
  AOI211_X1 U12467 ( .C1(n18852), .C2(n18867), .A(n16007), .B(n18378), .ZN(
        n19015) );
  INV_X1 U12468 ( .A(n19015), .ZN(n19012) );
  INV_X1 U12470 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18983) );
  AND2_X1 U12472 ( .A1(n13034), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20239)
         );
  NAND2_X1 U12474 ( .A1(n14576), .A2(n20099), .ZN(n14583) );
  OAI22_X1 U12475 ( .A1(n14913), .A2(n14727), .B1(n13058), .B2(n20153), .ZN(
        n13059) );
  AOI21_X1 U12476 ( .B1(n12396), .B2(n16367), .A(n12395), .ZN(n12397) );
  AOI21_X1 U12477 ( .B1(n14556), .B2(n16367), .A(n12343), .ZN(n12344) );
  NAND2_X1 U12478 ( .A1(n12366), .A2(n16360), .ZN(n12378) );
  OR2_X1 U12479 ( .A1(n14525), .A2(n19230), .ZN(n9959) );
  NAND2_X1 U12480 ( .A1(n9916), .A2(n19246), .ZN(n9915) );
  OAI211_X1 U12481 ( .C1(n12915), .C2(n16436), .A(n9870), .B(n9869), .ZN(
        P2_U2983) );
  NAND2_X1 U12482 ( .A1(n12912), .A2(n19400), .ZN(n9869) );
  OAI211_X1 U12483 ( .C1(n15513), .C2(n16435), .A(n9895), .B(n10912), .ZN(
        P2_U2984) );
  NAND2_X1 U12484 ( .A1(n15536), .A2(n19404), .ZN(n15302) );
  OAI211_X1 U12485 ( .C1(n15625), .C2(n16435), .A(n10085), .B(n10083), .ZN(
        P2_U2994) );
  AOI21_X1 U12486 ( .B1(n15628), .B2(n19403), .A(n15407), .ZN(n10085) );
  NAND2_X1 U12487 ( .A1(n10084), .A2(n19404), .ZN(n10083) );
  OR2_X1 U12488 ( .A1(n14525), .A2(n15834), .ZN(n12914) );
  OAI211_X1 U12489 ( .C1(n15834), .C2(n15524), .A(n15523), .B(n10089), .ZN(
        n15525) );
  AOI21_X1 U12490 ( .B1(n13352), .B2(n16723), .A(n9859), .ZN(n13386) );
  INV_X1 U12491 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12934) );
  AND3_X1 U12492 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10014), .A3(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n9772) );
  NAND2_X1 U12493 ( .A1(n14305), .A2(n10626), .ZN(n9773) );
  NAND2_X1 U12494 ( .A1(n12922), .A2(n9779), .ZN(n12920) );
  INV_X1 U12495 ( .A(n10626), .ZN(n10630) );
  NAND2_X1 U12496 ( .A1(n14482), .A2(n14484), .ZN(n14483) );
  AND2_X1 U12497 ( .A1(n14495), .A2(n10043), .ZN(n14656) );
  NAND2_X1 U12498 ( .A1(n13969), .A2(n13970), .ZN(n13968) );
  AND2_X1 U12499 ( .A1(n10022), .A2(n9814), .ZN(n9774) );
  AND2_X1 U12500 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12935) );
  AND2_X1 U12501 ( .A1(n14257), .A2(n9804), .ZN(n14384) );
  AND2_X1 U12502 ( .A1(n15151), .A2(n11231), .ZN(n11230) );
  AND3_X1 U12503 ( .A1(n17825), .A2(n13417), .A3(n17749), .ZN(n9775) );
  AND2_X1 U12504 ( .A1(n10026), .A2(n9812), .ZN(n9776) );
  INV_X1 U12505 ( .A(n10424), .ZN(n11177) );
  NAND2_X1 U12506 ( .A1(n12917), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12953) );
  NAND2_X1 U12507 ( .A1(n12922), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12921) );
  AND2_X1 U12508 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U12509 ( .A1(n13787), .A2(n11316), .ZN(n13854) );
  AND2_X1 U12510 ( .A1(n10016), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9778) );
  AND2_X1 U12511 ( .A1(n9902), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9779) );
  AND2_X1 U12512 ( .A1(n9830), .A2(n9990), .ZN(n9780) );
  NAND2_X1 U12513 ( .A1(n13969), .A2(n10004), .ZN(n10006) );
  OR3_X1 U12514 ( .A1(n12348), .A2(n15371), .A3(n9905), .ZN(n9781) );
  AND2_X1 U12515 ( .A1(n13199), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9782) );
  AND2_X1 U12516 ( .A1(n10019), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9783) );
  AND2_X1 U12517 ( .A1(n9907), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9784) );
  INV_X1 U12518 ( .A(n9863), .ZN(n18061) );
  OR2_X1 U12519 ( .A1(n17056), .A2(n13061), .ZN(n9785) );
  INV_X1 U12520 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19921) );
  OR2_X1 U12521 ( .A1(n14725), .A2(n14724), .ZN(n9786) );
  AND2_X1 U12522 ( .A1(n10081), .A2(n11288), .ZN(n10475) );
  NOR2_X1 U12523 ( .A1(n14641), .A2(n14643), .ZN(n14632) );
  AND2_X1 U12524 ( .A1(n14495), .A2(n10042), .ZN(n14700) );
  INV_X1 U12525 ( .A(n9994), .ZN(n11471) );
  NAND2_X1 U12526 ( .A1(n14378), .A2(n12095), .ZN(n14902) );
  NOR2_X1 U12527 ( .A1(n14641), .A2(n10040), .ZN(n14618) );
  AND4_X1 U12528 ( .A1(n11738), .A2(n11737), .A3(n11736), .A4(n11735), .ZN(
        n9788) );
  INV_X1 U12529 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12933) );
  INV_X1 U12530 ( .A(n10453), .ZN(n11178) );
  AND2_X1 U12531 ( .A1(n13921), .A2(n13930), .ZN(n9789) );
  NAND2_X1 U12532 ( .A1(n11853), .A2(n11887), .ZN(n11950) );
  NAND4_X1 U12533 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n9790) );
  NAND2_X2 U12534 ( .A1(n13068), .A2(n13067), .ZN(n13089) );
  AND2_X1 U12535 ( .A1(n14700), .A2(n14699), .ZN(n14701) );
  NAND2_X1 U12536 ( .A1(n9871), .A2(n14451), .ZN(n15500) );
  NAND2_X2 U12537 ( .A1(n10316), .A2(n10321), .ZN(n11277) );
  INV_X1 U12538 ( .A(n9878), .ZN(n18245) );
  OR2_X1 U12539 ( .A1(n17966), .A2(n13379), .ZN(n9878) );
  AND2_X1 U12540 ( .A1(n10636), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14305) );
  AND2_X1 U12541 ( .A1(n14470), .A2(n14496), .ZN(n14495) );
  XNOR2_X1 U12542 ( .A(n11886), .B(n11885), .ZN(n12425) );
  NAND2_X1 U12543 ( .A1(n13664), .A2(n11298), .ZN(n13737) );
  AND2_X2 U12544 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10370) );
  AND2_X1 U12545 ( .A1(n16236), .A2(n16235), .ZN(n9791) );
  AND2_X1 U12546 ( .A1(n13418), .A2(n17724), .ZN(n9792) );
  OR2_X1 U12547 ( .A1(n10334), .A2(n10333), .ZN(n10516) );
  AND4_X1 U12548 ( .A1(n13109), .A2(n13108), .A3(n13107), .A4(n10096), .ZN(
        n9793) );
  AND2_X1 U12549 ( .A1(n13184), .A2(n9918), .ZN(n9794) );
  INV_X1 U12550 ( .A(n10548), .ZN(n9845) );
  OR2_X1 U12551 ( .A1(n15098), .A2(n9971), .ZN(n9795) );
  AND2_X1 U12552 ( .A1(n10528), .A2(n10527), .ZN(n9796) );
  NOR2_X1 U12553 ( .A1(n15213), .A2(n15109), .ZN(n15110) );
  NAND4_X1 U12554 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n9797) );
  INV_X1 U12555 ( .A(n18818), .ZN(n18832) );
  NAND2_X1 U12556 ( .A1(n16003), .A2(n16001), .ZN(n18818) );
  AND2_X1 U12557 ( .A1(n9986), .A2(n9984), .ZN(n9798) );
  AND2_X1 U12558 ( .A1(n9789), .A2(n10007), .ZN(n9799) );
  AND2_X1 U12559 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9800) );
  AND2_X1 U12560 ( .A1(n10604), .A2(n10160), .ZN(n9801) );
  BUF_X1 U12561 ( .A(n11746), .Z(n11927) );
  NAND2_X1 U12562 ( .A1(n15204), .A2(n11519), .ZN(n11539) );
  INV_X1 U12563 ( .A(n14305), .ZN(n10547) );
  INV_X1 U12564 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18039) );
  AND2_X1 U12565 ( .A1(n10548), .A2(n9762), .ZN(n9802) );
  INV_X1 U12566 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9982) );
  INV_X2 U12567 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18986) );
  NAND2_X1 U12568 ( .A1(n11819), .A2(n12211), .ZN(n12217) );
  XNOR2_X2 U12569 ( .A(n12417), .B(n12416), .ZN(n13889) );
  NOR2_X1 U12570 ( .A1(n15711), .A2(n15712), .ZN(n15692) );
  NAND2_X1 U12571 ( .A1(n15765), .A2(n15750), .ZN(n15736) );
  AND2_X1 U12572 ( .A1(n12943), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12927) );
  NAND2_X1 U12573 ( .A1(n15151), .A2(n10010), .ZN(n15122) );
  NOR2_X1 U12574 ( .A1(n15233), .A2(n15234), .ZN(n14482) );
  AND2_X1 U12575 ( .A1(n9901), .A2(n9900), .ZN(n12931) );
  NAND2_X1 U12576 ( .A1(n14710), .A2(n14709), .ZN(n14704) );
  NOR2_X1 U12577 ( .A1(n12925), .A2(n21218), .ZN(n12922) );
  NAND2_X1 U12578 ( .A1(n14495), .A2(n14717), .ZN(n14655) );
  NOR2_X1 U12579 ( .A1(n14121), .A2(n14213), .ZN(n14126) );
  AND3_X1 U12580 ( .A1(n9880), .A2(n9881), .A3(n10652), .ZN(n10627) );
  AND2_X1 U12581 ( .A1(n11317), .A2(n10000), .ZN(n9803) );
  AND2_X1 U12582 ( .A1(n10862), .A2(n14386), .ZN(n9804) );
  NAND2_X1 U12583 ( .A1(n9968), .A2(n9966), .ZN(n14222) );
  AND2_X1 U12584 ( .A1(n11318), .A2(n9803), .ZN(n9805) );
  AND2_X1 U12585 ( .A1(n9936), .A2(n16241), .ZN(n9938) );
  AND2_X1 U12586 ( .A1(n12931), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12930) );
  AND2_X1 U12587 ( .A1(n14359), .A2(n14404), .ZN(n9806) );
  INV_X1 U12588 ( .A(n17847), .ZN(n17958) );
  NAND2_X1 U12589 ( .A1(n17548), .A2(n16566), .ZN(n17847) );
  NOR2_X1 U12590 ( .A1(n19435), .A2(n14261), .ZN(n9807) );
  AND2_X1 U12591 ( .A1(n10619), .A2(n10713), .ZN(n9808) );
  NOR2_X1 U12592 ( .A1(n14205), .A2(n14258), .ZN(n14257) );
  NAND2_X1 U12593 ( .A1(n12347), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12348) );
  INV_X1 U12594 ( .A(n18267), .ZN(n18851) );
  NAND2_X1 U12595 ( .A1(n16000), .A2(n19047), .ZN(n18267) );
  AND2_X1 U12596 ( .A1(n12036), .A2(n12064), .ZN(n9809) );
  NOR2_X1 U12597 ( .A1(n15210), .A2(n15209), .ZN(n9810) );
  INV_X1 U12598 ( .A(n10068), .ZN(n14627) );
  NOR2_X1 U12599 ( .A1(n14628), .A2(n14629), .ZN(n10068) );
  AND2_X1 U12600 ( .A1(n9804), .A2(n15239), .ZN(n9811) );
  AND2_X1 U12601 ( .A1(n10027), .A2(n17002), .ZN(n9812) );
  AND2_X1 U12602 ( .A1(n10059), .A2(n10056), .ZN(n9813) );
  AND2_X1 U12603 ( .A1(n10023), .A2(n17002), .ZN(n9814) );
  AND2_X1 U12604 ( .A1(n9777), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9815) );
  AND2_X1 U12605 ( .A1(n10061), .A2(n10060), .ZN(n9816) );
  INV_X1 U12606 ( .A(n15445), .ZN(n10079) );
  INV_X1 U12607 ( .A(n9882), .ZN(n10653) );
  OR2_X1 U12608 ( .A1(n10641), .A2(n10640), .ZN(n9882) );
  OR2_X1 U12609 ( .A1(n10466), .A2(n10465), .ZN(n11038) );
  AND2_X1 U12610 ( .A1(n14257), .A2(n10862), .ZN(n14385) );
  NAND2_X1 U12611 ( .A1(n14257), .A2(n9811), .ZN(n15161) );
  AOI211_X1 U12612 ( .C1(n16402), .C2(n19226), .A(n9914), .B(n15346), .ZN(
        n9913) );
  AND2_X1 U12613 ( .A1(n12922), .A2(n9902), .ZN(n9817) );
  AND2_X1 U12614 ( .A1(n13192), .A2(n13191), .ZN(n9818) );
  AND2_X1 U12615 ( .A1(n15110), .A2(n15199), .ZN(n15201) );
  AND2_X1 U12616 ( .A1(n10002), .A2(n10001), .ZN(n9819) );
  AND2_X1 U12617 ( .A1(n10028), .A2(n17002), .ZN(n9820) );
  OR2_X1 U12618 ( .A1(n20286), .A2(n21011), .ZN(n9821) );
  NOR2_X1 U12619 ( .A1(n16352), .A2(n16351), .ZN(n9822) );
  NOR2_X1 U12620 ( .A1(n12952), .A2(n15322), .ZN(n12917) );
  NOR2_X1 U12621 ( .A1(n12348), .A2(n15371), .ZN(n12919) );
  AND2_X1 U12622 ( .A1(n13808), .A2(n13895), .ZN(n13894) );
  NAND2_X1 U12623 ( .A1(n13632), .A2(n9960), .ZN(n14112) );
  NOR2_X1 U12624 ( .A1(n14262), .A2(n14264), .ZN(n14263) );
  INV_X1 U12625 ( .A(n10522), .ZN(n19641) );
  AND2_X1 U12626 ( .A1(n11318), .A2(n9999), .ZN(n9823) );
  NOR2_X1 U12627 ( .A1(n14262), .A2(n9979), .ZN(n15762) );
  AND2_X1 U12628 ( .A1(n11495), .A2(n11494), .ZN(n9824) );
  NAND2_X1 U12629 ( .A1(n14341), .A2(n11048), .ZN(n14458) );
  AND2_X1 U12630 ( .A1(n9976), .A2(n10102), .ZN(n9825) );
  AND2_X1 U12631 ( .A1(n14446), .A2(n14445), .ZN(n14361) );
  XNOR2_X1 U12632 ( .A(n9909), .B(n11267), .ZN(n12916) );
  NOR2_X1 U12633 ( .A1(n13631), .A2(n9962), .ZN(n14340) );
  AND2_X1 U12634 ( .A1(n9794), .A2(n17972), .ZN(n17957) );
  NOR2_X1 U12635 ( .A1(n15155), .A2(n19242), .ZN(n9826) );
  AND2_X1 U12636 ( .A1(n9825), .A2(n11228), .ZN(n9827) );
  AND2_X1 U12637 ( .A1(n12742), .A2(n12741), .ZN(n9828) );
  OR2_X1 U12638 ( .A1(n17730), .A2(n16774), .ZN(n9829) );
  AND2_X1 U12639 ( .A1(n9992), .A2(n14484), .ZN(n9830) );
  AND2_X1 U12640 ( .A1(n12917), .A2(n9907), .ZN(n9831) );
  AND2_X1 U12641 ( .A1(n14694), .A2(n16095), .ZN(n9832) );
  INV_X1 U12642 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10020) );
  INV_X1 U12643 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n9918) );
  NAND2_X1 U12644 ( .A1(n20049), .A2(n10606), .ZN(n16436) );
  OR2_X1 U12645 ( .A1(n19028), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n9833) );
  AND2_X2 U12646 ( .A1(n15855), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14321) );
  AND2_X1 U12647 ( .A1(n10835), .A2(n10834), .ZN(n9834) );
  INV_X1 U12648 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9897) );
  INV_X1 U12649 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9903) );
  INV_X1 U12650 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9905) );
  INV_X1 U12651 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10017) );
  INV_X1 U12652 ( .A(n19246), .ZN(n19928) );
  INV_X1 U12653 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9908) );
  NAND3_X2 U12654 ( .A1(n15855), .A2(n9982), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10178) );
  AND2_X1 U12655 ( .A1(n17836), .A2(n10016), .ZN(n9835) );
  INV_X1 U12656 ( .A(n13396), .ZN(n9922) );
  AND2_X1 U12657 ( .A1(n17725), .A2(n10019), .ZN(n9836) );
  AND2_X1 U12658 ( .A1(n10781), .A2(n15542), .ZN(n9837) );
  INV_X1 U12659 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10015) );
  INV_X1 U12660 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10021) );
  INV_X1 U12661 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9904) );
  INV_X1 U12662 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19763) );
  NAND2_X2 U12663 ( .A1(n19045), .A2(n18871), .ZN(n18358) );
  AOI22_X2 U12664 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20288), .B1(DATAI_21_), 
        .B2(n20240), .ZN(n20897) );
  AOI22_X2 U12665 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20288), .B1(DATAI_26_), 
        .B2(n20240), .ZN(n20739) );
  AOI22_X2 U12666 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20288), .B1(DATAI_28_), 
        .B2(n20240), .ZN(n20890) );
  AOI22_X2 U12667 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20288), .B1(DATAI_31_), 
        .B2(n20240), .ZN(n20919) );
  AOI22_X2 U12668 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20288), .B1(DATAI_27_), 
        .B2(n20240), .ZN(n20883) );
  NOR2_X4 U12669 ( .A1(n21022), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20980) );
  NOR2_X2 U12670 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18983), .ZN(n18747) );
  AND2_X2 U12671 ( .A1(n13739), .A2(n9712), .ZN(n14069) );
  NAND2_X1 U12672 ( .A1(n9761), .A2(n9762), .ZN(n10546) );
  NOR2_X1 U12673 ( .A1(n9762), .A2(n10548), .ZN(n9840) );
  NAND2_X1 U12674 ( .A1(n9764), .A2(n9802), .ZN(n9841) );
  NOR2_X1 U12675 ( .A1(n14305), .A2(n10548), .ZN(n9843) );
  INV_X1 U12676 ( .A(n9764), .ZN(n9844) );
  INV_X1 U12677 ( .A(n19698), .ZN(n9847) );
  INV_X4 U12678 ( .A(n11004), .ZN(n11007) );
  NAND2_X1 U12679 ( .A1(n10227), .A2(n10144), .ZN(n9848) );
  NAND2_X1 U12680 ( .A1(n10220), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9849) );
  NAND2_X2 U12681 ( .A1(n10441), .A2(n10442), .ZN(n10468) );
  NAND2_X1 U12682 ( .A1(n10086), .A2(n10443), .ZN(n9853) );
  OAI211_X1 U12683 ( .C1(n13392), .C2(n16723), .A(n13385), .B(n9860), .ZN(
        n9859) );
  NOR2_X1 U12684 ( .A1(n18379), .A2(n18398), .ZN(n9861) );
  NOR2_X2 U12685 ( .A1(n9864), .A2(n11288), .ZN(n10522) );
  NAND2_X1 U12686 ( .A1(n9865), .A2(n10785), .ZN(n9892) );
  XNOR2_X2 U12687 ( .A(n9868), .B(n9755), .ZN(n10636) );
  NAND3_X2 U12688 ( .A1(n10441), .A2(n11038), .A3(n10442), .ZN(n10635) );
  NAND2_X1 U12689 ( .A1(n15484), .A2(n10691), .ZN(n10071) );
  INV_X2 U12690 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19014) );
  NAND2_X2 U12691 ( .A1(n17044), .A2(n9800), .ZN(n17373) );
  INV_X1 U12692 ( .A(n15307), .ZN(n9891) );
  NOR2_X2 U12693 ( .A1(n10686), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10688) );
  INV_X1 U12694 ( .A(n9898), .ZN(n12924) );
  OAI21_X1 U12695 ( .B1(n14527), .B2(n9915), .A(n12980), .ZN(P2_U2825) );
  NAND2_X1 U12696 ( .A1(n12957), .A2(n12956), .ZN(n9916) );
  NOR2_X1 U12697 ( .A1(n12957), .A2(n12956), .ZN(n14527) );
  NOR2_X2 U12698 ( .A1(n17870), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17878) );
  NAND3_X1 U12699 ( .A1(n9794), .A2(n17847), .A3(n17972), .ZN(n17944) );
  NAND2_X2 U12700 ( .A1(n17973), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17972) );
  INV_X1 U12701 ( .A(n17794), .ZN(n9923) );
  NAND3_X1 U12702 ( .A1(n13192), .A2(n13191), .A3(n18082), .ZN(n17749) );
  NAND2_X2 U12703 ( .A1(n13064), .A2(n13065), .ZN(n15914) );
  NAND3_X1 U12704 ( .A1(n9928), .A2(n11833), .A3(n9926), .ZN(n9924) );
  INV_X1 U12705 ( .A(n11912), .ZN(n9927) );
  OAI211_X1 U12706 ( .C1(n12379), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12385), .B(n9931), .ZN(n9930) );
  OAI211_X1 U12707 ( .C1(n12385), .C2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n9930), .B(n9929), .ZN(n14515) );
  NAND2_X1 U12708 ( .A1(n12049), .A2(n9938), .ZN(n9935) );
  OAI21_X1 U12709 ( .B1(n12049), .B2(n9939), .A(n9938), .ZN(n16238) );
  NAND3_X1 U12710 ( .A1(n9945), .A2(n16191), .A3(n9944), .ZN(n12358) );
  NAND3_X1 U12711 ( .A1(n9945), .A2(n9942), .A3(n16191), .ZN(n12115) );
  NAND2_X1 U12712 ( .A1(n9956), .A2(n19425), .ZN(n10234) );
  NAND2_X1 U12713 ( .A1(n11284), .A2(n9734), .ZN(n15843) );
  OAI21_X1 U12714 ( .B1(n10961), .B2(n9736), .A(n10230), .ZN(n10962) );
  NAND3_X1 U12715 ( .A1(n14533), .A2(n14534), .A3(n9959), .ZN(P2_U2824) );
  NOR2_X1 U12716 ( .A1(n11031), .A2(n13631), .ZN(n14111) );
  NOR2_X1 U12717 ( .A1(n13630), .A2(n13629), .ZN(n13631) );
  INV_X1 U12718 ( .A(n11031), .ZN(n9965) );
  NOR2_X2 U12719 ( .A1(n14222), .A2(n14223), .ZN(n15651) );
  INV_X1 U12720 ( .A(n9973), .ZN(n12893) );
  NOR2_X2 U12721 ( .A1(n15127), .A2(n15126), .ZN(n15124) );
  NOR2_X2 U12722 ( .A1(n14262), .A2(n9977), .ZN(n15765) );
  NAND3_X1 U12723 ( .A1(n10246), .A2(n9722), .A3(n9981), .ZN(n10975) );
  NAND2_X1 U12724 ( .A1(n15196), .A2(n9986), .ZN(n9983) );
  NAND2_X1 U12725 ( .A1(n15196), .A2(n9798), .ZN(n9985) );
  INV_X1 U12726 ( .A(n11540), .ZN(n9987) );
  INV_X1 U12727 ( .A(n15234), .ZN(n9990) );
  INV_X1 U12728 ( .A(n9998), .ZN(n11518) );
  INV_X1 U12729 ( .A(n10006), .ZN(n14043) );
  NAND2_X1 U12730 ( .A1(n10901), .A2(n10900), .ZN(n15080) );
  OR2_X1 U12731 ( .A1(n14525), .A2(n15509), .ZN(n11276) );
  INV_X1 U12732 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10018) );
  INV_X1 U12733 ( .A(n10025), .ZN(n16808) );
  INV_X1 U12734 ( .A(n10028), .ZN(n16772) );
  NOR2_X4 U12735 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11694) );
  NAND2_X1 U12736 ( .A1(n12414), .A2(n12413), .ZN(n10034) );
  NAND2_X1 U12737 ( .A1(n10034), .A2(n10036), .ZN(n13822) );
  NAND2_X1 U12738 ( .A1(n10035), .A2(n12432), .ZN(n13825) );
  NAND2_X1 U12739 ( .A1(n12035), .A2(n12036), .ZN(n12062) );
  NAND2_X1 U12740 ( .A1(n12875), .A2(n10045), .ZN(n10048) );
  NAND2_X1 U12741 ( .A1(n12875), .A2(n12876), .ZN(n13012) );
  INV_X1 U12742 ( .A(n10048), .ZN(n13043) );
  INV_X1 U12743 ( .A(n13015), .ZN(n10047) );
  NOR2_X2 U12744 ( .A1(n14125), .A2(n10049), .ZN(n14367) );
  NAND2_X1 U12745 ( .A1(n12512), .A2(n12511), .ZN(n14125) );
  NAND3_X1 U12746 ( .A1(n13048), .A2(n13683), .A3(n13685), .ZN(n12216) );
  INV_X1 U12747 ( .A(n10055), .ZN(n14696) );
  INV_X1 U12748 ( .A(n10078), .ZN(n15423) );
  NAND2_X1 U12749 ( .A1(n10202), .A2(n10242), .ZN(n10186) );
  AND2_X1 U12750 ( .A1(n10081), .A2(n15835), .ZN(n19415) );
  NOR2_X1 U12751 ( .A1(n10352), .A2(n11277), .ZN(n10081) );
  NAND2_X1 U12752 ( .A1(n14449), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10082) );
  INV_X1 U12753 ( .A(n10442), .ZN(n10086) );
  NAND2_X1 U12754 ( .A1(n12910), .A2(n10088), .ZN(n12911) );
  OR2_X1 U12755 ( .A1(n13666), .A2(n13665), .ZN(n13667) );
  NAND2_X1 U12756 ( .A1(n13666), .A2(n13665), .ZN(n13664) );
  NAND2_X1 U12757 ( .A1(n12458), .A2(n12457), .ZN(n14087) );
  NAND2_X1 U12758 ( .A1(n15300), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11255) );
  NAND2_X1 U12759 ( .A1(n12346), .A2(n19404), .ZN(n12357) );
  NAND2_X1 U12760 ( .A1(n12346), .A2(n16461), .ZN(n11253) );
  XNOR2_X1 U12761 ( .A(n11255), .B(n11254), .ZN(n12915) );
  AOI21_X1 U12762 ( .B1(n12912), .B2(n16471), .A(n12911), .ZN(n12913) );
  AND2_X1 U12763 ( .A1(n12308), .A2(n13049), .ZN(n14556) );
  INV_X1 U12764 ( .A(n14330), .ZN(n15165) );
  NAND2_X1 U12765 ( .A1(n10243), .A2(n10805), .ZN(n10248) );
  AND2_X1 U12766 ( .A1(n10982), .A2(n10274), .ZN(n10275) );
  AND2_X1 U12767 ( .A1(n14126), .A2(n12510), .ZN(n12511) );
  INV_X1 U12768 ( .A(n14087), .ZN(n12512) );
  NAND2_X1 U12769 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11785) );
  CLKBUF_X1 U12770 ( .A(n12183), .Z(n13768) );
  NAND2_X1 U12771 ( .A1(n10985), .A2(n10262), .ZN(n10283) );
  INV_X1 U12772 ( .A(n12147), .ZN(n12207) );
  AOI22_X1 U12773 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10414) );
  OAI22_X1 U12774 ( .A1(n11521), .A2(n10480), .B1(n10516), .B2(n10409), .ZN(
        n10410) );
  OAI21_X2 U12775 ( .B1(n15700), .B2(n15380), .A(n15698), .ZN(n15444) );
  AOI21_X1 U12776 ( .B1(n10485), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n11007), .ZN(n10347) );
  NAND2_X1 U12777 ( .A1(n11913), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11835) );
  NAND2_X1 U12778 ( .A1(n20243), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12151) );
  OAI21_X1 U12779 ( .B1(n14171), .B2(n11262), .A(n14144), .ZN(n15815) );
  OR2_X1 U12780 ( .A1(n11912), .A2(n11911), .ZN(n11919) );
  OAI22_X1 U12781 ( .A1(n10297), .A2(n10282), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10292), .ZN(n10286) );
  AOI21_X1 U12782 ( .B1(n10814), .B2(n10813), .A(n10812), .ZN(n13791) );
  AOI22_X1 U12783 ( .A1(n10475), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n19698), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10422) );
  NAND2_X1 U12784 ( .A1(n11277), .A2(n11299), .ZN(n11283) );
  NAND2_X1 U12785 ( .A1(n11277), .A2(n10345), .ZN(n10333) );
  AOI22_X1 U12786 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U12787 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12992), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11745) );
  NAND2_X1 U12788 ( .A1(n11300), .A2(n10348), .ZN(n10355) );
  NAND2_X1 U12789 ( .A1(n11428), .A2(n10370), .ZN(n10087) );
  AND2_X1 U12790 ( .A1(n12909), .A2(n12908), .ZN(n10088) );
  OR3_X1 U12791 ( .A1(n15543), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15522), .ZN(n10089) );
  AND4_X1 U12792 ( .A1(n12193), .A2(n12398), .A3(n13019), .A4(n20286), .ZN(
        n10090) );
  AND2_X2 U12793 ( .A1(n11700), .A2(n13753), .ZN(n11997) );
  NOR2_X1 U12794 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12872) );
  NOR2_X1 U12795 ( .A1(n20998), .A2(n20851), .ZN(n10091) );
  AND3_X1 U12796 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .ZN(n10092) );
  AND2_X1 U12797 ( .A1(n9721), .A2(n12382), .ZN(n10093) );
  AND3_X1 U12798 ( .A1(n10726), .A2(n15409), .A3(n15383), .ZN(n10094) );
  OR3_X1 U12799 ( .A1(n15391), .A2(n15389), .A3(n10747), .ZN(n10095) );
  AND3_X1 U12800 ( .A1(n13106), .A2(n13105), .A3(n13104), .ZN(n10096) );
  INV_X1 U12801 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12380) );
  INV_X1 U12802 ( .A(n20230), .ZN(n20220) );
  AND2_X1 U12803 ( .A1(n15035), .A2(n12010), .ZN(n10097) );
  OR2_X1 U12804 ( .A1(n17210), .A2(n15929), .ZN(n10098) );
  OR2_X1 U12805 ( .A1(n17210), .A2(n17101), .ZN(n10099) );
  OR2_X1 U12806 ( .A1(n15392), .A2(n15391), .ZN(n10100) );
  NOR2_X1 U12807 ( .A1(n10733), .A2(n15392), .ZN(n10101) );
  NAND2_X1 U12808 ( .A1(n11223), .A2(n11222), .ZN(n10102) );
  INV_X1 U12809 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11254) );
  INV_X1 U12810 ( .A(n10392), .ZN(n11161) );
  AND2_X1 U12811 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .ZN(n10103) );
  AND3_X1 U12812 ( .A1(n13116), .A2(n13115), .A3(n13114), .ZN(n10104) );
  INV_X1 U12813 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20032) );
  AND2_X1 U12814 ( .A1(n17706), .A2(n17705), .ZN(n10105) );
  OR2_X1 U12815 ( .A1(n14535), .A2(n20238), .ZN(n10106) );
  AND3_X1 U12816 ( .A1(n11091), .A2(n11090), .A3(n11089), .ZN(n13855) );
  INV_X1 U12817 ( .A(n13855), .ZN(n11317) );
  AND3_X1 U12818 ( .A1(n17396), .A2(n17395), .A3(P3_EBX_REG_4__SCAN_IN), .ZN(
        n10107) );
  INV_X1 U12819 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10781) );
  NOR2_X1 U12820 ( .A1(n15488), .A2(n15491), .ZN(n10108) );
  INV_X1 U12821 ( .A(n10774), .ZN(n10775) );
  AND4_X1 U12822 ( .A1(n10202), .A2(n10257), .A3(n11013), .A4(n10240), .ZN(
        n10109) );
  NOR2_X1 U12823 ( .A1(n20720), .A2(n20851), .ZN(n10110) );
  OR2_X1 U12824 ( .A1(n18986), .A2(n13066), .ZN(n10111) );
  OR2_X1 U12825 ( .A1(n12353), .A2(n15800), .ZN(n10112) );
  XOR2_X1 U12826 ( .A(n12379), .B(n12121), .Z(n10113) );
  OR2_X1 U12827 ( .A1(n11379), .A2(n11378), .ZN(n10115) );
  AND2_X1 U12828 ( .A1(n9766), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10116) );
  AND2_X1 U12829 ( .A1(n13423), .A2(n13398), .ZN(n10117) );
  INV_X1 U12830 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13167) );
  AND2_X1 U12831 ( .A1(n15275), .A2(n15274), .ZN(n10118) );
  INV_X1 U12832 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n11002) );
  OR2_X1 U12833 ( .A1(n16077), .A2(n16076), .ZN(n10119) );
  OR2_X1 U12834 ( .A1(n17847), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10120) );
  INV_X1 U12835 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12426) );
  NOR2_X1 U12836 ( .A1(n12211), .A2(n20243), .ZN(n11836) );
  NAND2_X1 U12837 ( .A1(n11823), .A2(n20286), .ZN(n12190) );
  INV_X1 U12838 ( .A(n12190), .ZN(n11825) );
  NOR2_X1 U12839 ( .A1(n12147), .A2(n20243), .ZN(n10121) );
  INV_X1 U12840 ( .A(n12145), .ZN(n12164) );
  NOR2_X1 U12841 ( .A1(n11840), .A2(n20060), .ZN(n11845) );
  NOR2_X1 U12842 ( .A1(n10690), .A2(n15788), .ZN(n10691) );
  AND2_X1 U12843 ( .A1(n10475), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10349) );
  OR2_X1 U12844 ( .A1(n12032), .A2(n12031), .ZN(n12065) );
  INV_X1 U12845 ( .A(n15388), .ZN(n10729) );
  INV_X1 U12846 ( .A(n12146), .ZN(n12133) );
  INV_X1 U12847 ( .A(n13935), .ZN(n12458) );
  AND2_X1 U12848 ( .A1(n12009), .A2(n12008), .ZN(n12013) );
  BUF_X1 U12849 ( .A(n11828), .Z(n13744) );
  NOR2_X1 U12850 ( .A1(n11900), .A2(n11887), .ZN(n11938) );
  INV_X1 U12851 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U12852 ( .A1(n10094), .A2(n10729), .ZN(n10733) );
  NAND2_X1 U12853 ( .A1(n10972), .A2(n10970), .ZN(n10233) );
  AOI22_X1 U12854 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U12855 ( .A1(n13113), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13104) );
  INV_X1 U12856 ( .A(n14423), .ZN(n12529) );
  INV_X1 U12857 ( .A(n14713), .ZN(n12678) );
  INV_X1 U12858 ( .A(n14473), .ZN(n12609) );
  NAND2_X1 U12859 ( .A1(n12819), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11704) );
  OR2_X1 U12860 ( .A1(n12007), .A2(n12006), .ZN(n12041) );
  OR2_X1 U12861 ( .A1(n10610), .A2(n10611), .ZN(n10613) );
  INV_X1 U12862 ( .A(n10369), .ZN(n11410) );
  NAND2_X1 U12863 ( .A1(n10932), .A2(n10929), .ZN(n10591) );
  AND2_X1 U12864 ( .A1(n19143), .A2(n11262), .ZN(n10738) );
  AND2_X1 U12865 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11429) );
  NAND2_X1 U12866 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13228) );
  NAND2_X1 U12867 ( .A1(n11813), .A2(n10090), .ZN(n12183) );
  BUF_X1 U12868 ( .A(n12217), .Z(n12293) );
  INV_X1 U12869 ( .A(n11822), .ZN(n12143) );
  NAND2_X1 U12870 ( .A1(n10097), .A2(n12012), .ZN(n12038) );
  NOR2_X1 U12871 ( .A1(n12832), .A2(n14810), .ZN(n12833) );
  INV_X1 U12872 ( .A(n14633), .ZN(n12784) );
  OR2_X1 U12873 ( .A1(n12088), .A2(n12105), .ZN(n14889) );
  AND2_X1 U12874 ( .A1(n14879), .A2(n14881), .ZN(n12104) );
  OR2_X1 U12875 ( .A1(n12151), .A2(n13019), .ZN(n12167) );
  NAND2_X1 U12876 ( .A1(n10613), .A2(n10612), .ZN(n10640) );
  OR2_X1 U12877 ( .A1(n11469), .A2(n11468), .ZN(n11489) );
  INV_X1 U12878 ( .A(n10087), .ZN(n11402) );
  AND2_X1 U12879 ( .A1(n14388), .A2(n14219), .ZN(n11364) );
  NOR2_X1 U12880 ( .A1(n10509), .A2(n10508), .ZN(n11042) );
  AND2_X1 U12881 ( .A1(n10848), .A2(n10847), .ZN(n14243) );
  NOR2_X1 U12882 ( .A1(n13333), .A2(n13334), .ZN(n13209) );
  NAND3_X1 U12883 ( .A1(n9732), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13066) );
  INV_X1 U12884 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n21323) );
  NOR2_X1 U12885 ( .A1(n9719), .A2(n13326), .ZN(n13345) );
  AND2_X1 U12886 ( .A1(n17958), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13199) );
  INV_X1 U12887 ( .A(n13176), .ZN(n13174) );
  NOR2_X1 U12888 ( .A1(n15910), .A2(n18410), .ZN(n13314) );
  NAND2_X2 U12889 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13062), .ZN(
        n17298) );
  INV_X1 U12890 ( .A(n12196), .ZN(n13559) );
  NAND2_X1 U12891 ( .A1(n11975), .A2(n11974), .ZN(n20406) );
  NAND2_X1 U12892 ( .A1(n11820), .A2(n20243), .ZN(n11842) );
  AND4_X1 U12893 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11811) );
  NOR2_X1 U12894 ( .A1(n9721), .A2(n14833), .ZN(n12361) );
  AND2_X1 U12895 ( .A1(n12643), .A2(n12642), .ZN(n14717) );
  NOR2_X1 U12896 ( .A1(n12401), .A2(n12400), .ZN(n12438) );
  INV_X1 U12897 ( .A(n12558), .ZN(n12582) );
  AND2_X1 U12898 ( .A1(n12255), .A2(n12254), .ZN(n14131) );
  INV_X1 U12899 ( .A(n13937), .ZN(n12234) );
  INV_X1 U12900 ( .A(n13953), .ZN(n12225) );
  INV_X1 U12901 ( .A(n12313), .ZN(n15048) );
  AND2_X1 U12902 ( .A1(n20564), .A2(n20595), .ZN(n20572) );
  AND2_X1 U12903 ( .A1(n20680), .A2(n20714), .ZN(n20684) );
  INV_X1 U12904 ( .A(n20281), .ZN(n20287) );
  NAND2_X1 U12905 ( .A1(n10769), .A2(n10771), .ZN(n10783) );
  OR2_X1 U12906 ( .A1(n11069), .A2(n11068), .ZN(n11314) );
  OR2_X1 U12907 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  INV_X1 U12908 ( .A(n15124), .ZN(n15125) );
  AND2_X1 U12909 ( .A1(n19435), .A2(n11002), .ZN(n11008) );
  INV_X1 U12910 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10906) );
  AND2_X1 U12911 ( .A1(n10706), .A2(n10705), .ZN(n15453) );
  NOR2_X1 U12912 ( .A1(n11239), .A2(n16463), .ZN(n15794) );
  INV_X1 U12913 ( .A(n13627), .ZN(n15663) );
  AND2_X1 U12914 ( .A1(n12955), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11299) );
  INV_X1 U12915 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17354) );
  AOI21_X1 U12916 ( .B1(n17704), .B2(n17703), .A(n17971), .ZN(n17706) );
  INV_X1 U12917 ( .A(n13202), .ZN(n13200) );
  OAI21_X1 U12918 ( .B1(n13193), .B2(n13397), .A(n13190), .ZN(n13191) );
  NAND2_X1 U12919 ( .A1(n17901), .A2(n17904), .ZN(n17870) );
  NOR2_X1 U12920 ( .A1(n18814), .A2(n17548), .ZN(n18191) );
  NAND2_X1 U12921 ( .A1(n13314), .A2(n13313), .ZN(n13315) );
  NOR2_X1 U12922 ( .A1(n13231), .A2(n13230), .ZN(n13232) );
  NOR2_X1 U12923 ( .A1(n13267), .A2(n13266), .ZN(n13268) );
  AND2_X1 U12924 ( .A1(n12316), .A2(n12323), .ZN(n14562) );
  AND2_X1 U12925 ( .A1(n12274), .A2(n12273), .ZN(n14719) );
  INV_X1 U12926 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14413) );
  NOR2_X1 U12927 ( .A1(n14040), .A2(n14025), .ZN(n14038) );
  OR2_X1 U12928 ( .A1(n12875), .A2(n12876), .ZN(n12877) );
  NAND2_X1 U12929 ( .A1(n12804), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12832) );
  NAND2_X1 U12930 ( .A1(n12362), .A2(n12361), .ZN(n12363) );
  AND2_X1 U12931 ( .A1(n14210), .A2(n14128), .ZN(n14231) );
  AND2_X1 U12932 ( .A1(n12449), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12459) );
  AND2_X1 U12933 ( .A1(n12880), .A2(n14565), .ZN(n16040) );
  NAND2_X1 U12934 ( .A1(n12372), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12373) );
  AND2_X1 U12935 ( .A1(n14969), .A2(n12328), .ZN(n14979) );
  INV_X1 U12936 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n14021) );
  AND2_X1 U12937 ( .A1(n20300), .A2(n20299), .ZN(n20326) );
  AND2_X1 U12938 ( .A1(n20409), .A2(n20408), .ZN(n20434) );
  NOR2_X1 U12939 ( .A1(n20412), .A2(n20796), .ZN(n20643) );
  OR2_X1 U12940 ( .A1(n20241), .A2(n15036), .ZN(n20637) );
  INV_X1 U12941 ( .A(n20819), .ZN(n20871) );
  INV_X1 U12942 ( .A(n20840), .ZN(n20908) );
  AND2_X1 U12943 ( .A1(n13884), .A2(n13883), .ZN(n16043) );
  AND2_X1 U12944 ( .A1(n10861), .A2(n10860), .ZN(n14441) );
  AND3_X1 U12945 ( .A1(n11114), .A2(n11113), .A3(n11112), .ZN(n13979) );
  NAND2_X1 U12946 ( .A1(n19322), .A2(n11660), .ZN(n15284) );
  AND2_X1 U12947 ( .A1(n19322), .A2(n11677), .ZN(n13603) );
  OR2_X1 U12948 ( .A1(n15822), .A2(n15832), .ZN(n15708) );
  XNOR2_X1 U12949 ( .A(n10573), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16444) );
  OR2_X1 U12950 ( .A1(n11249), .A2(n10999), .ZN(n16474) );
  OR2_X1 U12951 ( .A1(n19848), .A2(n19841), .ZN(n19912) );
  AND2_X1 U12952 ( .A1(n10937), .A2(n10799), .ZN(n11635) );
  NAND2_X1 U12953 ( .A1(n17641), .A2(n15998), .ZN(n16696) );
  NOR2_X1 U12954 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16884), .ZN(n16870) );
  INV_X1 U12955 ( .A(n17068), .ZN(n17011) );
  INV_X1 U12956 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17029) );
  INV_X1 U12957 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n21214) );
  INV_X1 U12958 ( .A(n9720), .ZN(n13148) );
  INV_X1 U12959 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n21200) );
  NAND2_X1 U12960 ( .A1(n16078), .A2(n10119), .ZN(n16079) );
  INV_X1 U12961 ( .A(n17854), .ZN(n17813) );
  NOR2_X1 U12962 ( .A1(n13373), .A2(n13377), .ZN(n13379) );
  NAND2_X1 U12963 ( .A1(n13430), .A2(n10117), .ZN(n13431) );
  NOR2_X1 U12964 ( .A1(n18064), .A2(n16551), .ZN(n16536) );
  NOR2_X1 U12965 ( .A1(n18024), .A2(n18023), .ZN(n18022) );
  OAI221_X1 U12966 ( .B1(n16697), .B2(n17639), .C1(n16697), .C2(n17642), .A(
        n16004), .ZN(n16078) );
  INV_X1 U12967 ( .A(n18620), .ZN(n18721) );
  AND2_X1 U12968 ( .A1(n13256), .A2(n13255), .ZN(n13341) );
  NOR2_X1 U12969 ( .A1(n14537), .A2(n14414), .ZN(n16156) );
  AND2_X1 U12970 ( .A1(n20116), .A2(n14022), .ZN(n20099) );
  NOR2_X1 U12971 ( .A1(n20118), .A2(n14539), .ZN(n20106) );
  AND2_X1 U12972 ( .A1(n20116), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20128) );
  INV_X1 U12973 ( .A(n20153), .ZN(n14707) );
  NOR2_X1 U12974 ( .A1(n14771), .A2(n16581), .ZN(n13039) );
  NAND2_X1 U12975 ( .A1(n13023), .A2(n14575), .ZN(n14767) );
  INV_X1 U12976 ( .A(n13689), .ZN(n20201) );
  INV_X1 U12977 ( .A(n13712), .ZN(n20216) );
  NAND2_X1 U12978 ( .A1(n12675), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12710) );
  NAND2_X1 U12979 ( .A1(n12514), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12553) );
  AND2_X1 U12980 ( .A1(n16256), .A2(n20227), .ZN(n16252) );
  AND2_X1 U12981 ( .A1(n16040), .A2(n14575), .ZN(n20230) );
  NAND2_X1 U12982 ( .A1(n12342), .A2(n12341), .ZN(n12343) );
  NAND2_X1 U12983 ( .A1(n12374), .A2(n12373), .ZN(n12375) );
  OAI21_X1 U12984 ( .B1(n15002), .B2(n14954), .A(n14941), .ZN(n16304) );
  INV_X1 U12985 ( .A(n14979), .ZN(n16340) );
  INV_X1 U12986 ( .A(n16370), .ZN(n16360) );
  NAND2_X1 U12987 ( .A1(n12202), .A2(n14575), .ZN(n12331) );
  INV_X1 U12988 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21136) );
  INV_X1 U12989 ( .A(n16058), .ZN(n15064) );
  INV_X1 U12990 ( .A(n20366), .ZN(n20335) );
  OAI21_X1 U12991 ( .B1(n20341), .B2(n20339), .A(n20338), .ZN(n20363) );
  INV_X1 U12992 ( .A(n20399), .ZN(n20387) );
  INV_X1 U12993 ( .A(n20440), .ZN(n20419) );
  NAND2_X1 U12994 ( .A1(n12414), .A2(n20241), .ZN(n20370) );
  INV_X1 U12995 ( .A(n20463), .ZN(n20474) );
  NOR2_X1 U12996 ( .A1(n20532), .A2(n13889), .ZN(n20441) );
  INV_X1 U12997 ( .A(n20561), .ZN(n20551) );
  INV_X1 U12998 ( .A(n20554), .ZN(n20597) );
  OAI211_X1 U12999 ( .C1(n20591), .C2(n20726), .A(n20643), .B(n20574), .ZN(
        n20598) );
  INV_X1 U13000 ( .A(n20670), .ZN(n20632) );
  NOR2_X1 U13001 ( .A1(n20637), .A2(n13889), .ZN(n20609) );
  INV_X1 U13002 ( .A(n20702), .ZN(n20716) );
  OAI22_X1 U13003 ( .A1(n20731), .A2(n20730), .B1(n20729), .B2(n20728), .ZN(
        n20752) );
  AND2_X1 U13004 ( .A1(n20758), .A2(n12423), .ZN(n20790) );
  INV_X1 U13005 ( .A(n12423), .ZN(n20757) );
  NOR2_X1 U13006 ( .A1(n20272), .A2(n20412), .ZN(n20827) );
  NOR2_X1 U13007 ( .A1(n20291), .A2(n20412), .ZN(n20840) );
  NOR2_X1 U13008 ( .A1(n12414), .A2(n15038), .ZN(n20857) );
  INV_X1 U13009 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20932) );
  NAND2_X1 U13010 ( .A1(n12978), .A2(n12977), .ZN(n12979) );
  NOR2_X1 U13011 ( .A1(n16385), .A2(n19242), .ZN(n13443) );
  INV_X1 U13012 ( .A(n19252), .ZN(n19264) );
  INV_X1 U13013 ( .A(n11635), .ZN(n16502) );
  INV_X1 U13014 ( .A(n19250), .ZN(n19279) );
  NOR2_X1 U13015 ( .A1(n14248), .A2(n14249), .ZN(n14247) );
  INV_X1 U13016 ( .A(n15242), .ZN(n15235) );
  INV_X1 U13017 ( .A(n11626), .ZN(n11627) );
  AND2_X1 U13018 ( .A1(n13603), .A2(n15276), .ZN(n19290) );
  INV_X1 U13019 ( .A(n19324), .ZN(n19343) );
  INV_X1 U13020 ( .A(n13568), .ZN(n19393) );
  INV_X1 U13021 ( .A(n11670), .ZN(n14002) );
  OR2_X1 U13022 ( .A1(n12353), .A2(n16435), .ZN(n12354) );
  INV_X1 U13023 ( .A(n16428), .ZN(n16442) );
  NOR3_X1 U13024 ( .A1(n16482), .A2(n14164), .A3(n14163), .ZN(n15823) );
  INV_X1 U13025 ( .A(n16474), .ZN(n16457) );
  AOI21_X2 U13026 ( .B1(n15882), .B2(n13995), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19851) );
  INV_X1 U13027 ( .A(n19919), .ZN(n19442) );
  NOR2_X1 U13028 ( .A1(n19574), .A2(n20003), .ZN(n19524) );
  INV_X1 U13029 ( .A(n19527), .ZN(n19545) );
  INV_X1 U13030 ( .A(n19563), .ZN(n21345) );
  INV_X1 U13031 ( .A(n19592), .ZN(n19606) );
  NOR2_X1 U13032 ( .A1(n19846), .A2(n19574), .ZN(n19631) );
  NAND2_X1 U13033 ( .A1(n19503), .A2(n19277), .ZN(n19609) );
  NOR2_X1 U13034 ( .A1(n19690), .A2(n19455), .ZN(n19685) );
  NAND2_X1 U13035 ( .A1(n20020), .A2(n14061), .ZN(n19455) );
  NAND2_X1 U13036 ( .A1(n20020), .A2(n20026), .ZN(n20003) );
  INV_X1 U13037 ( .A(n19739), .ZN(n21346) );
  INV_X1 U13038 ( .A(n19758), .ZN(n19914) );
  AND3_X1 U13039 ( .A1(n19921), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19927) );
  INV_X1 U13040 ( .A(n19044), .ZN(n19046) );
  NOR2_X1 U13041 ( .A1(n17070), .A2(n16715), .ZN(n16758) );
  NOR2_X1 U13042 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16911), .ZN(n16891) );
  NOR4_X1 U13043 ( .A1(n17070), .A2(n18937), .A3(n18934), .A4(n16902), .ZN(
        n16883) );
  INV_X1 U13044 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17034) );
  INV_X1 U13045 ( .A(n17073), .ZN(n17058) );
  NAND2_X1 U13046 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17397), .ZN(n17389) );
  NAND2_X1 U13047 ( .A1(n17642), .A2(n17579), .ZN(n15912) );
  NOR2_X1 U13048 ( .A1(n17588), .A2(n17462), .ZN(n17457) );
  NOR3_X1 U13049 ( .A1(n17512), .A2(n17477), .A3(n17595), .ZN(n17473) );
  INV_X1 U13050 ( .A(n17565), .ZN(n17544) );
  AND2_X1 U13051 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13134) );
  INV_X1 U13052 ( .A(n13292), .ZN(n18410) );
  NOR2_X1 U13053 ( .A1(n18082), .A2(n18096), .ZN(n17737) );
  INV_X1 U13054 ( .A(n16563), .ZN(n18190) );
  NAND2_X1 U13055 ( .A1(n17837), .A2(n17864), .ZN(n18048) );
  INV_X1 U13056 ( .A(n19033), .ZN(n17642) );
  OAI21_X1 U13057 ( .B1(n18164), .B2(n17832), .A(n16564), .ZN(n18121) );
  INV_X1 U13058 ( .A(n17927), .ZN(n18240) );
  NOR2_X2 U13059 ( .A1(n18359), .A2(n18074), .ZN(n18263) );
  INV_X1 U13060 ( .A(n18343), .ZN(n18291) );
  INV_X1 U13061 ( .A(n18338), .ZN(n18359) );
  INV_X1 U13062 ( .A(n17060), .ZN(n18885) );
  INV_X1 U13063 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18871) );
  INV_X1 U13064 ( .A(U212), .ZN(n16629) );
  INV_X1 U13065 ( .A(n21016), .ZN(n14040) );
  INV_X1 U13066 ( .A(n20128), .ZN(n20094) );
  INV_X1 U13067 ( .A(n20127), .ZN(n16168) );
  INV_X1 U13068 ( .A(n16156), .ZN(n16174) );
  INV_X1 U13069 ( .A(n20154), .ZN(n20179) );
  NOR2_X1 U13070 ( .A1(n13593), .A2(n13592), .ZN(n13688) );
  AOI21_X1 U13071 ( .B1(n10113), .B2(n20230), .A(n12887), .ZN(n12888) );
  INV_X1 U13072 ( .A(n16252), .ZN(n20219) );
  INV_X1 U13073 ( .A(n13942), .ZN(n20238) );
  AOI21_X1 U13074 ( .B1(n12376), .B2(n16367), .A(n12375), .ZN(n12377) );
  OR2_X1 U13075 ( .A1(n12331), .A2(n12311), .ZN(n16341) );
  OR2_X1 U13076 ( .A1(n12331), .A2(n12210), .ZN(n16370) );
  INV_X1 U13077 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20236) );
  NAND2_X1 U13078 ( .A1(n20306), .A2(n12423), .ZN(n20332) );
  NAND2_X1 U13079 ( .A1(n20306), .A2(n20757), .ZN(n20366) );
  OR2_X1 U13080 ( .A1(n20370), .A2(n20638), .ZN(n20399) );
  OR2_X1 U13081 ( .A1(n20370), .A2(n20531), .ZN(n20440) );
  NAND2_X1 U13082 ( .A1(n20441), .A2(n20757), .ZN(n20513) );
  OR2_X1 U13083 ( .A1(n20532), .A2(n20531), .ZN(n20554) );
  NAND2_X1 U13084 ( .A1(n20480), .A2(n12423), .ZN(n20561) );
  NAND2_X1 U13085 ( .A1(n20609), .A2(n12423), .ZN(n20636) );
  NAND2_X1 U13086 ( .A1(n20609), .A2(n20757), .ZN(n20670) );
  NAND2_X1 U13087 ( .A1(n20691), .A2(n20794), .ZN(n20702) );
  NAND2_X1 U13088 ( .A1(n20691), .A2(n20690), .ZN(n20756) );
  NAND2_X1 U13089 ( .A1(n20758), .A2(n20757), .ZN(n20810) );
  NAND2_X1 U13090 ( .A1(n20857), .A2(n20690), .ZN(n20906) );
  NAND2_X1 U13091 ( .A1(n20857), .A2(n20794), .ZN(n20918) );
  INV_X1 U13092 ( .A(n20990), .ZN(n20923) );
  AND2_X1 U13093 ( .A1(n20932), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21009) );
  AOI21_X1 U13094 ( .B1(n15515), .B2(n19273), .A(n12979), .ZN(n12980) );
  INV_X1 U13095 ( .A(n19273), .ZN(n19230) );
  INV_X1 U13096 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19184) );
  NAND2_X1 U13097 ( .A1(n19222), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19250) );
  INV_X1 U13098 ( .A(n19266), .ZN(n19258) );
  AND2_X2 U13099 ( .A1(n11630), .A2(n19927), .ZN(n15229) );
  INV_X1 U13100 ( .A(n19339), .ZN(n19297) );
  NAND2_X1 U13101 ( .A1(n19385), .A2(n15074), .ZN(n19357) );
  AND2_X1 U13102 ( .A1(n13570), .A2(n13569), .ZN(n19385) );
  OR2_X1 U13103 ( .A1(n13463), .A2(n11284), .ZN(n13568) );
  INV_X1 U13104 ( .A(n19394), .ZN(n13541) );
  AND2_X1 U13105 ( .A1(n12355), .A2(n12354), .ZN(n12356) );
  INV_X1 U13106 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n21179) );
  INV_X1 U13107 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19209) );
  NAND2_X1 U13108 ( .A1(n19409), .A2(n20025), .ZN(n15509) );
  AOI211_X1 U13109 ( .C1(n15535), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15534), .B(n15533), .ZN(n15538) );
  AND2_X1 U13110 ( .A1(n11251), .A2(n10112), .ZN(n11252) );
  OR2_X1 U13111 ( .A1(n11249), .A2(n20048), .ZN(n16476) );
  INV_X1 U13112 ( .A(n16471), .ZN(n15800) );
  INV_X1 U13113 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20040) );
  INV_X1 U13114 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13556) );
  OR2_X1 U13115 ( .A1(n19455), .A2(n19574), .ZN(n19475) );
  OR2_X1 U13116 ( .A1(n19609), .A2(n20003), .ZN(n19527) );
  AOI21_X1 U13117 ( .B1(n15894), .B2(n15893), .A(n15892), .ZN(n19549) );
  AND2_X1 U13118 ( .A1(n19583), .A2(n19582), .ZN(n19592) );
  INV_X1 U13119 ( .A(n19599), .ZN(n21352) );
  INV_X1 U13120 ( .A(n19631), .ZN(n19638) );
  OR2_X1 U13121 ( .A1(n19609), .A2(n19846), .ZN(n19663) );
  INV_X1 U13122 ( .A(n19687), .ZN(n19678) );
  INV_X1 U13123 ( .A(n19685), .ZN(n19683) );
  OR2_X1 U13124 ( .A1(n19730), .A2(n19455), .ZN(n19723) );
  OR2_X1 U13125 ( .A1(n19690), .A2(n20003), .ZN(n19757) );
  INV_X1 U13126 ( .A(n19807), .ZN(n19801) );
  INV_X1 U13127 ( .A(n19798), .ZN(n19810) );
  OR2_X1 U13128 ( .A1(n19730), .A2(n19846), .ZN(n19919) );
  INV_X1 U13129 ( .A(n20002), .ZN(n19930) );
  INV_X1 U13130 ( .A(n17069), .ZN(n17062) );
  INV_X1 U13131 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17995) );
  NOR2_X1 U13132 ( .A1(n17084), .A2(n17083), .ZN(n17112) );
  NAND2_X1 U13133 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17134), .ZN(n17126) );
  AND2_X1 U13134 ( .A1(n17424), .A2(n17478), .ZN(n17422) );
  INV_X1 U13135 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17416) );
  INV_X1 U13136 ( .A(n17538), .ZN(n17542) );
  NAND2_X1 U13137 ( .A1(n17638), .A2(n17578), .ZN(n17636) );
  INV_X1 U13138 ( .A(n17691), .ZN(n17686) );
  INV_X1 U13139 ( .A(n18048), .ZN(n18034) );
  INV_X1 U13140 ( .A(n18047), .ZN(n18058) );
  OR2_X1 U13141 ( .A1(n18131), .A2(n18130), .ZN(n18154) );
  NAND2_X1 U13142 ( .A1(n18358), .A2(n18359), .ZN(n18343) );
  INV_X1 U13143 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18834) );
  INV_X1 U13144 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18418) );
  INV_X1 U13145 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18438) );
  INV_X1 U13146 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18614) );
  INV_X1 U13147 ( .A(n18598), .ZN(n18763) );
  INV_X1 U13148 ( .A(n18867), .ZN(n18883) );
  INV_X1 U13149 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18910) );
  INV_X1 U13150 ( .A(n16627), .ZN(n16632) );
  OAI21_X1 U13151 ( .B1(n14732), .B2(n14728), .A(n13060), .ZN(P1_U2842) );
  NAND2_X1 U13152 ( .A1(n12345), .A2(n12344), .ZN(P1_U3002) );
  OAI21_X1 U13153 ( .B1(n15368), .B2(n11253), .A(n11252), .ZN(P2_U3024) );
  AND2_X4 U13154 ( .A1(n14321), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11619) );
  AND2_X4 U13155 ( .A1(n14321), .A2(n10362), .ZN(n10221) );
  AND2_X4 U13156 ( .A1(n14323), .A2(n10362), .ZN(n10203) );
  AOI22_X1 U13157 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9726), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10124) );
  AND2_X4 U13158 ( .A1(n15852), .A2(n16484), .ZN(n11426) );
  AOI22_X1 U13159 ( .A1(n11426), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10123) );
  AND2_X4 U13160 ( .A1(n10370), .A2(n16484), .ZN(n10222) );
  AOI22_X1 U13161 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U13162 ( .A1(n10126), .A2(n15872), .ZN(n10133) );
  AOI22_X1 U13163 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9726), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U13164 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10221), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U13165 ( .A1(n11426), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U13166 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10127) );
  NAND4_X1 U13167 ( .A1(n10130), .A2(n10129), .A3(n10128), .A4(n10127), .ZN(
        n10131) );
  NAND2_X2 U13168 ( .A1(n10133), .A2(n10132), .ZN(n10240) );
  AOI22_X1 U13169 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10221), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U13170 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U13171 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10135) );
  NAND4_X1 U13172 ( .A1(n10138), .A2(n10137), .A3(n10136), .A4(n10135), .ZN(
        n10139) );
  NAND2_X1 U13173 ( .A1(n10139), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10147) );
  AOI22_X1 U13174 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10221), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U13175 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10142) );
  AOI22_X1 U13176 ( .A1(n11426), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U13177 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10140) );
  NAND4_X1 U13178 ( .A1(n10143), .A2(n10142), .A3(n10141), .A4(n10140), .ZN(
        n10145) );
  AOI22_X1 U13179 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11426), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U13180 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U13181 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U13182 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9726), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10148) );
  NAND4_X1 U13183 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n10152) );
  NAND2_X1 U13184 ( .A1(n10152), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10159) );
  AOI22_X1 U13185 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11426), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U13186 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9726), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U13187 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U13188 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10153) );
  NAND4_X1 U13189 ( .A1(n10156), .A2(n10155), .A3(n10154), .A4(n10153), .ZN(
        n10157) );
  NAND2_X1 U13190 ( .A1(n10157), .A2(n15872), .ZN(n10158) );
  NAND2_X1 U13191 ( .A1(n10257), .A2(n10242), .ZN(n10160) );
  AOI22_X1 U13192 ( .A1(n11426), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U13193 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U13194 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10221), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U13195 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10161) );
  NAND4_X1 U13196 ( .A1(n10164), .A2(n10163), .A3(n10162), .A4(n10161), .ZN(
        n10165) );
  NAND2_X1 U13197 ( .A1(n10165), .A2(n15872), .ZN(n10172) );
  AOI22_X1 U13198 ( .A1(n11426), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U13199 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10221), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U13200 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10166) );
  NAND4_X1 U13201 ( .A1(n10168), .A2(n10169), .A3(n10167), .A4(n10166), .ZN(
        n10170) );
  NAND2_X1 U13202 ( .A1(n10170), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10171) );
  AOI22_X1 U13203 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U13204 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U13205 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11426), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U13206 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10173) );
  NAND4_X1 U13207 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  AOI22_X1 U13208 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11426), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10182) );
  INV_X2 U13209 ( .A(n10178), .ZN(n11586) );
  AOI22_X1 U13210 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n11586), .ZN(n10181) );
  AOI22_X1 U13211 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13212 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10179) );
  NAND4_X1 U13213 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10183) );
  NAND2_X1 U13214 ( .A1(n10183), .A2(n15872), .ZN(n10184) );
  NAND2_X1 U13215 ( .A1(n10186), .A2(n10949), .ZN(n10201) );
  NAND2_X2 U13216 ( .A1(n10187), .A2(n10257), .ZN(n10231) );
  AOI22_X1 U13217 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13218 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13219 ( .A1(n11426), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U13220 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10188) );
  NAND4_X1 U13221 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n10192) );
  AOI22_X1 U13222 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13223 ( .A1(n11426), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U13224 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10194) );
  NAND2_X1 U13225 ( .A1(n10198), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10199) );
  NAND2_X1 U13226 ( .A1(n10231), .A2(n19425), .ZN(n10237) );
  AOI22_X1 U13227 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10206) );
  AOI22_X1 U13228 ( .A1(n11426), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U13229 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10204) );
  NAND4_X1 U13230 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n10208) );
  AOI22_X1 U13231 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U13232 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U13233 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10210) );
  NAND4_X1 U13234 ( .A1(n10213), .A2(n10212), .A3(n10211), .A4(n10210), .ZN(
        n10214) );
  AOI22_X1 U13235 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U13236 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11426), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10217) );
  AOI22_X1 U13237 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10216) );
  NAND4_X1 U13238 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10220) );
  AOI22_X1 U13239 ( .A1(n10203), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10226) );
  AOI22_X1 U13240 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11426), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U13241 ( .A1(n11619), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U13242 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10223) );
  NAND4_X1 U13243 ( .A1(n10226), .A2(n10225), .A3(n10224), .A4(n10223), .ZN(
        n10227) );
  AND2_X1 U13244 ( .A1(n10231), .A2(n11007), .ZN(n10228) );
  NAND2_X1 U13245 ( .A1(n10972), .A2(n10228), .ZN(n10272) );
  NAND2_X1 U13246 ( .A1(n10272), .A2(n9722), .ZN(n10229) );
  AND2_X1 U13247 ( .A1(n10955), .A2(n11013), .ZN(n10232) );
  NAND2_X1 U13248 ( .A1(n10607), .A2(n10242), .ZN(n10251) );
  NAND2_X1 U13249 ( .A1(n10251), .A2(n10231), .ZN(n10945) );
  NAND2_X1 U13250 ( .A1(n10945), .A2(n10202), .ZN(n10951) );
  NAND2_X1 U13251 ( .A1(n10234), .A2(n10233), .ZN(n10273) );
  NAND2_X1 U13252 ( .A1(n10273), .A2(n10263), .ZN(n10235) );
  NAND2_X1 U13253 ( .A1(n10274), .A2(n10235), .ZN(n10236) );
  NAND2_X1 U13254 ( .A1(n10236), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10245) );
  INV_X1 U13255 ( .A(n10237), .ZN(n10239) );
  AND2_X1 U13256 ( .A1(n10202), .A2(n10257), .ZN(n10238) );
  NAND2_X1 U13257 ( .A1(n10239), .A2(n10238), .ZN(n10944) );
  NOR2_X1 U13258 ( .A1(n11007), .A2(n10240), .ZN(n10241) );
  NAND2_X1 U13259 ( .A1(n10944), .A2(n10241), .ZN(n10244) );
  NAND2_X1 U13260 ( .A1(n10244), .A2(n10941), .ZN(n10998) );
  NAND2_X1 U13261 ( .A1(n9736), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13571) );
  NAND2_X2 U13262 ( .A1(n10245), .A2(n10270), .ZN(n10297) );
  NAND2_X1 U13263 ( .A1(n10297), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10256) );
  INV_X1 U13264 ( .A(n10246), .ZN(n10247) );
  NAND2_X1 U13265 ( .A1(n10247), .A2(n9722), .ZN(n10953) );
  NAND2_X1 U13266 ( .A1(n9742), .A2(n14076), .ZN(n10249) );
  NAND2_X1 U13267 ( .A1(n10262), .A2(n10250), .ZN(n10973) );
  INV_X1 U13268 ( .A(n10251), .ZN(n10252) );
  NOR2_X1 U13269 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10908) );
  AND2_X2 U13270 ( .A1(n10256), .A2(n10255), .ZN(n10288) );
  NAND2_X1 U13271 ( .A1(n10996), .A2(n10932), .ZN(n10261) );
  NOR2_X1 U13272 ( .A1(n10257), .A2(n11004), .ZN(n11001) );
  MUX2_X1 U13273 ( .A(n11001), .B(n10257), .S(n19425), .Z(n10259) );
  NOR2_X1 U13274 ( .A1(n9746), .A2(n10242), .ZN(n10258) );
  AND3_X2 U13275 ( .A1(n10259), .A2(n11634), .A3(n10258), .ZN(n10985) );
  INV_X1 U13276 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15833) );
  INV_X1 U13277 ( .A(n10972), .ZN(n10264) );
  NAND2_X1 U13278 ( .A1(n10292), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10266) );
  AND2_X4 U13279 ( .A1(n16515), .A2(n10280), .ZN(n11270) );
  AOI22_X1 U13280 ( .A1(n11270), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10265) );
  NAND2_X1 U13281 ( .A1(n10886), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10279) );
  INV_X1 U13282 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10643) );
  INV_X1 U13283 ( .A(n10908), .ZN(n10309) );
  NAND2_X1 U13284 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U13285 ( .A1(n10309), .A2(n10268), .ZN(n10269) );
  AOI21_X1 U13286 ( .B1(n11270), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10269), .ZN(
        n10271) );
  OAI211_X1 U13287 ( .C1(n10808), .C2(n10643), .A(n10271), .B(n10270), .ZN(
        n10277) );
  NAND2_X1 U13288 ( .A1(n10273), .A2(n10272), .ZN(n10982) );
  NOR2_X1 U13289 ( .A1(n10277), .A2(n10276), .ZN(n10278) );
  NAND2_X1 U13290 ( .A1(n10279), .A2(n10278), .ZN(n10324) );
  INV_X1 U13291 ( .A(n10280), .ZN(n10281) );
  NOR2_X1 U13292 ( .A1(n10281), .A2(n10981), .ZN(n10282) );
  INV_X1 U13293 ( .A(n14315), .ZN(n10284) );
  AOI22_X1 U13294 ( .A1(n10284), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n10908), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U13295 ( .A1(n10286), .A2(n10285), .ZN(n10323) );
  NAND2_X1 U13296 ( .A1(n10322), .A2(n10337), .ZN(n10291) );
  INV_X1 U13297 ( .A(n10287), .ZN(n10289) );
  NAND2_X1 U13298 ( .A1(n10289), .A2(n9737), .ZN(n10290) );
  NAND2_X1 U13299 ( .A1(n10291), .A2(n10290), .ZN(n10317) );
  NAND2_X1 U13300 ( .A1(n10292), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13301 ( .A1(n11270), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10293) );
  AND2_X1 U13302 ( .A1(n10294), .A2(n10293), .ZN(n10295) );
  AND2_X2 U13303 ( .A1(n10296), .A2(n10295), .ZN(n10302) );
  INV_X1 U13304 ( .A(n10302), .ZN(n10300) );
  OAI21_X1 U13305 ( .B1(n20024), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n19921), 
        .ZN(n10298) );
  INV_X1 U13306 ( .A(n10301), .ZN(n10299) );
  NAND2_X1 U13307 ( .A1(n10300), .A2(n10299), .ZN(n10303) );
  NAND2_X1 U13308 ( .A1(n10302), .A2(n10301), .ZN(n10304) );
  INV_X1 U13309 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14164) );
  INV_X1 U13310 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n14174) );
  OAI22_X1 U13311 ( .A1(n10896), .A2(n14174), .B1(n19921), .B2(n14176), .ZN(
        n10306) );
  AOI21_X1 U13312 ( .B1(n11271), .B2(P2_EBX_REG_3__SCAN_IN), .A(n10306), .ZN(
        n10307) );
  NOR2_X1 U13313 ( .A1(n10309), .A2(n20017), .ZN(n10310) );
  NAND2_X1 U13314 ( .A1(n10311), .A2(n10312), .ZN(n10811) );
  INV_X1 U13315 ( .A(n10311), .ZN(n10314) );
  INV_X1 U13316 ( .A(n10312), .ZN(n10313) );
  NAND2_X1 U13317 ( .A1(n10314), .A2(n10313), .ZN(n10315) );
  XNOR2_X2 U13318 ( .A(n10814), .B(n10813), .ZN(n11300) );
  BUF_X2 U13319 ( .A(n11300), .Z(n10334) );
  INV_X1 U13320 ( .A(n10317), .ZN(n10320) );
  INV_X1 U13321 ( .A(n10318), .ZN(n10319) );
  INV_X1 U13322 ( .A(n10323), .ZN(n10326) );
  INV_X1 U13323 ( .A(n10324), .ZN(n10325) );
  NAND2_X1 U13324 ( .A1(n10326), .A2(n10325), .ZN(n10327) );
  AND2_X1 U13325 ( .A1(n10322), .A2(n11289), .ZN(n10330) );
  NAND2_X1 U13326 ( .A1(n11277), .A2(n10330), .ZN(n10331) );
  INV_X1 U13327 ( .A(n10480), .ZN(n19612) );
  INV_X1 U13328 ( .A(n10322), .ZN(n10339) );
  AND2_X1 U13329 ( .A1(n10339), .A2(n11289), .ZN(n10345) );
  INV_X1 U13330 ( .A(n10333), .ZN(n10329) );
  AOI22_X1 U13331 ( .A1(n19612), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U13332 ( .A1(n13668), .A2(n10330), .ZN(n10335) );
  INV_X1 U13333 ( .A(n10481), .ZN(n10515) );
  INV_X1 U13334 ( .A(n10331), .ZN(n10332) );
  AND2_X2 U13335 ( .A1(n13739), .A2(n10332), .ZN(n19839) );
  AOI22_X1 U13336 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n19839), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10343) );
  INV_X1 U13337 ( .A(n10516), .ZN(n10484) );
  INV_X1 U13338 ( .A(n10335), .ZN(n10336) );
  AND2_X2 U13339 ( .A1(n13739), .A2(n10336), .ZN(n19725) );
  XNOR2_X2 U13340 ( .A(n10339), .B(n10338), .ZN(n11288) );
  INV_X1 U13341 ( .A(n10353), .ZN(n10340) );
  NAND2_X1 U13342 ( .A1(n10340), .A2(n10356), .ZN(n19759) );
  INV_X1 U13343 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11339) );
  NAND2_X1 U13344 ( .A1(n11277), .A2(n11288), .ZN(n10351) );
  OR2_X1 U13345 ( .A1(n10355), .A2(n10351), .ZN(n10524) );
  INV_X1 U13346 ( .A(n19451), .ZN(n10485) );
  INV_X1 U13347 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14074) );
  OAI211_X1 U13348 ( .C1(n10524), .C2(n19814), .A(n10347), .B(n10346), .ZN(
        n10350) );
  NOR2_X1 U13349 ( .A1(n10350), .A2(n10349), .ZN(n10359) );
  INV_X1 U13350 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11082) );
  OR2_X2 U13351 ( .A1(n10352), .A2(n10351), .ZN(n19584) );
  OR2_X2 U13352 ( .A1(n10353), .A2(n10352), .ZN(n15890) );
  INV_X1 U13353 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15902) );
  OAI22_X1 U13354 ( .A1(n11082), .A2(n19584), .B1(n15890), .B2(n15902), .ZN(
        n10354) );
  AOI21_X1 U13355 ( .B1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n19415), .A(
        n10354), .ZN(n10358) );
  AOI22_X1 U13356 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19698), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10357) );
  NAND4_X1 U13357 ( .A1(n10360), .A2(n10359), .A3(n10357), .A4(n10358), .ZN(
        n10408) );
  AOI22_X1 U13358 ( .A1(n11448), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11463), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10366) );
  AND2_X1 U13359 ( .A1(n11426), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10392) );
  AOI22_X1 U13360 ( .A1(n11451), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13361 ( .A1(n10116), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10364) );
  AND2_X2 U13362 ( .A1(n10801), .A2(n10362), .ZN(n11449) );
  AOI22_X1 U13363 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11449), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10363) );
  NAND4_X1 U13364 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n10377) );
  AND2_X1 U13365 ( .A1(n15855), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10367) );
  AND2_X1 U13366 ( .A1(n11428), .A2(n15852), .ZN(n10397) );
  AOI22_X1 U13367 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10375) );
  NOR2_X1 U13368 ( .A1(n15855), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10368) );
  AND2_X1 U13369 ( .A1(n11428), .A2(n10368), .ZN(n10369) );
  AOI22_X1 U13370 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13371 ( .A1(n11077), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10373) );
  AND2_X2 U13372 ( .A1(n11585), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11080) );
  AOI22_X1 U13373 ( .A1(n11080), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10372) );
  NAND4_X1 U13374 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(
        n10376) );
  NOR2_X1 U13375 ( .A1(n10377), .A2(n10376), .ZN(n11006) );
  OR2_X1 U13376 ( .A1(n11006), .A2(n11284), .ZN(n13620) );
  INV_X1 U13377 ( .A(n13620), .ZN(n10391) );
  AOI22_X1 U13378 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11080), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13379 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11448), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13380 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11450), .B1(
        n11449), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13381 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11451), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10378) );
  NAND4_X1 U13382 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10390) );
  AOI22_X1 U13383 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11077), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10388) );
  INV_X1 U13384 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U13385 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10383) );
  NAND2_X1 U13386 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10382) );
  OAI211_X1 U13387 ( .C1(n11461), .C2(n11081), .A(n10383), .B(n10382), .ZN(
        n10384) );
  INV_X1 U13388 ( .A(n10384), .ZN(n10387) );
  AOI22_X1 U13389 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11402), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10386) );
  NAND2_X1 U13390 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10385) );
  NAND4_X1 U13391 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10389) );
  NAND2_X1 U13392 ( .A1(n10391), .A2(n11017), .ZN(n10444) );
  AOI22_X1 U13393 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11448), .B1(
        n11451), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U13394 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n11080), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U13395 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11450), .B1(
        n11449), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13396 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10453), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10393) );
  NAND4_X1 U13397 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10406) );
  AOI22_X1 U13398 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11077), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10404) );
  INV_X1 U13399 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11104) );
  NAND2_X1 U13400 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10399) );
  NAND2_X1 U13401 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10398) );
  OAI211_X1 U13402 ( .C1(n11461), .C2(n11104), .A(n10399), .B(n10398), .ZN(
        n10400) );
  INV_X1 U13403 ( .A(n10400), .ZN(n10403) );
  AOI22_X1 U13404 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11402), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U13405 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10401) );
  NAND4_X1 U13406 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10405) );
  NAND2_X1 U13407 ( .A1(n10444), .A2(n11025), .ZN(n10407) );
  NAND2_X1 U13408 ( .A1(n10408), .A2(n10407), .ZN(n10443) );
  INV_X1 U13409 ( .A(n10443), .ZN(n10441) );
  AOI22_X1 U13410 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n19839), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13411 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19725), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10412) );
  INV_X1 U13412 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11521) );
  INV_X1 U13413 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10409) );
  INV_X1 U13414 ( .A(n10410), .ZN(n10411) );
  AOI22_X1 U13415 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19415), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10421) );
  INV_X1 U13416 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10416) );
  INV_X1 U13417 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10415) );
  OAI22_X1 U13418 ( .A1(n10416), .A2(n19584), .B1(n15890), .B2(n10415), .ZN(
        n10419) );
  INV_X1 U13419 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10417) );
  INV_X1 U13420 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11372) );
  OAI22_X1 U13421 ( .A1(n10417), .A2(n10524), .B1(n19759), .B2(n11372), .ZN(
        n10418) );
  NOR2_X1 U13422 ( .A1(n10419), .A2(n10418), .ZN(n10420) );
  NAND4_X1 U13423 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        n10440) );
  AOI22_X1 U13424 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n11080), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13425 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11448), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13426 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11450), .B1(
        n11449), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13427 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11451), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10425) );
  NAND4_X1 U13428 ( .A1(n10428), .A2(n10427), .A3(n10426), .A4(n10425), .ZN(
        n10437) );
  AOI22_X1 U13429 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11077), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10435) );
  INV_X1 U13430 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21198) );
  NAND2_X1 U13431 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10430) );
  NAND2_X1 U13432 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10429) );
  OAI211_X1 U13433 ( .C1(n11461), .C2(n21198), .A(n10430), .B(n10429), .ZN(
        n10431) );
  INV_X1 U13434 ( .A(n10431), .ZN(n10434) );
  AOI22_X1 U13435 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11402), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U13436 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10432) );
  NAND4_X1 U13437 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(
        n10436) );
  INV_X1 U13438 ( .A(n11033), .ZN(n10438) );
  NAND2_X1 U13439 ( .A1(n10438), .A2(n11007), .ZN(n10439) );
  AND2_X2 U13440 ( .A1(n10440), .A2(n10439), .ZN(n10442) );
  XOR2_X1 U13441 ( .A(n11025), .B(n10444), .Z(n13636) );
  NAND2_X1 U13442 ( .A1(n13620), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13619) );
  XOR2_X1 U13443 ( .A(n11006), .B(n11017), .Z(n10445) );
  NOR2_X1 U13444 ( .A1(n13619), .A2(n10445), .ZN(n10447) );
  INV_X1 U13445 ( .A(n13619), .ZN(n10446) );
  XOR2_X1 U13446 ( .A(n10446), .B(n10445), .Z(n13611) );
  NOR2_X1 U13447 ( .A1(n15833), .A2(n13611), .ZN(n13610) );
  NOR2_X1 U13448 ( .A1(n10447), .A2(n13610), .ZN(n10448) );
  XOR2_X1 U13449 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10448), .Z(
        n13635) );
  NOR2_X1 U13450 ( .A1(n13636), .A2(n13635), .ZN(n13634) );
  NOR2_X1 U13451 ( .A1(n10448), .A2(n9747), .ZN(n10449) );
  OR2_X1 U13452 ( .A1(n13634), .A2(n10449), .ZN(n10451) );
  XNOR2_X1 U13453 ( .A(n10451), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14170) );
  INV_X1 U13454 ( .A(n14170), .ZN(n10450) );
  NAND2_X1 U13455 ( .A1(n10451), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10452) );
  AOI22_X1 U13456 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11080), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13457 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11448), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13458 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11450), .B1(
        n11449), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U13459 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11451), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10454) );
  NAND4_X1 U13460 ( .A1(n10457), .A2(n10456), .A3(n10455), .A4(n10454), .ZN(
        n10466) );
  AOI22_X1 U13461 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11456), .B1(
        n11077), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10464) );
  NAND2_X1 U13462 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10459) );
  NAND2_X1 U13463 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10458) );
  OAI211_X1 U13464 ( .C1(n11461), .C2(n21251), .A(n10459), .B(n10458), .ZN(
        n10460) );
  INV_X1 U13465 ( .A(n10460), .ZN(n10463) );
  AOI22_X1 U13466 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11402), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U13467 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10461) );
  NAND4_X1 U13468 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10465) );
  INV_X1 U13469 ( .A(n11038), .ZN(n10467) );
  NAND2_X1 U13470 ( .A1(n10468), .A2(n10467), .ZN(n10469) );
  NAND2_X1 U13471 ( .A1(n10635), .A2(n10469), .ZN(n10471) );
  INV_X1 U13472 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15826) );
  NAND2_X1 U13473 ( .A1(n15825), .A2(n15826), .ZN(n10474) );
  INV_X1 U13474 ( .A(n10470), .ZN(n10472) );
  NAND2_X1 U13475 ( .A1(n10472), .A2(n10471), .ZN(n10473) );
  INV_X1 U13476 ( .A(n10475), .ZN(n19478) );
  INV_X1 U13477 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10476) );
  INV_X1 U13478 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11160) );
  INV_X1 U13479 ( .A(n10477), .ZN(n10496) );
  INV_X1 U13480 ( .A(n19415), .ZN(n10478) );
  INV_X1 U13481 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13901) );
  INV_X1 U13482 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11167) );
  OAI22_X1 U13483 ( .A1(n10478), .A2(n13901), .B1(n19641), .B2(n11167), .ZN(
        n10479) );
  INV_X1 U13484 ( .A(n10479), .ZN(n10495) );
  INV_X1 U13485 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10482) );
  INV_X1 U13486 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11563) );
  OAI22_X1 U13487 ( .A1(n10482), .A2(n10481), .B1(n10480), .B2(n11563), .ZN(
        n10483) );
  INV_X1 U13488 ( .A(n10483), .ZN(n10489) );
  AOI22_X1 U13489 ( .A1(n19555), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n19839), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13490 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19725), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13491 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10486) );
  INV_X1 U13492 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11162) );
  INV_X1 U13493 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10490) );
  OAI22_X1 U13494 ( .A1(n11162), .A2(n19584), .B1(n15890), .B2(n10490), .ZN(
        n10492) );
  INV_X1 U13495 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11400) );
  OAI22_X1 U13496 ( .A1(n19829), .A2(n10524), .B1(n19759), .B2(n11400), .ZN(
        n10491) );
  NOR2_X1 U13497 ( .A1(n10492), .A2(n10491), .ZN(n10493) );
  AOI22_X1 U13498 ( .A1(n11080), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13499 ( .A1(n11448), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13500 ( .A1(n11449), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13501 ( .A1(n11451), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10497) );
  NAND4_X1 U13502 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10509) );
  AOI22_X1 U13503 ( .A1(n11077), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10507) );
  NAND2_X1 U13504 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10502) );
  NAND2_X1 U13505 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10501) );
  OAI211_X1 U13506 ( .C1(n11461), .C2(n11160), .A(n10502), .B(n10501), .ZN(
        n10503) );
  INV_X1 U13507 ( .A(n10503), .ZN(n10506) );
  AOI22_X1 U13508 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10505) );
  NAND2_X1 U13509 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10504) );
  NAND4_X1 U13510 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10504), .ZN(
        n10508) );
  NAND2_X1 U13511 ( .A1(n11042), .A2(n11007), .ZN(n10510) );
  INV_X1 U13512 ( .A(n10636), .ZN(n10512) );
  INV_X1 U13513 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10513) );
  INV_X1 U13514 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11420) );
  INV_X1 U13515 ( .A(n10514), .ZN(n10530) );
  AOI22_X1 U13516 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n19839), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10521) );
  INV_X1 U13517 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11579) );
  INV_X1 U13518 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11409) );
  OAI22_X1 U13519 ( .A1(n11579), .A2(n10480), .B1(n10516), .B2(n11409), .ZN(
        n10517) );
  INV_X1 U13520 ( .A(n10517), .ZN(n10520) );
  AOI22_X1 U13521 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19725), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13522 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13523 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19415), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10528) );
  INV_X1 U13524 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11411) );
  INV_X1 U13525 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10523) );
  OAI22_X1 U13526 ( .A1(n11411), .A2(n19584), .B1(n15890), .B2(n10523), .ZN(
        n10526) );
  INV_X1 U13527 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11422) );
  INV_X1 U13528 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11415) );
  OAI22_X1 U13529 ( .A1(n11422), .A2(n10524), .B1(n19759), .B2(n11415), .ZN(
        n10525) );
  NOR2_X1 U13530 ( .A1(n10526), .A2(n10525), .ZN(n10527) );
  NAND3_X1 U13531 ( .A1(n10530), .A2(n10529), .A3(n9796), .ZN(n10545) );
  AOI22_X1 U13532 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11451), .B1(
        n11080), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13533 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10424), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13534 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11463), .B1(
        n11449), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13535 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11448), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10531) );
  NAND4_X1 U13536 ( .A1(n10534), .A2(n10533), .A3(n10532), .A4(n10531), .ZN(
        n10543) );
  AOI22_X1 U13537 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11077), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10541) );
  NAND2_X1 U13538 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10536) );
  NAND2_X1 U13539 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10535) );
  OAI211_X1 U13540 ( .C1(n11461), .C2(n11420), .A(n10536), .B(n10535), .ZN(
        n10537) );
  INV_X1 U13541 ( .A(n10537), .ZN(n10540) );
  AOI22_X1 U13542 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11402), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10539) );
  NAND2_X1 U13543 ( .A1(n11450), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10538) );
  NAND4_X1 U13544 ( .A1(n10541), .A2(n10540), .A3(n10539), .A4(n10538), .ZN(
        n10542) );
  NAND2_X1 U13545 ( .A1(n11046), .A2(n11007), .ZN(n10544) );
  NAND2_X1 U13546 ( .A1(n10545), .A2(n10544), .ZN(n10626) );
  XNOR2_X1 U13547 ( .A(n10551), .B(n10626), .ZN(n10548) );
  NAND2_X1 U13548 ( .A1(n10549), .A2(n9845), .ZN(n10550) );
  NAND2_X1 U13549 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10555) );
  NAND2_X1 U13550 ( .A1(n11448), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10554) );
  NAND2_X1 U13551 ( .A1(n11080), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10553) );
  NAND2_X1 U13552 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10552) );
  AOI22_X1 U13553 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10397), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10560) );
  NAND2_X1 U13554 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10559) );
  AOI22_X1 U13555 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11457), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10558) );
  INV_X1 U13556 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10556) );
  OR2_X1 U13557 ( .A1(n11461), .A2(n10556), .ZN(n10557) );
  NAND2_X1 U13558 ( .A1(n11451), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10564) );
  NAND2_X1 U13559 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10563) );
  NAND2_X1 U13560 ( .A1(n11449), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10562) );
  NAND2_X1 U13561 ( .A1(n11450), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10561) );
  AOI22_X1 U13562 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11456), .B1(
        n11077), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10565) );
  XNOR2_X1 U13563 ( .A(n10572), .B(n10615), .ZN(n10567) );
  NAND2_X1 U13564 ( .A1(n9729), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10571) );
  INV_X1 U13565 ( .A(n10567), .ZN(n10568) );
  NAND2_X1 U13566 ( .A1(n10569), .A2(n10568), .ZN(n10570) );
  NAND2_X1 U13567 ( .A1(n10574), .A2(n11262), .ZN(n10573) );
  NAND3_X1 U13568 ( .A1(n10574), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n11262), .ZN(n10575) );
  AND3_X1 U13569 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15647) );
  NAND2_X1 U13570 ( .A1(n15647), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11241) );
  INV_X1 U13571 ( .A(n11241), .ZN(n15627) );
  NAND2_X1 U13572 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15715) );
  INV_X1 U13573 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10705) );
  NOR2_X1 U13574 ( .A1(n15715), .A2(n10705), .ZN(n10576) );
  AND3_X1 U13575 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15707) );
  AND2_X1 U13576 ( .A1(n10576), .A2(n15707), .ZN(n11240) );
  NAND2_X1 U13577 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15618) );
  INV_X1 U13578 ( .A(n15618), .ZN(n10577) );
  NAND2_X1 U13579 ( .A1(n10577), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11242) );
  NAND2_X1 U13580 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15589) );
  NOR2_X1 U13581 ( .A1(n11242), .A2(n15589), .ZN(n10578) );
  AND3_X1 U13582 ( .A1(n15627), .A2(n11240), .A3(n10578), .ZN(n12901) );
  INV_X1 U13583 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12897) );
  INV_X1 U13584 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21297) );
  INV_X1 U13585 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15301) );
  NAND2_X1 U13586 ( .A1(n20040), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10797) );
  OAI21_X1 U13587 ( .B1(n20040), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10797), .ZN(n10920) );
  MUX2_X1 U13588 ( .A(n10920), .B(n11006), .S(n10263), .Z(n10644) );
  MUX2_X1 U13589 ( .A(n20032), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10919) );
  INV_X1 U13590 ( .A(n10919), .ZN(n10585) );
  INV_X1 U13591 ( .A(n10797), .ZN(n10579) );
  NAND2_X1 U13592 ( .A1(n10919), .A2(n10579), .ZN(n10581) );
  NAND2_X1 U13593 ( .A1(n20032), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10580) );
  NAND2_X1 U13594 ( .A1(n10581), .A2(n10580), .ZN(n10587) );
  XNOR2_X1 U13595 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10586) );
  INV_X1 U13596 ( .A(n10586), .ZN(n10582) );
  XNOR2_X1 U13597 ( .A(n10587), .B(n10582), .ZN(n10918) );
  MUX2_X1 U13598 ( .A(n10918), .B(n10583), .S(n10263), .Z(n10608) );
  INV_X1 U13599 ( .A(n10608), .ZN(n10584) );
  OAI21_X1 U13600 ( .B1(n10644), .B2(n10585), .A(n10584), .ZN(n10603) );
  NAND2_X1 U13601 ( .A1(n10587), .A2(n10586), .ZN(n10589) );
  NAND2_X1 U13602 ( .A1(n20024), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10588) );
  XNOR2_X1 U13603 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10594) );
  INV_X1 U13604 ( .A(n10594), .ZN(n10590) );
  XNOR2_X1 U13605 ( .A(n10595), .B(n10590), .ZN(n10929) );
  NOR2_X1 U13606 ( .A1(n15872), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10593) );
  NOR2_X1 U13607 ( .A1(n16493), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10596) );
  NAND2_X1 U13608 ( .A1(n10598), .A2(n10596), .ZN(n10931) );
  MUX2_X1 U13609 ( .A(n11038), .B(n10931), .S(n10932), .Z(n10614) );
  NAND2_X1 U13610 ( .A1(n10610), .A2(n10614), .ZN(n10916) );
  INV_X1 U13611 ( .A(n10916), .ZN(n10602) );
  NAND2_X1 U13612 ( .A1(n16493), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10597) );
  NAND2_X1 U13613 ( .A1(n10598), .A2(n10597), .ZN(n10600) );
  NAND2_X1 U13614 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13556), .ZN(
        n10599) );
  INV_X1 U13615 ( .A(n10937), .ZN(n10601) );
  AOI21_X1 U13616 ( .B1(n10603), .B2(n10602), .A(n10601), .ZN(n20049) );
  AND2_X1 U13617 ( .A1(n9736), .A2(n11013), .ZN(n10947) );
  NAND2_X1 U13618 ( .A1(n10947), .A2(n10604), .ZN(n10605) );
  NOR2_X1 U13619 ( .A1(n10944), .A2(n10605), .ZN(n16497) );
  NAND2_X1 U13620 ( .A1(n16497), .A2(n11007), .ZN(n20048) );
  INV_X1 U13621 ( .A(n19927), .ZN(n13464) );
  NOR2_X1 U13622 ( .A1(n20048), .A2(n13464), .ZN(n10606) );
  INV_X1 U13623 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14154) );
  NOR2_X1 U13624 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10609) );
  MUX2_X1 U13625 ( .A(n10609), .B(n11017), .S(n19435), .Z(n10648) );
  NAND2_X1 U13626 ( .A1(n10649), .A2(n10648), .ZN(n10641) );
  NAND2_X1 U13627 ( .A1(n10611), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10612) );
  INV_X1 U13628 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13793) );
  MUX2_X1 U13629 ( .A(n10614), .B(n13793), .S(n10611), .Z(n10652) );
  MUX2_X1 U13630 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n11042), .S(n19435), .Z(
        n10637) );
  MUX2_X1 U13631 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n11046), .S(n19435), .Z(
        n10628) );
  INV_X1 U13632 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10831) );
  NOR2_X1 U13633 ( .A1(n19435), .A2(n10831), .ZN(n10662) );
  INV_X1 U13634 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19192) );
  INV_X1 U13635 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13974) );
  NAND2_X1 U13636 ( .A1(n10694), .A2(n10774), .ZN(n10681) );
  NAND2_X1 U13637 ( .A1(n10611), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10618) );
  NAND2_X1 U13638 ( .A1(n10611), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10713) );
  OAI21_X1 U13639 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n10611), .ZN(n10619) );
  INV_X1 U13640 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14261) );
  NAND2_X1 U13641 ( .A1(n10611), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10723) );
  INV_X1 U13642 ( .A(n10723), .ZN(n10620) );
  NOR2_X2 U13643 ( .A1(n10724), .A2(n10620), .ZN(n10697) );
  NAND2_X1 U13644 ( .A1(n10611), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10698) );
  NAND2_X1 U13645 ( .A1(n10697), .A2(n10698), .ZN(n10721) );
  INV_X1 U13646 ( .A(n10721), .ZN(n10623) );
  INV_X1 U13647 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10621) );
  NOR2_X1 U13648 ( .A1(n19435), .A2(n10621), .ZN(n10720) );
  INV_X1 U13649 ( .A(n10720), .ZN(n10622) );
  INV_X1 U13650 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15167) );
  NOR2_X1 U13651 ( .A1(n10748), .A2(n10775), .ZN(n10732) );
  INV_X1 U13652 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n10624) );
  NOR2_X1 U13653 ( .A1(n19435), .A2(n10624), .ZN(n10749) );
  NAND2_X1 U13654 ( .A1(n10611), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10752) );
  INV_X1 U13655 ( .A(n10752), .ZN(n10625) );
  XNOR2_X1 U13656 ( .A(n10753), .B(n10625), .ZN(n15136) );
  NAND3_X1 U13657 ( .A1(n9710), .A2(n10615), .A3(n10626), .ZN(n10634) );
  NAND3_X1 U13658 ( .A1(n10630), .A2(n9754), .A3(n10615), .ZN(n10629) );
  INV_X1 U13659 ( .A(n10628), .ZN(n10665) );
  XNOR2_X1 U13660 ( .A(n10627), .B(n10665), .ZN(n19223) );
  XNOR2_X1 U13661 ( .A(n10661), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14450) );
  AND2_X1 U13662 ( .A1(n10651), .A2(n10637), .ZN(n10638) );
  OR2_X1 U13663 ( .A1(n10638), .A2(n10627), .ZN(n19238) );
  NAND2_X1 U13664 ( .A1(n10639), .A2(n19238), .ZN(n14300) );
  NAND2_X1 U13665 ( .A1(n14300), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10660) );
  NAND2_X1 U13666 ( .A1(n10641), .A2(n10640), .ZN(n10642) );
  NAND2_X1 U13667 ( .A1(n9882), .A2(n10642), .ZN(n14144) );
  MUX2_X1 U13668 ( .A(n10644), .B(n10643), .S(n10611), .Z(n19271) );
  INV_X1 U13669 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10645) );
  NOR2_X1 U13670 ( .A1(n19271), .A2(n10645), .ZN(n13613) );
  INV_X1 U13671 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n19251) );
  NOR3_X1 U13672 ( .A1(n19435), .A2(n10643), .A3(n19251), .ZN(n10646) );
  NOR2_X1 U13673 ( .A1(n10648), .A2(n10646), .ZN(n19254) );
  NAND2_X1 U13674 ( .A1(n13613), .A2(n19254), .ZN(n10647) );
  NOR2_X1 U13675 ( .A1(n13613), .A2(n19254), .ZN(n13612) );
  AOI21_X1 U13676 ( .B1(n15833), .B2(n10647), .A(n13612), .ZN(n13639) );
  XNOR2_X1 U13677 ( .A(n10649), .B(n10648), .ZN(n14158) );
  XNOR2_X1 U13678 ( .A(n14158), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13638) );
  NOR2_X1 U13679 ( .A1(n14158), .A2(n9747), .ZN(n10650) );
  AOI21_X1 U13680 ( .B1(n13639), .B2(n13638), .A(n10650), .ZN(n10654) );
  OAI21_X1 U13681 ( .B1(n10653), .B2(n10652), .A(n10651), .ZN(n15818) );
  AND2_X1 U13682 ( .A1(n15818), .A2(n15826), .ZN(n10655) );
  AOI21_X1 U13683 ( .B1(n10654), .B2(n14164), .A(n10655), .ZN(n10659) );
  INV_X1 U13684 ( .A(n10654), .ZN(n15816) );
  INV_X1 U13685 ( .A(n10655), .ZN(n10656) );
  NAND3_X1 U13686 ( .A1(n15816), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n10656), .ZN(n10657) );
  OAI21_X1 U13687 ( .B1(n15818), .B2(n15826), .A(n10657), .ZN(n10658) );
  AOI21_X1 U13688 ( .B1(n15815), .B2(n10659), .A(n10658), .ZN(n14301) );
  NAND2_X1 U13689 ( .A1(n10661), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15502) );
  NAND2_X1 U13690 ( .A1(n10663), .A2(n10662), .ZN(n10664) );
  NAND2_X1 U13691 ( .A1(n10686), .A2(n10664), .ZN(n14274) );
  NOR2_X1 U13692 ( .A1(n14274), .A2(n10615), .ZN(n10682) );
  AND2_X1 U13693 ( .A1(n10682), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16448) );
  INV_X1 U13694 ( .A(n16448), .ZN(n10669) );
  NAND2_X1 U13695 ( .A1(n10627), .A2(n10665), .ZN(n10668) );
  INV_X1 U13696 ( .A(n10666), .ZN(n10667) );
  XNOR2_X1 U13697 ( .A(n10668), .B(n10667), .ZN(n19213) );
  NAND2_X1 U13698 ( .A1(n19213), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15503) );
  AND2_X1 U13699 ( .A1(n10669), .A2(n15503), .ZN(n10670) );
  AND2_X1 U13700 ( .A1(n15502), .A2(n10670), .ZN(n10671) );
  NAND2_X1 U13701 ( .A1(n10688), .A2(n19192), .ZN(n10675) );
  NOR2_X1 U13702 ( .A1(n10688), .A2(n19192), .ZN(n10672) );
  NAND2_X1 U13703 ( .A1(n10611), .A2(n10672), .ZN(n10673) );
  AND2_X1 U13704 ( .A1(n10774), .A2(n10673), .ZN(n10674) );
  NAND2_X1 U13705 ( .A1(n10675), .A2(n10674), .ZN(n19189) );
  OR2_X1 U13706 ( .A1(n19189), .A2(n10615), .ZN(n10676) );
  INV_X1 U13707 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15777) );
  NAND2_X1 U13708 ( .A1(n10676), .A2(n15777), .ZN(n15774) );
  INV_X1 U13709 ( .A(n19213), .ZN(n10678) );
  INV_X1 U13710 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10677) );
  NAND2_X1 U13711 ( .A1(n10678), .A2(n10677), .ZN(n16445) );
  NAND2_X1 U13712 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n10675), .ZN(n10679) );
  NOR2_X1 U13713 ( .A1(n19435), .A2(n10679), .ZN(n10680) );
  OR2_X1 U13714 ( .A1(n10681), .A2(n10680), .ZN(n19174) );
  INV_X1 U13715 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15749) );
  OAI21_X1 U13716 ( .B1(n19174), .B2(n10615), .A(n15749), .ZN(n15490) );
  INV_X1 U13717 ( .A(n10682), .ZN(n10684) );
  INV_X1 U13718 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10683) );
  NAND2_X1 U13719 ( .A1(n10684), .A2(n10683), .ZN(n16447) );
  NAND4_X1 U13720 ( .A1(n15774), .A2(n16445), .A3(n15490), .A4(n16447), .ZN(
        n10690) );
  INV_X1 U13721 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10685) );
  NOR2_X1 U13722 ( .A1(n19435), .A2(n10685), .ZN(n10687) );
  MUX2_X1 U13723 ( .A(n19435), .B(n10687), .S(n10686), .Z(n10689) );
  NOR2_X1 U13724 ( .A1(n10689), .A2(n10688), .ZN(n19198) );
  AOI21_X1 U13725 ( .B1(n19198), .B2(n11262), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15788) );
  AND2_X1 U13726 ( .A1(n11262), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10692) );
  NAND2_X1 U13727 ( .A1(n19198), .A2(n10692), .ZN(n15786) );
  OR3_X1 U13728 ( .A1(n19189), .A2(n10615), .A3(n15777), .ZN(n15773) );
  NAND2_X1 U13729 ( .A1(n15786), .A2(n15773), .ZN(n15488) );
  NAND2_X1 U13730 ( .A1(n11262), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10693) );
  NOR2_X1 U13731 ( .A1(n19174), .A2(n10693), .ZN(n15491) );
  NAND2_X1 U13732 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n10694), .ZN(n10695) );
  NOR2_X1 U13733 ( .A1(n19435), .A2(n10695), .ZN(n10696) );
  OR2_X1 U13734 ( .A1(n10714), .A2(n10696), .ZN(n19165) );
  INV_X1 U13735 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15742) );
  NOR3_X1 U13736 ( .A1(n19165), .A2(n10615), .A3(n15742), .ZN(n15475) );
  INV_X1 U13737 ( .A(n10697), .ZN(n10700) );
  INV_X1 U13738 ( .A(n10698), .ZN(n10699) );
  NAND2_X1 U13739 ( .A1(n10700), .A2(n10699), .ZN(n10701) );
  NAND2_X1 U13740 ( .A1(n10721), .A2(n10701), .ZN(n19098) );
  OR2_X1 U13741 ( .A1(n19098), .A2(n10615), .ZN(n10737) );
  INV_X1 U13742 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10863) );
  NAND3_X1 U13743 ( .A1(n10710), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n10611), 
        .ZN(n10702) );
  OAI211_X1 U13744 ( .C1(n10710), .C2(P2_EBX_REG_16__SCAN_IN), .A(n10702), .B(
        n10774), .ZN(n19122) );
  OR2_X1 U13745 ( .A1(n19122), .A2(n10615), .ZN(n10739) );
  INV_X1 U13746 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15687) );
  XNOR2_X1 U13747 ( .A(n10739), .B(n15687), .ZN(n15445) );
  NAND2_X1 U13748 ( .A1(n10611), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10703) );
  MUX2_X1 U13749 ( .A(n10703), .B(n10611), .S(n10716), .Z(n10704) );
  INV_X1 U13750 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n14242) );
  NAND2_X1 U13751 ( .A1(n10716), .A2(n14242), .ZN(n10709) );
  INV_X1 U13752 ( .A(n10738), .ZN(n10706) );
  INV_X1 U13753 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10707) );
  NOR2_X1 U13754 ( .A1(n19435), .A2(n10707), .ZN(n10708) );
  NAND2_X1 U13755 ( .A1(n10709), .A2(n10708), .ZN(n10711) );
  NAND2_X1 U13756 ( .A1(n10711), .A2(n10710), .ZN(n19132) );
  OR2_X1 U13757 ( .A1(n19132), .A2(n10615), .ZN(n10712) );
  INV_X1 U13758 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15704) );
  NAND2_X1 U13759 ( .A1(n10712), .A2(n15704), .ZN(n15698) );
  NOR2_X1 U13760 ( .A1(n10714), .A2(n10713), .ZN(n10715) );
  OR2_X1 U13761 ( .A1(n10716), .A2(n10715), .ZN(n19151) );
  INV_X1 U13762 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15723) );
  OAI21_X1 U13763 ( .B1(n19151), .B2(n10615), .A(n15723), .ZN(n15462) );
  INV_X1 U13764 ( .A(n19165), .ZN(n10717) );
  AOI21_X1 U13765 ( .B1(n10717), .B2(n11262), .A(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15477) );
  INV_X1 U13766 ( .A(n15477), .ZN(n10718) );
  NAND3_X1 U13767 ( .A1(n15698), .A2(n15462), .A3(n10718), .ZN(n10719) );
  NOR4_X1 U13768 ( .A1(n15420), .A2(n15445), .A3(n15453), .A4(n10719), .ZN(
        n10726) );
  NAND2_X1 U13769 ( .A1(n10721), .A2(n10720), .ZN(n10722) );
  AND2_X1 U13770 ( .A1(n10728), .A2(n10722), .ZN(n19084) );
  AOI21_X1 U13771 ( .B1(n19084), .B2(n11262), .A(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15385) );
  INV_X1 U13772 ( .A(n15385), .ZN(n15409) );
  XNOR2_X1 U13773 ( .A(n10724), .B(n10723), .ZN(n19110) );
  NAND2_X1 U13774 ( .A1(n19110), .A2(n11262), .ZN(n10725) );
  INV_X1 U13775 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15675) );
  NAND2_X1 U13776 ( .A1(n10725), .A2(n15675), .ZN(n15383) );
  NAND2_X1 U13777 ( .A1(n10611), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10727) );
  XNOR2_X1 U13778 ( .A(n10728), .B(n10727), .ZN(n15177) );
  AOI21_X1 U13779 ( .B1(n15177), .B2(n11262), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15388) );
  NAND3_X1 U13780 ( .A1(n10730), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n10611), 
        .ZN(n10731) );
  AND2_X1 U13781 ( .A1(n10732), .A2(n10731), .ZN(n15159) );
  AOI21_X1 U13782 ( .B1(n15159), .B2(n11262), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15392) );
  INV_X1 U13783 ( .A(n15159), .ZN(n10735) );
  NAND2_X1 U13784 ( .A1(n11262), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10734) );
  NOR2_X1 U13785 ( .A1(n10735), .A2(n10734), .ZN(n15391) );
  AND2_X1 U13786 ( .A1(n11262), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10736) );
  NOR2_X1 U13787 ( .A1(n10737), .A2(n10863), .ZN(n15421) );
  INV_X1 U13788 ( .A(n15421), .ZN(n10746) );
  NAND2_X1 U13789 ( .A1(n10738), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15452) );
  INV_X1 U13790 ( .A(n10739), .ZN(n10740) );
  NAND2_X1 U13791 ( .A1(n10740), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15381) );
  NAND2_X1 U13792 ( .A1(n11262), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10741) );
  NOR2_X1 U13793 ( .A1(n19132), .A2(n10741), .ZN(n15380) );
  INV_X1 U13794 ( .A(n15380), .ZN(n15699) );
  NAND2_X1 U13795 ( .A1(n11262), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10742) );
  NOR2_X1 U13796 ( .A1(n19151), .A2(n10742), .ZN(n15379) );
  INV_X1 U13797 ( .A(n15379), .ZN(n15463) );
  AND4_X1 U13798 ( .A1(n15452), .A2(n15381), .A3(n15699), .A4(n15463), .ZN(
        n10745) );
  AND2_X1 U13799 ( .A1(n11262), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10743) );
  NAND2_X1 U13800 ( .A1(n19110), .A2(n10743), .ZN(n15382) );
  AND2_X1 U13801 ( .A1(n11262), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10744) );
  NAND2_X1 U13802 ( .A1(n19084), .A2(n10744), .ZN(n15408) );
  NAND4_X1 U13803 ( .A1(n10746), .A2(n10745), .A3(n15382), .A4(n15408), .ZN(
        n10747) );
  INV_X1 U13804 ( .A(n10748), .ZN(n10750) );
  AND2_X1 U13805 ( .A1(n10750), .A2(n10749), .ZN(n10751) );
  OR2_X1 U13806 ( .A1(n10753), .A2(n10751), .ZN(n15139) );
  NOR2_X1 U13807 ( .A1(n15139), .A2(n10615), .ZN(n10758) );
  NOR2_X1 U13808 ( .A1(n10758), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11246) );
  NOR2_X2 U13809 ( .A1(n11247), .A2(n11246), .ZN(n15355) );
  OAI21_X1 U13810 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15356), .A(
        n15355), .ZN(n10763) );
  INV_X1 U13811 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15216) );
  NAND2_X1 U13812 ( .A1(n10611), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10754) );
  OAI21_X1 U13813 ( .B1(n10755), .B2(n10754), .A(n10774), .ZN(n10756) );
  OR2_X1 U13814 ( .A1(n10776), .A2(n10756), .ZN(n16405) );
  INV_X1 U13815 ( .A(n16405), .ZN(n10757) );
  NAND2_X1 U13816 ( .A1(n10757), .A2(n11262), .ZN(n10760) );
  NOR2_X1 U13817 ( .A1(n10760), .A2(n12897), .ZN(n15352) );
  NAND2_X1 U13818 ( .A1(n10758), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11245) );
  INV_X1 U13819 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15359) );
  INV_X1 U13820 ( .A(n15356), .ZN(n15360) );
  AOI21_X1 U13821 ( .B1(n11245), .B2(n15359), .A(n15360), .ZN(n10759) );
  NOR2_X1 U13822 ( .A1(n15352), .A2(n10759), .ZN(n10762) );
  INV_X1 U13823 ( .A(n10760), .ZN(n10761) );
  NOR2_X1 U13824 ( .A1(n10761), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15353) );
  INV_X1 U13825 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15207) );
  NAND2_X1 U13826 ( .A1(n10764), .A2(n10774), .ZN(n10769) );
  INV_X1 U13827 ( .A(n10769), .ZN(n11261) );
  NAND3_X1 U13828 ( .A1(n10611), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10765), 
        .ZN(n10766) );
  INV_X1 U13829 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21158) );
  NOR3_X1 U13830 ( .A1(n16395), .A2(n10615), .A3(n21158), .ZN(n10788) );
  INV_X1 U13831 ( .A(n16395), .ZN(n10767) );
  AOI21_X1 U13832 ( .B1(n10767), .B2(n11262), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10768) );
  NAND2_X1 U13833 ( .A1(n10611), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10771) );
  OR2_X1 U13834 ( .A1(n10771), .A2(n10770), .ZN(n10772) );
  AND2_X1 U13835 ( .A1(n10783), .A2(n10772), .ZN(n13444) );
  NAND2_X1 U13836 ( .A1(n13444), .A2(n11262), .ZN(n15308) );
  INV_X1 U13837 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15542) );
  NOR2_X1 U13838 ( .A1(n10776), .A2(n15207), .ZN(n10773) );
  NAND2_X1 U13839 ( .A1(n10611), .A2(n10773), .ZN(n10778) );
  AOI21_X1 U13840 ( .B1(n10776), .B2(n15207), .A(n10775), .ZN(n10777) );
  NOR2_X1 U13841 ( .A1(n10786), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15340) );
  AOI21_X1 U13842 ( .B1(n15308), .B2(n15542), .A(n15340), .ZN(n10779) );
  INV_X1 U13843 ( .A(n10779), .ZN(n10780) );
  INV_X1 U13844 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15102) );
  NOR2_X1 U13845 ( .A1(n10257), .A2(n15102), .ZN(n10782) );
  AND2_X1 U13846 ( .A1(n10783), .A2(n10782), .ZN(n10784) );
  NOR2_X1 U13847 ( .A1(n10791), .A2(n10784), .ZN(n15106) );
  NAND2_X1 U13848 ( .A1(n15106), .A2(n11262), .ZN(n15311) );
  INV_X1 U13849 ( .A(n15311), .ZN(n10785) );
  INV_X1 U13850 ( .A(n10786), .ZN(n10787) );
  NOR2_X1 U13851 ( .A1(n10787), .A2(n21297), .ZN(n15339) );
  NOR2_X1 U13852 ( .A1(n15339), .A2(n10788), .ZN(n15306) );
  NAND2_X1 U13853 ( .A1(n10611), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10790) );
  XNOR2_X1 U13854 ( .A(n10791), .B(n10790), .ZN(n10789) );
  OAI21_X1 U13855 ( .B1(n10789), .B2(n10615), .A(n15301), .ZN(n15292) );
  NAND2_X1 U13856 ( .A1(n15294), .A2(n15292), .ZN(n11258) );
  INV_X1 U13857 ( .A(n10789), .ZN(n15083) );
  NAND3_X1 U13858 ( .A1(n15083), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11262), .ZN(n15293) );
  NAND2_X1 U13859 ( .A1(n11258), .A2(n15293), .ZN(n10796) );
  NAND2_X1 U13860 ( .A1(n10791), .A2(n10790), .ZN(n11259) );
  INV_X1 U13861 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12972) );
  NOR2_X1 U13862 ( .A1(n10257), .A2(n12972), .ZN(n10792) );
  XNOR2_X1 U13863 ( .A(n11259), .B(n10792), .ZN(n12975) );
  INV_X1 U13864 ( .A(n12975), .ZN(n10793) );
  AOI21_X1 U13865 ( .B1(n10793), .B2(n11262), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11257) );
  INV_X1 U13866 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15519) );
  INV_X1 U13867 ( .A(n11256), .ZN(n10794) );
  NOR2_X1 U13868 ( .A1(n11257), .A2(n10794), .ZN(n10795) );
  NAND3_X1 U13869 ( .A1(n10931), .A2(n10929), .A3(n10918), .ZN(n10800) );
  XNOR2_X1 U13870 ( .A(n10919), .B(n10797), .ZN(n10921) );
  INV_X1 U13871 ( .A(n10800), .ZN(n10798) );
  NAND2_X1 U13872 ( .A1(n10921), .A2(n10798), .ZN(n10799) );
  OAI211_X1 U13873 ( .C1(n10920), .C2(n10800), .A(n19921), .B(n11635), .ZN(
        n10804) );
  INV_X1 U13874 ( .A(n10801), .ZN(n15869) );
  NAND2_X1 U13875 ( .A1(n15869), .A2(n13556), .ZN(n13553) );
  INV_X1 U13876 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13551) );
  OAI21_X1 U13877 ( .B1(n11080), .B2(n13553), .A(n13551), .ZN(n10802) );
  AND2_X1 U13878 ( .A1(n10802), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20037) );
  INV_X1 U13879 ( .A(n20037), .ZN(n10803) );
  NAND3_X1 U13880 ( .A1(n10805), .A2(n10263), .A3(n19927), .ZN(n10806) );
  OR2_X1 U13881 ( .A1(n10944), .A2(n10806), .ZN(n10807) );
  AOI22_X1 U13882 ( .A1(n11270), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10809) );
  OAI21_X1 U13883 ( .B1(n10808), .B2(n12972), .A(n10809), .ZN(n10810) );
  AOI21_X1 U13884 ( .B1(n10886), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10810), .ZN(n10902) );
  INV_X1 U13885 ( .A(n10811), .ZN(n10812) );
  OR2_X1 U13886 ( .A1(n9771), .A2(n15826), .ZN(n10816) );
  AOI22_X1 U13887 ( .A1(n11270), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10815) );
  OAI211_X1 U13888 ( .C1(n13793), .C2(n10808), .A(n10816), .B(n10815), .ZN(
        n13790) );
  NAND2_X1 U13889 ( .A1(n13791), .A2(n13790), .ZN(n13809) );
  INV_X1 U13890 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10990) );
  OR2_X1 U13891 ( .A1(n9771), .A2(n10990), .ZN(n10820) );
  NAND2_X1 U13892 ( .A1(n10292), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13893 ( .A1(n11270), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10817) );
  AND2_X1 U13894 ( .A1(n10818), .A2(n10817), .ZN(n10819) );
  INV_X1 U13895 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16464) );
  OR2_X1 U13896 ( .A1(n9771), .A2(n16464), .ZN(n10824) );
  NAND2_X1 U13897 ( .A1(n11271), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13898 ( .A1(n11270), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10821) );
  AND2_X1 U13899 ( .A1(n10822), .A2(n10821), .ZN(n10823) );
  NAND2_X1 U13900 ( .A1(n10824), .A2(n10823), .ZN(n13895) );
  OR2_X1 U13901 ( .A1(n9771), .A2(n10677), .ZN(n10828) );
  NAND2_X1 U13902 ( .A1(n10292), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13903 ( .A1(n11270), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10825) );
  AND2_X1 U13904 ( .A1(n10826), .A2(n10825), .ZN(n10827) );
  NAND2_X1 U13905 ( .A1(n10828), .A2(n10827), .ZN(n13930) );
  NAND2_X1 U13906 ( .A1(n10886), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10830) );
  AOI22_X1 U13907 ( .A1(n11270), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10829) );
  OAI211_X1 U13908 ( .C1(n10831), .C2(n10808), .A(n10830), .B(n10829), .ZN(
        n13921) );
  INV_X1 U13909 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15793) );
  OR2_X1 U13910 ( .A1(n9771), .A2(n15793), .ZN(n10835) );
  NAND2_X1 U13911 ( .A1(n11271), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13912 ( .A1(n11270), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10832) );
  AND2_X1 U13913 ( .A1(n10833), .A2(n10832), .ZN(n10834) );
  OR2_X1 U13914 ( .A1(n9771), .A2(n15777), .ZN(n10838) );
  INV_X1 U13915 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19188) );
  OAI22_X1 U13916 ( .A1(n10896), .A2(n19188), .B1(n19921), .B2(n10906), .ZN(
        n10836) );
  AOI21_X1 U13917 ( .B1(n11271), .B2(P2_EBX_REG_10__SCAN_IN), .A(n10836), .ZN(
        n10837) );
  OR2_X1 U13918 ( .A1(n9771), .A2(n15749), .ZN(n10841) );
  INV_X1 U13919 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19965) );
  OAI22_X1 U13920 ( .A1(n10896), .A2(n19965), .B1(n19921), .B2(n19184), .ZN(
        n10839) );
  AOI21_X1 U13921 ( .B1(n10292), .B2(P2_EBX_REG_11__SCAN_IN), .A(n10839), .ZN(
        n10840) );
  NAND2_X1 U13922 ( .A1(n10841), .A2(n10840), .ZN(n13970) );
  OR2_X1 U13923 ( .A1(n9771), .A2(n15742), .ZN(n10845) );
  INV_X1 U13924 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19967) );
  INV_X1 U13925 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10842) );
  OAI22_X1 U13926 ( .A1(n10896), .A2(n19967), .B1(n19921), .B2(n10842), .ZN(
        n10843) );
  AOI21_X1 U13927 ( .B1(n11271), .B2(P2_EBX_REG_12__SCAN_IN), .A(n10843), .ZN(
        n10844) );
  OR2_X1 U13928 ( .A1(n9771), .A2(n15723), .ZN(n10848) );
  INV_X1 U13929 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n21161) );
  INV_X1 U13930 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19161) );
  OAI22_X1 U13931 ( .A1(n10896), .A2(n21161), .B1(n19921), .B2(n19161), .ZN(
        n10846) );
  AOI21_X1 U13932 ( .B1(n11271), .B2(P2_EBX_REG_13__SCAN_IN), .A(n10846), .ZN(
        n10847) );
  AOI22_X1 U13933 ( .A1(n11270), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10849) );
  OAI21_X1 U13934 ( .B1(n10808), .B2(n14242), .A(n10849), .ZN(n10850) );
  AOI21_X1 U13935 ( .B1(n10886), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10850), .ZN(n14239) );
  OR2_X1 U13936 ( .A1(n9771), .A2(n15704), .ZN(n10854) );
  NAND2_X1 U13937 ( .A1(n11271), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13938 ( .A1(n11270), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10851) );
  AND2_X1 U13939 ( .A1(n10852), .A2(n10851), .ZN(n10853) );
  NAND2_X1 U13940 ( .A1(n10854), .A2(n10853), .ZN(n14206) );
  NAND2_X1 U13941 ( .A1(n14204), .A2(n14206), .ZN(n14205) );
  OR2_X1 U13942 ( .A1(n9771), .A2(n15687), .ZN(n10858) );
  INV_X1 U13943 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n10855) );
  OAI22_X1 U13944 ( .A1(n10896), .A2(n10855), .B1(n19921), .B2(n9897), .ZN(
        n10856) );
  AOI21_X1 U13945 ( .B1(n11271), .B2(P2_EBX_REG_16__SCAN_IN), .A(n10856), .ZN(
        n10857) );
  OR2_X1 U13946 ( .A1(n9771), .A2(n15675), .ZN(n10861) );
  INV_X1 U13947 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n15436) );
  INV_X1 U13948 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n21218) );
  OAI22_X1 U13949 ( .A1(n10896), .A2(n15436), .B1(n19921), .B2(n21218), .ZN(
        n10859) );
  AOI21_X1 U13950 ( .B1(n11271), .B2(P2_EBX_REG_17__SCAN_IN), .A(n10859), .ZN(
        n10860) );
  OR2_X1 U13951 ( .A1(n9771), .A2(n10863), .ZN(n10866) );
  INV_X1 U13952 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19974) );
  OAI22_X1 U13953 ( .A1(n10896), .A2(n19974), .B1(n19921), .B2(n9903), .ZN(
        n10864) );
  AOI21_X1 U13954 ( .B1(n11271), .B2(P2_EBX_REG_18__SCAN_IN), .A(n10864), .ZN(
        n10865) );
  NAND2_X1 U13955 ( .A1(n10866), .A2(n10865), .ZN(n14386) );
  INV_X1 U13956 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21279) );
  OR2_X1 U13957 ( .A1(n9771), .A2(n21279), .ZN(n10869) );
  INV_X1 U13958 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19976) );
  INV_X1 U13959 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15413) );
  OAI22_X1 U13960 ( .A1(n10896), .A2(n19976), .B1(n19921), .B2(n15413), .ZN(
        n10867) );
  AOI21_X1 U13961 ( .B1(n11271), .B2(P2_EBX_REG_19__SCAN_IN), .A(n10867), .ZN(
        n10868) );
  NAND2_X1 U13962 ( .A1(n10869), .A2(n10868), .ZN(n15239) );
  AOI22_X1 U13963 ( .A1(n11270), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10870) );
  OAI21_X1 U13964 ( .B1(n10808), .B2(n15167), .A(n10870), .ZN(n10871) );
  AOI21_X1 U13965 ( .B1(n10886), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10871), .ZN(n15162) );
  INV_X1 U13966 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10914) );
  OR2_X1 U13967 ( .A1(n9771), .A2(n10914), .ZN(n10874) );
  INV_X1 U13968 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19979) );
  INV_X1 U13969 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15396) );
  OAI22_X1 U13970 ( .A1(n10896), .A2(n19979), .B1(n19921), .B2(n15396), .ZN(
        n10872) );
  AOI21_X1 U13971 ( .B1(n11271), .B2(P2_EBX_REG_21__SCAN_IN), .A(n10872), .ZN(
        n10873) );
  INV_X1 U13972 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10915) );
  OR2_X1 U13973 ( .A1(n9771), .A2(n10915), .ZN(n10877) );
  INV_X1 U13974 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19980) );
  INV_X1 U13975 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15138) );
  OAI22_X1 U13976 ( .A1(n10896), .A2(n19980), .B1(n19921), .B2(n15138), .ZN(
        n10875) );
  AOI21_X1 U13977 ( .B1(n11271), .B2(P2_EBX_REG_22__SCAN_IN), .A(n10875), .ZN(
        n10876) );
  NAND2_X1 U13978 ( .A1(n10877), .A2(n10876), .ZN(n11231) );
  OR2_X1 U13979 ( .A1(n9771), .A2(n15359), .ZN(n10880) );
  INV_X1 U13980 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19982) );
  INV_X1 U13981 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15371) );
  OAI22_X1 U13982 ( .A1(n10896), .A2(n19982), .B1(n19921), .B2(n15371), .ZN(
        n10878) );
  AOI21_X1 U13983 ( .B1(n11271), .B2(P2_EBX_REG_23__SCAN_IN), .A(n10878), .ZN(
        n10879) );
  NAND2_X1 U13984 ( .A1(n10880), .A2(n10879), .ZN(n15123) );
  OR2_X1 U13985 ( .A1(n9771), .A2(n12897), .ZN(n10883) );
  INV_X1 U13986 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19984) );
  OAI22_X1 U13987 ( .A1(n10896), .A2(n19984), .B1(n19921), .B2(n9905), .ZN(
        n10881) );
  AOI21_X1 U13988 ( .B1(n11271), .B2(P2_EBX_REG_24__SCAN_IN), .A(n10881), .ZN(
        n10882) );
  AND2_X1 U13989 ( .A1(n10883), .A2(n10882), .ZN(n15215) );
  AOI22_X1 U13990 ( .A1(n11270), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10884) );
  OAI21_X1 U13991 ( .B1(n10808), .B2(n15207), .A(n10884), .ZN(n10885) );
  AOI21_X1 U13992 ( .B1(n10886), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10885), .ZN(n15109) );
  OR2_X1 U13993 ( .A1(n9771), .A2(n21158), .ZN(n10889) );
  INV_X1 U13994 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n15333) );
  INV_X1 U13995 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16390) );
  OAI22_X1 U13996 ( .A1(n10896), .A2(n15333), .B1(n19921), .B2(n16390), .ZN(
        n10887) );
  AOI21_X1 U13997 ( .B1(n11271), .B2(P2_EBX_REG_26__SCAN_IN), .A(n10887), .ZN(
        n10888) );
  NAND2_X1 U13998 ( .A1(n10889), .A2(n10888), .ZN(n15199) );
  OR2_X1 U13999 ( .A1(n9771), .A2(n15542), .ZN(n10892) );
  INV_X1 U14000 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19989) );
  INV_X1 U14001 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15322) );
  OAI22_X1 U14002 ( .A1(n10896), .A2(n19989), .B1(n19921), .B2(n15322), .ZN(
        n10890) );
  AOI21_X1 U14003 ( .B1(n11271), .B2(P2_EBX_REG_27__SCAN_IN), .A(n10890), .ZN(
        n10891) );
  NAND2_X1 U14004 ( .A1(n10892), .A2(n10891), .ZN(n13447) );
  NAND2_X1 U14005 ( .A1(n15201), .A2(n13447), .ZN(n13446) );
  OR2_X1 U14006 ( .A1(n9771), .A2(n10781), .ZN(n10895) );
  INV_X1 U14007 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n21168) );
  OAI22_X1 U14008 ( .A1(n10896), .A2(n21168), .B1(n19921), .B2(n9908), .ZN(
        n10893) );
  AOI21_X1 U14009 ( .B1(n11271), .B2(P2_EBX_REG_28__SCAN_IN), .A(n10893), .ZN(
        n10894) );
  AND2_X1 U14010 ( .A1(n10895), .A2(n10894), .ZN(n15091) );
  OR2_X1 U14011 ( .A1(n9771), .A2(n15301), .ZN(n10899) );
  INV_X1 U14012 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19991) );
  INV_X1 U14013 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15296) );
  OAI22_X1 U14014 ( .A1(n10896), .A2(n19991), .B1(n19921), .B2(n15296), .ZN(
        n10897) );
  AOI21_X1 U14015 ( .B1(n11271), .B2(P2_EBX_REG_29__SCAN_IN), .A(n10897), .ZN(
        n10898) );
  AND2_X1 U14016 ( .A1(n10899), .A2(n10898), .ZN(n15078) );
  INV_X1 U14017 ( .A(n15078), .ZN(n10900) );
  NOR2_X2 U14018 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20004) );
  NAND2_X1 U14019 ( .A1(n19921), .A2(n20033), .ZN(n20006) );
  INV_X1 U14020 ( .A(n20006), .ZN(n15858) );
  OR2_X1 U14021 ( .A1(n20004), .A2(n15858), .ZN(n20007) );
  INV_X1 U14022 ( .A(n20007), .ZN(n20034) );
  INV_X1 U14023 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19691) );
  NOR2_X1 U14024 ( .A1(n19921), .A2(n19691), .ZN(n20025) );
  INV_X1 U14025 ( .A(n11299), .ZN(n10904) );
  NAND2_X1 U14026 ( .A1(n19691), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10903) );
  NAND2_X1 U14027 ( .A1(n10904), .A2(n10903), .ZN(n13621) );
  NAND2_X1 U14028 ( .A1(n12930), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12929) );
  INV_X1 U14029 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15343) );
  XOR2_X1 U14030 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n9831), .Z(n12956) );
  INV_X1 U14031 ( .A(n12956), .ZN(n10910) );
  INV_X2 U14032 ( .A(n19214), .ZN(n19399) );
  NAND2_X1 U14033 ( .A1(n19399), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15518) );
  NAND2_X1 U14034 ( .A1(n16442), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10909) );
  OAI211_X1 U14035 ( .C1(n16455), .C2(n10910), .A(n15518), .B(n10909), .ZN(
        n10911) );
  AOI21_X1 U14036 ( .B1(n15515), .B2(n19403), .A(n10911), .ZN(n10912) );
  NAND2_X1 U14037 ( .A1(n15377), .A2(n10915), .ZN(n12346) );
  NAND2_X1 U14038 ( .A1(n10916), .A2(n10932), .ZN(n10935) );
  INV_X1 U14039 ( .A(n13571), .ZN(n10917) );
  MUX2_X1 U14040 ( .A(n10917), .B(n10932), .S(n10918), .Z(n10928) );
  INV_X1 U14041 ( .A(n10918), .ZN(n10925) );
  OAI21_X1 U14042 ( .B1(n10920), .B2(n10585), .A(n10263), .ZN(n10924) );
  INV_X1 U14043 ( .A(n10920), .ZN(n10922) );
  OAI211_X1 U14044 ( .C1(n11284), .C2(n10922), .A(n9722), .B(n10921), .ZN(
        n10923) );
  OAI211_X1 U14045 ( .C1(n10926), .C2(n10925), .A(n10924), .B(n10923), .ZN(
        n10927) );
  OAI21_X1 U14046 ( .B1(n10928), .B2(n11007), .A(n10927), .ZN(n10930) );
  NAND2_X1 U14047 ( .A1(n10930), .A2(n10929), .ZN(n10934) );
  OAI21_X1 U14048 ( .B1(n10932), .B2(n10931), .A(n10937), .ZN(n10933) );
  AOI21_X1 U14049 ( .B1(n10935), .B2(n10934), .A(n10933), .ZN(n10936) );
  MUX2_X1 U14050 ( .A(n13556), .B(n10936), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n10961) );
  INV_X1 U14051 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19052) );
  INV_X1 U14052 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19950) );
  NOR2_X1 U14053 ( .A1(n19052), .A2(n19950), .ZN(n19941) );
  NOR2_X1 U14054 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19943) );
  NOR3_X1 U14055 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19941), .A3(n19943), 
        .ZN(n19935) );
  NAND2_X1 U14056 ( .A1(n19935), .A2(n11284), .ZN(n10939) );
  OR2_X1 U14057 ( .A1(n16501), .A2(n10939), .ZN(n13548) );
  NAND2_X1 U14058 ( .A1(n11635), .A2(n11007), .ZN(n10940) );
  AOI21_X1 U14059 ( .B1(n13548), .B2(n10940), .A(n10604), .ZN(n10943) );
  NOR2_X1 U14060 ( .A1(n16502), .A2(n10941), .ZN(n13467) );
  AND2_X1 U14061 ( .A1(n13467), .A2(n11284), .ZN(n10942) );
  NAND2_X1 U14062 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19922) );
  OAI21_X1 U14063 ( .B1(n10943), .B2(n10942), .A(n19922), .ZN(n10968) );
  INV_X1 U14064 ( .A(n20045), .ZN(n10960) );
  NOR2_X1 U14065 ( .A1(n10944), .A2(n11007), .ZN(n10959) );
  INV_X1 U14066 ( .A(n19922), .ZN(n19942) );
  INV_X1 U14067 ( .A(n19935), .ZN(n15068) );
  NOR2_X1 U14068 ( .A1(n19942), .A2(n15068), .ZN(n13458) );
  INV_X1 U14069 ( .A(n11013), .ZN(n11676) );
  OR2_X1 U14070 ( .A1(n10945), .A2(n11676), .ZN(n10946) );
  NAND2_X1 U14071 ( .A1(n11007), .A2(n9736), .ZN(n12961) );
  INV_X1 U14072 ( .A(n12961), .ZN(n15067) );
  NAND2_X1 U14073 ( .A1(n10946), .A2(n15067), .ZN(n10971) );
  INV_X1 U14074 ( .A(n10947), .ZN(n10948) );
  OAI211_X1 U14075 ( .C1(n9746), .C2(n11284), .A(n10948), .B(n10604), .ZN(
        n10950) );
  NAND4_X1 U14076 ( .A1(n10971), .A2(n10981), .A3(n10951), .A4(n10950), .ZN(
        n10952) );
  AOI21_X1 U14077 ( .B1(n13467), .B2(n13458), .A(n10952), .ZN(n10958) );
  NAND2_X1 U14078 ( .A1(n10955), .A2(n10604), .ZN(n10956) );
  NAND2_X1 U14079 ( .A1(n10954), .A2(n10956), .ZN(n10957) );
  NAND2_X1 U14080 ( .A1(n10958), .A2(n10957), .ZN(n13543) );
  AOI21_X1 U14081 ( .B1(n10960), .B2(n10959), .A(n13543), .ZN(n10967) );
  INV_X1 U14082 ( .A(n10962), .ZN(n10963) );
  OAI21_X1 U14083 ( .B1(n16501), .B2(n11007), .A(n10963), .ZN(n10966) );
  INV_X1 U14084 ( .A(n20048), .ZN(n10964) );
  NAND2_X1 U14085 ( .A1(n20049), .A2(n10964), .ZN(n10965) );
  NAND4_X1 U14086 ( .A1(n10968), .A2(n10967), .A3(n10966), .A4(n10965), .ZN(
        n10969) );
  AOI21_X1 U14087 ( .B1(n15843), .B2(n10971), .A(n10970), .ZN(n10979) );
  NOR2_X1 U14088 ( .A1(n10973), .A2(n10972), .ZN(n11637) );
  INV_X1 U14089 ( .A(n11637), .ZN(n10977) );
  NAND2_X1 U14090 ( .A1(n10981), .A2(n10202), .ZN(n10974) );
  INV_X1 U14091 ( .A(n9750), .ZN(n13462) );
  AOI22_X1 U14092 ( .A1(n10974), .A2(n13462), .B1(n9736), .B2(n10240), .ZN(
        n10976) );
  NAND3_X1 U14093 ( .A1(n10977), .A2(n10976), .A3(n10975), .ZN(n10978) );
  NOR2_X1 U14094 ( .A1(n10979), .A2(n10978), .ZN(n10980) );
  OAI21_X1 U14095 ( .B1(n10982), .B2(n10981), .A(n10980), .ZN(n15863) );
  NOR2_X1 U14096 ( .A1(n15863), .A2(n11629), .ZN(n10983) );
  NAND2_X1 U14097 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15831) );
  NOR2_X1 U14098 ( .A1(n9747), .A2(n15831), .ZN(n11237) );
  NAND2_X1 U14099 ( .A1(n11249), .A2(n19214), .ZN(n16469) );
  OAI21_X1 U14100 ( .B1(n15667), .B2(n11237), .A(n16469), .ZN(n10984) );
  INV_X1 U14101 ( .A(n10984), .ZN(n10988) );
  AND3_X1 U14102 ( .A1(n10604), .A2(n11007), .A3(n19435), .ZN(n10986) );
  NAND2_X1 U14103 ( .A1(n9749), .A2(n10986), .ZN(n16505) );
  AND2_X1 U14104 ( .A1(n15831), .A2(n9747), .ZN(n10987) );
  NAND2_X1 U14105 ( .A1(n15663), .A2(n10987), .ZN(n13643) );
  AND2_X1 U14106 ( .A1(n10988), .A2(n13643), .ZN(n14162) );
  NAND2_X1 U14107 ( .A1(n15832), .A2(n14164), .ZN(n10989) );
  NAND2_X1 U14108 ( .A1(n14162), .A2(n10989), .ZN(n15822) );
  NOR2_X1 U14109 ( .A1(n10990), .A2(n15826), .ZN(n11238) );
  INV_X1 U14110 ( .A(n11238), .ZN(n14343) );
  OR2_X1 U14111 ( .A1(n15822), .A2(n14343), .ZN(n10991) );
  NAND2_X1 U14112 ( .A1(n15708), .A2(n10991), .ZN(n16456) );
  NAND3_X1 U14113 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U14114 ( .A1(n15832), .A2(n11239), .ZN(n10992) );
  NAND2_X1 U14115 ( .A1(n16456), .A2(n10992), .ZN(n15792) );
  INV_X1 U14116 ( .A(n11240), .ZN(n10993) );
  NOR2_X1 U14117 ( .A1(n15792), .A2(n10993), .ZN(n15664) );
  NOR2_X1 U14118 ( .A1(n11241), .A2(n11242), .ZN(n10995) );
  INV_X1 U14119 ( .A(n15792), .ZN(n10994) );
  AOI22_X1 U14120 ( .A1(n15664), .A2(n10995), .B1(n16482), .B2(n10994), .ZN(
        n15621) );
  AND2_X1 U14121 ( .A1(n10998), .A2(n9749), .ZN(n16503) );
  AOI21_X1 U14122 ( .B1(n11284), .B2(n10997), .A(n16503), .ZN(n10999) );
  AND2_X1 U14123 ( .A1(n11013), .A2(n11002), .ZN(n11000) );
  NAND2_X1 U14124 ( .A1(n11001), .A2(n11000), .ZN(n11133) );
  INV_X2 U14125 ( .A(n11133), .ZN(n11053) );
  NAND2_X1 U14126 ( .A1(n11053), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11003) );
  INV_X1 U14127 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13499) );
  MUX2_X1 U14128 ( .A(n11013), .B(n20040), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11005) );
  NAND2_X1 U14129 ( .A1(n11639), .A2(n11032), .ZN(n11024) );
  AND2_X1 U14130 ( .A1(n11005), .A2(n11024), .ZN(n11012) );
  INV_X1 U14131 ( .A(n11006), .ZN(n11010) );
  NAND2_X2 U14132 ( .A1(n11008), .A2(n11007), .ZN(n11212) );
  NAND2_X1 U14133 ( .A1(n11010), .A2(n11009), .ZN(n11011) );
  NAND2_X1 U14134 ( .A1(n11012), .A2(n11011), .ZN(n13605) );
  AND2_X2 U14135 ( .A1(n13604), .A2(n13605), .ZN(n13607) );
  NAND2_X1 U14136 ( .A1(n11053), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11015) );
  NOR2_X1 U14137 ( .A1(n11013), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U14138 ( .A1(n11026), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11014) );
  NAND2_X1 U14139 ( .A1(n11015), .A2(n11014), .ZN(n11020) );
  NAND2_X1 U14140 ( .A1(n10231), .A2(n11013), .ZN(n11016) );
  MUX2_X1 U14141 ( .A(n11016), .B(n20032), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11019) );
  NAND2_X1 U14142 ( .A1(n11009), .A2(n11017), .ZN(n11018) );
  NAND2_X1 U14143 ( .A1(n11019), .A2(n11018), .ZN(n13827) );
  NOR2_X1 U14144 ( .A1(n13828), .A2(n13827), .ZN(n11022) );
  NOR2_X1 U14145 ( .A1(n13607), .A2(n11020), .ZN(n11021) );
  NAND2_X1 U14146 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11023) );
  OAI211_X1 U14147 ( .C1(n11212), .C2(n11025), .A(n11024), .B(n11023), .ZN(
        n11030) );
  NAND2_X1 U14148 ( .A1(n11053), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U14149 ( .A1(n12889), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11027) );
  NAND2_X1 U14150 ( .A1(n11028), .A2(n11027), .ZN(n13629) );
  NOR2_X1 U14151 ( .A1(n11029), .A2(n11030), .ZN(n11031) );
  NAND2_X1 U14152 ( .A1(n11053), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U14153 ( .A1(n11032), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11036) );
  NAND2_X1 U14154 ( .A1(n11009), .A2(n11033), .ZN(n11035) );
  NAND2_X1 U14155 ( .A1(n12889), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11034) );
  NAND4_X1 U14156 ( .A1(n11037), .A2(n11036), .A3(n11035), .A4(n11034), .ZN(
        n14110) );
  NAND2_X1 U14157 ( .A1(n11053), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U14158 ( .A1(n12889), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11040) );
  NAND2_X1 U14159 ( .A1(n11009), .A2(n11038), .ZN(n11039) );
  INV_X1 U14160 ( .A(n11042), .ZN(n11043) );
  AOI22_X1 U14161 ( .A1(n11053), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11009), 
        .B2(n11043), .ZN(n11045) );
  AOI22_X1 U14162 ( .A1(n12889), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11044) );
  NAND2_X1 U14163 ( .A1(n11045), .A2(n11044), .ZN(n14342) );
  NAND2_X1 U14164 ( .A1(n14340), .A2(n14342), .ZN(n14341) );
  INV_X1 U14165 ( .A(n11046), .ZN(n11047) );
  NAND2_X1 U14166 ( .A1(n11009), .A2(n11047), .ZN(n11048) );
  NAND2_X1 U14167 ( .A1(n11053), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U14168 ( .A1(n12889), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11049) );
  NAND2_X1 U14169 ( .A1(n11050), .A2(n11049), .ZN(n14459) );
  NAND2_X1 U14170 ( .A1(n14458), .A2(n14459), .ZN(n11052) );
  NAND2_X1 U14171 ( .A1(n11009), .A2(n11262), .ZN(n11051) );
  NAND2_X1 U14172 ( .A1(n11053), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14173 ( .A1(n12889), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11054) );
  NAND2_X1 U14174 ( .A1(n11055), .A2(n11054), .ZN(n15803) );
  AOI22_X1 U14175 ( .A1(n11451), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14176 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11449), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14177 ( .A1(n11080), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U14178 ( .A1(n11448), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11056) );
  NAND4_X1 U14179 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n11069) );
  AOI22_X1 U14180 ( .A1(n11077), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11067) );
  INV_X1 U14181 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11062) );
  NAND2_X1 U14182 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11061) );
  NAND2_X1 U14183 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11060) );
  OAI211_X1 U14184 ( .C1(n11461), .C2(n11062), .A(n11061), .B(n11060), .ZN(
        n11063) );
  INV_X1 U14185 ( .A(n11063), .ZN(n11066) );
  AOI22_X1 U14186 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11065) );
  NAND2_X1 U14187 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11064) );
  NAND4_X1 U14188 ( .A1(n11067), .A2(n11066), .A3(n11065), .A4(n11064), .ZN(
        n11068) );
  INV_X1 U14189 ( .A(n11314), .ZN(n13922) );
  AOI22_X1 U14190 ( .A1(n12889), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11070) );
  OAI21_X1 U14191 ( .B1(n13922), .B2(n11212), .A(n11070), .ZN(n11071) );
  AOI21_X1 U14192 ( .B1(n11053), .B2(P2_REIP_REG_8__SCAN_IN), .A(n11071), .ZN(
        n14264) );
  AOI22_X1 U14193 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10397), .B1(
        n11457), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14194 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10369), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11075) );
  INV_X1 U14195 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11072) );
  OR2_X1 U14196 ( .A1(n11461), .A2(n11072), .ZN(n11074) );
  NAND2_X1 U14197 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11073) );
  NAND4_X1 U14198 ( .A1(n11076), .A2(n11075), .A3(n11074), .A4(n11073), .ZN(
        n11079) );
  INV_X1 U14199 ( .A(n11456), .ZN(n15871) );
  INV_X1 U14200 ( .A(n11077), .ZN(n11421) );
  INV_X1 U14201 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14009) );
  OAI22_X1 U14202 ( .A1(n14074), .A2(n15871), .B1(n11421), .B2(n14009), .ZN(
        n11078) );
  NOR2_X1 U14203 ( .A1(n11079), .A2(n11078), .ZN(n11091) );
  INV_X1 U14204 ( .A(n11080), .ZN(n11159) );
  INV_X1 U14205 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11481) );
  OAI22_X1 U14206 ( .A1(n19814), .A2(n11177), .B1(n11159), .B2(n11481), .ZN(
        n11084) );
  INV_X1 U14207 ( .A(n11451), .ZN(n11163) );
  OAI22_X1 U14208 ( .A1(n11163), .A2(n11082), .B1(n11161), .B2(n11081), .ZN(
        n11083) );
  NOR2_X1 U14209 ( .A1(n11084), .A2(n11083), .ZN(n11090) );
  INV_X1 U14210 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11474) );
  INV_X1 U14211 ( .A(n11448), .ZN(n11166) );
  OAI22_X1 U14212 ( .A1(n11474), .A2(n11166), .B1(n11178), .B2(n11339), .ZN(
        n11088) );
  INV_X1 U14213 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11086) );
  INV_X1 U14214 ( .A(n11449), .ZN(n11169) );
  INV_X1 U14215 ( .A(n11450), .ZN(n11168) );
  INV_X1 U14216 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11085) );
  OAI22_X1 U14217 ( .A1(n11086), .A2(n11169), .B1(n11168), .B2(n11085), .ZN(
        n11087) );
  NOR2_X1 U14218 ( .A1(n11088), .A2(n11087), .ZN(n11089) );
  NAND2_X1 U14219 ( .A1(n11053), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U14220 ( .A1(n12889), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11092) );
  OAI211_X1 U14221 ( .C1(n13855), .C2(n11212), .A(n11093), .B(n11092), .ZN(
        n15795) );
  AOI22_X1 U14222 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10397), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14223 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10369), .B1(
        n11457), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11097) );
  INV_X1 U14224 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11094) );
  OR2_X1 U14225 ( .A1(n11461), .A2(n11094), .ZN(n11096) );
  NAND2_X1 U14226 ( .A1(n11449), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11095) );
  NAND4_X1 U14227 ( .A1(n11098), .A2(n11097), .A3(n11096), .A4(n11095), .ZN(
        n11102) );
  INV_X1 U14228 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11100) );
  INV_X1 U14229 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11099) );
  OAI22_X1 U14230 ( .A1(n11100), .A2(n15871), .B1(n11421), .B2(n11099), .ZN(
        n11101) );
  NOR2_X1 U14231 ( .A1(n11102), .A2(n11101), .ZN(n11114) );
  INV_X1 U14232 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11103) );
  INV_X1 U14233 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11499) );
  OAI22_X1 U14234 ( .A1(n11103), .A2(n11163), .B1(n11166), .B2(n11499), .ZN(
        n11106) );
  INV_X1 U14235 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11506) );
  OAI22_X1 U14236 ( .A1(n11159), .A2(n11506), .B1(n11161), .B2(n11104), .ZN(
        n11105) );
  NOR2_X1 U14237 ( .A1(n11106), .A2(n11105), .ZN(n11113) );
  INV_X1 U14238 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11325) );
  OAI22_X1 U14239 ( .A1(n19818), .A2(n11177), .B1(n11178), .B2(n11325), .ZN(
        n11111) );
  INV_X1 U14240 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11109) );
  INV_X1 U14241 ( .A(n11463), .ZN(n11108) );
  INV_X1 U14242 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11107) );
  OAI22_X1 U14243 ( .A1(n11109), .A2(n11108), .B1(n11168), .B2(n11107), .ZN(
        n11110) );
  NOR2_X1 U14244 ( .A1(n11111), .A2(n11110), .ZN(n11112) );
  NAND2_X1 U14245 ( .A1(n11053), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U14246 ( .A1(n12889), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11115) );
  OAI211_X1 U14247 ( .C1(n13979), .C2(n11212), .A(n11116), .B(n11115), .ZN(
        n15763) );
  AOI22_X1 U14248 ( .A1(n12889), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11132) );
  AOI22_X1 U14249 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10424), .B1(
        n11080), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11120) );
  AOI22_X1 U14250 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11448), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14251 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11449), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14252 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11451), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11117) );
  NAND4_X1 U14253 ( .A1(n11120), .A2(n11119), .A3(n11118), .A4(n11117), .ZN(
        n11130) );
  AOI22_X1 U14254 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11456), .B1(
        n11077), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11128) );
  INV_X1 U14255 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11123) );
  NAND2_X1 U14256 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11122) );
  NAND2_X1 U14257 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11121) );
  OAI211_X1 U14258 ( .C1(n11461), .C2(n11123), .A(n11122), .B(n11121), .ZN(
        n11124) );
  INV_X1 U14259 ( .A(n11124), .ZN(n11127) );
  AOI22_X1 U14260 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10369), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11126) );
  NAND2_X1 U14261 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11125) );
  NAND4_X1 U14262 ( .A1(n11128), .A2(n11127), .A3(n11126), .A4(n11125), .ZN(
        n11129) );
  NAND2_X1 U14263 ( .A1(n11009), .A2(n13967), .ZN(n11131) );
  OAI211_X1 U14264 ( .C1(n11133), .C2(n19965), .A(n11132), .B(n11131), .ZN(
        n15750) );
  AOI22_X1 U14265 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11448), .B1(
        n11080), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11137) );
  AOI22_X1 U14266 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11451), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11136) );
  AOI22_X1 U14267 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11449), .B1(
        n11463), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11135) );
  AOI22_X1 U14268 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10453), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11134) );
  NAND4_X1 U14269 ( .A1(n11137), .A2(n11136), .A3(n11135), .A4(n11134), .ZN(
        n11147) );
  AOI22_X1 U14270 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11077), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11145) );
  INV_X1 U14271 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11140) );
  NAND2_X1 U14272 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11139) );
  NAND2_X1 U14273 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11138) );
  OAI211_X1 U14274 ( .C1(n11461), .C2(n11140), .A(n11139), .B(n11138), .ZN(
        n11141) );
  INV_X1 U14275 ( .A(n11141), .ZN(n11144) );
  AOI22_X1 U14276 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10369), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11143) );
  NAND2_X1 U14277 ( .A1(n11450), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11142) );
  NAND4_X1 U14278 ( .A1(n11145), .A2(n11144), .A3(n11143), .A4(n11142), .ZN(
        n11146) );
  NOR2_X1 U14279 ( .A1(n11147), .A2(n11146), .ZN(n14045) );
  AOI22_X1 U14280 ( .A1(n12889), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11148) );
  OAI21_X1 U14281 ( .B1(n14045), .B2(n11212), .A(n11148), .ZN(n11149) );
  AOI21_X1 U14282 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n11053), .A(n11149), 
        .ZN(n15737) );
  NOR2_X2 U14283 ( .A1(n15736), .A2(n15737), .ZN(n15724) );
  AOI22_X1 U14284 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11154) );
  AOI22_X1 U14285 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11153) );
  INV_X1 U14286 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11150) );
  OR2_X1 U14287 ( .A1(n11461), .A2(n11150), .ZN(n11152) );
  NAND2_X1 U14288 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11151) );
  NAND4_X1 U14289 ( .A1(n11154), .A2(n11153), .A3(n11152), .A4(n11151), .ZN(
        n11158) );
  INV_X1 U14290 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11156) );
  INV_X1 U14291 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11155) );
  OAI22_X1 U14292 ( .A1(n11421), .A2(n11156), .B1(n15871), .B2(n11155), .ZN(
        n11157) );
  NOR2_X1 U14293 ( .A1(n11158), .A2(n11157), .ZN(n11174) );
  INV_X1 U14294 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11570) );
  OAI22_X1 U14295 ( .A1(n11159), .A2(n11570), .B1(n11177), .B2(n19829), .ZN(
        n11165) );
  OAI22_X1 U14296 ( .A1(n11163), .A2(n11162), .B1(n11161), .B2(n11160), .ZN(
        n11164) );
  NOR2_X1 U14297 ( .A1(n11165), .A2(n11164), .ZN(n11173) );
  OAI22_X1 U14298 ( .A1(n11166), .A2(n11563), .B1(n11178), .B2(n11400), .ZN(
        n11171) );
  OAI22_X1 U14299 ( .A1(n11169), .A2(n13901), .B1(n11168), .B2(n11167), .ZN(
        n11170) );
  NOR2_X1 U14300 ( .A1(n11171), .A2(n11170), .ZN(n11172) );
  NAND2_X1 U14301 ( .A1(n11053), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U14302 ( .A1(n12889), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11175) );
  OAI211_X1 U14303 ( .C1(n14249), .C2(n11212), .A(n11176), .B(n11175), .ZN(
        n15725) );
  NAND2_X1 U14304 ( .A1(n11053), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14305 ( .A1(n12889), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14306 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11448), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11182) );
  AOI22_X1 U14307 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11449), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14308 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n11080), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11180) );
  AOI22_X1 U14309 ( .A1(n11451), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11179) );
  NAND4_X1 U14310 ( .A1(n11182), .A2(n11181), .A3(n11180), .A4(n11179), .ZN(
        n11192) );
  AOI22_X1 U14311 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11456), .B1(
        n11077), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11190) );
  INV_X1 U14312 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U14313 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11184) );
  NAND2_X1 U14314 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11183) );
  OAI211_X1 U14315 ( .C1(n11461), .C2(n11185), .A(n11184), .B(n11183), .ZN(
        n11186) );
  INV_X1 U14316 ( .A(n11186), .ZN(n11189) );
  AOI22_X1 U14317 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10369), .B1(
        n11457), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11188) );
  NAND2_X1 U14318 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11187) );
  NAND4_X1 U14319 ( .A1(n11190), .A2(n11189), .A3(n11188), .A4(n11187), .ZN(
        n11191) );
  OR2_X1 U14320 ( .A1(n11192), .A2(n11191), .ZN(n14238) );
  NAND2_X1 U14321 ( .A1(n11009), .A2(n14238), .ZN(n11193) );
  AOI22_X1 U14322 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10424), .B1(
        n11080), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11199) );
  AOI22_X1 U14323 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11448), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14324 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11449), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14325 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11451), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11196) );
  NAND4_X1 U14326 ( .A1(n11199), .A2(n11198), .A3(n11197), .A4(n11196), .ZN(
        n11209) );
  AOI22_X1 U14327 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11456), .B1(
        n11077), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11207) );
  INV_X1 U14328 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11202) );
  NAND2_X1 U14329 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11201) );
  NAND2_X1 U14330 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11200) );
  OAI211_X1 U14331 ( .C1(n11461), .C2(n11202), .A(n11201), .B(n11200), .ZN(
        n11203) );
  INV_X1 U14332 ( .A(n11203), .ZN(n11206) );
  AOI22_X1 U14333 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10369), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11205) );
  NAND2_X1 U14334 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11204) );
  NAND4_X1 U14335 ( .A1(n11207), .A2(n11206), .A3(n11205), .A4(n11204), .ZN(
        n11208) );
  OR2_X1 U14336 ( .A1(n11209), .A2(n11208), .ZN(n14203) );
  INV_X1 U14337 ( .A(n14203), .ZN(n11213) );
  NAND2_X1 U14338 ( .A1(n11053), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14339 ( .A1(n12889), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11210) );
  OAI211_X1 U14340 ( .C1(n11213), .C2(n11212), .A(n11211), .B(n11210), .ZN(
        n15693) );
  NAND2_X1 U14341 ( .A1(n11053), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14342 ( .A1(n12889), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11214) );
  NAND2_X1 U14343 ( .A1(n11215), .A2(n11214), .ZN(n15679) );
  NAND2_X1 U14344 ( .A1(n11053), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14345 ( .A1(n12889), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11216) );
  NAND2_X1 U14346 ( .A1(n11053), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14347 ( .A1(n12889), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11218) );
  NAND2_X1 U14348 ( .A1(n11219), .A2(n11218), .ZN(n15650) );
  NAND2_X1 U14349 ( .A1(n11053), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14350 ( .A1(n12889), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11220) );
  AND2_X1 U14351 ( .A1(n11221), .A2(n11220), .ZN(n14332) );
  NAND2_X1 U14352 ( .A1(n11053), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14353 ( .A1(n12889), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11222) );
  NAND2_X1 U14354 ( .A1(n11053), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14355 ( .A1(n12889), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11224) );
  AND2_X1 U14356 ( .A1(n11225), .A2(n11224), .ZN(n14485) );
  NAND2_X1 U14357 ( .A1(n11053), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14358 ( .A1(n12889), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11226) );
  NAND2_X1 U14359 ( .A1(n11227), .A2(n11226), .ZN(n11228) );
  OR2_X1 U14360 ( .A1(n14486), .A2(n11228), .ZN(n11229) );
  NAND2_X1 U14361 ( .A1(n15127), .A2(n11229), .ZN(n15143) );
  NOR2_X1 U14362 ( .A1(n15151), .A2(n11231), .ZN(n11232) );
  OR2_X1 U14363 ( .A1(n11230), .A2(n11232), .ZN(n15225) );
  INV_X1 U14364 ( .A(n15225), .ZN(n11235) );
  NAND2_X1 U14365 ( .A1(n11233), .A2(n11007), .ZN(n11234) );
  NAND2_X1 U14366 ( .A1(n11235), .A2(n16479), .ZN(n11236) );
  NAND2_X1 U14367 ( .A1(n19399), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12350) );
  OAI211_X1 U14368 ( .C1(n16474), .C2(n15143), .A(n11236), .B(n12350), .ZN(
        n11244) );
  INV_X1 U14369 ( .A(n15831), .ZN(n13640) );
  OAI22_X1 U14370 ( .A1(n15663), .A2(n11237), .B1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13640), .ZN(n14163) );
  NAND2_X1 U14371 ( .A1(n15794), .A2(n11240), .ZN(n15691) );
  NOR2_X1 U14372 ( .A1(n15639), .A2(n11242), .ZN(n12899) );
  INV_X1 U14373 ( .A(n12899), .ZN(n15607) );
  NOR2_X1 U14374 ( .A1(n15607), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11243) );
  AOI211_X1 U14375 ( .C1(n15621), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11244), .B(n11243), .ZN(n11251) );
  INV_X1 U14376 ( .A(n11245), .ZN(n15354) );
  NOR2_X1 U14377 ( .A1(n11246), .A2(n15354), .ZN(n11248) );
  XOR2_X1 U14378 ( .A(n11248), .B(n11247), .Z(n12353) );
  INV_X1 U14379 ( .A(n11249), .ZN(n11250) );
  AND2_X1 U14380 ( .A1(n16497), .A2(n11284), .ZN(n20044) );
  OAI211_X2 U14381 ( .C1(n11258), .C2(n11257), .A(n11256), .B(n15293), .ZN(
        n11265) );
  NOR2_X1 U14382 ( .A1(n11259), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11260) );
  MUX2_X1 U14383 ( .A(n11261), .B(n11260), .S(n10611), .Z(n14532) );
  NAND2_X1 U14384 ( .A1(n14532), .A2(n11262), .ZN(n11263) );
  XOR2_X1 U14385 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11263), .Z(
        n11264) );
  INV_X1 U14386 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n11266) );
  NOR2_X1 U14387 ( .A1(n19214), .A2(n11266), .ZN(n12894) );
  INV_X1 U14388 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11267) );
  NOR2_X1 U14389 ( .A1(n16455), .A2(n12916), .ZN(n11268) );
  AOI211_X1 U14390 ( .C1(n16442), .C2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12894), .B(n11268), .ZN(n11269) );
  AOI22_X1 U14391 ( .A1(n11270), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11273) );
  NAND2_X1 U14392 ( .A1(n11271), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11272) );
  OAI211_X1 U14393 ( .C1(n9771), .C2(n11254), .A(n11273), .B(n11272), .ZN(
        n11274) );
  NAND2_X1 U14394 ( .A1(n10242), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11278) );
  NAND2_X1 U14395 ( .A1(n11278), .A2(n20033), .ZN(n11304) );
  NOR2_X1 U14396 ( .A1(n20024), .A2(n20032), .ZN(n19579) );
  AND2_X1 U14397 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19579), .ZN(
        n11301) );
  INV_X1 U14398 ( .A(n11301), .ZN(n11280) );
  NAND2_X1 U14399 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19611) );
  NAND2_X1 U14400 ( .A1(n19611), .A2(n20024), .ZN(n11279) );
  NAND2_X1 U14401 ( .A1(n11280), .A2(n11279), .ZN(n15886) );
  NOR2_X1 U14402 ( .A1(n20013), .A2(n15886), .ZN(n11281) );
  AOI21_X1 U14403 ( .B1(n11304), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11281), .ZN(n11282) );
  NAND2_X1 U14404 ( .A1(n11536), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11295) );
  NAND2_X1 U14405 ( .A1(n11304), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11286) );
  NAND2_X1 U14406 ( .A1(n20032), .A2(n20040), .ZN(n19410) );
  AND2_X1 U14407 ( .A1(n19611), .A2(n19410), .ZN(n19694) );
  NAND2_X1 U14408 ( .A1(n19694), .A2(n20004), .ZN(n19587) );
  NAND2_X1 U14409 ( .A1(n11286), .A2(n19587), .ZN(n11287) );
  AOI22_X1 U14410 ( .A1(n11304), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20004), .B2(n20040), .ZN(n11290) );
  NAND2_X1 U14411 ( .A1(n11536), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11292) );
  NAND2_X1 U14412 ( .A1(n13599), .A2(n13600), .ZN(n13598) );
  INV_X1 U14413 ( .A(n11292), .ZN(n11293) );
  OR2_X1 U14414 ( .A1(n15849), .A2(n11293), .ZN(n11294) );
  INV_X1 U14415 ( .A(n11295), .ZN(n11296) );
  NAND2_X1 U14416 ( .A1(n11297), .A2(n11296), .ZN(n11298) );
  NAND2_X1 U14417 ( .A1(n11300), .A2(n11299), .ZN(n11306) );
  OAI21_X1 U14418 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11301), .A(
        n20004), .ZN(n11302) );
  AND2_X1 U14419 ( .A1(n11301), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19853) );
  NOR2_X1 U14420 ( .A1(n11302), .A2(n19853), .ZN(n11303) );
  AOI21_X1 U14421 ( .B1(n11304), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11303), .ZN(n11305) );
  NAND2_X1 U14422 ( .A1(n11306), .A2(n11305), .ZN(n11312) );
  INV_X1 U14423 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11307) );
  NOR2_X1 U14424 ( .A1(n13783), .A2(n11307), .ZN(n11308) );
  OR2_X1 U14425 ( .A1(n11312), .A2(n11308), .ZN(n11309) );
  NAND2_X1 U14426 ( .A1(n11312), .A2(n11308), .ZN(n13785) );
  NAND2_X1 U14427 ( .A1(n13737), .A2(n13738), .ZN(n11311) );
  NAND2_X1 U14428 ( .A1(n10242), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11310) );
  AND2_X1 U14429 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11313) );
  AND2_X1 U14430 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13903) );
  NAND4_X1 U14431 ( .A1(n11314), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .A4(n13903), .ZN(n11315) );
  NOR2_X1 U14432 ( .A1(n13783), .A2(n11315), .ZN(n11316) );
  INV_X1 U14433 ( .A(n13854), .ZN(n11318) );
  AOI22_X1 U14434 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11080), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11322) );
  AOI22_X1 U14435 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n11448), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14436 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11449), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14437 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11451), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11319) );
  NAND4_X1 U14438 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(
        n11332) );
  AOI22_X1 U14439 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n11077), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U14440 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11324) );
  NAND2_X1 U14441 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11323) );
  OAI211_X1 U14442 ( .C1(n11461), .C2(n11325), .A(n11324), .B(n11323), .ZN(
        n11326) );
  INV_X1 U14443 ( .A(n11326), .ZN(n11329) );
  AOI22_X1 U14444 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11402), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11328) );
  NAND2_X1 U14445 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11327) );
  NAND4_X1 U14446 ( .A1(n11330), .A2(n11329), .A3(n11328), .A4(n11327), .ZN(
        n11331) );
  OR2_X1 U14447 ( .A1(n11332), .A2(n11331), .ZN(n14388) );
  AOI22_X1 U14448 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11080), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14449 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11448), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14450 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11449), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14451 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11451), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11333) );
  NAND4_X1 U14452 ( .A1(n11336), .A2(n11335), .A3(n11334), .A4(n11333), .ZN(
        n11346) );
  AOI22_X1 U14453 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11077), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11344) );
  NAND2_X1 U14454 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11338) );
  NAND2_X1 U14455 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11337) );
  OAI211_X1 U14456 ( .C1(n11461), .C2(n11339), .A(n11338), .B(n11337), .ZN(
        n11340) );
  INV_X1 U14457 ( .A(n11340), .ZN(n11343) );
  AOI22_X1 U14458 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11402), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U14459 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11341) );
  NAND4_X1 U14460 ( .A1(n11344), .A2(n11343), .A3(n11342), .A4(n11341), .ZN(
        n11345) );
  OR2_X1 U14461 ( .A1(n11346), .A2(n11345), .ZN(n14221) );
  AOI22_X1 U14462 ( .A1(n11080), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14463 ( .A1(n11448), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14464 ( .A1(n11449), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14465 ( .A1(n11451), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11347) );
  NAND4_X1 U14466 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n11360) );
  AOI22_X1 U14467 ( .A1(n11077), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11358) );
  INV_X1 U14468 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11353) );
  NAND2_X1 U14469 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11352) );
  NAND2_X1 U14470 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11351) );
  OAI211_X1 U14471 ( .C1(n11461), .C2(n11353), .A(n11352), .B(n11351), .ZN(
        n11354) );
  INV_X1 U14472 ( .A(n11354), .ZN(n11357) );
  AOI22_X1 U14473 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11356) );
  NAND2_X1 U14474 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11355) );
  NAND4_X1 U14475 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(
        n11359) );
  NOR2_X1 U14476 ( .A1(n11360), .A2(n11359), .ZN(n14256) );
  INV_X1 U14477 ( .A(n14256), .ZN(n11361) );
  AND2_X1 U14478 ( .A1(n14203), .A2(n14238), .ZN(n14202) );
  AND2_X1 U14479 ( .A1(n11361), .A2(n14202), .ZN(n14218) );
  NAND2_X1 U14480 ( .A1(n14221), .A2(n14218), .ZN(n11362) );
  OR2_X1 U14481 ( .A1(n11362), .A2(n14249), .ZN(n11363) );
  NOR2_X1 U14482 ( .A1(n11363), .A2(n14045), .ZN(n14219) );
  AOI22_X1 U14483 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11080), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14484 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11448), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14485 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11449), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14486 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11451), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11366) );
  NAND4_X1 U14487 ( .A1(n11369), .A2(n11368), .A3(n11367), .A4(n11366), .ZN(
        n11379) );
  AOI22_X1 U14488 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n11077), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11377) );
  NAND2_X1 U14489 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11371) );
  NAND2_X1 U14490 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11370) );
  OAI211_X1 U14491 ( .C1(n11461), .C2(n11372), .A(n11371), .B(n11370), .ZN(
        n11373) );
  INV_X1 U14492 ( .A(n11373), .ZN(n11376) );
  AOI22_X1 U14493 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11402), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11375) );
  NAND2_X1 U14494 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11374) );
  NAND4_X1 U14495 ( .A1(n11377), .A2(n11376), .A3(n11375), .A4(n11374), .ZN(
        n11378) );
  AOI22_X1 U14496 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11080), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14497 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11448), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14498 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11449), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14499 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11451), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11380) );
  NAND4_X1 U14500 ( .A1(n11383), .A2(n11382), .A3(n11381), .A4(n11380), .ZN(
        n11393) );
  AOI22_X1 U14501 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11077), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11391) );
  INV_X1 U14502 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11386) );
  NAND2_X1 U14503 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11385) );
  NAND2_X1 U14504 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11384) );
  OAI211_X1 U14505 ( .C1(n11461), .C2(n11386), .A(n11385), .B(n11384), .ZN(
        n11387) );
  INV_X1 U14506 ( .A(n11387), .ZN(n11390) );
  AOI22_X1 U14507 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11402), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11389) );
  NAND2_X1 U14508 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11388) );
  NAND4_X1 U14509 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n11392) );
  NOR2_X1 U14510 ( .A1(n11393), .A2(n11392), .ZN(n15234) );
  AOI22_X1 U14511 ( .A1(n11080), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14512 ( .A1(n11448), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14513 ( .A1(n11449), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14514 ( .A1(n11451), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11394) );
  NAND4_X1 U14515 ( .A1(n11397), .A2(n11396), .A3(n11395), .A4(n11394), .ZN(
        n11408) );
  AOI22_X1 U14516 ( .A1(n11077), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11456), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11406) );
  NAND2_X1 U14517 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11399) );
  NAND2_X1 U14518 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11398) );
  OAI211_X1 U14519 ( .C1(n11461), .C2(n11400), .A(n11399), .B(n11398), .ZN(
        n11401) );
  INV_X1 U14520 ( .A(n11401), .ZN(n11405) );
  AOI22_X1 U14521 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11404) );
  NAND2_X1 U14522 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11403) );
  NAND4_X1 U14523 ( .A1(n11406), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(
        n11407) );
  OR2_X1 U14524 ( .A1(n11408), .A2(n11407), .ZN(n14484) );
  OAI22_X1 U14525 ( .A1(n11411), .A2(n10087), .B1(n11410), .B2(n11409), .ZN(
        n11412) );
  AOI21_X1 U14526 ( .B1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n11463), .A(
        n11412), .ZN(n11414) );
  AOI22_X1 U14527 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11457), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11413) );
  OAI211_X1 U14528 ( .C1(n11415), .C2(n11461), .A(n11414), .B(n11413), .ZN(
        n11425) );
  AOI22_X1 U14529 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11080), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14530 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11448), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14531 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11449), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14532 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11451), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11416) );
  NAND4_X1 U14533 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n11424) );
  OAI22_X1 U14534 ( .A1(n11422), .A2(n11421), .B1(n15871), .B2(n11420), .ZN(
        n11423) );
  NOR3_X1 U14535 ( .A1(n11425), .A2(n11424), .A3(n11423), .ZN(n14501) );
  INV_X1 U14536 ( .A(n11426), .ZN(n11615) );
  INV_X1 U14537 ( .A(n11615), .ZN(n11603) );
  AOI22_X1 U14538 ( .A1(n10361), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14539 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14540 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10222), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11436) );
  INV_X1 U14541 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11433) );
  NAND2_X1 U14542 ( .A1(n9766), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11432) );
  INV_X1 U14543 ( .A(n11428), .ZN(n11431) );
  INV_X1 U14544 ( .A(n11429), .ZN(n11430) );
  NAND2_X1 U14545 ( .A1(n11431), .A2(n11430), .ZN(n11612) );
  OAI211_X1 U14546 ( .C1(n9725), .C2(n11433), .A(n11432), .B(n11612), .ZN(
        n11434) );
  INV_X1 U14547 ( .A(n11434), .ZN(n11435) );
  NAND4_X1 U14548 ( .A1(n11438), .A2(n11437), .A3(n11436), .A4(n11435), .ZN(
        n11447) );
  AOI22_X1 U14549 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14550 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14551 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11443) );
  INV_X1 U14552 ( .A(n10222), .ZN(n11611) );
  INV_X1 U14553 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11440) );
  NAND2_X1 U14554 ( .A1(n11586), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11439) );
  INV_X1 U14555 ( .A(n11612), .ZN(n11587) );
  OAI211_X1 U14556 ( .C1(n11611), .C2(n11440), .A(n11439), .B(n11587), .ZN(
        n11441) );
  INV_X1 U14557 ( .A(n11441), .ZN(n11442) );
  NAND4_X1 U14558 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11446) );
  AND2_X1 U14559 ( .A1(n11447), .A2(n11446), .ZN(n11492) );
  NAND2_X1 U14560 ( .A1(n11284), .A2(n11492), .ZN(n11470) );
  AOI22_X1 U14561 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11448), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U14562 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11449), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14563 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11080), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14564 ( .A1(n11451), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11450), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11452) );
  NAND4_X1 U14565 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n11469) );
  AOI22_X1 U14566 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n11456), .B1(
        n11077), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11467) );
  INV_X1 U14567 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11460) );
  NAND2_X1 U14568 ( .A1(n11457), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11459) );
  NAND2_X1 U14569 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11458) );
  OAI211_X1 U14570 ( .C1(n11461), .C2(n11460), .A(n11459), .B(n11458), .ZN(
        n11462) );
  INV_X1 U14571 ( .A(n11462), .ZN(n11466) );
  AOI22_X1 U14572 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11402), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11465) );
  NAND2_X1 U14573 ( .A1(n11463), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11464) );
  NAND4_X1 U14574 ( .A1(n11467), .A2(n11466), .A3(n11465), .A4(n11464), .ZN(
        n11468) );
  XNOR2_X1 U14575 ( .A(n11470), .B(n11489), .ZN(n11495) );
  NAND2_X1 U14576 ( .A1(n11007), .A2(n11492), .ZN(n15220) );
  AOI22_X1 U14577 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14578 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14579 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11477) );
  NAND2_X1 U14580 ( .A1(n11586), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11473) );
  OAI211_X1 U14581 ( .C1(n11611), .C2(n11474), .A(n11473), .B(n11612), .ZN(
        n11475) );
  INV_X1 U14582 ( .A(n11475), .ZN(n11476) );
  NAND4_X1 U14583 ( .A1(n11479), .A2(n11478), .A3(n11477), .A4(n11476), .ZN(
        n11488) );
  AOI22_X1 U14584 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14585 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14586 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11484) );
  NAND2_X1 U14587 ( .A1(n9766), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11480) );
  OAI211_X1 U14588 ( .C1(n11611), .C2(n11481), .A(n11480), .B(n11587), .ZN(
        n11482) );
  INV_X1 U14589 ( .A(n11482), .ZN(n11483) );
  NAND4_X1 U14590 ( .A1(n11486), .A2(n11485), .A3(n11484), .A4(n11483), .ZN(
        n11487) );
  NAND2_X1 U14591 ( .A1(n11488), .A2(n11487), .ZN(n11496) );
  NAND2_X1 U14592 ( .A1(n11489), .A2(n11492), .ZN(n11497) );
  XOR2_X1 U14593 ( .A(n11496), .B(n11497), .Z(n11490) );
  NAND2_X1 U14594 ( .A1(n11490), .A2(n11536), .ZN(n15209) );
  INV_X1 U14595 ( .A(n11496), .ZN(n11491) );
  NAND2_X1 U14596 ( .A1(n11007), .A2(n11491), .ZN(n15212) );
  INV_X1 U14597 ( .A(n11492), .ZN(n11493) );
  NOR2_X1 U14598 ( .A1(n15212), .A2(n11493), .ZN(n11494) );
  NOR2_X1 U14599 ( .A1(n11497), .A2(n11496), .ZN(n11514) );
  AOI22_X1 U14600 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14601 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14602 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11502) );
  NAND2_X1 U14603 ( .A1(n9766), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11498) );
  OAI211_X1 U14604 ( .C1(n11611), .C2(n11499), .A(n11498), .B(n11612), .ZN(
        n11500) );
  INV_X1 U14605 ( .A(n11500), .ZN(n11501) );
  NAND4_X1 U14606 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11513) );
  AOI22_X1 U14607 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14608 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14609 ( .A1(n10361), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11509) );
  NAND2_X1 U14610 ( .A1(n11586), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11505) );
  OAI211_X1 U14611 ( .C1(n11611), .C2(n11506), .A(n11505), .B(n11587), .ZN(
        n11507) );
  INV_X1 U14612 ( .A(n11507), .ZN(n11508) );
  NAND4_X1 U14613 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(
        n11512) );
  AND2_X1 U14614 ( .A1(n11513), .A2(n11512), .ZN(n11515) );
  NAND2_X1 U14615 ( .A1(n11514), .A2(n11515), .ZN(n11558) );
  OAI211_X1 U14616 ( .C1(n11514), .C2(n11515), .A(n11536), .B(n11558), .ZN(
        n11517) );
  INV_X1 U14617 ( .A(n11515), .ZN(n11516) );
  NOR2_X1 U14618 ( .A1(n11284), .A2(n11516), .ZN(n15205) );
  AOI22_X1 U14619 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14620 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14621 ( .A1(n10361), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U14622 ( .A1(n11586), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11520) );
  OAI211_X1 U14623 ( .C1(n11611), .C2(n11521), .A(n11520), .B(n11612), .ZN(
        n11522) );
  INV_X1 U14624 ( .A(n11522), .ZN(n11523) );
  NAND4_X1 U14625 ( .A1(n11526), .A2(n11525), .A3(n11524), .A4(n11523), .ZN(
        n11535) );
  AOI22_X1 U14626 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14627 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14628 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11531) );
  INV_X1 U14629 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11528) );
  NAND2_X1 U14630 ( .A1(n11586), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11527) );
  OAI211_X1 U14631 ( .C1(n11611), .C2(n11528), .A(n11527), .B(n11587), .ZN(
        n11529) );
  INV_X1 U14632 ( .A(n11529), .ZN(n11530) );
  NAND4_X1 U14633 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11534) );
  AND2_X1 U14634 ( .A1(n11535), .A2(n11534), .ZN(n11538) );
  XNOR2_X1 U14635 ( .A(n11558), .B(n11538), .ZN(n11537) );
  NAND2_X1 U14636 ( .A1(n11537), .A2(n11536), .ZN(n11540) );
  INV_X1 U14637 ( .A(n11538), .ZN(n11557) );
  NOR2_X1 U14638 ( .A1(n11284), .A2(n11557), .ZN(n15197) );
  AOI22_X1 U14639 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14640 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14641 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11545) );
  INV_X1 U14642 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11542) );
  NAND2_X1 U14643 ( .A1(n9726), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11541) );
  OAI211_X1 U14644 ( .C1(n11611), .C2(n11542), .A(n11541), .B(n11612), .ZN(
        n11543) );
  INV_X1 U14645 ( .A(n11543), .ZN(n11544) );
  NAND4_X1 U14646 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11556) );
  AOI22_X1 U14647 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11554) );
  INV_X1 U14648 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n21251) );
  AOI22_X1 U14649 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11553) );
  INV_X1 U14650 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n19677) );
  AOI22_X1 U14651 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11552) );
  INV_X1 U14652 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U14653 ( .A1(n9726), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11548) );
  OAI211_X1 U14654 ( .C1(n11611), .C2(n11549), .A(n11548), .B(n11587), .ZN(
        n11550) );
  INV_X1 U14655 ( .A(n11550), .ZN(n11551) );
  NAND4_X1 U14656 ( .A1(n11554), .A2(n11553), .A3(n11552), .A4(n11551), .ZN(
        n11555) );
  NAND2_X1 U14657 ( .A1(n11556), .A2(n11555), .ZN(n11561) );
  OR2_X1 U14658 ( .A1(n11558), .A2(n11557), .ZN(n11559) );
  NOR2_X1 U14659 ( .A1(n11559), .A2(n11561), .ZN(n15184) );
  NOR2_X1 U14660 ( .A1(n11284), .A2(n11561), .ZN(n15192) );
  NAND2_X1 U14661 ( .A1(n15193), .A2(n15192), .ZN(n15191) );
  AOI22_X1 U14662 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14663 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14664 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11566) );
  NAND2_X1 U14665 ( .A1(n11586), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11562) );
  OAI211_X1 U14666 ( .C1(n11611), .C2(n11563), .A(n11562), .B(n11612), .ZN(
        n11564) );
  INV_X1 U14667 ( .A(n11564), .ZN(n11565) );
  NAND4_X1 U14668 ( .A1(n11568), .A2(n11567), .A3(n11566), .A4(n11565), .ZN(
        n11577) );
  AOI22_X1 U14669 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14670 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14671 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11573) );
  NAND2_X1 U14672 ( .A1(n9766), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11569) );
  OAI211_X1 U14673 ( .C1(n11611), .C2(n11570), .A(n11569), .B(n11587), .ZN(
        n11571) );
  INV_X1 U14674 ( .A(n11571), .ZN(n11572) );
  NAND4_X1 U14675 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11576) );
  NAND2_X1 U14676 ( .A1(n11577), .A2(n11576), .ZN(n11597) );
  AOI21_X1 U14677 ( .B1(n15191), .B2(n15186), .A(n11597), .ZN(n15180) );
  AOI22_X1 U14678 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14679 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14680 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11582) );
  NAND2_X1 U14681 ( .A1(n9726), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11578) );
  OAI211_X1 U14682 ( .C1(n11611), .C2(n11579), .A(n11578), .B(n11612), .ZN(
        n11580) );
  INV_X1 U14683 ( .A(n11580), .ZN(n11581) );
  NAND4_X1 U14684 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11596) );
  AOI22_X1 U14685 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14686 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14687 ( .A1(n10361), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11592) );
  INV_X1 U14688 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11589) );
  NAND2_X1 U14689 ( .A1(n9726), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11588) );
  OAI211_X1 U14690 ( .C1(n11611), .C2(n11589), .A(n11588), .B(n11587), .ZN(
        n11590) );
  INV_X1 U14691 ( .A(n11590), .ZN(n11591) );
  NAND4_X1 U14692 ( .A1(n11594), .A2(n11593), .A3(n11592), .A4(n11591), .ZN(
        n11595) );
  NAND2_X1 U14693 ( .A1(n11596), .A2(n11595), .ZN(n11600) );
  INV_X1 U14694 ( .A(n11597), .ZN(n15187) );
  AND2_X1 U14695 ( .A1(n11284), .A2(n15187), .ZN(n11598) );
  NAND2_X1 U14696 ( .A1(n15184), .A2(n11598), .ZN(n11599) );
  NOR2_X1 U14697 ( .A1(n11599), .A2(n11600), .ZN(n11601) );
  AOI21_X1 U14698 ( .B1(n11600), .B2(n11599), .A(n11601), .ZN(n15179) );
  NAND2_X1 U14699 ( .A1(n15180), .A2(n15179), .ZN(n15181) );
  INV_X1 U14700 ( .A(n11601), .ZN(n11602) );
  NAND2_X1 U14701 ( .A1(n15181), .A2(n11602), .ZN(n11628) );
  AOI22_X1 U14702 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11603), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14703 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11606) );
  NAND2_X1 U14704 ( .A1(n11607), .A2(n11606), .ZN(n11625) );
  INV_X1 U14705 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14706 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10193), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11609) );
  AOI21_X1 U14707 ( .B1(n9766), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n11612), .ZN(n11608) );
  OAI211_X1 U14708 ( .C1(n11611), .C2(n11610), .A(n11609), .B(n11608), .ZN(
        n11624) );
  INV_X1 U14709 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11613) );
  OAI21_X1 U14710 ( .B1(n10178), .B2(n11613), .A(n11612), .ZN(n11617) );
  INV_X1 U14711 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15907) );
  INV_X1 U14712 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11614) );
  OAI22_X1 U14713 ( .A1(n11615), .A2(n15907), .B1(n9725), .B2(n11614), .ZN(
        n11616) );
  AOI211_X1 U14714 ( .C1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .C2(n10222), .A(
        n11617), .B(n11616), .ZN(n11622) );
  AOI22_X1 U14715 ( .A1(n11605), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14716 ( .A1(n11585), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11620) );
  NAND3_X1 U14717 ( .A1(n11622), .A2(n11621), .A3(n11620), .ZN(n11623) );
  OAI21_X1 U14718 ( .B1(n11625), .B2(n11624), .A(n11623), .ZN(n11626) );
  XNOR2_X1 U14719 ( .A(n11628), .B(n11627), .ZN(n11681) );
  NAND2_X1 U14720 ( .A1(n16501), .A2(n16503), .ZN(n13545) );
  INV_X1 U14721 ( .A(n11629), .ZN(n14314) );
  NAND2_X1 U14722 ( .A1(n13545), .A2(n14314), .ZN(n11630) );
  NAND2_X1 U14723 ( .A1(n15515), .A2(n15229), .ZN(n11632) );
  NAND2_X1 U14724 ( .A1(n13900), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11631) );
  OAI21_X1 U14725 ( .B1(n11681), .B2(n15242), .A(n11633), .ZN(P2_U2857) );
  AND2_X1 U14726 ( .A1(n9750), .A2(n19922), .ZN(n13459) );
  NAND3_X1 U14727 ( .A1(n10997), .A2(n11635), .A3(n13459), .ZN(n11636) );
  OAI21_X1 U14728 ( .B1(n16501), .B2(n16505), .A(n11636), .ZN(n13547) );
  NAND2_X1 U14729 ( .A1(n11053), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14730 ( .A1(n12889), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11640) );
  AND2_X1 U14731 ( .A1(n11641), .A2(n11640), .ZN(n15126) );
  NAND2_X1 U14732 ( .A1(n11053), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14733 ( .A1(n12889), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11642) );
  AND2_X1 U14734 ( .A1(n11643), .A2(n11642), .ZN(n15273) );
  INV_X1 U14735 ( .A(n15273), .ZN(n11644) );
  NAND2_X1 U14736 ( .A1(n11053), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14737 ( .A1(n12889), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11645) );
  AND2_X1 U14738 ( .A1(n11646), .A2(n11645), .ZN(n15113) );
  NAND2_X1 U14739 ( .A1(n11053), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14740 ( .A1(n12889), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U14741 ( .A1(n11648), .A2(n11647), .ZN(n15261) );
  NAND2_X1 U14742 ( .A1(n15112), .A2(n15261), .ZN(n13448) );
  NAND2_X1 U14743 ( .A1(n11053), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14744 ( .A1(n12889), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11649) );
  AND2_X1 U14745 ( .A1(n11650), .A2(n11649), .ZN(n13449) );
  INV_X1 U14746 ( .A(n11651), .ZN(n15098) );
  NAND2_X1 U14747 ( .A1(n11053), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14748 ( .A1(n12889), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11652) );
  AND2_X1 U14749 ( .A1(n11653), .A2(n11652), .ZN(n15097) );
  NAND2_X1 U14750 ( .A1(n11053), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14751 ( .A1(n12889), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U14752 ( .A1(n11655), .A2(n11654), .ZN(n15081) );
  NAND2_X1 U14753 ( .A1(n11053), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14754 ( .A1(n12889), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11656) );
  AND2_X1 U14755 ( .A1(n11657), .A2(n11656), .ZN(n11658) );
  NAND2_X1 U14756 ( .A1(n9795), .A2(n11658), .ZN(n11659) );
  NOR2_X1 U14757 ( .A1(n11676), .A2(n10257), .ZN(n11660) );
  NOR4_X1 U14758 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n11664) );
  NOR4_X1 U14759 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n11663) );
  NOR4_X1 U14760 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n11662) );
  NOR4_X1 U14761 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_8__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_9__SCAN_IN), .ZN(n11661) );
  NAND4_X1 U14762 ( .A1(n11664), .A2(n11663), .A3(n11662), .A4(n11661), .ZN(
        n11669) );
  NOR4_X1 U14763 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_2__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n11667) );
  NOR4_X1 U14764 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n11666) );
  NOR4_X1 U14765 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n11665) );
  INV_X1 U14766 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19952) );
  NAND4_X1 U14767 ( .A1(n11667), .A2(n11666), .A3(n11665), .A4(n19952), .ZN(
        n11668) );
  OAI21_X1 U14768 ( .B1(n11669), .B2(n11668), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n11670) );
  NAND2_X1 U14769 ( .A1(n15276), .A2(BUF2_REG_14__SCAN_IN), .ZN(n11672) );
  INV_X1 U14770 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14371) );
  OR2_X1 U14771 ( .A1(n15276), .A2(n14371), .ZN(n11671) );
  NAND2_X1 U14772 ( .A1(n11672), .A2(n11671), .ZN(n19388) );
  INV_X1 U14773 ( .A(n19388), .ZN(n11674) );
  INV_X1 U14774 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n11673) );
  OAI22_X1 U14775 ( .A1(n15284), .A2(n11674), .B1(n19322), .B2(n11673), .ZN(
        n11675) );
  AOI21_X1 U14776 ( .B1(n15516), .B2(n19339), .A(n11675), .ZN(n11679) );
  NOR2_X1 U14777 ( .A1(n11676), .A2(n10187), .ZN(n11677) );
  AOI22_X1 U14778 ( .A1(n19291), .A2(BUF1_REG_30__SCAN_IN), .B1(n19290), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n11678) );
  OAI21_X1 U14779 ( .B1(n11681), .B2(n19324), .A(n11680), .ZN(P2_U2889) );
  AND2_X4 U14780 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15044) );
  NAND2_X1 U14781 ( .A1(n11854), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11689) );
  INV_X1 U14782 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11683) );
  AND2_X2 U14783 ( .A1(n11700), .A2(n11701), .ZN(n12589) );
  NAND2_X1 U14784 ( .A1(n12839), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11688) );
  AND2_X2 U14785 ( .A1(n11684), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13755) );
  INV_X1 U14786 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11685) );
  AND2_X2 U14787 ( .A1(n11685), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11699) );
  NAND2_X1 U14788 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11687) );
  AND2_X2 U14789 ( .A1(n13755), .A2(n15044), .ZN(n11754) );
  NAND2_X1 U14791 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11686) );
  AND2_X4 U14792 ( .A1(n13753), .A2(n11699), .ZN(n12992) );
  NAND2_X1 U14793 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11693) );
  NOR2_X4 U14794 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15045) );
  NAND2_X1 U14795 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11692) );
  NAND2_X1 U14796 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11691) );
  NAND2_X1 U14797 ( .A1(n11747), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11690) );
  NAND2_X1 U14798 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11698) );
  NAND2_X1 U14799 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11697) );
  AND2_X2 U14800 ( .A1(n11694), .A2(n15045), .ZN(n11740) );
  NAND2_X1 U14801 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11696) );
  NAND2_X1 U14802 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11695) );
  AND2_X2 U14803 ( .A1(n11699), .A2(n11701), .ZN(n11746) );
  NAND2_X1 U14804 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11705) );
  AND2_X2 U14805 ( .A1(n11700), .A2(n13755), .ZN(n11867) );
  BUF_X2 U14806 ( .A(n11867), .Z(n12819) );
  BUF_X2 U14807 ( .A(n11859), .Z(n12862) );
  NAND2_X1 U14808 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11703) );
  NAND2_X1 U14809 ( .A1(n11741), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11702) );
  AOI22_X1 U14810 ( .A1(n11854), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14811 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14812 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14813 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11710) );
  NAND4_X1 U14814 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n11719) );
  AOI22_X1 U14815 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11717) );
  BUF_X2 U14816 ( .A(n11867), .Z(n12995) );
  AOI22_X1 U14817 ( .A1(n12995), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11724), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14818 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11747), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14819 ( .A1(n12987), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11714) );
  NAND4_X1 U14820 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11718) );
  NAND2_X1 U14821 ( .A1(n12206), .A2(n20286), .ZN(n11826) );
  AOI22_X1 U14822 ( .A1(n11854), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11723) );
  AOI22_X1 U14823 ( .A1(n12995), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11746), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U14824 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14825 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11747), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11720) );
  NAND4_X1 U14826 ( .A1(n11723), .A2(n11722), .A3(n11721), .A4(n11720), .ZN(
        n11730) );
  AOI22_X1 U14827 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11724), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14828 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14829 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14830 ( .A1(n12987), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11725) );
  NAND4_X1 U14831 ( .A1(n11728), .A2(n11727), .A3(n11726), .A4(n11725), .ZN(
        n11729) );
  NAND2_X2 U14832 ( .A1(n11837), .A2(n20286), .ZN(n12184) );
  NAND2_X1 U14833 ( .A1(n11826), .A2(n12184), .ZN(n11769) );
  AOI22_X1 U14834 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14835 ( .A1(n11854), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12839), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14836 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11724), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14837 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11747), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14838 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14839 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14840 ( .A1(n12995), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14841 ( .A1(n12987), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14842 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14843 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11743) );
  BUF_X2 U14844 ( .A(n11867), .Z(n12856) );
  AOI22_X1 U14845 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11742) );
  NAND4_X1 U14846 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11753) );
  BUF_X2 U14847 ( .A(n11746), .Z(n12812) );
  AOI22_X1 U14848 ( .A1(n12812), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12862), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14849 ( .A1(n11854), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11747), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14850 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11748) );
  NAND4_X1 U14851 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11752) );
  AOI22_X1 U14853 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14854 ( .A1(n11854), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12839), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14855 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11724), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14856 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11747), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11755) );
  NAND4_X1 U14857 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n11755), .ZN(
        n11764) );
  AOI22_X1 U14858 ( .A1(n12995), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14859 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U14860 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14861 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11759) );
  NAND4_X1 U14862 ( .A1(n11762), .A2(n11761), .A3(n11760), .A4(n11759), .ZN(
        n11763) );
  OR2_X2 U14863 ( .A1(n11764), .A2(n11763), .ZN(n11819) );
  NAND2_X1 U14864 ( .A1(n11880), .A2(n20266), .ZN(n11766) );
  NAND2_X2 U14865 ( .A1(n12398), .A2(n11822), .ZN(n12189) );
  NAND2_X1 U14866 ( .A1(n11766), .A2(n12189), .ZN(n11768) );
  NAND2_X4 U14867 ( .A1(n11822), .A2(n13019), .ZN(n12147) );
  NAND2_X1 U14868 ( .A1(n20261), .A2(n12147), .ZN(n11767) );
  NAND3_X1 U14869 ( .A1(n11769), .A2(n11768), .A3(n11767), .ZN(n11828) );
  INV_X1 U14870 ( .A(n11828), .ZN(n11791) );
  NAND2_X1 U14871 ( .A1(n11854), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11773) );
  NAND2_X1 U14872 ( .A1(n12839), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11772) );
  NAND2_X1 U14873 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11771) );
  NAND2_X1 U14874 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11770) );
  NAND2_X1 U14875 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U14876 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11776) );
  NAND2_X1 U14877 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11775) );
  NAND2_X1 U14878 ( .A1(n11747), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11774) );
  NAND2_X1 U14879 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U14880 ( .A1(n12819), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11780) );
  NAND2_X1 U14881 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11779) );
  NAND2_X1 U14882 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11786) );
  NAND2_X1 U14883 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11784) );
  NAND2_X1 U14884 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11783) );
  NAND2_X1 U14885 ( .A1(n11854), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11795) );
  NAND2_X1 U14886 ( .A1(n12839), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11794) );
  NAND2_X1 U14887 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11793) );
  NAND2_X1 U14888 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11792) );
  NAND2_X1 U14889 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11799) );
  NAND2_X1 U14890 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11798) );
  NAND2_X1 U14891 ( .A1(n12819), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11797) );
  NAND2_X1 U14892 ( .A1(n11741), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11796) );
  NAND2_X1 U14893 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11804) );
  NAND2_X1 U14894 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11802) );
  NAND2_X1 U14895 ( .A1(n11747), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11801) );
  NAND2_X1 U14896 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11807) );
  NAND2_X1 U14897 ( .A1(n12812), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11806) );
  NAND2_X1 U14898 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11805) );
  NAND2_X1 U14899 ( .A1(n12189), .A2(n12192), .ZN(n11841) );
  INV_X1 U14900 ( .A(n11841), .ZN(n11813) );
  NAND2_X1 U14901 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20928) );
  OAI21_X1 U14902 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20928), .ZN(n12139) );
  NAND2_X1 U14903 ( .A1(n20257), .A2(n12139), .ZN(n11816) );
  NOR2_X1 U14904 ( .A1(n12184), .A2(n20275), .ZN(n11815) );
  NAND2_X1 U14905 ( .A1(n12203), .A2(n11817), .ZN(n11818) );
  NAND2_X1 U14906 ( .A1(n20261), .A2(n20243), .ZN(n12314) );
  NAND2_X1 U14907 ( .A1(n12143), .A2(n11837), .ZN(n11823) );
  OR2_X2 U14908 ( .A1(n11826), .A2(n12189), .ZN(n12313) );
  INV_X1 U14909 ( .A(n13863), .ZN(n12320) );
  NAND3_X1 U14910 ( .A1(n11839), .A2(n11846), .A3(n12320), .ZN(n11827) );
  NAND2_X1 U14911 ( .A1(n11827), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11830) );
  INV_X2 U14912 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n11887) );
  INV_X1 U14913 ( .A(n11976), .ZN(n11945) );
  OAI21_X1 U14914 ( .B1(n13744), .B2(n14026), .A(n11945), .ZN(n11829) );
  AND2_X2 U14915 ( .A1(n11830), .A2(n11829), .ZN(n11831) );
  NAND2_X2 U14916 ( .A1(n11912), .A2(n11831), .ZN(n11913) );
  NAND2_X1 U14917 ( .A1(n15060), .A2(n11887), .ZN(n12881) );
  NAND2_X1 U14918 ( .A1(n20998), .A2(n20759), .ZN(n20720) );
  NAND2_X1 U14919 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20368) );
  NAND2_X1 U14920 ( .A1(n20720), .A2(n20368), .ZN(n20642) );
  OR2_X1 U14921 ( .A1(n16054), .A2(n20998), .ZN(n11910) );
  OAI21_X1 U14922 ( .B1(n12881), .B2(n20642), .A(n11910), .ZN(n11832) );
  INV_X1 U14923 ( .A(n11832), .ZN(n11833) );
  MUX2_X1 U14924 ( .A(n12881), .B(n16054), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11834) );
  NOR2_X1 U14925 ( .A1(n12320), .A2(n11837), .ZN(n11838) );
  AOI21_X1 U14926 ( .B1(n13744), .B2(n14023), .A(n11838), .ZN(n12317) );
  INV_X1 U14927 ( .A(n11839), .ZN(n11840) );
  NAND2_X1 U14928 ( .A1(n15060), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20060) );
  INV_X1 U14929 ( .A(n11836), .ZN(n14573) );
  NAND2_X1 U14930 ( .A1(n13566), .A2(n11841), .ZN(n11844) );
  INV_X1 U14931 ( .A(n13591), .ZN(n21013) );
  NAND2_X1 U14932 ( .A1(n12190), .A2(n21013), .ZN(n11843) );
  NAND2_X1 U14933 ( .A1(n11846), .A2(n20243), .ZN(n11847) );
  NAND2_X1 U14934 ( .A1(n11847), .A2(n14026), .ZN(n11848) );
  NAND3_X1 U14935 ( .A1(n12317), .A2(n11849), .A3(n11848), .ZN(n11884) );
  NAND2_X2 U14936 ( .A1(n20371), .A2(n11850), .ZN(n11921) );
  INV_X1 U14937 ( .A(n11850), .ZN(n11851) );
  NAND2_X1 U14938 ( .A1(n11852), .A2(n11851), .ZN(n20297) );
  NAND2_X1 U14939 ( .A1(n11921), .A2(n20297), .ZN(n14100) );
  INV_X1 U14940 ( .A(n14100), .ZN(n11853) );
  AOI22_X1 U14941 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U14942 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12992), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U14943 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14944 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11855) );
  NAND4_X1 U14945 ( .A1(n11858), .A2(n11857), .A3(n11856), .A4(n11855), .ZN(
        n11865) );
  AOI22_X1 U14947 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12771), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14948 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U14949 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14950 ( .A1(n12818), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11860) );
  NAND4_X1 U14951 ( .A1(n11863), .A2(n11862), .A3(n11861), .A4(n11860), .ZN(
        n11864) );
  INV_X1 U14952 ( .A(n11960), .ZN(n11866) );
  OR2_X1 U14953 ( .A1(n11866), .A2(n11977), .ZN(n11951) );
  AOI22_X1 U14954 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12856), .B1(
        n9715), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14955 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12715), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14956 ( .A1(n12861), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14957 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n12812), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11869) );
  NAND4_X1 U14958 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11878) );
  AOI22_X1 U14959 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12992), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14960 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14961 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14962 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12771), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11873) );
  NAND4_X1 U14963 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11877) );
  INV_X1 U14964 ( .A(n11959), .ZN(n11879) );
  XNOR2_X1 U14965 ( .A(n11879), .B(n11960), .ZN(n11881) );
  AOI21_X1 U14966 ( .B1(n11881), .B2(n21013), .A(n11880), .ZN(n11882) );
  NAND2_X1 U14967 ( .A1(n11883), .A2(n11882), .ZN(n11906) );
  INV_X1 U14968 ( .A(n11884), .ZN(n11885) );
  NAND2_X1 U14969 ( .A1(n12425), .A2(n11887), .ZN(n11943) );
  BUF_X1 U14970 ( .A(n12589), .Z(n12679) );
  AOI22_X1 U14971 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14972 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12985), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14973 ( .A1(n12995), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12812), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U14974 ( .A1(n12714), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11888) );
  NAND4_X1 U14975 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11897) );
  AOI22_X1 U14976 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14977 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U14978 ( .A1(n12771), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U14979 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11892) );
  NAND4_X1 U14980 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11896) );
  NAND2_X1 U14981 ( .A1(n13019), .A2(n12090), .ZN(n11900) );
  NOR2_X1 U14982 ( .A1(n11977), .A2(n12090), .ZN(n11944) );
  MUX2_X1 U14983 ( .A(n11938), .B(n11944), .S(n11959), .Z(n11898) );
  INV_X1 U14984 ( .A(n11898), .ZN(n11939) );
  NAND2_X1 U14985 ( .A1(n11943), .A2(n11939), .ZN(n11902) );
  INV_X1 U14986 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11901) );
  OAI21_X1 U14987 ( .B1(n11887), .B2(n11959), .A(n12151), .ZN(n11899) );
  OAI211_X1 U14988 ( .C1(n12167), .C2(n11901), .A(n11900), .B(n11899), .ZN(
        n11937) );
  NAND2_X1 U14989 ( .A1(n20275), .A2(n14026), .ZN(n12141) );
  NAND2_X1 U14990 ( .A1(n14025), .A2(n12192), .ZN(n11964) );
  OAI21_X1 U14991 ( .B1(n13591), .B2(n11959), .A(n11964), .ZN(n11903) );
  INV_X1 U14992 ( .A(n11903), .ZN(n11904) );
  NAND2_X1 U14993 ( .A1(n13912), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11909) );
  INV_X1 U14994 ( .A(n11906), .ZN(n11907) );
  OR2_X1 U14995 ( .A1(n11907), .A2(n13814), .ZN(n11908) );
  NAND2_X1 U14996 ( .A1(n11909), .A2(n11908), .ZN(n11967) );
  XNOR2_X1 U14997 ( .A(n11967), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13948) );
  AND2_X1 U14998 ( .A1(n11910), .A2(n13867), .ZN(n11911) );
  NAND2_X1 U14999 ( .A1(n11921), .A2(n11919), .ZN(n11917) );
  NOR2_X1 U15000 ( .A1(n16054), .A2(n20562), .ZN(n11915) );
  INV_X1 U15001 ( .A(n12881), .ZN(n11973) );
  XNOR2_X1 U15002 ( .A(n20368), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20252) );
  NAND2_X1 U15003 ( .A1(n11973), .A2(n20252), .ZN(n11918) );
  NAND2_X1 U15004 ( .A1(n11920), .A2(n11918), .ZN(n11916) );
  NAND2_X1 U15005 ( .A1(n11917), .A2(n11916), .ZN(n11969) );
  NAND4_X1 U15006 ( .A1(n11921), .A2(n11920), .A3(n11919), .A4(n11918), .ZN(
        n11922) );
  NAND2_X1 U15007 ( .A1(n11969), .A2(n11922), .ZN(n13860) );
  AOI22_X1 U15008 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15009 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12839), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U15010 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15011 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11923) );
  NAND4_X1 U15012 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11933) );
  AOI22_X1 U15013 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11931) );
  INV_X1 U15014 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21195) );
  AOI22_X1 U15015 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15016 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15017 ( .A1(n12987), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11928) );
  NAND4_X1 U15018 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(
        n11932) );
  INV_X1 U15019 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11934) );
  OAI22_X1 U15020 ( .A1(n12167), .A2(n11934), .B1(n11961), .B2(n11976), .ZN(
        n11935) );
  XNOR2_X1 U15021 ( .A(n11936), .B(n11935), .ZN(n11956) );
  INV_X1 U15022 ( .A(n11937), .ZN(n11941) );
  AND2_X1 U15023 ( .A1(n11939), .A2(n12085), .ZN(n11940) );
  NAND2_X1 U15024 ( .A1(n11943), .A2(n11942), .ZN(n11953) );
  INV_X1 U15025 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11948) );
  INV_X1 U15026 ( .A(n11944), .ZN(n11947) );
  NAND2_X1 U15027 ( .A1(n11945), .A2(n11960), .ZN(n11946) );
  OAI211_X1 U15028 ( .C1(n12167), .C2(n11948), .A(n11947), .B(n11946), .ZN(
        n11952) );
  INV_X1 U15029 ( .A(n11952), .ZN(n11949) );
  NAND3_X1 U15030 ( .A1(n12415), .A2(n11951), .A3(n11950), .ZN(n11955) );
  NAND2_X1 U15031 ( .A1(n11955), .A2(n11954), .ZN(n11957) );
  OR2_X2 U15032 ( .A1(n11956), .A2(n11957), .ZN(n12011) );
  NAND2_X1 U15033 ( .A1(n11956), .A2(n11957), .ZN(n11958) );
  INV_X1 U15034 ( .A(n12414), .ZN(n15036) );
  INV_X1 U15035 ( .A(n12141), .ZN(n12081) );
  NAND2_X1 U15036 ( .A1(n11960), .A2(n11959), .ZN(n11962) );
  AND2_X1 U15037 ( .A1(n11962), .A2(n11961), .ZN(n12017) );
  NOR2_X1 U15038 ( .A1(n11962), .A2(n11961), .ZN(n11963) );
  OAI21_X1 U15039 ( .B1(n12017), .B2(n11963), .A(n21013), .ZN(n11965) );
  NAND2_X1 U15040 ( .A1(n11965), .A2(n11964), .ZN(n11966) );
  NAND2_X1 U15041 ( .A1(n11967), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11968) );
  INV_X1 U15042 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14187) );
  NAND2_X1 U15043 ( .A1(n11914), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11975) );
  INV_X1 U15044 ( .A(n20368), .ZN(n20678) );
  NAND2_X1 U15045 ( .A1(n21136), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20478) );
  INV_X1 U15046 ( .A(n20478), .ZN(n11970) );
  NAND2_X1 U15047 ( .A1(n20678), .A2(n11970), .ZN(n20556) );
  NAND2_X1 U15048 ( .A1(n20556), .A2(n21136), .ZN(n11972) );
  NAND2_X1 U15049 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20851) );
  INV_X1 U15050 ( .A(n20851), .ZN(n11971) );
  NAND2_X1 U15051 ( .A1(n20678), .A2(n11971), .ZN(n20910) );
  INV_X1 U15052 ( .A(n16054), .ZN(n16047) );
  AOI22_X1 U15053 ( .A1(n20565), .A2(n11973), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16047), .ZN(n11974) );
  AOI22_X1 U15054 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U15055 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12839), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U15056 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15057 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11978) );
  NAND4_X1 U15058 ( .A1(n11981), .A2(n11980), .A3(n11979), .A4(n11978), .ZN(
        n11987) );
  AOI22_X1 U15059 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U15060 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15061 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15062 ( .A1(n12987), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11982) );
  NAND4_X1 U15063 ( .A1(n11985), .A2(n11984), .A3(n11983), .A4(n11982), .ZN(
        n11986) );
  AOI22_X1 U15064 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12173), .B1(
        n12145), .B2(n12016), .ZN(n11988) );
  NAND2_X1 U15065 ( .A1(n12011), .A2(n15038), .ZN(n11990) );
  OR2_X1 U15066 ( .A1(n20241), .A2(n12141), .ZN(n11993) );
  XNOR2_X1 U15067 ( .A(n12017), .B(n12016), .ZN(n11991) );
  NAND2_X1 U15068 ( .A1(n11991), .A2(n21013), .ZN(n11992) );
  NAND2_X1 U15069 ( .A1(n11993), .A2(n11992), .ZN(n13941) );
  NAND2_X1 U15070 ( .A1(n13940), .A2(n13941), .ZN(n11996) );
  NAND2_X1 U15071 ( .A1(n11994), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11995) );
  NAND2_X1 U15072 ( .A1(n11996), .A2(n11995), .ZN(n14080) );
  NAND2_X1 U15073 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12009) );
  AOI22_X1 U15074 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15075 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12819), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15076 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15077 ( .A1(n12812), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12862), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11998) );
  NAND4_X1 U15078 ( .A1(n12001), .A2(n12000), .A3(n11999), .A4(n11998), .ZN(
        n12007) );
  AOI22_X1 U15079 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U15080 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15081 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15082 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12002) );
  NAND4_X1 U15083 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n12006) );
  NAND2_X1 U15084 ( .A1(n12145), .A2(n12041), .ZN(n12008) );
  INV_X1 U15085 ( .A(n12011), .ZN(n12012) );
  NAND2_X1 U15086 ( .A1(n12014), .A2(n12013), .ZN(n12015) );
  NAND2_X1 U15087 ( .A1(n12038), .A2(n12015), .ZN(n12434) );
  INV_X1 U15088 ( .A(n12016), .ZN(n12018) );
  NOR2_X1 U15089 ( .A1(n12018), .A2(n12017), .ZN(n12042) );
  XNOR2_X1 U15090 ( .A(n12041), .B(n12042), .ZN(n12019) );
  OAI22_X1 U15091 ( .A1(n12434), .A2(n12141), .B1(n12019), .B2(n13591), .ZN(
        n12020) );
  INV_X1 U15092 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12228) );
  XNOR2_X1 U15093 ( .A(n12020), .B(n12228), .ZN(n14081) );
  NAND2_X1 U15094 ( .A1(n14080), .A2(n14081), .ZN(n12022) );
  NAND2_X1 U15095 ( .A1(n12020), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12021) );
  NAND2_X1 U15096 ( .A1(n12022), .A2(n12021), .ZN(n16250) );
  INV_X1 U15097 ( .A(n12038), .ZN(n12035) );
  NAND2_X1 U15098 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12034) );
  AOI22_X1 U15099 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15100 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12839), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U15101 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15102 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12023) );
  NAND4_X1 U15103 ( .A1(n12026), .A2(n12025), .A3(n12024), .A4(n12023), .ZN(
        n12032) );
  AOI22_X1 U15104 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15105 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15106 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15107 ( .A1(n12987), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12027) );
  NAND4_X1 U15108 ( .A1(n12030), .A2(n12029), .A3(n12028), .A4(n12027), .ZN(
        n12031) );
  NAND2_X1 U15109 ( .A1(n12145), .A2(n12065), .ZN(n12033) );
  NAND2_X1 U15110 ( .A1(n12034), .A2(n12033), .ZN(n12036) );
  INV_X1 U15111 ( .A(n12036), .ZN(n12037) );
  NAND2_X1 U15112 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  NAND2_X1 U15113 ( .A1(n12062), .A2(n12039), .ZN(n12448) );
  INV_X1 U15114 ( .A(n12448), .ZN(n12040) );
  NAND2_X1 U15115 ( .A1(n12040), .A2(n12081), .ZN(n12045) );
  NAND2_X1 U15116 ( .A1(n12042), .A2(n12041), .ZN(n12066) );
  XNOR2_X1 U15117 ( .A(n12065), .B(n12066), .ZN(n12043) );
  NAND2_X1 U15118 ( .A1(n21013), .A2(n12043), .ZN(n12044) );
  NAND2_X1 U15119 ( .A1(n12045), .A2(n12044), .ZN(n12047) );
  INV_X1 U15120 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12046) );
  XNOR2_X1 U15121 ( .A(n12047), .B(n12046), .ZN(n16249) );
  NAND2_X1 U15122 ( .A1(n16250), .A2(n16249), .ZN(n12049) );
  NAND2_X1 U15123 ( .A1(n12047), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12048) );
  AOI22_X1 U15124 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15125 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12839), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15126 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15127 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12050) );
  NAND4_X1 U15128 ( .A1(n12053), .A2(n12052), .A3(n12051), .A4(n12050), .ZN(
        n12059) );
  AOI22_X1 U15129 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15130 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15131 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15132 ( .A1(n12987), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12054) );
  NAND4_X1 U15133 ( .A1(n12057), .A2(n12056), .A3(n12055), .A4(n12054), .ZN(
        n12058) );
  NAND2_X1 U15134 ( .A1(n12145), .A2(n12077), .ZN(n12063) );
  NAND2_X1 U15135 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12060) );
  AND2_X1 U15136 ( .A1(n12063), .A2(n12060), .ZN(n12061) );
  NAND2_X1 U15137 ( .A1(n12062), .A2(n12061), .ZN(n12456) );
  INV_X1 U15138 ( .A(n12063), .ZN(n12064) );
  NAND3_X1 U15139 ( .A1(n12456), .A2(n12087), .A3(n12081), .ZN(n12071) );
  INV_X1 U15140 ( .A(n12065), .ZN(n12067) );
  NOR2_X1 U15141 ( .A1(n12067), .A2(n12066), .ZN(n12078) );
  INV_X1 U15142 ( .A(n12078), .ZN(n12068) );
  XNOR2_X1 U15143 ( .A(n12077), .B(n12068), .ZN(n12069) );
  NAND2_X1 U15144 ( .A1(n21013), .A2(n12069), .ZN(n12070) );
  NAND2_X1 U15145 ( .A1(n12071), .A2(n12070), .ZN(n12072) );
  OR2_X1 U15146 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16242) );
  NAND2_X1 U15147 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16241) );
  INV_X1 U15148 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12074) );
  NAND2_X1 U15149 ( .A1(n12145), .A2(n12090), .ZN(n12073) );
  OAI21_X1 U15150 ( .B1(n12074), .B2(n12167), .A(n12073), .ZN(n12075) );
  AND2_X1 U15151 ( .A1(n12078), .A2(n12077), .ZN(n12089) );
  XNOR2_X1 U15152 ( .A(n12090), .B(n12089), .ZN(n12079) );
  NOR2_X1 U15153 ( .A1(n13591), .A2(n12079), .ZN(n12080) );
  AOI21_X1 U15154 ( .B1(n12465), .B2(n12081), .A(n12080), .ZN(n16236) );
  INV_X1 U15155 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16235) );
  INV_X1 U15156 ( .A(n16236), .ZN(n12082) );
  NAND2_X1 U15157 ( .A1(n12082), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12083) );
  NOR2_X1 U15158 ( .A1(n12085), .A2(n12141), .ZN(n12086) );
  NAND2_X4 U15159 ( .A1(n12087), .A2(n12086), .ZN(n12088) );
  NAND2_X1 U15160 ( .A1(n12090), .A2(n12089), .ZN(n12091) );
  OR2_X1 U15161 ( .A1(n12091), .A2(n13591), .ZN(n12092) );
  NAND2_X1 U15162 ( .A1(n12088), .A2(n12092), .ZN(n14292) );
  AND2_X1 U15163 ( .A1(n14292), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12094) );
  INV_X1 U15164 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15030) );
  NAND2_X1 U15165 ( .A1(n12088), .A2(n15030), .ZN(n12096) );
  INV_X1 U15166 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15002) );
  NAND2_X1 U15167 ( .A1(n12088), .A2(n15002), .ZN(n12097) );
  NAND2_X1 U15168 ( .A1(n16212), .A2(n12097), .ZN(n14895) );
  INV_X1 U15169 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15017) );
  NAND2_X1 U15170 ( .A1(n12088), .A2(n15017), .ZN(n14893) );
  NAND2_X1 U15171 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U15172 ( .A1(n12088), .A2(n12098), .ZN(n14891) );
  NAND2_X1 U15173 ( .A1(n14893), .A2(n14891), .ZN(n12099) );
  NOR2_X1 U15174 ( .A1(n14895), .A2(n12099), .ZN(n16214) );
  INV_X1 U15175 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16317) );
  NAND2_X1 U15176 ( .A1(n12088), .A2(n16317), .ZN(n12100) );
  NAND2_X1 U15177 ( .A1(n16214), .A2(n12100), .ZN(n14877) );
  OR2_X1 U15178 ( .A1(n12088), .A2(n16317), .ZN(n12101) );
  INV_X1 U15179 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12102) );
  NAND2_X1 U15180 ( .A1(n12088), .A2(n12102), .ZN(n14964) );
  NAND2_X1 U15181 ( .A1(n14967), .A2(n14964), .ZN(n12103) );
  AOI21_X1 U15182 ( .B1(n14877), .B2(n12104), .A(n12103), .ZN(n14868) );
  NAND2_X1 U15183 ( .A1(n14868), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12107) );
  NOR2_X1 U15184 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12105) );
  NAND2_X1 U15185 ( .A1(n14892), .A2(n14889), .ZN(n14866) );
  OAI21_X1 U15186 ( .B1(n14865), .B2(n12107), .A(n12106), .ZN(n12108) );
  INV_X1 U15187 ( .A(n12108), .ZN(n12112) );
  NOR2_X1 U15188 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12109) );
  INV_X1 U15189 ( .A(n12110), .ZN(n12111) );
  INV_X1 U15190 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21294) );
  INV_X1 U15191 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16292) );
  NAND2_X1 U15192 ( .A1(n21294), .A2(n16292), .ZN(n12113) );
  INV_X1 U15193 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16063) );
  INV_X1 U15194 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16069) );
  XNOR2_X1 U15195 ( .A(n12088), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14860) );
  NAND2_X1 U15196 ( .A1(n14861), .A2(n14860), .ZN(n14851) );
  AND3_X1 U15197 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12339) );
  INV_X1 U15198 ( .A(n12339), .ZN(n12114) );
  INV_X1 U15199 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14833) );
  INV_X1 U15200 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14845) );
  INV_X1 U15201 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12371) );
  NAND3_X1 U15202 ( .A1(n14833), .A2(n14845), .A3(n12371), .ZN(n14797) );
  NAND2_X1 U15203 ( .A1(n12115), .A2(n9721), .ZN(n14820) );
  NAND2_X1 U15204 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12369) );
  INV_X1 U15205 ( .A(n12369), .ZN(n12116) );
  NAND2_X1 U15206 ( .A1(n12116), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14796) );
  NAND2_X1 U15207 ( .A1(n12358), .A2(n14796), .ZN(n12118) );
  NAND2_X1 U15208 ( .A1(n12117), .A2(n12088), .ZN(n12360) );
  NAND3_X1 U15209 ( .A1(n12118), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n12360), .ZN(n14808) );
  NAND2_X1 U15210 ( .A1(n14820), .A2(n14808), .ZN(n14807) );
  NOR2_X1 U15211 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14923) );
  INV_X1 U15212 ( .A(n14923), .ZN(n12119) );
  AND2_X1 U15213 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14924) );
  NAND2_X1 U15214 ( .A1(n14807), .A2(n14924), .ZN(n12381) );
  INV_X1 U15215 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12382) );
  XNOR2_X1 U15216 ( .A(n12088), .B(n12382), .ZN(n12121) );
  XNOR2_X1 U15217 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12132) );
  NAND2_X1 U15218 ( .A1(n20759), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12146) );
  NAND2_X1 U15219 ( .A1(n12132), .A2(n12133), .ZN(n12123) );
  NAND2_X1 U15220 ( .A1(n20998), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12122) );
  NAND2_X1 U15221 ( .A1(n12123), .A2(n12122), .ZN(n12137) );
  XNOR2_X1 U15222 ( .A(n21244), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12136) );
  NAND2_X1 U15223 ( .A1(n12137), .A2(n12136), .ZN(n12125) );
  NAND2_X1 U15224 ( .A1(n20562), .A2(n21244), .ZN(n12124) );
  NAND2_X1 U15225 ( .A1(n12125), .A2(n12124), .ZN(n12135) );
  MUX2_X1 U15226 ( .A(n21136), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12134) );
  NAND2_X1 U15227 ( .A1(n12135), .A2(n12134), .ZN(n12127) );
  NAND2_X1 U15228 ( .A1(n21136), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12126) );
  NAND2_X1 U15229 ( .A1(n12127), .A2(n12126), .ZN(n12131) );
  INV_X1 U15230 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13878) );
  NOR2_X1 U15231 ( .A1(n13878), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12128) );
  XNOR2_X1 U15232 ( .A(n12133), .B(n12132), .ZN(n12155) );
  XNOR2_X1 U15233 ( .A(n12135), .B(n12134), .ZN(n12169) );
  XNOR2_X1 U15234 ( .A(n12137), .B(n12136), .ZN(n12162) );
  NOR4_X1 U15235 ( .A1(n12172), .A2(n12155), .A3(n12169), .A4(n12162), .ZN(
        n12138) );
  NOR2_X1 U15236 ( .A1(n12142), .A2(n12138), .ZN(n13558) );
  OR2_X1 U15237 ( .A1(n12139), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n16073) );
  NAND2_X1 U15238 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21018) );
  INV_X1 U15239 ( .A(n21018), .ZN(n20924) );
  AOI21_X1 U15240 ( .B1(n14026), .B2(n16073), .A(n20924), .ZN(n12140) );
  NAND2_X1 U15241 ( .A1(n13558), .A2(n12140), .ZN(n12188) );
  NAND2_X1 U15242 ( .A1(n12170), .A2(n12142), .ZN(n12182) );
  NAND2_X1 U15243 ( .A1(n12142), .A2(n12145), .ZN(n12180) );
  AOI22_X1 U15244 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12143), .B1(n12145), 
        .B2(n14026), .ZN(n12157) );
  INV_X1 U15245 ( .A(n12157), .ZN(n12144) );
  NOR2_X1 U15246 ( .A1(n12155), .A2(n12144), .ZN(n12154) );
  OAI21_X1 U15247 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20759), .A(
        n12146), .ZN(n12148) );
  NOR2_X1 U15248 ( .A1(n12164), .A2(n12148), .ZN(n12153) );
  INV_X1 U15249 ( .A(n12148), .ZN(n12150) );
  NAND2_X1 U15250 ( .A1(n12143), .A2(n20243), .ZN(n12149) );
  NAND2_X1 U15251 ( .A1(n12149), .A2(n20257), .ZN(n12163) );
  OAI211_X1 U15252 ( .C1(n12147), .C2(n12151), .A(n12150), .B(n12163), .ZN(
        n12152) );
  OAI21_X1 U15253 ( .B1(n12170), .B2(n12153), .A(n12152), .ZN(n12156) );
  NAND2_X1 U15254 ( .A1(n12154), .A2(n12156), .ZN(n12161) );
  NAND2_X1 U15255 ( .A1(n12157), .A2(n14026), .ZN(n12175) );
  OAI211_X1 U15256 ( .C1(n12157), .C2(n12156), .A(n12155), .B(n12175), .ZN(
        n12160) );
  NAND2_X1 U15257 ( .A1(n12173), .A2(n12162), .ZN(n12158) );
  OAI211_X1 U15258 ( .C1(n12164), .C2(n12162), .A(n12158), .B(n12163), .ZN(
        n12159) );
  NAND3_X1 U15259 ( .A1(n12161), .A2(n12160), .A3(n12159), .ZN(n12166) );
  AOI22_X1 U15260 ( .A1(n12167), .A2(n12169), .B1(n12166), .B2(n12165), .ZN(
        n12168) );
  AOI21_X1 U15261 ( .B1(n12170), .B2(n12169), .A(n12168), .ZN(n12177) );
  INV_X1 U15262 ( .A(n12172), .ZN(n12171) );
  NOR2_X1 U15263 ( .A1(n12173), .A2(n12171), .ZN(n12176) );
  NAND2_X1 U15264 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  OAI22_X1 U15265 ( .A1(n12177), .A2(n12176), .B1(n12175), .B2(n12174), .ZN(
        n12178) );
  AOI21_X1 U15266 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n11887), .A(
        n12178), .ZN(n12179) );
  NAND2_X1 U15267 ( .A1(n12180), .A2(n12179), .ZN(n12181) );
  NAND2_X1 U15268 ( .A1(n20257), .A2(n16073), .ZN(n14028) );
  NAND2_X1 U15269 ( .A1(n14028), .A2(n21018), .ZN(n12185) );
  OAI211_X1 U15270 ( .C1(n13768), .C2(n12185), .A(n20243), .B(n12184), .ZN(
        n12186) );
  NAND2_X1 U15271 ( .A1(n14565), .A2(n12186), .ZN(n12187) );
  MUX2_X1 U15272 ( .A(n12188), .B(n12187), .S(n12193), .Z(n12201) );
  INV_X1 U15273 ( .A(n12189), .ZN(n12197) );
  NAND2_X1 U15274 ( .A1(n12197), .A2(n13019), .ZN(n12191) );
  AND2_X1 U15275 ( .A1(n12191), .A2(n11825), .ZN(n12321) );
  NAND2_X1 U15276 ( .A1(n12313), .A2(n14025), .ZN(n12194) );
  NAND4_X1 U15277 ( .A1(n12321), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n12879) );
  AOI21_X1 U15278 ( .B1(n12197), .B2(n14026), .A(n14025), .ZN(n12198) );
  AND2_X1 U15279 ( .A1(n12199), .A2(n12198), .ZN(n12318) );
  AOI21_X1 U15280 ( .B1(n12879), .B2(n13559), .A(n12318), .ZN(n13766) );
  NAND3_X1 U15281 ( .A1(n14569), .A2(n15048), .A3(n14026), .ZN(n12200) );
  NAND3_X1 U15282 ( .A1(n12201), .A2(n13766), .A3(n12200), .ZN(n12202) );
  NAND2_X1 U15283 ( .A1(n16054), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20057) );
  AOI22_X1 U15284 ( .A1(n14567), .A2(n14026), .B1(n12309), .B2(n20270), .ZN(
        n12209) );
  INV_X1 U15285 ( .A(n12879), .ZN(n13016) );
  OR2_X1 U15286 ( .A1(n12207), .A2(n14023), .ZN(n12208) );
  NAND2_X1 U15287 ( .A1(n13016), .A2(n12208), .ZN(n14566) );
  AND3_X1 U15288 ( .A1(n12204), .A2(n12209), .A3(n14566), .ZN(n12210) );
  NAND2_X1 U15289 ( .A1(n10113), .A2(n16360), .ZN(n12345) );
  INV_X1 U15290 ( .A(n12217), .ZN(n13048) );
  INV_X1 U15291 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U15292 ( .A1(n12300), .A2(n12212), .ZN(n12214) );
  INV_X1 U15293 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13685) );
  NAND2_X1 U15294 ( .A1(n13683), .A2(n13685), .ZN(n12213) );
  NAND3_X1 U15295 ( .A1(n12214), .A2(n12293), .A3(n12213), .ZN(n12215) );
  NAND2_X1 U15296 ( .A1(n12300), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12219) );
  INV_X1 U15297 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14034) );
  NAND2_X1 U15298 ( .A1(n12293), .A2(n14034), .ZN(n12218) );
  NAND2_X1 U15299 ( .A1(n12219), .A2(n12218), .ZN(n13805) );
  XNOR2_X1 U15300 ( .A(n12220), .B(n13805), .ZN(n13684) );
  NAND2_X1 U15301 ( .A1(n13684), .A2(n13683), .ZN(n13682) );
  NAND2_X1 U15302 ( .A1(n13682), .A2(n12220), .ZN(n13954) );
  OR2_X1 U15303 ( .A1(n12306), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12224) );
  INV_X1 U15304 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13951) );
  NAND2_X1 U15305 ( .A1(n12300), .A2(n13951), .ZN(n12222) );
  INV_X1 U15306 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14522) );
  NAND2_X1 U15307 ( .A1(n13683), .A2(n14522), .ZN(n12221) );
  NAND3_X1 U15308 ( .A1(n12222), .A2(n12293), .A3(n12221), .ZN(n12223) );
  MUX2_X1 U15309 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12227) );
  OAI21_X1 U15310 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13804), .A(
        n12227), .ZN(n13989) );
  OR2_X1 U15311 ( .A1(n12306), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n12232) );
  NAND2_X1 U15312 ( .A1(n12300), .A2(n12228), .ZN(n12230) );
  INV_X1 U15313 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14054) );
  NAND2_X1 U15314 ( .A1(n13683), .A2(n14054), .ZN(n12229) );
  NAND3_X1 U15315 ( .A1(n12230), .A2(n12293), .A3(n12229), .ZN(n12231) );
  NAND2_X1 U15316 ( .A1(n12232), .A2(n12231), .ZN(n13962) );
  MUX2_X1 U15317 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12233) );
  OAI21_X1 U15318 ( .B1(n13804), .B2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12233), .ZN(n13937) );
  OR2_X1 U15319 ( .A1(n12306), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n12238) );
  INV_X1 U15320 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16345) );
  NAND2_X1 U15321 ( .A1(n12300), .A2(n16345), .ZN(n12236) );
  INV_X1 U15322 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14093) );
  NAND2_X1 U15323 ( .A1(n13683), .A2(n14093), .ZN(n12235) );
  NAND3_X1 U15324 ( .A1(n12236), .A2(n12293), .A3(n12235), .ZN(n12237) );
  INV_X1 U15325 ( .A(n12298), .ZN(n12239) );
  INV_X1 U15326 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20152) );
  NAND2_X1 U15327 ( .A1(n12239), .A2(n20152), .ZN(n12243) );
  NAND2_X1 U15328 ( .A1(n13683), .A2(n20152), .ZN(n12241) );
  NAND2_X1 U15329 ( .A1(n12293), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12240) );
  NAND3_X1 U15330 ( .A1(n12241), .A2(n12300), .A3(n12240), .ZN(n12242) );
  MUX2_X1 U15331 ( .A(n12306), .B(n12300), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12247) );
  INV_X1 U15332 ( .A(n12300), .ZN(n12244) );
  NAND2_X1 U15333 ( .A1(n12244), .A2(n14572), .ZN(n12278) );
  NAND2_X1 U15334 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n14572), .ZN(
        n12245) );
  AND2_X1 U15335 ( .A1(n12278), .A2(n12245), .ZN(n12246) );
  NAND2_X1 U15336 ( .A1(n12247), .A2(n12246), .ZN(n14216) );
  INV_X1 U15337 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20147) );
  NAND2_X1 U15338 ( .A1(n13683), .A2(n20147), .ZN(n12249) );
  NAND2_X1 U15339 ( .A1(n12293), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12248) );
  NAND3_X1 U15340 ( .A1(n12249), .A2(n12300), .A3(n12248), .ZN(n12250) );
  OAI21_X1 U15341 ( .B1(n12298), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12250), .ZN(
        n14396) );
  OR2_X1 U15342 ( .A1(n12306), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n12255) );
  INV_X1 U15343 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14906) );
  NAND2_X1 U15344 ( .A1(n12300), .A2(n14906), .ZN(n12253) );
  INV_X1 U15345 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n12251) );
  NAND2_X1 U15346 ( .A1(n13683), .A2(n12251), .ZN(n12252) );
  NAND3_X1 U15347 ( .A1(n12253), .A2(n12293), .A3(n12252), .ZN(n12254) );
  MUX2_X1 U15348 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12257) );
  OR2_X1 U15349 ( .A1(n13804), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12256) );
  MUX2_X1 U15350 ( .A(n12306), .B(n12300), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12260) );
  NAND2_X1 U15351 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14572), .ZN(
        n12258) );
  AND2_X1 U15352 ( .A1(n12278), .A2(n12258), .ZN(n12259) );
  NAND2_X1 U15353 ( .A1(n12260), .A2(n12259), .ZN(n14362) );
  MUX2_X1 U15354 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12261) );
  OAI21_X1 U15355 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13804), .A(
        n12261), .ZN(n14407) );
  MUX2_X1 U15356 ( .A(n12306), .B(n12300), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12263) );
  NAND2_X1 U15357 ( .A1(n14572), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12262) );
  MUX2_X1 U15358 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12264) );
  OAI21_X1 U15359 ( .B1(n13804), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12264), .ZN(n14435) );
  OR2_X1 U15360 ( .A1(n12306), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n12269) );
  INV_X1 U15361 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16303) );
  NAND2_X1 U15362 ( .A1(n12300), .A2(n16303), .ZN(n12267) );
  INV_X1 U15363 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n12265) );
  NAND2_X1 U15364 ( .A1(n13683), .A2(n12265), .ZN(n12266) );
  NAND3_X1 U15365 ( .A1(n12267), .A2(n12293), .A3(n12266), .ZN(n12268) );
  NAND2_X1 U15366 ( .A1(n12269), .A2(n12268), .ZN(n14474) );
  MUX2_X1 U15367 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12270) );
  OAI21_X1 U15368 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13804), .A(
        n12270), .ZN(n14724) );
  OR2_X1 U15369 ( .A1(n12306), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n12274) );
  NAND2_X1 U15370 ( .A1(n12300), .A2(n21294), .ZN(n12272) );
  INV_X1 U15371 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16119) );
  NAND2_X1 U15372 ( .A1(n13683), .A2(n16119), .ZN(n12271) );
  NAND3_X1 U15373 ( .A1(n12272), .A2(n12217), .A3(n12271), .ZN(n12273) );
  MUX2_X1 U15374 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12276) );
  OR2_X1 U15375 ( .A1(n13804), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12275) );
  AND2_X1 U15376 ( .A1(n12276), .A2(n12275), .ZN(n14658) );
  MUX2_X1 U15377 ( .A(n12306), .B(n12300), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12280) );
  NAND2_X1 U15378 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n14572), .ZN(
        n12277) );
  AND2_X1 U15379 ( .A1(n12278), .A2(n12277), .ZN(n12279) );
  NAND2_X1 U15380 ( .A1(n12280), .A2(n12279), .ZN(n14709) );
  MUX2_X1 U15381 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12281) );
  OAI21_X1 U15382 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13804), .A(
        n12281), .ZN(n14705) );
  MUX2_X1 U15383 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12282) );
  OAI21_X1 U15384 ( .B1(n13804), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12282), .ZN(n12283) );
  INV_X1 U15385 ( .A(n12283), .ZN(n14694) );
  OR2_X1 U15386 ( .A1(n12306), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n12288) );
  INV_X1 U15387 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12284) );
  NAND2_X1 U15388 ( .A1(n12300), .A2(n12284), .ZN(n12286) );
  INV_X1 U15389 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16189) );
  NAND2_X1 U15390 ( .A1(n13683), .A2(n16189), .ZN(n12285) );
  NAND3_X1 U15391 ( .A1(n12286), .A2(n12293), .A3(n12285), .ZN(n12287) );
  NAND2_X1 U15392 ( .A1(n12288), .A2(n12287), .ZN(n16095) );
  OR2_X1 U15393 ( .A1(n12306), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U15394 ( .A1(n12300), .A2(n14833), .ZN(n12290) );
  INV_X1 U15395 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14691) );
  NAND2_X1 U15396 ( .A1(n13683), .A2(n14691), .ZN(n12289) );
  NAND3_X1 U15397 ( .A1(n12290), .A2(n12293), .A3(n12289), .ZN(n12291) );
  NAND2_X1 U15398 ( .A1(n12292), .A2(n12291), .ZN(n14651) );
  MUX2_X1 U15399 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12295) );
  OR2_X1 U15400 ( .A1(n13804), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12294) );
  AND2_X1 U15401 ( .A1(n12295), .A2(n12294), .ZN(n12367) );
  MUX2_X1 U15402 ( .A(n12306), .B(n12300), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12297) );
  NAND2_X1 U15403 ( .A1(n14572), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12296) );
  AND2_X1 U15404 ( .A1(n12297), .A2(n12296), .ZN(n14629) );
  MUX2_X1 U15405 ( .A(n12298), .B(n12293), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12299) );
  OAI21_X1 U15406 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13804), .A(
        n12299), .ZN(n14611) );
  MUX2_X1 U15407 ( .A(n12306), .B(n12300), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12302) );
  NAND2_X1 U15408 ( .A1(n14572), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12301) );
  AND2_X1 U15409 ( .A1(n12302), .A2(n12301), .ZN(n14595) );
  OR2_X1 U15410 ( .A1(n13804), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12305) );
  INV_X1 U15411 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n12303) );
  NAND2_X1 U15412 ( .A1(n13683), .A2(n12303), .ZN(n12304) );
  NAND2_X1 U15413 ( .A1(n12305), .A2(n12304), .ZN(n13050) );
  OAI22_X1 U15414 ( .A1(n13050), .A2(n13048), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12306), .ZN(n12307) );
  OR2_X1 U15415 ( .A1(n14597), .A2(n12307), .ZN(n12308) );
  NAND2_X1 U15416 ( .A1(n14567), .A2(n20257), .ZN(n16051) );
  NAND2_X1 U15417 ( .A1(n12309), .A2(n13019), .ZN(n12310) );
  AND2_X1 U15418 ( .A1(n16051), .A2(n12310), .ZN(n12311) );
  NAND2_X1 U15419 ( .A1(n12147), .A2(n14025), .ZN(n12319) );
  NAND2_X1 U15420 ( .A1(n12319), .A2(n14026), .ZN(n12312) );
  NOR2_X1 U15421 ( .A1(n12313), .A2(n12312), .ZN(n12316) );
  INV_X1 U15422 ( .A(n12314), .ZN(n12315) );
  AOI21_X1 U15423 ( .B1(n13804), .B2(n20266), .A(n12315), .ZN(n12323) );
  INV_X1 U15424 ( .A(n14562), .ZN(n13751) );
  NAND2_X1 U15425 ( .A1(n12196), .A2(n14026), .ZN(n13868) );
  OAI21_X1 U15426 ( .B1(n20243), .B2(n13745), .A(n12317), .ZN(n12326) );
  INV_X1 U15427 ( .A(n12318), .ZN(n12325) );
  NAND3_X1 U15428 ( .A1(n12321), .A2(n12320), .A3(n12319), .ZN(n12322) );
  NAND2_X1 U15429 ( .A1(n12322), .A2(n14026), .ZN(n12324) );
  NAND3_X1 U15430 ( .A1(n12325), .A2(n12324), .A3(n12323), .ZN(n13748) );
  NOR2_X1 U15431 ( .A1(n12326), .A2(n13748), .ZN(n12327) );
  NAND2_X1 U15432 ( .A1(n16333), .A2(n14974), .ZN(n13817) );
  INV_X1 U15433 ( .A(n13817), .ZN(n12328) );
  NAND2_X1 U15434 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16280) );
  NOR2_X1 U15435 ( .A1(n16063), .A2(n16292), .ZN(n16068) );
  NAND2_X1 U15436 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13984) );
  NAND2_X1 U15437 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16337) );
  INV_X1 U15438 ( .A(n16337), .ZN(n16332) );
  NAND2_X1 U15439 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16332), .ZN(
        n12329) );
  OR2_X1 U15440 ( .A1(n13984), .A2(n12329), .ZN(n15014) );
  INV_X1 U15441 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16322) );
  NOR2_X1 U15442 ( .A1(n14906), .A2(n15030), .ZN(n16323) );
  NAND4_X1 U15443 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n16323), .ZN(n15013) );
  NOR2_X1 U15444 ( .A1(n16322), .A2(n15013), .ZN(n15020) );
  NAND2_X1 U15445 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15020), .ZN(
        n12330) );
  NOR2_X1 U15446 ( .A1(n15014), .A2(n12330), .ZN(n14998) );
  NAND4_X1 U15447 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16296) );
  NOR2_X1 U15448 ( .A1(n21294), .A2(n16296), .ZN(n12338) );
  AND2_X1 U15449 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12338), .ZN(
        n14955) );
  NAND2_X1 U15450 ( .A1(n14998), .A2(n14955), .ZN(n14956) );
  INV_X1 U15451 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15051) );
  OAI21_X1 U15452 ( .B1(n15051), .B2(n12212), .A(n13951), .ZN(n13985) );
  NAND3_X1 U15453 ( .A1(n16332), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n13985), .ZN(n15007) );
  NOR2_X1 U15454 ( .A1(n12330), .A2(n15007), .ZN(n16318) );
  AOI21_X1 U15455 ( .B1(n14955), .B2(n16318), .A(n16333), .ZN(n12332) );
  OR2_X2 U15456 ( .A1(n12881), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20100) );
  NAND2_X1 U15457 ( .A1(n12331), .A2(n20100), .ZN(n14971) );
  OAI21_X1 U15458 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14974), .A(
        n14971), .ZN(n15012) );
  AOI211_X1 U15459 ( .C1(n16338), .C2(n14956), .A(n12332), .B(n15012), .ZN(
        n16289) );
  NOR2_X1 U15460 ( .A1(n16340), .A2(n15012), .ZN(n15025) );
  AOI21_X1 U15461 ( .B1(n16068), .B2(n16289), .A(n15025), .ZN(n16278) );
  AOI21_X1 U15462 ( .B1(n16340), .B2(n16280), .A(n16278), .ZN(n16276) );
  OAI21_X1 U15463 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16333), .A(
        n16276), .ZN(n14942) );
  NAND2_X1 U15464 ( .A1(n12369), .A2(n16338), .ZN(n12334) );
  OR2_X1 U15465 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n16333), .ZN(
        n12333) );
  NAND2_X1 U15466 ( .A1(n12334), .A2(n12333), .ZN(n12335) );
  NOR2_X1 U15467 ( .A1(n14942), .A2(n12335), .ZN(n12370) );
  NAND2_X1 U15468 ( .A1(n12370), .A2(n14979), .ZN(n12392) );
  INV_X1 U15469 ( .A(n14924), .ZN(n12340) );
  NAND2_X1 U15470 ( .A1(n12392), .A2(n12340), .ZN(n12336) );
  NAND2_X1 U15471 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n12370), .ZN(
        n14933) );
  OAI21_X1 U15472 ( .B1(n12371), .B2(n14933), .A(n12392), .ZN(n14922) );
  AND2_X1 U15473 ( .A1(n12336), .A2(n14922), .ZN(n12391) );
  OR2_X1 U15474 ( .A1(n12391), .A2(n12382), .ZN(n12342) );
  INV_X2 U15475 ( .A(n20100), .ZN(n20232) );
  NAND2_X1 U15476 ( .A1(n13958), .A2(n16318), .ZN(n14954) );
  AND2_X1 U15477 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14998), .ZN(
        n14970) );
  NAND2_X1 U15478 ( .A1(n15016), .A2(n14970), .ZN(n14941) );
  NAND4_X1 U15479 ( .A1(n12339), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n12338), .A4(n16304), .ZN(n16269) );
  NOR2_X1 U15480 ( .A1(n14796), .A2(n16269), .ZN(n14935) );
  NAND2_X1 U15481 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n14935), .ZN(
        n16261) );
  NOR2_X1 U15482 ( .A1(n12340), .A2(n16261), .ZN(n12388) );
  AOI22_X1 U15483 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n20232), .B1(n12388), 
        .B2(n12382), .ZN(n12341) );
  INV_X1 U15484 ( .A(n16436), .ZN(n19404) );
  OAI21_X1 U15485 ( .B1(n12347), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n12348), .ZN(n12349) );
  INV_X1 U15486 ( .A(n12349), .ZN(n15145) );
  OAI21_X1 U15487 ( .B1(n19409), .B2(n15138), .A(n12350), .ZN(n12352) );
  NOR2_X1 U15488 ( .A1(n15225), .A2(n15509), .ZN(n12351) );
  AOI211_X1 U15489 ( .C1(n19398), .C2(n15145), .A(n12352), .B(n12351), .ZN(
        n12355) );
  OAI21_X1 U15490 ( .B1(n15368), .B2(n12357), .A(n12356), .ZN(P2_U2992) );
  INV_X1 U15491 ( .A(n14841), .ZN(n12359) );
  NAND2_X1 U15492 ( .A1(n12359), .A2(n9721), .ZN(n14840) );
  OR2_X2 U15493 ( .A1(n14840), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12364) );
  NAND2_X1 U15494 ( .A1(n12360), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14832) );
  OAI21_X2 U15495 ( .B1(n12364), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12363), .ZN(n12365) );
  INV_X1 U15496 ( .A(n14831), .ZN(n12366) );
  OR2_X1 U15497 ( .A1(n14649), .A2(n12367), .ZN(n12368) );
  NAND2_X1 U15498 ( .A1(n14628), .A2(n12368), .ZN(n14689) );
  INV_X1 U15499 ( .A(n14689), .ZN(n12376) );
  NOR3_X1 U15500 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n12369), .A3(
        n16269), .ZN(n14934) );
  AOI21_X1 U15501 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n20232), .A(n14934), 
        .ZN(n12374) );
  INV_X1 U15502 ( .A(n12370), .ZN(n12372) );
  NAND2_X1 U15503 ( .A1(n12378), .A2(n12377), .ZN(P1_U3006) );
  INV_X1 U15504 ( .A(n12381), .ZN(n12384) );
  INV_X1 U15505 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15052) );
  AOI22_X1 U15506 ( .A1(n13804), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14572), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13054) );
  MUX2_X1 U15507 ( .A(n13054), .B(n12217), .S(n13049), .Z(n12387) );
  AOI22_X1 U15508 ( .A1(n13804), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14572), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12386) );
  XNOR2_X2 U15509 ( .A(n12387), .B(n12386), .ZN(n14685) );
  INV_X1 U15510 ( .A(n14685), .ZN(n12396) );
  NAND2_X1 U15511 ( .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n12388), .ZN(
        n14916) );
  NAND2_X1 U15512 ( .A1(n15052), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12394) );
  OAI21_X1 U15513 ( .B1(n14979), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12389) );
  INV_X1 U15514 ( .A(n12389), .ZN(n12390) );
  NAND2_X1 U15515 ( .A1(n12391), .A2(n12390), .ZN(n14918) );
  NAND3_X1 U15516 ( .A1(n14918), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12392), .ZN(n12393) );
  NAND2_X1 U15517 ( .A1(n20232), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14511) );
  OAI211_X1 U15518 ( .C1(n14916), .C2(n12394), .A(n12393), .B(n14511), .ZN(
        n12395) );
  OAI21_X1 U15519 ( .B1(n14515), .B2(n16370), .A(n12397), .ZN(P1_U3000) );
  INV_X1 U15520 ( .A(n20241), .ZN(n12399) );
  NAND2_X1 U15521 ( .A1(n20280), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12558) );
  INV_X1 U15522 ( .A(n12184), .ZN(n13024) );
  NAND2_X1 U15523 ( .A1(n13024), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12435) );
  INV_X1 U15524 ( .A(n12872), .ZN(n12409) );
  INV_X1 U15525 ( .A(n12409), .ZN(n13006) );
  NAND2_X1 U15526 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12401) );
  INV_X1 U15527 ( .A(n12401), .ZN(n12403) );
  INV_X1 U15528 ( .A(n12438), .ZN(n12402) );
  OAI21_X1 U15529 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12403), .A(
        n12402), .ZN(n20114) );
  AOI22_X1 U15530 ( .A1(n13006), .A2(n20114), .B1(n13013), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12405) );
  INV_X2 U15531 ( .A(n9821), .ZN(n13014) );
  NAND2_X1 U15532 ( .A1(n13014), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12404) );
  OAI211_X1 U15533 ( .C1(n12435), .C2(n13752), .A(n12405), .B(n12404), .ZN(
        n12406) );
  INV_X1 U15534 ( .A(n12406), .ZN(n12407) );
  INV_X1 U15535 ( .A(n21244), .ZN(n13862) );
  XNOR2_X1 U15536 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20130) );
  AOI21_X1 U15537 ( .B1(n12872), .B2(n20130), .A(n13013), .ZN(n12411) );
  NAND2_X1 U15538 ( .A1(n13014), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12410) );
  OAI211_X1 U15539 ( .C1(n12435), .C2(n13862), .A(n12411), .B(n12410), .ZN(
        n12412) );
  INV_X1 U15540 ( .A(n12412), .ZN(n12413) );
  NAND2_X1 U15541 ( .A1(n13013), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12433) );
  INV_X1 U15542 ( .A(n12415), .ZN(n12416) );
  NAND2_X1 U15543 ( .A1(n13889), .A2(n12582), .ZN(n12422) );
  NAND2_X1 U15544 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n21011), .ZN(
        n12419) );
  NAND2_X1 U15545 ( .A1(n13014), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n12418) );
  OAI211_X1 U15546 ( .C1(n12435), .C2(n13867), .A(n12419), .B(n12418), .ZN(
        n12420) );
  INV_X1 U15547 ( .A(n12420), .ZN(n12421) );
  NAND2_X1 U15548 ( .A1(n12422), .A2(n12421), .ZN(n13681) );
  NAND2_X1 U15549 ( .A1(n12423), .A2(n20280), .ZN(n12424) );
  NAND2_X1 U15550 ( .A1(n12424), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13800) );
  NAND2_X1 U15551 ( .A1(n21011), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12428) );
  NAND2_X1 U15552 ( .A1(n13014), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12427) );
  OAI211_X1 U15553 ( .C1(n12435), .C2(n12426), .A(n12428), .B(n12427), .ZN(
        n12429) );
  AOI21_X1 U15554 ( .B1(n20372), .B2(n12582), .A(n12429), .ZN(n12430) );
  OR2_X1 U15555 ( .A1(n13800), .A2(n12430), .ZN(n13801) );
  INV_X1 U15556 ( .A(n12430), .ZN(n13802) );
  OR2_X1 U15557 ( .A1(n13802), .A2(n12409), .ZN(n12431) );
  NAND2_X1 U15558 ( .A1(n13801), .A2(n12431), .ZN(n13680) );
  NAND2_X1 U15559 ( .A1(n13681), .A2(n13680), .ZN(n13823) );
  INV_X1 U15560 ( .A(n13823), .ZN(n12432) );
  NAND2_X1 U15561 ( .A1(n13837), .A2(n13838), .ZN(n13836) );
  INV_X1 U15562 ( .A(n12434), .ZN(n12443) );
  INV_X1 U15563 ( .A(n12435), .ZN(n12436) );
  NAND2_X1 U15564 ( .A1(n12436), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12441) );
  INV_X1 U15565 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21293) );
  AOI21_X1 U15566 ( .B1(n21293), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12437) );
  AOI21_X1 U15567 ( .B1(n13014), .B2(P1_EAX_REG_4__SCAN_IN), .A(n12437), .ZN(
        n12440) );
  NOR2_X1 U15568 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12438), .ZN(
        n12439) );
  NOR2_X1 U15569 ( .A1(n12444), .A2(n12439), .ZN(n14083) );
  AOI22_X1 U15570 ( .A1(n12441), .A2(n12440), .B1(n12872), .B2(n14083), .ZN(
        n12442) );
  NOR2_X2 U15571 ( .A1(n13836), .A2(n13961), .ZN(n13933) );
  NOR2_X1 U15572 ( .A1(n12444), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12445) );
  NOR2_X1 U15573 ( .A1(n12449), .A2(n12445), .ZN(n20105) );
  INV_X1 U15574 ( .A(n13013), .ZN(n12623) );
  INV_X1 U15575 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16257) );
  OAI22_X1 U15576 ( .A1(n20105), .A2(n12409), .B1(n12623), .B2(n16257), .ZN(
        n12446) );
  AOI21_X1 U15577 ( .B1(n13014), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12446), .ZN(
        n12447) );
  NAND2_X1 U15578 ( .A1(n13933), .A2(n13936), .ZN(n13935) );
  INV_X1 U15579 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12454) );
  INV_X1 U15580 ( .A(n12459), .ZN(n12460) );
  INV_X1 U15581 ( .A(n12449), .ZN(n12451) );
  INV_X1 U15582 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U15583 ( .A1(n12451), .A2(n12450), .ZN(n12452) );
  NAND2_X1 U15584 ( .A1(n12460), .A2(n12452), .ZN(n16248) );
  AOI22_X1 U15585 ( .A1(n16248), .A2(n13006), .B1(n13013), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12453) );
  OAI21_X1 U15586 ( .B1(n9821), .B2(n12454), .A(n12453), .ZN(n12455) );
  INV_X1 U15587 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n14123) );
  INV_X1 U15588 ( .A(n12490), .ZN(n12462) );
  INV_X1 U15589 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20093) );
  NAND2_X1 U15590 ( .A1(n12460), .A2(n20093), .ZN(n12461) );
  NAND2_X1 U15591 ( .A1(n12462), .A2(n12461), .ZN(n20089) );
  AOI22_X1 U15592 ( .A1(n20089), .A2(n13006), .B1(n13013), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12463) );
  OAI21_X1 U15593 ( .B1(n9821), .B2(n14123), .A(n12463), .ZN(n12464) );
  AOI21_X1 U15594 ( .B1(n12465), .B2(n12582), .A(n12464), .ZN(n14121) );
  AOI22_X1 U15595 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12983), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U15596 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12819), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U15597 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n12812), .B1(
        n12771), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U15598 ( .A1(n12861), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12466) );
  NAND4_X1 U15599 ( .A1(n12469), .A2(n12468), .A3(n12467), .A4(n12466), .ZN(
        n12475) );
  AOI22_X1 U15600 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9715), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15601 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15602 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15603 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n12659), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12470) );
  NAND4_X1 U15604 ( .A1(n12473), .A2(n12472), .A3(n12471), .A4(n12470), .ZN(
        n12474) );
  OAI21_X1 U15605 ( .B1(n12475), .B2(n12474), .A(n12582), .ZN(n12479) );
  NAND2_X1 U15606 ( .A1(n13014), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12478) );
  XNOR2_X1 U15607 ( .A(n12490), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14676) );
  NAND2_X1 U15608 ( .A1(n14676), .A2(n13006), .ZN(n12477) );
  NAND2_X1 U15609 ( .A1(n13013), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12476) );
  AOI22_X1 U15610 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12992), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15611 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12819), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15612 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15613 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12771), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12480) );
  NAND4_X1 U15614 ( .A1(n12483), .A2(n12482), .A3(n12481), .A4(n12480), .ZN(
        n12489) );
  AOI22_X1 U15615 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15616 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15617 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15618 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12484) );
  NAND4_X1 U15619 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12488) );
  NOR2_X1 U15620 ( .A1(n12489), .A2(n12488), .ZN(n12493) );
  XNOR2_X1 U15621 ( .A(n12513), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16177) );
  NAND2_X1 U15622 ( .A1(n16177), .A2(n13006), .ZN(n12492) );
  AOI22_X1 U15623 ( .A1(n13014), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n13013), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12491) );
  OAI211_X1 U15624 ( .C1(n12493), .C2(n12558), .A(n12492), .B(n12491), .ZN(
        n14129) );
  XOR2_X1 U15625 ( .A(n20083), .B(n12494), .Z(n20081) );
  INV_X1 U15626 ( .A(n20081), .ZN(n12509) );
  AOI22_X1 U15627 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12839), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15628 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12715), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U15629 ( .A1(n12995), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15630 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12495) );
  NAND4_X1 U15631 ( .A1(n12498), .A2(n12497), .A3(n12496), .A4(n12495), .ZN(
        n12504) );
  AOI22_X1 U15632 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15633 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12771), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15634 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15635 ( .A1(n12861), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12499) );
  NAND4_X1 U15636 ( .A1(n12502), .A2(n12501), .A3(n12500), .A4(n12499), .ZN(
        n12503) );
  OAI21_X1 U15637 ( .B1(n12504), .B2(n12503), .A(n12582), .ZN(n12507) );
  NAND2_X1 U15638 ( .A1(n13014), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12506) );
  NAND2_X1 U15639 ( .A1(n13013), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12505) );
  NAND3_X1 U15640 ( .A1(n12507), .A2(n12506), .A3(n12505), .ZN(n12508) );
  AOI21_X1 U15641 ( .B1(n12509), .B2(n13006), .A(n12508), .ZN(n14228) );
  INV_X1 U15642 ( .A(n14228), .ZN(n14127) );
  AND2_X1 U15643 ( .A1(n14129), .A2(n14127), .ZN(n12510) );
  INV_X1 U15644 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12516) );
  OAI21_X1 U15645 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12514), .A(
        n12553), .ZN(n16234) );
  NAND2_X1 U15646 ( .A1(n16234), .A2(n12872), .ZN(n12515) );
  OAI21_X1 U15647 ( .B1(n12516), .B2(n12623), .A(n12515), .ZN(n12517) );
  AOI21_X1 U15648 ( .B1(n13014), .B2(P1_EAX_REG_11__SCAN_IN), .A(n12517), .ZN(
        n14355) );
  AOI22_X1 U15649 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12521) );
  AOI22_X1 U15650 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12715), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12520) );
  AOI22_X1 U15651 ( .A1(n12995), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12771), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U15652 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12518) );
  NAND4_X1 U15653 ( .A1(n12521), .A2(n12520), .A3(n12519), .A4(n12518), .ZN(
        n12527) );
  AOI22_X1 U15654 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U15655 ( .A1(n12861), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U15656 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9714), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U15657 ( .A1(n12812), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12522) );
  NAND4_X1 U15658 ( .A1(n12525), .A2(n12524), .A3(n12523), .A4(n12522), .ZN(
        n12526) );
  OR2_X1 U15659 ( .A1(n12527), .A2(n12526), .ZN(n12528) );
  NAND2_X1 U15660 ( .A1(n12582), .A2(n12528), .ZN(n14423) );
  INV_X1 U15661 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14366) );
  AOI22_X1 U15662 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U15663 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12992), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U15664 ( .A1(n12995), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12812), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15665 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12530) );
  NAND4_X1 U15666 ( .A1(n12533), .A2(n12532), .A3(n12531), .A4(n12530), .ZN(
        n12539) );
  AOI22_X1 U15667 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15668 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U15669 ( .A1(n12987), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12535) );
  AOI22_X1 U15670 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12534) );
  NAND4_X1 U15671 ( .A1(n12537), .A2(n12536), .A3(n12535), .A4(n12534), .ZN(
        n12538) );
  OAI21_X1 U15672 ( .B1(n12539), .B2(n12538), .A(n12582), .ZN(n12542) );
  XNOR2_X1 U15673 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12553), .ZN(
        n16223) );
  OAI22_X1 U15674 ( .A1(n16223), .A2(n12409), .B1(n12623), .B2(n16159), .ZN(
        n12540) );
  INV_X1 U15675 ( .A(n12540), .ZN(n12541) );
  OAI211_X1 U15676 ( .C1(n9821), .C2(n14366), .A(n12542), .B(n12541), .ZN(
        n14359) );
  AOI22_X1 U15677 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12839), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15678 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12715), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U15679 ( .A1(n12861), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U15680 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12543) );
  NAND4_X1 U15681 ( .A1(n12546), .A2(n12545), .A3(n12544), .A4(n12543), .ZN(
        n12552) );
  AOI22_X1 U15682 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15683 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12771), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15684 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15685 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12547) );
  NAND4_X1 U15686 ( .A1(n12550), .A2(n12549), .A3(n12548), .A4(n12547), .ZN(
        n12551) );
  NOR2_X1 U15687 ( .A1(n12552), .A2(n12551), .ZN(n12557) );
  INV_X1 U15688 ( .A(n12559), .ZN(n12554) );
  XNOR2_X1 U15689 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12554), .ZN(
        n14897) );
  AOI22_X1 U15690 ( .A1(n13006), .A2(n14897), .B1(n13013), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12556) );
  NAND2_X1 U15691 ( .A1(n13014), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12555) );
  OAI211_X1 U15692 ( .C1(n12558), .C2(n12557), .A(n12556), .B(n12555), .ZN(
        n14404) );
  XOR2_X1 U15693 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n12573), .Z(
        n16218) );
  AOI22_X1 U15694 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15695 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9715), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U15696 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U15697 ( .A1(n12791), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12560) );
  NAND4_X1 U15698 ( .A1(n12563), .A2(n12562), .A3(n12561), .A4(n12560), .ZN(
        n12569) );
  AOI22_X1 U15699 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12715), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U15700 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U15701 ( .A1(n12714), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15702 ( .A1(n12771), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12564) );
  NAND4_X1 U15703 ( .A1(n12567), .A2(n12566), .A3(n12565), .A4(n12564), .ZN(
        n12568) );
  OR2_X1 U15704 ( .A1(n12569), .A2(n12568), .ZN(n12570) );
  AOI22_X1 U15705 ( .A1(n12582), .A2(n12570), .B1(n13013), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12572) );
  NAND2_X1 U15706 ( .A1(n13014), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12571) );
  OAI211_X1 U15707 ( .C1(n16218), .C2(n12409), .A(n12572), .B(n12571), .ZN(
        n14370) );
  NAND2_X1 U15708 ( .A1(n14367), .A2(n14370), .ZN(n14369) );
  XNOR2_X1 U15709 ( .A(n12605), .B(n12604), .ZN(n14884) );
  AOI22_X1 U15710 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U15711 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U15712 ( .A1(n12985), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U15713 ( .A1(n12771), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12574) );
  NAND4_X1 U15714 ( .A1(n12577), .A2(n12576), .A3(n12575), .A4(n12574), .ZN(
        n12584) );
  AOI22_X1 U15715 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12992), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15716 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15717 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12812), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15718 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12578) );
  NAND4_X1 U15719 ( .A1(n12581), .A2(n12580), .A3(n12579), .A4(n12578), .ZN(
        n12583) );
  OAI21_X1 U15720 ( .B1(n12584), .B2(n12583), .A(n12582), .ZN(n12587) );
  NAND2_X1 U15721 ( .A1(n13014), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U15722 ( .A1(n13013), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12585) );
  NAND3_X1 U15723 ( .A1(n12587), .A2(n12586), .A3(n12585), .ZN(n12588) );
  AOI21_X1 U15724 ( .B1(n14884), .B2(n13006), .A(n12588), .ZN(n14433) );
  AOI22_X1 U15725 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12679), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15726 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12715), .B1(
        n12992), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15727 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12994), .B1(
        n12812), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15728 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n9715), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12590) );
  NAND4_X1 U15729 ( .A1(n12593), .A2(n12592), .A3(n12591), .A4(n12590), .ZN(
        n12599) );
  AOI22_X1 U15730 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15731 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n12856), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15732 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12771), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15733 ( .A1(n12714), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12594) );
  NAND4_X1 U15734 ( .A1(n12597), .A2(n12596), .A3(n12595), .A4(n12594), .ZN(
        n12598) );
  NOR2_X1 U15735 ( .A1(n12599), .A2(n12598), .ZN(n12603) );
  NAND2_X1 U15736 ( .A1(n21011), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12600) );
  NAND2_X1 U15737 ( .A1(n12409), .A2(n12600), .ZN(n12601) );
  AOI21_X1 U15738 ( .B1(n13014), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12601), .ZN(
        n12602) );
  OAI21_X1 U15739 ( .B1(n13009), .B2(n12603), .A(n12602), .ZN(n12608) );
  OAI21_X1 U15740 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12606), .A(
        n12622), .ZN(n16211) );
  OR2_X1 U15741 ( .A1(n12409), .A2(n16211), .ZN(n12607) );
  NAND2_X1 U15742 ( .A1(n12608), .A2(n12607), .ZN(n14473) );
  AOI22_X1 U15743 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12715), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15744 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U15745 ( .A1(n12861), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U15746 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12611) );
  NAND4_X1 U15747 ( .A1(n12614), .A2(n12613), .A3(n12612), .A4(n12611), .ZN(
        n12620) );
  AOI22_X1 U15748 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15749 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15750 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U15751 ( .A1(n12771), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12615) );
  NAND4_X1 U15752 ( .A1(n12618), .A2(n12617), .A3(n12616), .A4(n12615), .ZN(
        n12619) );
  OR2_X1 U15753 ( .A1(n12620), .A2(n12619), .ZN(n12621) );
  NAND2_X1 U15754 ( .A1(n12869), .A2(n12621), .ZN(n12626) );
  AOI21_X1 U15755 ( .B1(n21087), .B2(n12622), .A(n12641), .ZN(n16128) );
  OAI22_X1 U15756 ( .A1(n16128), .A2(n12409), .B1(n21087), .B2(n12623), .ZN(
        n12624) );
  AOI21_X1 U15757 ( .B1(n13014), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12624), .ZN(
        n12625) );
  NAND2_X1 U15758 ( .A1(n12626), .A2(n12625), .ZN(n14496) );
  AOI22_X1 U15759 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15760 ( .A1(n12985), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12714), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15761 ( .A1(n12819), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U15762 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12627) );
  NAND4_X1 U15763 ( .A1(n12630), .A2(n12629), .A3(n12628), .A4(n12627), .ZN(
        n12636) );
  AOI22_X1 U15764 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U15765 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U15766 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U15767 ( .A1(n12771), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12631) );
  NAND4_X1 U15768 ( .A1(n12634), .A2(n12633), .A3(n12632), .A4(n12631), .ZN(
        n12635) );
  NOR2_X1 U15769 ( .A1(n12636), .A2(n12635), .ZN(n12640) );
  INV_X1 U15770 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21012) );
  OAI21_X1 U15771 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21012), .A(
        n21011), .ZN(n12637) );
  INV_X1 U15772 ( .A(n12637), .ZN(n12638) );
  AOI21_X1 U15773 ( .B1(n13014), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12638), .ZN(
        n12639) );
  OAI21_X1 U15774 ( .B1(n13009), .B2(n12640), .A(n12639), .ZN(n12643) );
  OAI21_X1 U15775 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12641), .A(
        n12674), .ZN(n16118) );
  OR2_X1 U15776 ( .A1(n12409), .A2(n16118), .ZN(n12642) );
  AOI22_X1 U15777 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U15778 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12714), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U15779 ( .A1(n12812), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12771), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12645) );
  AOI22_X1 U15780 ( .A1(n12791), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12644) );
  NAND4_X1 U15781 ( .A1(n12647), .A2(n12646), .A3(n12645), .A4(n12644), .ZN(
        n12653) );
  AOI22_X1 U15782 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12985), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U15783 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15784 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U15785 ( .A1(n12819), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12648) );
  NAND4_X1 U15786 ( .A1(n12651), .A2(n12650), .A3(n12649), .A4(n12648), .ZN(
        n12652) );
  NOR2_X1 U15787 ( .A1(n12653), .A2(n12652), .ZN(n12656) );
  INV_X1 U15788 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14855) );
  OAI21_X1 U15789 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14855), .A(n12409), 
        .ZN(n12654) );
  AOI21_X1 U15790 ( .B1(n13014), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12654), .ZN(
        n12655) );
  OAI21_X1 U15791 ( .B1(n13009), .B2(n12656), .A(n12655), .ZN(n12658) );
  XNOR2_X1 U15792 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12674), .ZN(
        n14857) );
  NAND2_X1 U15793 ( .A1(n12872), .A2(n14857), .ZN(n12657) );
  NAND2_X1 U15794 ( .A1(n12658), .A2(n12657), .ZN(n14657) );
  AOI22_X1 U15795 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12715), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15796 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12819), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U15797 ( .A1(n12985), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12714), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U15798 ( .A1(n12771), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12660) );
  NAND4_X1 U15799 ( .A1(n12663), .A2(n12662), .A3(n12661), .A4(n12660), .ZN(
        n12669) );
  AOI22_X1 U15800 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12992), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U15801 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U15802 ( .A1(n12791), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U15803 ( .A1(n12812), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12664) );
  NAND4_X1 U15804 ( .A1(n12667), .A2(n12666), .A3(n12665), .A4(n12664), .ZN(
        n12668) );
  NOR2_X1 U15805 ( .A1(n12669), .A2(n12668), .ZN(n12673) );
  NAND2_X1 U15806 ( .A1(n21011), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12670) );
  NAND2_X1 U15807 ( .A1(n12409), .A2(n12670), .ZN(n12671) );
  AOI21_X1 U15808 ( .B1(n13014), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12671), .ZN(
        n12672) );
  OAI21_X1 U15809 ( .B1(n13009), .B2(n12673), .A(n12672), .ZN(n12677) );
  OAI21_X1 U15810 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12675), .A(
        n12710), .ZN(n16206) );
  OR2_X1 U15811 ( .A1(n12409), .A2(n16206), .ZN(n12676) );
  NAND2_X1 U15812 ( .A1(n12677), .A2(n12676), .ZN(n14713) );
  AOI22_X1 U15813 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U15814 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12715), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U15815 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12771), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U15816 ( .A1(n12714), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12680) );
  NAND4_X1 U15817 ( .A1(n12683), .A2(n12682), .A3(n12681), .A4(n12680), .ZN(
        n12689) );
  AOI22_X1 U15818 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U15819 ( .A1(n12819), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15820 ( .A1(n12812), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U15821 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12684) );
  NAND4_X1 U15822 ( .A1(n12687), .A2(n12686), .A3(n12685), .A4(n12684), .ZN(
        n12688) );
  NOR2_X1 U15823 ( .A1(n12689), .A2(n12688), .ZN(n12692) );
  INV_X1 U15824 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12709) );
  OAI21_X1 U15825 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n12709), .A(n12409), 
        .ZN(n12690) );
  AOI21_X1 U15826 ( .B1(n13014), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12690), .ZN(
        n12691) );
  OAI21_X1 U15827 ( .B1(n13009), .B2(n12692), .A(n12691), .ZN(n12694) );
  XNOR2_X1 U15828 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12710), .ZN(
        n16197) );
  NAND2_X1 U15829 ( .A1(n16197), .A2(n12872), .ZN(n12693) );
  AOI22_X1 U15830 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U15831 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12714), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U15832 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12771), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U15833 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12695) );
  NAND4_X1 U15834 ( .A1(n12698), .A2(n12697), .A3(n12696), .A4(n12695), .ZN(
        n12704) );
  AOI22_X1 U15835 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15836 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15837 ( .A1(n12995), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U15838 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12699) );
  NAND4_X1 U15839 ( .A1(n12702), .A2(n12701), .A3(n12700), .A4(n12699), .ZN(
        n12703) );
  NOR2_X1 U15840 ( .A1(n12704), .A2(n12703), .ZN(n12708) );
  OAI21_X1 U15841 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21012), .A(
        n21011), .ZN(n12705) );
  INV_X1 U15842 ( .A(n12705), .ZN(n12706) );
  AOI21_X1 U15843 ( .B1(n13014), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12706), .ZN(
        n12707) );
  OAI21_X1 U15844 ( .B1(n13009), .B2(n12708), .A(n12707), .ZN(n12713) );
  OAI21_X1 U15845 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12711), .A(
        n12761), .ZN(n16196) );
  OR2_X1 U15846 ( .A1(n12409), .A2(n16196), .ZN(n12712) );
  NAND2_X1 U15847 ( .A1(n14701), .A2(n14756), .ZN(n14692) );
  INV_X1 U15848 ( .A(n14692), .ZN(n12743) );
  AOI22_X1 U15849 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U15850 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12679), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15851 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12714), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15852 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12716) );
  NAND4_X1 U15853 ( .A1(n12719), .A2(n12718), .A3(n12717), .A4(n12716), .ZN(
        n12725) );
  AOI22_X1 U15854 ( .A1(n12819), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12812), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U15855 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15856 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15857 ( .A1(n12771), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12720) );
  NAND4_X1 U15858 ( .A1(n12723), .A2(n12722), .A3(n12721), .A4(n12720), .ZN(
        n12724) );
  NOR2_X1 U15859 ( .A1(n12725), .A2(n12724), .ZN(n12744) );
  AOI22_X1 U15860 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15861 ( .A1(n12985), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15862 ( .A1(n12818), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U15863 ( .A1(n12987), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12727) );
  NAND4_X1 U15864 ( .A1(n12730), .A2(n12729), .A3(n12728), .A4(n12727), .ZN(
        n12736) );
  AOI22_X1 U15865 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12992), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U15866 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U15867 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U15868 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12731) );
  NAND4_X1 U15869 ( .A1(n12734), .A2(n12733), .A3(n12732), .A4(n12731), .ZN(
        n12735) );
  NOR2_X1 U15870 ( .A1(n12736), .A2(n12735), .ZN(n12745) );
  XOR2_X1 U15871 ( .A(n12744), .B(n12745), .Z(n12737) );
  NAND2_X1 U15872 ( .A1(n12869), .A2(n12737), .ZN(n12740) );
  INV_X1 U15873 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16092) );
  OAI21_X1 U15874 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n16092), .A(n12409), 
        .ZN(n12738) );
  AOI21_X1 U15875 ( .B1(n13014), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12738), .ZN(
        n12739) );
  NAND2_X1 U15876 ( .A1(n12740), .A2(n12739), .ZN(n12742) );
  XNOR2_X1 U15877 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12761), .ZN(
        n16082) );
  NAND2_X1 U15878 ( .A1(n12872), .A2(n16082), .ZN(n12741) );
  NAND2_X1 U15879 ( .A1(n12743), .A2(n9828), .ZN(n14641) );
  NOR2_X1 U15880 ( .A1(n12745), .A2(n12744), .ZN(n12766) );
  AOI22_X1 U15881 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15882 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12679), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U15883 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U15884 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12813), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12747) );
  NAND4_X1 U15885 ( .A1(n12750), .A2(n12749), .A3(n12748), .A4(n12747), .ZN(
        n12756) );
  AOI22_X1 U15886 ( .A1(n12819), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15887 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U15888 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U15889 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12751) );
  NAND4_X1 U15890 ( .A1(n12754), .A2(n12753), .A3(n12752), .A4(n12751), .ZN(
        n12755) );
  OR2_X1 U15891 ( .A1(n12756), .A2(n12755), .ZN(n12765) );
  INV_X1 U15892 ( .A(n12765), .ZN(n12757) );
  XNOR2_X1 U15893 ( .A(n12766), .B(n12757), .ZN(n12760) );
  INV_X1 U15894 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14747) );
  NAND2_X1 U15895 ( .A1(n21011), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12758) );
  OAI211_X1 U15896 ( .C1(n9821), .C2(n14747), .A(n12409), .B(n12758), .ZN(
        n12759) );
  AOI21_X1 U15897 ( .B1(n12760), .B2(n12869), .A(n12759), .ZN(n12764) );
  OAI21_X1 U15898 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12762), .A(
        n12802), .ZN(n14836) );
  NOR2_X1 U15899 ( .A1(n14836), .A2(n12409), .ZN(n12763) );
  NAND2_X1 U15900 ( .A1(n12766), .A2(n12765), .ZN(n12785) );
  AOI22_X1 U15901 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U15902 ( .A1(n12819), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U15903 ( .A1(n12812), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U15904 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12767) );
  NAND4_X1 U15905 ( .A1(n12770), .A2(n12769), .A3(n12768), .A4(n12767), .ZN(
        n12777) );
  AOI22_X1 U15906 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U15907 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U15908 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12771), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U15909 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12772) );
  NAND4_X1 U15910 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n12776) );
  NOR2_X1 U15911 ( .A1(n12777), .A2(n12776), .ZN(n12786) );
  XOR2_X1 U15912 ( .A(n12785), .B(n12786), .Z(n12778) );
  NAND2_X1 U15913 ( .A1(n12778), .A2(n12869), .ZN(n12781) );
  INV_X1 U15914 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14826) );
  AOI21_X1 U15915 ( .B1(n14826), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12779) );
  AOI21_X1 U15916 ( .B1(n13014), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12779), .ZN(
        n12780) );
  NAND2_X1 U15917 ( .A1(n12781), .A2(n12780), .ZN(n12783) );
  XNOR2_X1 U15918 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n12802), .ZN(
        n14828) );
  NAND2_X1 U15919 ( .A1(n12872), .A2(n14828), .ZN(n12782) );
  NAND2_X1 U15920 ( .A1(n12783), .A2(n12782), .ZN(n14633) );
  NOR2_X1 U15921 ( .A1(n12786), .A2(n12785), .ZN(n12811) );
  AOI22_X1 U15922 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U15923 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12679), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12789) );
  INV_X1 U15924 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n21127) );
  AOI22_X1 U15925 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12714), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U15926 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12787) );
  NAND4_X1 U15927 ( .A1(n12790), .A2(n12789), .A3(n12788), .A4(n12787), .ZN(
        n12797) );
  AOI22_X1 U15928 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U15929 ( .A1(n12985), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12794) );
  AOI22_X1 U15930 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U15931 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12792) );
  NAND4_X1 U15932 ( .A1(n12795), .A2(n12794), .A3(n12793), .A4(n12792), .ZN(
        n12796) );
  OR2_X1 U15933 ( .A1(n12797), .A2(n12796), .ZN(n12810) );
  INV_X1 U15934 ( .A(n12810), .ZN(n12798) );
  XNOR2_X1 U15935 ( .A(n12811), .B(n12798), .ZN(n12799) );
  NAND2_X1 U15936 ( .A1(n12799), .A2(n12869), .ZN(n12809) );
  NAND2_X1 U15937 ( .A1(n21011), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12800) );
  NAND2_X1 U15938 ( .A1(n12409), .A2(n12800), .ZN(n12801) );
  AOI21_X1 U15939 ( .B1(n13014), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12801), .ZN(
        n12808) );
  INV_X1 U15940 ( .A(n12802), .ZN(n12803) );
  INV_X1 U15941 ( .A(n12804), .ZN(n12805) );
  INV_X1 U15942 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14621) );
  NAND2_X1 U15943 ( .A1(n12805), .A2(n14621), .ZN(n12806) );
  NAND2_X1 U15944 ( .A1(n12832), .A2(n12806), .ZN(n14817) );
  NOR2_X1 U15945 ( .A1(n14817), .A2(n12409), .ZN(n12807) );
  AOI21_X1 U15946 ( .B1(n12809), .B2(n12808), .A(n12807), .ZN(n14620) );
  NAND2_X1 U15947 ( .A1(n12811), .A2(n12810), .ZN(n12836) );
  AOI22_X1 U15948 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12985), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U15949 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12816) );
  AOI22_X1 U15950 ( .A1(n12812), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U15951 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12814) );
  NAND4_X1 U15952 ( .A1(n12817), .A2(n12816), .A3(n12815), .A4(n12814), .ZN(
        n12825) );
  AOI22_X1 U15953 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U15954 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12992), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12822) );
  AOI22_X1 U15955 ( .A1(n12819), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U15956 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12820) );
  NAND4_X1 U15957 ( .A1(n12823), .A2(n12822), .A3(n12821), .A4(n12820), .ZN(
        n12824) );
  NOR2_X1 U15958 ( .A1(n12825), .A2(n12824), .ZN(n12837) );
  XOR2_X1 U15959 ( .A(n12836), .B(n12837), .Z(n12826) );
  NAND2_X1 U15960 ( .A1(n12826), .A2(n12869), .ZN(n12831) );
  NAND2_X1 U15961 ( .A1(n21011), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12827) );
  NAND2_X1 U15962 ( .A1(n12409), .A2(n12827), .ZN(n12828) );
  AOI21_X1 U15963 ( .B1(n13014), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12828), .ZN(
        n12830) );
  XNOR2_X1 U15964 ( .A(n12832), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14814) );
  AOI21_X1 U15965 ( .B1(n12831), .B2(n12830), .A(n12829), .ZN(n14608) );
  INV_X1 U15966 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14810) );
  NAND2_X1 U15967 ( .A1(n12833), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12981) );
  INV_X1 U15968 ( .A(n12833), .ZN(n12834) );
  INV_X1 U15969 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n21091) );
  NAND2_X1 U15970 ( .A1(n12834), .A2(n21091), .ZN(n12835) );
  NAND2_X1 U15971 ( .A1(n12981), .A2(n12835), .ZN(n14803) );
  NOR2_X1 U15972 ( .A1(n12837), .A2(n12836), .ZN(n12855) );
  AOI22_X1 U15973 ( .A1(n12838), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12843) );
  AOI22_X1 U15974 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12839), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U15975 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U15976 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12840) );
  NAND4_X1 U15977 ( .A1(n12843), .A2(n12842), .A3(n12841), .A4(n12840), .ZN(
        n12849) );
  INV_X1 U15978 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n21221) );
  AOI22_X1 U15979 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U15980 ( .A1(n12985), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U15981 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U15982 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12844) );
  NAND4_X1 U15983 ( .A1(n12847), .A2(n12846), .A3(n12845), .A4(n12844), .ZN(
        n12848) );
  OR2_X1 U15984 ( .A1(n12849), .A2(n12848), .ZN(n12854) );
  XNOR2_X1 U15985 ( .A(n12855), .B(n12854), .ZN(n12852) );
  NOR2_X1 U15986 ( .A1(n21091), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12850) );
  AOI211_X1 U15987 ( .C1(n13014), .C2(P1_EAX_REG_28__SCAN_IN), .A(n13006), .B(
        n12850), .ZN(n12851) );
  OAI21_X1 U15988 ( .B1(n12852), .B2(n13009), .A(n12851), .ZN(n12853) );
  OAI21_X1 U15989 ( .B1(n12409), .B2(n14803), .A(n12853), .ZN(n14594) );
  NAND2_X1 U15990 ( .A1(n12855), .A2(n12854), .ZN(n13002) );
  AOI22_X1 U15991 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12860) );
  AOI22_X1 U15992 ( .A1(n12715), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12859) );
  AOI22_X1 U15993 ( .A1(n12856), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9714), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U15994 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12857) );
  NAND4_X1 U15995 ( .A1(n12860), .A2(n12859), .A3(n12858), .A4(n12857), .ZN(
        n12868) );
  AOI22_X1 U15996 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U15997 ( .A1(n12985), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12714), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12865) );
  AOI22_X1 U15998 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U15999 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12863) );
  NAND4_X1 U16000 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n12863), .ZN(
        n12867) );
  NOR2_X1 U16001 ( .A1(n12868), .A2(n12867), .ZN(n13003) );
  XOR2_X1 U16002 ( .A(n13002), .B(n13003), .Z(n12870) );
  NAND2_X1 U16003 ( .A1(n12870), .A2(n12869), .ZN(n12874) );
  INV_X1 U16004 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12884) );
  NOR2_X1 U16005 ( .A1(n12884), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12871) );
  AOI211_X1 U16006 ( .C1(n13014), .C2(P1_EAX_REG_29__SCAN_IN), .A(n13006), .B(
        n12871), .ZN(n12873) );
  XNOR2_X1 U16007 ( .A(n12981), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14550) );
  AOI22_X1 U16008 ( .A1(n12874), .A2(n12873), .B1(n12872), .B2(n14550), .ZN(
        n12876) );
  NAND2_X1 U16009 ( .A1(n13012), .A2(n12877), .ZN(n14535) );
  NAND3_X1 U16010 ( .A1(n11887), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16377) );
  INV_X1 U16011 ( .A(n16377), .ZN(n12878) );
  AND2_X1 U16012 ( .A1(n12878), .A2(n20689), .ZN(n13942) );
  NOR2_X1 U16013 ( .A1(n12879), .A2(n12147), .ZN(n12880) );
  INV_X1 U16014 ( .A(n20689), .ZN(n20760) );
  NAND2_X1 U16015 ( .A1(n20760), .A2(n12881), .ZN(n21017) );
  AND2_X1 U16016 ( .A1(n21017), .A2(n11887), .ZN(n12882) );
  NAND2_X1 U16017 ( .A1(n11887), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16048) );
  NAND2_X1 U16018 ( .A1(n21012), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12883) );
  NAND2_X1 U16019 ( .A1(n16048), .A2(n12883), .ZN(n20227) );
  INV_X1 U16020 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14546) );
  OAI22_X1 U16021 ( .A1(n16256), .A2(n12884), .B1(n20100), .B2(n14546), .ZN(
        n12885) );
  AOI21_X1 U16022 ( .B1(n16252), .B2(n14550), .A(n12885), .ZN(n12886) );
  INV_X1 U16023 ( .A(n12886), .ZN(n12887) );
  NAND2_X1 U16024 ( .A1(n10106), .A2(n12888), .ZN(P1_U2970) );
  NAND2_X1 U16025 ( .A1(n11053), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U16026 ( .A1(n12889), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12890) );
  AND2_X1 U16027 ( .A1(n12891), .A2(n12890), .ZN(n12892) );
  INV_X1 U16028 ( .A(n12894), .ZN(n12895) );
  OAI21_X1 U16029 ( .B1(n14528), .B2(n16474), .A(n12895), .ZN(n12896) );
  INV_X1 U16030 ( .A(n12896), .ZN(n12910) );
  NOR2_X1 U16031 ( .A1(n15589), .A2(n12897), .ZN(n12898) );
  NAND2_X1 U16032 ( .A1(n12899), .A2(n12898), .ZN(n15575) );
  NAND2_X1 U16033 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12903) );
  INV_X1 U16034 ( .A(n15543), .ZN(n12900) );
  NAND3_X1 U16035 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15522) );
  INV_X1 U16036 ( .A(n15522), .ZN(n12905) );
  NAND4_X1 U16037 ( .A1(n12900), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n11254), .A4(n12905), .ZN(n12909) );
  OAI21_X1 U16038 ( .B1(n16482), .B2(n12901), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12902) );
  OR2_X1 U16039 ( .A1(n15792), .A2(n12902), .ZN(n15590) );
  NAND2_X1 U16040 ( .A1(n15590), .A2(n15708), .ZN(n15576) );
  NAND2_X1 U16041 ( .A1(n15708), .A2(n12903), .ZN(n12904) );
  NAND2_X1 U16042 ( .A1(n15576), .A2(n12904), .ZN(n15561) );
  NOR2_X1 U16043 ( .A1(n16482), .A2(n12905), .ZN(n12906) );
  NOR2_X1 U16044 ( .A1(n15561), .A2(n12906), .ZN(n15520) );
  OAI21_X1 U16045 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16482), .A(
        n15520), .ZN(n12907) );
  NAND2_X1 U16046 ( .A1(n12907), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12908) );
  OAI211_X1 U16047 ( .C1(n12915), .C2(n16476), .A(n12914), .B(n12913), .ZN(
        P2_U3015) );
  AND2_X1 U16048 ( .A1(n12952), .A2(n15322), .ZN(n12918) );
  NOR2_X1 U16049 ( .A1(n12917), .A2(n12918), .ZN(n15324) );
  OAI21_X1 U16050 ( .B1(n12919), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n9781), .ZN(n15365) );
  INV_X1 U16051 ( .A(n15365), .ZN(n16403) );
  OAI21_X1 U16052 ( .B1(n9817), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n12920), .ZN(n15404) );
  INV_X1 U16053 ( .A(n15404), .ZN(n15172) );
  OR2_X1 U16054 ( .A1(n12922), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12923) );
  NAND2_X1 U16055 ( .A1(n12921), .A2(n12923), .ZN(n15427) );
  INV_X1 U16056 ( .A(n15427), .ZN(n19096) );
  OAI21_X1 U16057 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12924), .A(
        n12925), .ZN(n12926) );
  INV_X1 U16058 ( .A(n12926), .ZN(n19120) );
  OAI21_X1 U16059 ( .B1(n12948), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n12949), .ZN(n15459) );
  INV_X1 U16060 ( .A(n15459), .ZN(n19142) );
  INV_X1 U16061 ( .A(n12927), .ZN(n12928) );
  OAI21_X1 U16062 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12943), .A(
        n12928), .ZN(n19163) );
  INV_X1 U16063 ( .A(n19163), .ZN(n12946) );
  NOR2_X1 U16064 ( .A1(n19209), .A2(n12929), .ZN(n12940) );
  OAI21_X1 U16065 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12940), .A(
        n12944), .ZN(n19186) );
  INV_X1 U16066 ( .A(n19186), .ZN(n12942) );
  OAI21_X1 U16067 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12930), .A(
        n12929), .ZN(n16454) );
  INV_X1 U16068 ( .A(n16454), .ZN(n12939) );
  AOI21_X1 U16069 ( .B1(n19235), .B2(n12936), .A(n12931), .ZN(n19228) );
  NOR2_X1 U16070 ( .A1(n19408), .A2(n12932), .ZN(n12937) );
  AOI21_X1 U16071 ( .B1(n19408), .B2(n12932), .A(n12937), .ZN(n19397) );
  AOI21_X1 U16072 ( .B1(n12933), .B2(n12934), .A(n12935), .ZN(n14151) );
  INV_X1 U16073 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U16074 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n12955), .ZN(n14313) );
  AOI22_X1 U16075 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n12933), .B2(n12955), .ZN(
        n14312) );
  NAND2_X1 U16076 ( .A1(n14313), .A2(n14312), .ZN(n14311) );
  NOR2_X1 U16077 ( .A1(n14151), .A2(n14311), .ZN(n14138) );
  OAI21_X1 U16078 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12935), .A(
        n12932), .ZN(n14175) );
  NAND2_X1 U16079 ( .A1(n14138), .A2(n14175), .ZN(n14192) );
  NOR2_X1 U16080 ( .A1(n19397), .A2(n14192), .ZN(n19241) );
  OAI21_X1 U16081 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12937), .A(
        n12936), .ZN(n19243) );
  NAND2_X1 U16082 ( .A1(n19241), .A2(n19243), .ZN(n19225) );
  NOR2_X1 U16083 ( .A1(n19228), .A2(n19225), .ZN(n19210) );
  INV_X1 U16084 ( .A(n12930), .ZN(n12938) );
  OAI21_X1 U16085 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12931), .A(
        n12938), .ZN(n19212) );
  NAND2_X1 U16086 ( .A1(n19210), .A2(n19212), .ZN(n14265) );
  NOR2_X1 U16087 ( .A1(n12939), .A2(n14265), .ZN(n19201) );
  AOI21_X1 U16088 ( .B1(n19209), .B2(n12929), .A(n12940), .ZN(n19203) );
  INV_X1 U16089 ( .A(n19203), .ZN(n12941) );
  NAND2_X1 U16090 ( .A1(n19201), .A2(n12941), .ZN(n19185) );
  NOR2_X1 U16091 ( .A1(n12942), .A2(n19185), .ZN(n19176) );
  AOI21_X1 U16092 ( .B1(n12944), .B2(n19184), .A(n12943), .ZN(n19178) );
  INV_X1 U16093 ( .A(n19178), .ZN(n12945) );
  NAND2_X1 U16094 ( .A1(n19176), .A2(n12945), .ZN(n19162) );
  NOR2_X1 U16095 ( .A1(n12946), .A2(n19162), .ZN(n19153) );
  NOR2_X1 U16096 ( .A1(n12927), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12947) );
  OR2_X1 U16097 ( .A1(n12948), .A2(n12947), .ZN(n15468) );
  NAND2_X1 U16098 ( .A1(n19153), .A2(n15468), .ZN(n19140) );
  NOR2_X1 U16099 ( .A1(n19142), .A2(n19140), .ZN(n19129) );
  AOI21_X1 U16100 ( .B1(n21179), .B2(n12949), .A(n12924), .ZN(n16422) );
  INV_X1 U16101 ( .A(n16422), .ZN(n19131) );
  NAND2_X1 U16102 ( .A1(n19129), .A2(n19131), .ZN(n19118) );
  NOR2_X1 U16103 ( .A1(n19120), .A2(n19118), .ZN(n19107) );
  AOI21_X1 U16104 ( .B1(n12925), .B2(n21218), .A(n12922), .ZN(n15438) );
  INV_X1 U16105 ( .A(n15438), .ZN(n19109) );
  NAND2_X1 U16106 ( .A1(n19107), .A2(n19109), .ZN(n19094) );
  NOR2_X1 U16107 ( .A1(n19096), .A2(n19094), .ZN(n19081) );
  AOI21_X1 U16108 ( .B1(n15413), .B2(n12921), .A(n9817), .ZN(n15416) );
  INV_X1 U16109 ( .A(n15416), .ZN(n19083) );
  NAND2_X1 U16110 ( .A1(n19081), .A2(n19083), .ZN(n15171) );
  NOR2_X1 U16111 ( .A1(n15172), .A2(n15171), .ZN(n15170) );
  AOI21_X1 U16112 ( .B1(n12920), .B2(n15396), .A(n12347), .ZN(n15394) );
  AND2_X1 U16113 ( .A1(n12348), .A2(n15371), .ZN(n12950) );
  NOR2_X1 U16114 ( .A1(n12919), .A2(n12950), .ZN(n15374) );
  NOR2_X1 U16115 ( .A1(n15133), .A2(n15374), .ZN(n15132) );
  NOR2_X1 U16116 ( .A1(n19242), .A2(n15132), .ZN(n16402) );
  AOI21_X1 U16117 ( .B1(n15343), .B2(n9781), .A(n12951), .ZN(n15346) );
  OAI21_X1 U16118 ( .B1(n12951), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n12952), .ZN(n15334) );
  INV_X1 U16119 ( .A(n15334), .ZN(n16387) );
  NOR2_X1 U16120 ( .A1(n16386), .A2(n16387), .ZN(n16385) );
  NOR2_X1 U16121 ( .A1(n15324), .A2(n13443), .ZN(n13442) );
  NOR2_X1 U16122 ( .A1(n19242), .A2(n13442), .ZN(n15094) );
  OAI21_X1 U16123 ( .B1(n12917), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n12953), .ZN(n12954) );
  INV_X1 U16124 ( .A(n12954), .ZN(n15316) );
  NOR2_X1 U16125 ( .A1(n15094), .A2(n15316), .ZN(n15095) );
  NOR2_X1 U16126 ( .A1(n19242), .A2(n15095), .ZN(n15086) );
  AOI21_X1 U16127 ( .B1(n15296), .B2(n12953), .A(n9831), .ZN(n15299) );
  NOR2_X1 U16128 ( .A1(n15086), .A2(n15299), .ZN(n15087) );
  NOR2_X1 U16129 ( .A1(n19242), .A2(n15087), .ZN(n12957) );
  AND4_X1 U16130 ( .A1(n12955), .A2(n19763), .A3(n19691), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19246) );
  OR3_X1 U16131 ( .A1(n10954), .A2(n13464), .A3(n16502), .ZN(n14201) );
  AND2_X1 U16132 ( .A1(n9736), .A2(n19927), .ZN(n12958) );
  NAND2_X1 U16133 ( .A1(n13467), .A2(n12958), .ZN(n13463) );
  NAND2_X1 U16134 ( .A1(n14201), .A2(n13463), .ZN(n19057) );
  NAND2_X1 U16135 ( .A1(n19691), .A2(n19922), .ZN(n12967) );
  INV_X1 U16136 ( .A(n12967), .ZN(n12959) );
  AND2_X1 U16137 ( .A1(n10263), .A2(n12959), .ZN(n12960) );
  NAND2_X1 U16138 ( .A1(n19691), .A2(n13458), .ZN(n12965) );
  NOR2_X1 U16139 ( .A1(n12961), .A2(n12965), .ZN(n16517) );
  NAND2_X1 U16140 ( .A1(n15516), .A2(n19266), .ZN(n12978) );
  AND3_X1 U16141 ( .A1(n10263), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n12967), .ZN(
        n12962) );
  NAND2_X1 U16142 ( .A1(n19057), .A2(n12962), .ZN(n19270) );
  NAND2_X1 U16143 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19763), .ZN(n19923) );
  NOR3_X1 U16144 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n20033), .A3(n19923), 
        .ZN(n16514) );
  NAND2_X1 U16145 ( .A1(n19214), .A2(n19928), .ZN(n12963) );
  OR2_X1 U16146 ( .A1(n16514), .A2(n12963), .ZN(n12964) );
  INV_X1 U16147 ( .A(n12965), .ZN(n12970) );
  INV_X1 U16148 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12966) );
  NAND2_X1 U16149 ( .A1(n12967), .A2(n12966), .ZN(n12968) );
  AND2_X1 U16150 ( .A1(n11284), .A2(n12968), .ZN(n12969) );
  NAND2_X1 U16151 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19279), .ZN(
        n12971) );
  OAI21_X1 U16152 ( .B1(n19252), .B2(n12972), .A(n12971), .ZN(n12973) );
  AOI21_X1 U16153 ( .B1(n19265), .B2(P2_REIP_REG_30__SCAN_IN), .A(n12973), 
        .ZN(n12974) );
  OAI21_X1 U16154 ( .B1(n12975), .B2(n19270), .A(n12974), .ZN(n12976) );
  INV_X1 U16155 ( .A(n12976), .ZN(n12977) );
  INV_X1 U16156 ( .A(n12981), .ZN(n12982) );
  XNOR2_X1 U16157 ( .A(n14018), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14792) );
  AOI22_X1 U16158 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12838), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16159 ( .A1(n9715), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U16160 ( .A1(n12861), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12986), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12989) );
  AOI22_X1 U16161 ( .A1(n12987), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12659), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12988) );
  NAND4_X1 U16162 ( .A1(n12991), .A2(n12990), .A3(n12989), .A4(n12988), .ZN(
        n13001) );
  AOI22_X1 U16163 ( .A1(n12992), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12715), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U16164 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U16165 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12791), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U16166 ( .A1(n12995), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12996) );
  NAND4_X1 U16167 ( .A1(n12999), .A2(n12998), .A3(n12997), .A4(n12996), .ZN(
        n13000) );
  NOR2_X1 U16168 ( .A1(n13001), .A2(n13000), .ZN(n13005) );
  NOR2_X1 U16169 ( .A1(n13003), .A2(n13002), .ZN(n13004) );
  XOR2_X1 U16170 ( .A(n13005), .B(n13004), .Z(n13010) );
  AOI21_X1 U16171 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21011), .A(
        n13006), .ZN(n13008) );
  NAND2_X1 U16172 ( .A1(n13014), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n13007) );
  OAI211_X1 U16173 ( .C1(n13010), .C2(n13009), .A(n13008), .B(n13007), .ZN(
        n13011) );
  OAI21_X1 U16174 ( .B1(n12409), .B2(n14792), .A(n13011), .ZN(n13044) );
  AOI22_X1 U16175 ( .A1(n13014), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13013), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13015) );
  INV_X1 U16176 ( .A(n20286), .ZN(n13057) );
  INV_X1 U16177 ( .A(n12204), .ZN(n13778) );
  NAND3_X1 U16178 ( .A1(n13778), .A2(n13558), .A3(n21018), .ZN(n13767) );
  NAND2_X1 U16179 ( .A1(n13016), .A2(n14023), .ZN(n13769) );
  INV_X1 U16180 ( .A(n13768), .ZN(n13017) );
  NAND3_X1 U16181 ( .A1(n13017), .A2(n13683), .A3(n21018), .ZN(n13018) );
  NAND2_X1 U16182 ( .A1(n13769), .A2(n13018), .ZN(n13772) );
  NAND2_X1 U16183 ( .A1(n13772), .A2(n14565), .ZN(n13022) );
  AND4_X1 U16184 ( .A1(n12143), .A2(n13057), .A3(n13019), .A4(n11837), .ZN(
        n13020) );
  AND2_X1 U16185 ( .A1(n13020), .A2(n13863), .ZN(n13045) );
  NAND2_X1 U16186 ( .A1(n13045), .A2(n14023), .ZN(n13021) );
  NAND3_X1 U16187 ( .A1(n13767), .A2(n13022), .A3(n13021), .ZN(n13023) );
  INV_X2 U16188 ( .A(n14767), .ZN(n14748) );
  NAND3_X1 U16189 ( .A1(n14576), .A2(n13057), .A3(n14748), .ZN(n13042) );
  NAND2_X1 U16190 ( .A1(n14748), .A2(n13024), .ZN(n13037) );
  NOR4_X1 U16191 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n13028) );
  NOR4_X1 U16192 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(
        P1_ADDRESS_REG_20__SCAN_IN), .A3(P1_ADDRESS_REG_19__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13027) );
  NOR4_X1 U16193 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13026) );
  NOR4_X1 U16194 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n13025) );
  AND4_X1 U16195 ( .A1(n13028), .A2(n13027), .A3(n13026), .A4(n13025), .ZN(
        n13033) );
  NOR4_X1 U16196 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_6__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n13031) );
  NOR4_X1 U16197 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_22__SCAN_IN), .ZN(n13030) );
  NOR4_X1 U16198 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_3__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13029) );
  INV_X1 U16199 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20943) );
  AND4_X1 U16200 ( .A1(n13031), .A2(n13030), .A3(n13029), .A4(n20943), .ZN(
        n13032) );
  NAND2_X1 U16201 ( .A1(n13033), .A2(n13032), .ZN(n13034) );
  AOI22_X1 U16202 ( .A1(n13035), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14767), .ZN(n13036) );
  INV_X1 U16203 ( .A(n13036), .ZN(n13040) );
  INV_X1 U16204 ( .A(n13037), .ZN(n13038) );
  NAND2_X1 U16205 ( .A1(n13038), .A2(n20239), .ZN(n14771) );
  INV_X1 U16206 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16581) );
  NOR2_X1 U16207 ( .A1(n13040), .A2(n13039), .ZN(n13041) );
  NAND2_X1 U16208 ( .A1(n13042), .A2(n13041), .ZN(P1_U2873) );
  INV_X1 U16209 ( .A(n14794), .ZN(n14732) );
  NAND2_X1 U16210 ( .A1(n14562), .A2(n14569), .ZN(n13765) );
  NAND2_X1 U16211 ( .A1(n13045), .A2(n13683), .ZN(n13046) );
  NAND2_X1 U16212 ( .A1(n13765), .A2(n13046), .ZN(n13047) );
  NAND2_X1 U16213 ( .A1(n13049), .A2(n13048), .ZN(n13053) );
  INV_X1 U16214 ( .A(n13050), .ZN(n13051) );
  NAND2_X1 U16215 ( .A1(n14597), .A2(n13051), .ZN(n13052) );
  NAND2_X1 U16216 ( .A1(n13053), .A2(n13052), .ZN(n13056) );
  INV_X1 U16217 ( .A(n13054), .ZN(n13055) );
  INV_X1 U16218 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13058) );
  INV_X1 U16219 ( .A(n13059), .ZN(n13060) );
  NAND2_X1 U16220 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13061) );
  INV_X2 U16221 ( .A(n9785), .ZN(n17376) );
  AOI22_X1 U16222 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13078) );
  AOI22_X1 U16223 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9720), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13077) );
  OR2_X2 U16224 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n16008), .ZN(
        n17317) );
  INV_X2 U16225 ( .A(n17317), .ZN(n17375) );
  NAND4_X2 U16226 ( .A1(n13063), .A2(n18986), .A3(n13208), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U16227 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13076) );
  NOR3_X1 U16228 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n19014), .ZN(n13062) );
  INV_X1 U16229 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17106) );
  OAI22_X1 U16230 ( .A1(n17373), .A2(n21122), .B1(n17298), .B2(n17106), .ZN(
        n13074) );
  NAND2_X1 U16231 ( .A1(n13065), .A2(n17044), .ZN(n13250) );
  AOI22_X1 U16232 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13072) );
  NAND2_X1 U16233 ( .A1(n17044), .A2(n13067), .ZN(n17205) );
  AOI22_X1 U16234 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16235 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13070) );
  NAND2_X1 U16236 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n13069) );
  NAND4_X1 U16237 ( .A1(n13072), .A2(n13071), .A3(n13070), .A4(n13069), .ZN(
        n13073) );
  AOI211_X1 U16238 ( .C1(n17368), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n13074), .B(n13073), .ZN(n13075) );
  INV_X1 U16239 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U16240 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13088) );
  INV_X1 U16241 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U16242 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U16243 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13079) );
  OAI211_X1 U16244 ( .C1(n17298), .C2(n17286), .A(n13080), .B(n13079), .ZN(
        n13086) );
  AOI22_X1 U16245 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U16246 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U16247 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13082) );
  NAND2_X1 U16248 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13081) );
  NAND4_X1 U16249 ( .A1(n13084), .A2(n13083), .A3(n13082), .A4(n13081), .ZN(
        n13085) );
  AOI211_X1 U16250 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n13086), .B(n13085), .ZN(n13087) );
  OAI211_X1 U16251 ( .C1(n17371), .C2(n17277), .A(n13088), .B(n13087), .ZN(
        n13365) );
  INV_X1 U16252 ( .A(n13365), .ZN(n17556) );
  AOI22_X1 U16253 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13100) );
  INV_X1 U16254 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15922) );
  AOI22_X1 U16255 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16256 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13091) );
  OAI211_X1 U16257 ( .C1(n17298), .C2(n15922), .A(n13092), .B(n13091), .ZN(
        n13098) );
  AOI22_X1 U16258 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9720), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U16259 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16260 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13094) );
  NAND2_X1 U16261 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13093) );
  NAND4_X1 U16262 ( .A1(n13096), .A2(n13095), .A3(n13094), .A4(n13093), .ZN(
        n13097) );
  AOI211_X1 U16263 ( .C1(n13113), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n13098), .B(n13097), .ZN(n13099) );
  INV_X1 U16264 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U16265 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9720), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17332), .ZN(n13102) );
  AOI22_X1 U16266 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17376), .ZN(n13101) );
  OAI211_X1 U16267 ( .C1(n17298), .C2(n17353), .A(n13102), .B(n13101), .ZN(
        n13103) );
  INV_X1 U16268 ( .A(n13103), .ZN(n13109) );
  NAND2_X1 U16269 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13108) );
  AOI22_X1 U16270 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n9767), .ZN(n13107) );
  AOI22_X1 U16271 ( .A1(n13140), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U16272 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n9716), .ZN(n13105) );
  AOI22_X1 U16273 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17199), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13111) );
  INV_X1 U16274 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18421) );
  INV_X1 U16275 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17346) );
  OAI22_X1 U16276 ( .A1(n17210), .A2(n21323), .B1(n17298), .B2(n17346), .ZN(
        n13112) );
  INV_X1 U16277 ( .A(n13112), .ZN(n13120) );
  AOI22_X1 U16278 ( .A1(n13140), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16279 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16280 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9767), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U16281 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13114) );
  NAND4_X1 U16282 ( .A1(n13120), .A2(n13119), .A3(n10104), .A4(n13118), .ZN(
        n13124) );
  INV_X1 U16283 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15958) );
  AOI22_X1 U16284 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13121) );
  OAI21_X1 U16285 ( .B1(n9785), .B2(n15958), .A(n13121), .ZN(n13123) );
  INV_X1 U16286 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U16287 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13132) );
  INV_X1 U16288 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15967) );
  AOI22_X1 U16289 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13126) );
  OAI21_X1 U16290 ( .B1(n13089), .B2(n15967), .A(n13126), .ZN(n13130) );
  INV_X1 U16291 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17306) );
  AOI22_X1 U16292 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16293 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9720), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13127) );
  OAI211_X1 U16294 ( .C1(n17298), .C2(n17306), .A(n13128), .B(n13127), .ZN(
        n13129) );
  AOI211_X1 U16295 ( .C1(n13113), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n13130), .B(n13129), .ZN(n13131) );
  OAI211_X1 U16296 ( .C1(n17371), .C2(n17301), .A(n13132), .B(n13131), .ZN(
        n13136) );
  AOI22_X1 U16297 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13133) );
  OAI21_X1 U16298 ( .B1(n17373), .B2(n17407), .A(n13133), .ZN(n13135) );
  INV_X1 U16299 ( .A(n9718), .ZN(n13137) );
  NAND2_X1 U16300 ( .A1(n13170), .A2(n13137), .ZN(n13173) );
  AOI22_X1 U16301 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17377), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13138) );
  INV_X1 U16302 ( .A(n13138), .ZN(n13150) );
  INV_X1 U16303 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U16304 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13147) );
  INV_X1 U16305 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U16306 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13139) );
  OAI21_X1 U16307 ( .B1(n17373), .B2(n17400), .A(n13139), .ZN(n13145) );
  AOI22_X1 U16308 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17314), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13143) );
  AOI22_X1 U16309 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13142) );
  AOI22_X1 U16310 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13141) );
  NAND3_X1 U16311 ( .A1(n13143), .A2(n13142), .A3(n13141), .ZN(n13144) );
  AOI211_X1 U16312 ( .C1(n17199), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n13145), .B(n13144), .ZN(n13146) );
  OAI211_X1 U16313 ( .C1(n13148), .C2(n17146), .A(n13147), .B(n13146), .ZN(
        n13149) );
  NOR2_X1 U16314 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17958), .ZN(
        n13151) );
  AOI21_X1 U16315 ( .B1(n17958), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n13151), .ZN(n13207) );
  NAND2_X1 U16316 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17796) );
  INV_X1 U16317 ( .A(n17796), .ZN(n18137) );
  NAND3_X1 U16318 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n18137), .ZN(n17782) );
  INV_X1 U16319 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18129) );
  NOR2_X1 U16320 ( .A1(n17782), .A2(n18129), .ZN(n18109) );
  NAND2_X1 U16321 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18109), .ZN(
        n18103) );
  INV_X1 U16322 ( .A(n18103), .ZN(n13417) );
  NAND2_X1 U16323 ( .A1(n13163), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13162) );
  INV_X1 U16324 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18597) );
  AOI22_X1 U16325 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9716), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13161) );
  INV_X1 U16326 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n21155) );
  AOI22_X1 U16327 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13152) );
  OAI211_X1 U16328 ( .C1(n17298), .C2(n21155), .A(n13153), .B(n13152), .ZN(
        n13159) );
  AOI22_X1 U16329 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U16330 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U16331 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U16332 ( .A1(n13113), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13154) );
  NAND4_X1 U16333 ( .A1(n13157), .A2(n13156), .A3(n13155), .A4(n13154), .ZN(
        n13158) );
  AOI211_X1 U16334 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n13159), .B(n13158), .ZN(n13160) );
  OAI211_X1 U16335 ( .C1(n13089), .C2(n18597), .A(n13161), .B(n13160), .ZN(
        n16080) );
  INV_X1 U16336 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19011) );
  NOR2_X1 U16337 ( .A1(n18053), .A2(n19011), .ZN(n18052) );
  INV_X1 U16338 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18994) );
  NAND2_X1 U16339 ( .A1(n18052), .A2(n18045), .ZN(n18044) );
  NAND2_X1 U16340 ( .A1(n13162), .A2(n18044), .ZN(n18036) );
  XNOR2_X1 U16341 ( .A(n17567), .B(n13163), .ZN(n13164) );
  INV_X1 U16342 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18341) );
  XNOR2_X1 U16343 ( .A(n13164), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18037) );
  NAND2_X1 U16344 ( .A1(n18036), .A2(n18037), .ZN(n18035) );
  OR2_X1 U16345 ( .A1(n18341), .A2(n13164), .ZN(n13165) );
  NAND2_X1 U16346 ( .A1(n18035), .A2(n13165), .ZN(n18026) );
  NAND2_X1 U16347 ( .A1(n18026), .A2(n18027), .ZN(n18025) );
  NAND2_X1 U16348 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13168), .ZN(
        n13169) );
  NAND2_X1 U16349 ( .A1(n18025), .A2(n13169), .ZN(n18010) );
  XNOR2_X1 U16350 ( .A(n13170), .B(n9718), .ZN(n13171) );
  XOR2_X1 U16351 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n13171), .Z(
        n18011) );
  NAND2_X1 U16352 ( .A1(n18010), .A2(n18011), .ZN(n18009) );
  NAND2_X1 U16353 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13171), .ZN(
        n13172) );
  NAND2_X2 U16354 ( .A1(n18009), .A2(n13172), .ZN(n13175) );
  XOR2_X1 U16355 ( .A(n17556), .B(n13173), .Z(n13176) );
  XNOR2_X2 U16356 ( .A(n13175), .B(n13174), .ZN(n18003) );
  NAND2_X1 U16357 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  XOR2_X1 U16358 ( .A(n17552), .B(n13178), .Z(n13179) );
  XOR2_X1 U16359 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13179), .Z(
        n17986) );
  NAND2_X1 U16360 ( .A1(n17985), .A2(n17986), .ZN(n17984) );
  NAND2_X1 U16361 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13179), .ZN(
        n13180) );
  NAND2_X1 U16362 ( .A1(n17984), .A2(n13180), .ZN(n13182) );
  OAI21_X1 U16363 ( .B1(n17548), .B2(n16566), .A(n17847), .ZN(n13181) );
  INV_X1 U16364 ( .A(n13181), .ZN(n13183) );
  XNOR2_X1 U16365 ( .A(n13182), .B(n13181), .ZN(n17973) );
  NAND2_X1 U16366 ( .A1(n13183), .A2(n13182), .ZN(n13184) );
  INV_X1 U16367 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17943) );
  NAND2_X1 U16368 ( .A1(n17931), .A2(n17943), .ZN(n17919) );
  NOR2_X2 U16369 ( .A1(n17919), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17901) );
  INV_X1 U16370 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17904) );
  NOR2_X1 U16371 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18195) );
  INV_X1 U16372 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18203) );
  NAND2_X1 U16373 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17920) );
  INV_X1 U16374 ( .A(n17920), .ZN(n18247) );
  NAND2_X1 U16375 ( .A1(n18247), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18228) );
  INV_X1 U16376 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18227) );
  NOR2_X1 U16377 ( .A1(n18228), .A2(n18227), .ZN(n18202) );
  NAND2_X1 U16378 ( .A1(n18202), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18204) );
  NOR2_X1 U16379 ( .A1(n18203), .A2(n18204), .ZN(n18180) );
  NAND2_X1 U16380 ( .A1(n18180), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18163) );
  INV_X1 U16381 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18182) );
  NOR2_X2 U16382 ( .A1(n17839), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17838) );
  NAND2_X1 U16383 ( .A1(n18190), .A2(n13188), .ZN(n17848) );
  INV_X1 U16384 ( .A(n17848), .ZN(n13193) );
  INV_X1 U16385 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18171) );
  NOR2_X1 U16386 ( .A1(n18182), .A2(n18171), .ZN(n18158) );
  NAND2_X1 U16387 ( .A1(n18158), .A2(n13417), .ZN(n13397) );
  INV_X1 U16388 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18131) );
  NAND2_X1 U16389 ( .A1(n18131), .A2(n17847), .ZN(n17824) );
  NOR2_X1 U16390 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17824), .ZN(
        n13189) );
  INV_X1 U16391 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21224) );
  NAND2_X1 U16392 ( .A1(n13189), .A2(n21224), .ZN(n17795) );
  INV_X1 U16393 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18113) );
  NAND3_X1 U16394 ( .A1(n17783), .A2(n18113), .A3(n18129), .ZN(n13190) );
  INV_X1 U16395 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18082) );
  INV_X1 U16396 ( .A(n18158), .ZN(n17832) );
  INV_X1 U16397 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21220) );
  NOR2_X2 U16398 ( .A1(n17732), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17731) );
  NAND2_X1 U16399 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13396) );
  NOR2_X1 U16400 ( .A1(n17731), .A2(n13196), .ZN(n13198) );
  NOR2_X1 U16401 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17958), .ZN(
        n13197) );
  NAND2_X1 U16402 ( .A1(n16561), .A2(n13197), .ZN(n16014) );
  NAND2_X1 U16403 ( .A1(n13198), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16560) );
  INV_X1 U16404 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16537) );
  OAI22_X1 U16405 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n13200), .B1(
        n13389), .B2(n17847), .ZN(n13206) );
  NAND2_X1 U16406 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17958), .ZN(
        n13201) );
  INV_X1 U16407 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13398) );
  OAI22_X1 U16408 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17958), .B1(
        n13201), .B2(n13398), .ZN(n13205) );
  OAI211_X1 U16409 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n13398), .A(
        n13203), .B(n13202), .ZN(n13204) );
  AOI22_X1 U16410 ( .A1(n13207), .A2(n13206), .B1(n13205), .B2(n13204), .ZN(
        n16555) );
  INV_X1 U16411 ( .A(n17548), .ZN(n13347) );
  AOI21_X1 U16412 ( .B1(n18833), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13209), .ZN(n13215) );
  OAI21_X1 U16413 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13063), .A(
        n13210), .ZN(n13211) );
  OAI22_X1 U16414 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18859), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13211), .ZN(n13216) );
  NOR2_X1 U16415 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18859), .ZN(
        n13212) );
  NAND2_X1 U16416 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13211), .ZN(
        n13217) );
  AOI22_X1 U16417 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13216), .B1(
        n13212), .B2(n13217), .ZN(n13221) );
  OAI21_X1 U16418 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18834), .A(
        n13334), .ZN(n13338) );
  NOR2_X1 U16419 ( .A1(n13333), .A2(n13338), .ZN(n13220) );
  OAI21_X1 U16420 ( .B1(n13215), .B2(n13214), .A(n13221), .ZN(n13213) );
  AOI21_X1 U16421 ( .B1(n13217), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n13216), .ZN(n13218) );
  AOI21_X1 U16422 ( .B1(n18859), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13218), .ZN(n13219) );
  INV_X1 U16423 ( .A(n13219), .ZN(n13335) );
  AOI22_X1 U16424 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13222) );
  OAI21_X1 U16425 ( .B1(n17373), .B2(n17354), .A(n13222), .ZN(n13226) );
  INV_X1 U16426 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18601) );
  AOI22_X1 U16427 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13224) );
  AOI22_X1 U16428 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13223) );
  OAI211_X1 U16429 ( .C1(n17298), .C2(n18601), .A(n13224), .B(n13223), .ZN(
        n13225) );
  AOI211_X1 U16430 ( .C1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .C2(n13113), .A(
        n13226), .B(n13225), .ZN(n13233) );
  INV_X1 U16431 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U16432 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17314), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13227) );
  OAI21_X1 U16433 ( .B1(n17229), .B2(n17214), .A(n13227), .ZN(n13231) );
  AOI22_X1 U16434 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13229) );
  INV_X1 U16435 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15929) );
  NAND3_X1 U16436 ( .A1(n13229), .A2(n10098), .A3(n13228), .ZN(n13230) );
  AND2_X2 U16437 ( .A1(n13233), .A2(n13232), .ZN(n19033) );
  AOI22_X1 U16438 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13243) );
  INV_X1 U16439 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17278) );
  AOI22_X1 U16440 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U16441 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13234) );
  OAI211_X1 U16442 ( .C1(n17298), .C2(n17278), .A(n13235), .B(n13234), .ZN(
        n13241) );
  AOI22_X1 U16443 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13239) );
  AOI22_X1 U16444 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13238) );
  AOI22_X1 U16445 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13237) );
  NAND2_X1 U16446 ( .A1(n13113), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13236) );
  NAND4_X1 U16447 ( .A1(n13239), .A2(n13238), .A3(n13237), .A4(n13236), .ZN(
        n13240) );
  OAI22_X1 U16448 ( .A1(n17298), .A2(n15967), .B1(n17322), .B2(n17407), .ZN(
        n13248) );
  AOI22_X1 U16449 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U16450 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9767), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U16451 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13244) );
  NAND3_X1 U16452 ( .A1(n13246), .A2(n13245), .A3(n13244), .ZN(n13247) );
  AOI211_X1 U16453 ( .C1(n17368), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n13248), .B(n13247), .ZN(n13256) );
  INV_X1 U16454 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17294) );
  AOI22_X1 U16455 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13249) );
  OAI21_X1 U16456 ( .B1(n9785), .B2(n17294), .A(n13249), .ZN(n13254) );
  AOI22_X1 U16457 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13252) );
  INV_X1 U16458 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15968) );
  AOI22_X1 U16459 ( .A1(n13113), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13257) );
  OAI21_X1 U16460 ( .B1(n17210), .B2(n21214), .A(n13257), .ZN(n13261) );
  AOI22_X1 U16461 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13259) );
  AOI22_X1 U16462 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13258) );
  OAI211_X1 U16463 ( .C1(n17298), .C2(n18614), .A(n13259), .B(n13258), .ZN(
        n13260) );
  AOI211_X1 U16464 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n13261), .B(n13260), .ZN(n13269) );
  INV_X1 U16465 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U16466 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13262) );
  OAI21_X1 U16467 ( .B1(n13148), .B2(n17263), .A(n13262), .ZN(n13267) );
  AOI22_X1 U16468 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13265) );
  INV_X1 U16469 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U16470 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13279) );
  AOI22_X1 U16471 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13271) );
  AOI22_X1 U16472 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13270) );
  OAI211_X1 U16473 ( .C1(n17317), .C2(n21323), .A(n13271), .B(n13270), .ZN(
        n13277) );
  AOI22_X1 U16474 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9720), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13275) );
  AOI22_X1 U16475 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U16476 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13273) );
  NAND2_X1 U16477 ( .A1(n17377), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13272) );
  NAND4_X1 U16478 ( .A1(n13275), .A2(n13274), .A3(n13273), .A4(n13272), .ZN(
        n13276) );
  INV_X2 U16479 ( .A(n13340), .ZN(n18386) );
  NAND3_X1 U16480 ( .A1(n18822), .A2(n13342), .A3(n18386), .ZN(n13324) );
  NAND2_X1 U16481 ( .A1(n18398), .A2(n18386), .ZN(n13404) );
  INV_X1 U16482 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n21093) );
  OAI22_X1 U16483 ( .A1(n13090), .A2(n21093), .B1(n17338), .B2(n18438), .ZN(
        n13284) );
  AOI22_X1 U16484 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U16485 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17332), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16486 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17377), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13280) );
  NAND3_X1 U16487 ( .A1(n13282), .A2(n13281), .A3(n13280), .ZN(n13283) );
  AOI211_X1 U16488 ( .C1(n9765), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n13284), .B(n13283), .ZN(n13291) );
  AOI22_X1 U16489 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13290) );
  AOI22_X1 U16490 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13285) );
  OAI21_X1 U16491 ( .B1(n17322), .B2(n21122), .A(n13285), .ZN(n13288) );
  INV_X1 U16492 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17101) );
  NAND3_X1 U16493 ( .A1(n13291), .A2(n13290), .A3(n13289), .ZN(n13292) );
  AOI22_X1 U16494 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13302) );
  AOI22_X1 U16495 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13294) );
  AOI22_X1 U16496 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13293) );
  OAI211_X1 U16497 ( .C1(n17298), .C2(n21200), .A(n13294), .B(n13293), .ZN(
        n13300) );
  AOI22_X1 U16498 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13298) );
  AOI22_X1 U16499 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U16500 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13296) );
  NAND2_X1 U16501 ( .A1(n13113), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13295) );
  NAND4_X1 U16502 ( .A1(n13298), .A2(n13297), .A3(n13296), .A4(n13295), .ZN(
        n13299) );
  AOI22_X1 U16503 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U16504 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13303) );
  OAI211_X1 U16505 ( .C1(n17338), .C2(n18418), .A(n13304), .B(n13303), .ZN(
        n13310) );
  AOI22_X1 U16506 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9767), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13308) );
  AOI22_X1 U16507 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13307) );
  AOI22_X1 U16508 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13306) );
  NAND2_X1 U16509 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13305) );
  NAND4_X1 U16510 ( .A1(n13308), .A2(n13307), .A3(n13306), .A4(n13305), .ZN(
        n13309) );
  NAND2_X1 U16511 ( .A1(n13292), .A2(n18379), .ZN(n13317) );
  NAND2_X1 U16512 ( .A1(n17432), .A2(n18398), .ZN(n13319) );
  AND2_X1 U16513 ( .A1(n13340), .A2(n13329), .ZN(n16672) );
  INV_X1 U16514 ( .A(n16696), .ZN(n13316) );
  NAND2_X1 U16515 ( .A1(n18386), .A2(n13326), .ZN(n18821) );
  NAND2_X1 U16516 ( .A1(n19033), .A2(n18379), .ZN(n16076) );
  INV_X1 U16517 ( .A(n16076), .ZN(n13313) );
  OAI211_X1 U16518 ( .C1(n18410), .C2(n18829), .A(n17579), .B(n19033), .ZN(
        n13409) );
  AOI22_X1 U16519 ( .A1(n13341), .A2(n18829), .B1(n13326), .B2(n13317), .ZN(
        n13323) );
  NAND2_X1 U16520 ( .A1(n13292), .A2(n13319), .ZN(n13321) );
  INV_X1 U16521 ( .A(n13346), .ZN(n13320) );
  AOI22_X1 U16522 ( .A1(n13321), .A2(n18393), .B1(n13320), .B2(n13319), .ZN(
        n13322) );
  OAI211_X1 U16523 ( .C1(n17579), .C2(n13324), .A(n13323), .B(n13322), .ZN(
        n13407) );
  INV_X1 U16524 ( .A(n13407), .ZN(n13325) );
  OAI211_X1 U16525 ( .C1(n13327), .C2(n13326), .A(n13409), .B(n13325), .ZN(
        n13330) );
  INV_X1 U16526 ( .A(n13330), .ZN(n13328) );
  NAND2_X1 U16527 ( .A1(n13329), .A2(n13328), .ZN(n16001) );
  NOR2_X1 U16528 ( .A1(n13345), .A2(n16696), .ZN(n13331) );
  AOI21_X1 U16529 ( .B1(n13331), .B2(n17642), .A(n13330), .ZN(n18820) );
  NOR2_X2 U16530 ( .A1(n18822), .A2(n13332), .ZN(n16000) );
  NAND2_X1 U16531 ( .A1(n16076), .A2(n15912), .ZN(n19047) );
  INV_X1 U16532 ( .A(n13337), .ZN(n13339) );
  XOR2_X1 U16533 ( .A(n13334), .B(n13333), .Z(n13336) );
  OAI21_X1 U16534 ( .B1(n13339), .B2(n13338), .A(n18812), .ZN(n13415) );
  INV_X1 U16535 ( .A(n13415), .ZN(n18813) );
  NOR2_X1 U16536 ( .A1(n19033), .A2(n13340), .ZN(n13406) );
  NAND2_X1 U16537 ( .A1(n13406), .A2(n17432), .ZN(n13413) );
  AOI21_X1 U16538 ( .B1(n13342), .B2(n13341), .A(n18829), .ZN(n13343) );
  INV_X1 U16539 ( .A(n13343), .ZN(n13344) );
  NAND3_X1 U16540 ( .A1(n13346), .A2(n13345), .A3(n13344), .ZN(n13408) );
  NOR3_X1 U16541 ( .A1(n18871), .A2(n18866), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18867) );
  NAND2_X1 U16542 ( .A1(n16555), .A2(n17953), .ZN(n13387) );
  INV_X1 U16543 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18887) );
  NAND2_X1 U16544 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18363) );
  NAND2_X1 U16545 ( .A1(n18983), .A2(n18363), .ZN(n19028) );
  INV_X1 U16546 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19032) );
  NOR2_X1 U16547 ( .A1(n18887), .A2(n19032), .ZN(n17851) );
  INV_X1 U16548 ( .A(n17851), .ZN(n18017) );
  INV_X1 U16549 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16723) );
  INV_X1 U16550 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21104) );
  NAND2_X1 U16551 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17960) );
  NAND2_X1 U16552 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17922) );
  NOR2_X1 U16553 ( .A1(n17960), .A2(n17922), .ZN(n16929) );
  NAND2_X1 U16554 ( .A1(n16929), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16888) );
  INV_X1 U16555 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17910) );
  NOR2_X1 U16556 ( .A1(n17910), .A2(n17896), .ZN(n17891) );
  NAND3_X1 U16557 ( .A1(n17892), .A2(n17891), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17850) );
  NAND2_X1 U16558 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17856) );
  NAND2_X1 U16559 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17814) );
  INV_X1 U16560 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21288) );
  INV_X1 U16561 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17792) );
  NOR2_X1 U16562 ( .A1(n21288), .A2(n17792), .ZN(n17780) );
  INV_X1 U16563 ( .A(n17780), .ZN(n16709) );
  NAND2_X1 U16564 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17740) );
  NAND2_X1 U16565 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17710) );
  NAND2_X1 U16566 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n13391), .ZN(
        n13349) );
  XOR2_X2 U16567 ( .A(n16723), .B(n13349), .Z(n17002) );
  INV_X1 U16568 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18970) );
  NOR2_X1 U16569 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19010) );
  INV_X1 U16570 ( .A(n19010), .ZN(n18996) );
  NOR2_X1 U16571 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18996), .ZN(n19045) );
  NOR2_X1 U16572 ( .A1(n18970), .A2(n18358), .ZN(n16553) );
  INV_X1 U16573 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16727) );
  NOR2_X1 U16574 ( .A1(n18866), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n17895) );
  NOR2_X1 U16575 ( .A1(n18983), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19008) );
  INV_X1 U16576 ( .A(n19008), .ZN(n19002) );
  OAI21_X1 U16577 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n18363), .ZN(n18890) );
  NAND2_X1 U16578 ( .A1(n19002), .A2(n18890), .ZN(n18377) );
  NOR3_X1 U16579 ( .A1(n19032), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n15997) );
  OAI21_X1 U16580 ( .B1(n21104), .B2(n17837), .A(n18693), .ZN(n17854) );
  NOR2_X1 U16581 ( .A1(n17813), .A2(n13350), .ZN(n13351) );
  INV_X1 U16582 ( .A(n13351), .ZN(n13393) );
  NOR2_X1 U16583 ( .A1(n16727), .A2(n13393), .ZN(n13352) );
  NOR2_X1 U16584 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17837), .ZN(
        n16543) );
  NOR2_X1 U16585 ( .A1(n21104), .A2(n17739), .ZN(n16710) );
  NAND3_X1 U16586 ( .A1(n16710), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17695) );
  NOR2_X1 U16587 ( .A1(n10020), .A2(n17695), .ZN(n16706) );
  NAND2_X1 U16588 ( .A1(n16706), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16705) );
  INV_X1 U16589 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16704) );
  NOR2_X1 U16590 ( .A1(n16705), .A2(n16704), .ZN(n16703) );
  INV_X1 U16591 ( .A(n17895), .ZN(n18891) );
  NAND2_X1 U16592 ( .A1(n18753), .A2(n13350), .ZN(n16530) );
  OAI211_X1 U16593 ( .C1(n16703), .C2(n18891), .A(n18054), .B(n16530), .ZN(
        n16532) );
  AOI211_X1 U16594 ( .C1(n13351), .C2(n16727), .A(n16543), .B(n16532), .ZN(
        n13392) );
  INV_X1 U16595 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18993) );
  NAND2_X1 U16596 ( .A1(n17567), .A2(n13355), .ZN(n13354) );
  NAND2_X1 U16597 ( .A1(n13354), .A2(n13353), .ZN(n13362) );
  NOR2_X1 U16598 ( .A1(n9718), .A2(n13362), .ZN(n13366) );
  NAND2_X1 U16599 ( .A1(n13366), .A2(n13365), .ZN(n13368) );
  NOR2_X1 U16600 ( .A1(n17552), .A2(n13368), .ZN(n13372) );
  NAND2_X1 U16601 ( .A1(n13372), .A2(n17548), .ZN(n13373) );
  XNOR2_X1 U16602 ( .A(n13354), .B(n17562), .ZN(n13360) );
  NOR2_X1 U16603 ( .A1(n13358), .A2(n18341), .ZN(n13359) );
  NOR2_X1 U16604 ( .A1(n13163), .A2(n19011), .ZN(n13357) );
  NAND3_X1 U16605 ( .A1(n18053), .A2(n13163), .A3(n19011), .ZN(n13356) );
  OAI221_X1 U16606 ( .B1(n13357), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18053), .C2(n13163), .A(n13356), .ZN(n18335) );
  XOR2_X1 U16607 ( .A(n13167), .B(n13360), .Z(n18023) );
  INV_X1 U16608 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18313) );
  NOR2_X1 U16609 ( .A1(n13363), .A2(n18313), .ZN(n13364) );
  XNOR2_X1 U16610 ( .A(n13362), .B(n9718), .ZN(n18014) );
  XNOR2_X1 U16611 ( .A(n13366), .B(n13365), .ZN(n18000) );
  NOR2_X1 U16612 ( .A1(n17999), .A2(n18000), .ZN(n13367) );
  NAND2_X1 U16613 ( .A1(n17999), .A2(n18000), .ZN(n17998) );
  XNOR2_X1 U16614 ( .A(n13368), .B(n17552), .ZN(n13369) );
  NOR2_X1 U16615 ( .A1(n13370), .A2(n13369), .ZN(n13371) );
  INV_X1 U16616 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18297) );
  XNOR2_X1 U16617 ( .A(n13372), .B(n17548), .ZN(n13375) );
  INV_X1 U16618 ( .A(n13373), .ZN(n13378) );
  OR2_X1 U16619 ( .A1(n13375), .A2(n13374), .ZN(n17979) );
  OAI21_X1 U16620 ( .B1(n13378), .B2(n13377), .A(n17979), .ZN(n13376) );
  INV_X1 U16621 ( .A(n13397), .ZN(n13381) );
  NAND2_X1 U16622 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16533) );
  NOR2_X1 U16623 ( .A1(n16533), .A2(n16537), .ZN(n13423) );
  INV_X1 U16624 ( .A(n13423), .ZN(n16551) );
  NAND2_X1 U16625 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16536), .ZN(
        n13380) );
  XNOR2_X1 U16626 ( .A(n18993), .B(n13380), .ZN(n16559) );
  NAND2_X1 U16627 ( .A1(n13381), .A2(n16563), .ZN(n18096) );
  NAND2_X1 U16628 ( .A1(n9922), .A2(n17737), .ZN(n18063) );
  NAND2_X1 U16629 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16534), .ZN(
        n13382) );
  XOR2_X1 U16630 ( .A(n18993), .B(n13382), .Z(n16556) );
  NAND2_X1 U16631 ( .A1(n16556), .A2(n17968), .ZN(n13383) );
  OAI21_X1 U16632 ( .B1(n16559), .B2(n18058), .A(n13383), .ZN(n13384) );
  INV_X1 U16633 ( .A(n13384), .ZN(n13385) );
  NAND2_X1 U16634 ( .A1(n13387), .A2(n13386), .ZN(P3_U2799) );
  NOR2_X1 U16635 ( .A1(n13389), .A2(n13388), .ZN(n13390) );
  XOR2_X1 U16636 ( .A(n13390), .B(n13398), .Z(n13435) );
  INV_X1 U16637 ( .A(n13391), .ZN(n16541) );
  AOI22_X1 U16638 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n13391), .B1(
        n16541), .B2(n16727), .ZN(n16726) );
  AOI21_X1 U16639 ( .B1(n16727), .B2(n13393), .A(n13392), .ZN(n13394) );
  INV_X1 U16640 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18972) );
  NOR2_X1 U16641 ( .A1(n18358), .A2(n18972), .ZN(n13427) );
  AOI211_X1 U16642 ( .C1(n17914), .C2(n16726), .A(n13394), .B(n13427), .ZN(
        n13401) );
  INV_X1 U16643 ( .A(n17968), .ZN(n17887) );
  OAI22_X1 U16644 ( .A1(n16536), .A2(n18058), .B1(n16534), .B2(n17887), .ZN(
        n13395) );
  NAND2_X1 U16645 ( .A1(n13395), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13400) );
  NOR2_X1 U16646 ( .A1(n18082), .A2(n13396), .ZN(n13418) );
  NAND2_X1 U16647 ( .A1(n9792), .A2(n10117), .ZN(n13399) );
  NAND3_X1 U16648 ( .A1(n13401), .A2(n13400), .A3(n13399), .ZN(n13402) );
  AOI21_X1 U16649 ( .B1(n13435), .B2(n17953), .A(n13402), .ZN(n13403) );
  INV_X1 U16650 ( .A(n13403), .ZN(P3_U2800) );
  INV_X1 U16651 ( .A(n13404), .ZN(n13412) );
  INV_X1 U16652 ( .A(n18812), .ZN(n16677) );
  NAND2_X1 U16653 ( .A1(n18910), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19042) );
  INV_X2 U16654 ( .A(n19042), .ZN(n19041) );
  NAND2_X1 U16655 ( .A1(n19041), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18973) );
  OAI211_X1 U16656 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18910), .B(n18967), .ZN(n19031) );
  OAI21_X1 U16657 ( .B1(n18386), .B2(n17642), .A(n19031), .ZN(n13405) );
  NAND2_X1 U16658 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19034) );
  OAI21_X1 U16659 ( .B1(n13406), .B2(n13405), .A(n19034), .ZN(n16676) );
  NOR3_X1 U16660 ( .A1(n13412), .A2(n16677), .A3(n16676), .ZN(n13411) );
  NOR2_X1 U16661 ( .A1(n13408), .A2(n13407), .ZN(n13410) );
  OAI21_X1 U16662 ( .B1(n13410), .B2(n16672), .A(n13409), .ZN(n15999) );
  AOI211_X1 U16663 ( .C1(n13412), .C2(n18809), .A(n13411), .B(n15999), .ZN(
        n13414) );
  AOI221_X4 U16664 ( .B1(n13415), .B2(n13414), .C1(n13413), .C2(n13414), .A(
        n18883), .ZN(n18338) );
  NAND2_X1 U16665 ( .A1(n13425), .A2(n17548), .ZN(n18074) );
  NOR2_X1 U16666 ( .A1(n18341), .A2(n18994), .ZN(n18308) );
  INV_X1 U16667 ( .A(n18308), .ZN(n13416) );
  NAND3_X1 U16668 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18162) );
  NOR2_X1 U16669 ( .A1(n13416), .A2(n18162), .ZN(n18266) );
  INV_X1 U16670 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18285) );
  NOR3_X1 U16671 ( .A1(n18285), .A2(n18297), .A3(n9918), .ZN(n18217) );
  NAND2_X1 U16672 ( .A1(n18266), .A2(n18217), .ZN(n18201) );
  NOR2_X1 U16673 ( .A1(n18163), .A2(n18201), .ZN(n18155) );
  NAND2_X1 U16674 ( .A1(n18158), .A2(n18155), .ZN(n13422) );
  NAND2_X1 U16675 ( .A1(n13417), .A2(n13418), .ZN(n16565) );
  INV_X1 U16676 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18059) );
  NAND2_X1 U16677 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n13418), .ZN(
        n13419) );
  NOR3_X1 U16678 ( .A1(n18129), .A2(n18059), .A3(n13419), .ZN(n13420) );
  INV_X1 U16679 ( .A(n17782), .ZN(n18122) );
  INV_X1 U16680 ( .A(n13422), .ZN(n13428) );
  NAND2_X1 U16681 ( .A1(n18122), .A2(n13428), .ZN(n18062) );
  OAI21_X1 U16682 ( .B1(n19011), .B2(n18062), .A(n18828), .ZN(n18060) );
  OAI21_X1 U16683 ( .B1(n19011), .B2(n18994), .A(n18341), .ZN(n18161) );
  INV_X1 U16684 ( .A(n18161), .ZN(n18328) );
  NOR2_X1 U16685 ( .A1(n18328), .A2(n18162), .ZN(n18268) );
  NAND2_X1 U16686 ( .A1(n18217), .A2(n18268), .ZN(n18176) );
  NOR3_X1 U16687 ( .A1(n18163), .A2(n17832), .A3(n18176), .ZN(n18116) );
  NAND2_X1 U16688 ( .A1(n18109), .A2(n18116), .ZN(n18100) );
  OAI21_X1 U16689 ( .B1(n18100), .B2(n13419), .A(n18851), .ZN(n18065) );
  OAI211_X1 U16690 ( .C1(n18843), .C2(n13420), .A(n18060), .B(n18065), .ZN(
        n13421) );
  AOI221_X1 U16691 ( .B1(n13422), .B2(n18818), .C1(n16565), .C2(n18818), .A(
        n13421), .ZN(n16010) );
  OAI21_X1 U16692 ( .B1(n16011), .B2(n13423), .A(n16010), .ZN(n13424) );
  AOI21_X1 U16693 ( .B1(n18338), .B2(n13424), .A(n18291), .ZN(n16548) );
  INV_X1 U16694 ( .A(n16548), .ZN(n13426) );
  INV_X1 U16695 ( .A(n13425), .ZN(n18814) );
  NAND2_X1 U16696 ( .A1(n18338), .A2(n18191), .ZN(n18210) );
  NAND2_X1 U16697 ( .A1(n18808), .A2(n18338), .ZN(n18317) );
  OAI22_X1 U16698 ( .A1(n16534), .A2(n18210), .B1(n16536), .B2(n18317), .ZN(
        n16012) );
  OAI21_X1 U16699 ( .B1(n13426), .B2(n16012), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13433) );
  INV_X1 U16700 ( .A(n13427), .ZN(n13432) );
  INV_X1 U16701 ( .A(n18064), .ZN(n17700) );
  INV_X1 U16702 ( .A(n18191), .ZN(n18239) );
  AOI21_X1 U16703 ( .B1(n18832), .B2(n19011), .A(n9863), .ZN(n18329) );
  AOI22_X1 U16704 ( .A1(n18851), .A2(n18116), .B1(n13428), .B2(n18329), .ZN(
        n16564) );
  NOR3_X1 U16705 ( .A1(n16564), .A2(n18082), .A3(n18103), .ZN(n18081) );
  NAND2_X1 U16706 ( .A1(n9922), .A2(n18081), .ZN(n16549) );
  OAI21_X1 U16707 ( .B1(n18239), .B2(n18063), .A(n16549), .ZN(n13429) );
  AOI22_X1 U16708 ( .A1(n17700), .A2(n18355), .B1(n18338), .B2(n13429), .ZN(
        n16017) );
  INV_X1 U16709 ( .A(n16017), .ZN(n13430) );
  NAND3_X1 U16710 ( .A1(n13433), .A2(n13432), .A3(n13431), .ZN(n13434) );
  AOI21_X1 U16711 ( .B1(n13435), .B2(n18263), .A(n13434), .ZN(n13436) );
  INV_X1 U16712 ( .A(n13436), .ZN(P3_U2832) );
  INV_X1 U16713 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21008) );
  NOR3_X1 U16714 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21008), .ZN(n13438) );
  NOR4_X1 U16715 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13437) );
  NAND4_X1 U16716 ( .A1(n20239), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13438), .A4(
        n13437), .ZN(U214) );
  NOR2_X1 U16717 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13440) );
  NOR4_X1 U16718 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13439) );
  NAND4_X1 U16719 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13440), .A4(n13439), .ZN(n13441) );
  NOR2_X1 U16720 ( .A1(n15276), .A2(n13441), .ZN(n16580) );
  NAND2_X1 U16721 ( .A1(n16580), .A2(U214), .ZN(U212) );
  NOR2_X1 U16722 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13441), .ZN(n16653)
         );
  AOI211_X1 U16723 ( .C1(n15324), .C2(n13443), .A(n13442), .B(n19928), .ZN(
        n13455) );
  INV_X1 U16724 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n21112) );
  OAI22_X1 U16725 ( .A1(n21112), .A2(n19252), .B1(n19989), .B2(n19222), .ZN(
        n13454) );
  INV_X1 U16726 ( .A(n13444), .ZN(n13445) );
  OAI22_X1 U16727 ( .A1(n13445), .A2(n19270), .B1(n19250), .B2(n15322), .ZN(
        n13453) );
  OAI21_X1 U16728 ( .B1(n15201), .B2(n13447), .A(n13446), .ZN(n15558) );
  NAND2_X1 U16729 ( .A1(n13448), .A2(n13449), .ZN(n13450) );
  AND2_X1 U16730 ( .A1(n15098), .A2(n13450), .ZN(n15555) );
  INV_X1 U16731 ( .A(n15555), .ZN(n13451) );
  OAI22_X1 U16732 ( .A1(n15558), .A2(n19230), .B1(n13451), .B2(n19258), .ZN(
        n13452) );
  OR4_X1 U16733 ( .A1(n13455), .A2(n13454), .A3(n13453), .A4(n13452), .ZN(
        P2_U2828) );
  INV_X1 U16734 ( .A(n14201), .ZN(n19276) );
  INV_X1 U16735 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13457) );
  NOR2_X1 U16736 ( .A1(n20013), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13460) );
  INV_X1 U16737 ( .A(n13460), .ZN(n13456) );
  OAI211_X1 U16738 ( .C1(n19276), .C2(n13457), .A(n13463), .B(n13456), .ZN(
        P2_U2814) );
  NOR4_X1 U16739 ( .A1(n10253), .A2(n13459), .A3(n13458), .A4(n16502), .ZN(
        n16496) );
  NOR2_X1 U16740 ( .A1(n16496), .A2(n13464), .ZN(n20050) );
  OAI211_X1 U16741 ( .C1(n20050), .C2(n13551), .A(n16436), .B(n16435), .ZN(
        P2_U2819) );
  INV_X1 U16742 ( .A(n19057), .ZN(n15073) );
  OAI21_X1 U16743 ( .B1(n13460), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n15073), 
        .ZN(n13461) );
  OAI21_X1 U16744 ( .B1(n13462), .B2(n15073), .A(n13461), .ZN(P2_U3612) );
  INV_X1 U16745 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19363) );
  NOR2_X1 U16746 ( .A1(n13464), .A2(n19942), .ZN(n13465) );
  AND2_X1 U16747 ( .A1(n10263), .A2(n13465), .ZN(n13466) );
  NAND2_X1 U16748 ( .A1(n13467), .A2(n13466), .ZN(n13540) );
  NAND2_X1 U16749 ( .A1(n19394), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13470) );
  INV_X1 U16750 ( .A(n13540), .ZN(n19389) );
  NAND2_X1 U16751 ( .A1(n15276), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13469) );
  INV_X1 U16752 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16611) );
  OR2_X1 U16753 ( .A1(n15276), .A2(n16611), .ZN(n13468) );
  NAND2_X1 U16754 ( .A1(n13469), .A2(n13468), .ZN(n19304) );
  NAND2_X1 U16755 ( .A1(n19389), .A2(n19304), .ZN(n13500) );
  OAI211_X1 U16756 ( .C1(n19363), .C2(n13568), .A(n13470), .B(n13500), .ZN(
        P2_U2979) );
  INV_X1 U16757 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19366) );
  NAND2_X1 U16758 ( .A1(n19394), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13473) );
  NAND2_X1 U16759 ( .A1(n15276), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13472) );
  INV_X1 U16760 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16615) );
  OR2_X1 U16761 ( .A1(n15276), .A2(n16615), .ZN(n13471) );
  NAND2_X1 U16762 ( .A1(n13472), .A2(n13471), .ZN(n19309) );
  NAND2_X1 U16763 ( .A1(n19389), .A2(n19309), .ZN(n13502) );
  OAI211_X1 U16764 ( .C1(n19366), .C2(n13568), .A(n13473), .B(n13502), .ZN(
        P2_U2977) );
  INV_X1 U16765 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15268) );
  NAND2_X1 U16766 ( .A1(n19394), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13477) );
  INV_X1 U16767 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14232) );
  OR2_X1 U16768 ( .A1(n15276), .A2(n14232), .ZN(n13475) );
  NAND2_X1 U16769 ( .A1(n15276), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13474) );
  AND2_X1 U16770 ( .A1(n13475), .A2(n13474), .ZN(n19312) );
  INV_X1 U16771 ( .A(n19312), .ZN(n13476) );
  NAND2_X1 U16772 ( .A1(n19389), .A2(n13476), .ZN(n13482) );
  OAI211_X1 U16773 ( .C1(n13568), .C2(n15268), .A(n13477), .B(n13482), .ZN(
        P2_U2961) );
  INV_X1 U16774 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15256) );
  NAND2_X1 U16775 ( .A1(n19394), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13481) );
  INV_X1 U16776 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14424) );
  OR2_X1 U16777 ( .A1(n15276), .A2(n14424), .ZN(n13479) );
  NAND2_X1 U16778 ( .A1(n15276), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13478) );
  AND2_X1 U16779 ( .A1(n13479), .A2(n13478), .ZN(n19307) );
  INV_X1 U16780 ( .A(n19307), .ZN(n13480) );
  NAND2_X1 U16781 ( .A1(n19389), .A2(n13480), .ZN(n13494) );
  OAI211_X1 U16782 ( .C1(n13568), .C2(n15256), .A(n13481), .B(n13494), .ZN(
        P2_U2963) );
  INV_X1 U16783 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n13484) );
  NAND2_X1 U16784 ( .A1(n19394), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13483) );
  OAI211_X1 U16785 ( .C1(n13568), .C2(n13484), .A(n13483), .B(n13482), .ZN(
        P2_U2976) );
  INV_X1 U16786 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13486) );
  NAND2_X1 U16787 ( .A1(n19394), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13485) );
  OAI22_X1 U16788 ( .A1(n15276), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14002), .ZN(n14075) );
  INV_X1 U16789 ( .A(n14075), .ZN(n19288) );
  NAND2_X1 U16790 ( .A1(n19389), .A2(n19288), .ZN(n13497) );
  OAI211_X1 U16791 ( .C1(n13568), .C2(n13486), .A(n13485), .B(n13497), .ZN(
        P2_U2952) );
  INV_X1 U16792 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n13491) );
  NAND2_X1 U16793 ( .A1(n19394), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13490) );
  INV_X1 U16794 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14427) );
  OR2_X1 U16795 ( .A1(n15276), .A2(n14427), .ZN(n13488) );
  NAND2_X1 U16796 ( .A1(n15276), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13487) );
  AND2_X1 U16797 ( .A1(n13488), .A2(n13487), .ZN(n19302) );
  INV_X1 U16798 ( .A(n19302), .ZN(n13489) );
  NAND2_X1 U16799 ( .A1(n19389), .A2(n13489), .ZN(n13492) );
  OAI211_X1 U16800 ( .C1(n13568), .C2(n13491), .A(n13490), .B(n13492), .ZN(
        P2_U2980) );
  INV_X1 U16801 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15245) );
  NAND2_X1 U16802 ( .A1(n19394), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13493) );
  OAI211_X1 U16803 ( .C1(n13568), .C2(n15245), .A(n13493), .B(n13492), .ZN(
        P2_U2965) );
  INV_X1 U16804 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n13496) );
  NAND2_X1 U16805 ( .A1(n19394), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13495) );
  OAI211_X1 U16806 ( .C1(n13568), .C2(n13496), .A(n13495), .B(n13494), .ZN(
        P2_U2978) );
  NAND2_X1 U16807 ( .A1(n19394), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n13498) );
  OAI211_X1 U16808 ( .C1(n13568), .C2(n13499), .A(n13498), .B(n13497), .ZN(
        P2_U2967) );
  INV_X1 U16809 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13584) );
  NAND2_X1 U16810 ( .A1(n19394), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13501) );
  OAI211_X1 U16811 ( .C1(n13584), .C2(n13568), .A(n13501), .B(n13500), .ZN(
        P2_U2964) );
  INV_X1 U16812 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13573) );
  NAND2_X1 U16813 ( .A1(n19394), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13503) );
  OAI211_X1 U16814 ( .C1(n13573), .C2(n13568), .A(n13503), .B(n13502), .ZN(
        P2_U2962) );
  INV_X1 U16815 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13505) );
  AOI22_X1 U16816 ( .A1(n14002), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15276), .ZN(n19348) );
  NOR2_X1 U16817 ( .A1(n13540), .A2(n19348), .ZN(n13533) );
  AOI21_X1 U16818 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n19393), .A(n13533), .ZN(
        n13504) );
  OAI21_X1 U16819 ( .B1(n13541), .B2(n13505), .A(n13504), .ZN(P2_U2968) );
  INV_X1 U16820 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n13507) );
  AOI22_X1 U16821 ( .A1(n14002), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15276), .ZN(n19320) );
  NOR2_X1 U16822 ( .A1(n13540), .A2(n19320), .ZN(n13524) );
  AOI21_X1 U16823 ( .B1(n19393), .B2(P2_EAX_REG_6__SCAN_IN), .A(n13524), .ZN(
        n13506) );
  OAI21_X1 U16824 ( .B1(n13541), .B2(n13507), .A(n13506), .ZN(P2_U2973) );
  INV_X1 U16825 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13509) );
  OAI22_X1 U16826 ( .A1(n15276), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14002), .ZN(n19422) );
  NOR2_X1 U16827 ( .A1(n13540), .A2(n19422), .ZN(n13518) );
  AOI21_X1 U16828 ( .B1(n19393), .B2(P2_EAX_REG_2__SCAN_IN), .A(n13518), .ZN(
        n13508) );
  OAI21_X1 U16829 ( .B1(n13541), .B2(n13509), .A(n13508), .ZN(P2_U2969) );
  INV_X1 U16830 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13511) );
  OAI22_X1 U16831 ( .A1(n15276), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14002), .ZN(n19429) );
  NOR2_X1 U16832 ( .A1(n13540), .A2(n19429), .ZN(n13521) );
  AOI21_X1 U16833 ( .B1(n19393), .B2(P2_EAX_REG_20__SCAN_IN), .A(n13521), .ZN(
        n13510) );
  OAI21_X1 U16834 ( .B1(n13541), .B2(n13511), .A(n13510), .ZN(P2_U2956) );
  INV_X1 U16835 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13513) );
  AOI22_X1 U16836 ( .A1(n14002), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15276), .ZN(n19436) );
  NOR2_X1 U16837 ( .A1(n13540), .A2(n19436), .ZN(n13530) );
  AOI21_X1 U16838 ( .B1(n19393), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13530), .ZN(
        n13512) );
  OAI21_X1 U16839 ( .B1(n13541), .B2(n13513), .A(n13512), .ZN(P2_U2957) );
  INV_X1 U16840 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13515) );
  AOI22_X1 U16841 ( .A1(n14002), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15276), .ZN(n19318) );
  NOR2_X1 U16842 ( .A1(n13540), .A2(n19318), .ZN(n13527) );
  AOI21_X1 U16843 ( .B1(n19393), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13527), .ZN(
        n13514) );
  OAI21_X1 U16844 ( .B1(n13541), .B2(n13515), .A(n13514), .ZN(P2_U2959) );
  INV_X1 U16845 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U16846 ( .A1(n14002), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15276), .ZN(n19426) );
  NOR2_X1 U16847 ( .A1(n13540), .A2(n19426), .ZN(n13536) );
  AOI21_X1 U16848 ( .B1(n19393), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13536), .ZN(
        n13516) );
  OAI21_X1 U16849 ( .B1(n13541), .B2(n13517), .A(n13516), .ZN(P2_U2955) );
  INV_X1 U16850 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13520) );
  AOI21_X1 U16851 ( .B1(n19393), .B2(P2_EAX_REG_18__SCAN_IN), .A(n13518), .ZN(
        n13519) );
  OAI21_X1 U16852 ( .B1(n13541), .B2(n13520), .A(n13519), .ZN(P2_U2954) );
  INV_X1 U16853 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n13523) );
  AOI21_X1 U16854 ( .B1(n19393), .B2(P2_EAX_REG_4__SCAN_IN), .A(n13521), .ZN(
        n13522) );
  OAI21_X1 U16855 ( .B1(n13541), .B2(n13523), .A(n13522), .ZN(P2_U2971) );
  INV_X1 U16856 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13526) );
  AOI21_X1 U16857 ( .B1(n19393), .B2(P2_EAX_REG_22__SCAN_IN), .A(n13524), .ZN(
        n13525) );
  OAI21_X1 U16858 ( .B1(n13541), .B2(n13526), .A(n13525), .ZN(P2_U2958) );
  INV_X1 U16859 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13529) );
  AOI21_X1 U16860 ( .B1(n19393), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13527), .ZN(
        n13528) );
  OAI21_X1 U16861 ( .B1(n13541), .B2(n13529), .A(n13528), .ZN(P2_U2974) );
  INV_X1 U16862 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13532) );
  AOI21_X1 U16863 ( .B1(n19393), .B2(P2_EAX_REG_5__SCAN_IN), .A(n13530), .ZN(
        n13531) );
  OAI21_X1 U16864 ( .B1(n13541), .B2(n13532), .A(n13531), .ZN(P2_U2972) );
  INV_X1 U16865 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13535) );
  AOI21_X1 U16866 ( .B1(n19393), .B2(P2_EAX_REG_17__SCAN_IN), .A(n13533), .ZN(
        n13534) );
  OAI21_X1 U16867 ( .B1(n13541), .B2(n13535), .A(n13534), .ZN(P2_U2953) );
  INV_X1 U16868 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13538) );
  AOI21_X1 U16869 ( .B1(n19393), .B2(P2_EAX_REG_3__SCAN_IN), .A(n13536), .ZN(
        n13537) );
  OAI21_X1 U16870 ( .B1(n13541), .B2(n13538), .A(n13537), .ZN(P2_U2970) );
  INV_X1 U16871 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13542) );
  AOI22_X1 U16872 ( .A1(n14002), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15276), .ZN(n19298) );
  INV_X1 U16873 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13539) );
  OAI222_X1 U16874 ( .A1(n13542), .A2(n13541), .B1(n13540), .B2(n19298), .C1(
        n13539), .C2(n13568), .ZN(P2_U2982) );
  INV_X1 U16875 ( .A(n13543), .ZN(n13544) );
  NAND2_X1 U16876 ( .A1(n13545), .A2(n13544), .ZN(n13546) );
  NOR2_X1 U16877 ( .A1(n13547), .A2(n13546), .ZN(n13550) );
  NOR2_X1 U16878 ( .A1(n13548), .A2(n10954), .ZN(n13567) );
  NAND2_X1 U16879 ( .A1(n13567), .A2(n19922), .ZN(n13549) );
  NAND2_X1 U16880 ( .A1(n13550), .A2(n13549), .ZN(n16486) );
  NAND2_X1 U16881 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n13994) );
  NOR2_X1 U16882 ( .A1(n12955), .A2(n13994), .ZN(n16527) );
  INV_X1 U16883 ( .A(n16527), .ZN(n16526) );
  OAI22_X1 U16884 ( .A1(n16526), .A2(n13551), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n20033), .ZN(n13552) );
  AOI21_X1 U16885 ( .B1(n16486), .B2(n19927), .A(n13552), .ZN(n15883) );
  INV_X1 U16886 ( .A(n15883), .ZN(n13557) );
  INV_X1 U16887 ( .A(n10954), .ZN(n13554) );
  NAND3_X1 U16888 ( .A1(n13554), .A2(n11007), .A3(n13553), .ZN(n16498) );
  OR3_X1 U16889 ( .A1(n15883), .A2(n20006), .A3(n16498), .ZN(n13555) );
  OAI21_X1 U16890 ( .B1(n13557), .B2(n13556), .A(n13555), .ZN(P2_U3595) );
  INV_X1 U16891 ( .A(n13558), .ZN(n14561) );
  NOR2_X1 U16892 ( .A1(n13559), .A2(n14561), .ZN(n14568) );
  NAND2_X1 U16893 ( .A1(n14568), .A2(n14575), .ZN(n13563) );
  AND2_X1 U16894 ( .A1(n20689), .A2(n14021), .ZN(n13564) );
  NAND2_X1 U16895 ( .A1(n14567), .A2(n14575), .ZN(n13560) );
  INV_X1 U16896 ( .A(n13593), .ZN(n13561) );
  AOI211_X1 U16897 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n13563), .A(n13564), 
        .B(n13561), .ZN(n13562) );
  INV_X1 U16898 ( .A(n13562), .ZN(P1_U2801) );
  OAI21_X1 U16899 ( .B1(n13564), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n14040), 
        .ZN(n13565) );
  OAI21_X1 U16900 ( .B1(n13566), .B2(n14040), .A(n13565), .ZN(P1_U3487) );
  NAND2_X1 U16901 ( .A1(n13567), .A2(n19927), .ZN(n13570) );
  OR2_X1 U16902 ( .A1(n13568), .A2(n15068), .ZN(n13569) );
  OR2_X1 U16903 ( .A1(n19385), .A2(n13571), .ZN(n19350) );
  OR2_X1 U16904 ( .A1(n13994), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15074) );
  INV_X2 U16905 ( .A(n15074), .ZN(n19383) );
  AOI22_X1 U16906 ( .A1(P2_UWORD_REG_10__SCAN_IN), .A2(n19383), .B1(n19382), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13572) );
  OAI21_X1 U16907 ( .B1(n13573), .B2(n19350), .A(n13572), .ZN(P2_U2925) );
  INV_X1 U16908 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13575) );
  AOI22_X1 U16909 ( .A1(n19383), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13574) );
  OAI21_X1 U16910 ( .B1(n13575), .B2(n19350), .A(n13574), .ZN(P2_U2931) );
  INV_X1 U16911 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14334) );
  AOI22_X1 U16912 ( .A1(n19383), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13576) );
  OAI21_X1 U16913 ( .B1(n14334), .B2(n19350), .A(n13576), .ZN(P2_U2932) );
  INV_X1 U16914 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14503) );
  AOI22_X1 U16915 ( .A1(n19383), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13577) );
  OAI21_X1 U16916 ( .B1(n14503), .B2(n19350), .A(n13577), .ZN(P2_U2929) );
  INV_X1 U16917 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15283) );
  AOI22_X1 U16918 ( .A1(n19383), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13578) );
  OAI21_X1 U16919 ( .B1(n15283), .B2(n19350), .A(n13578), .ZN(P2_U2928) );
  INV_X1 U16920 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n21309) );
  AOI22_X1 U16921 ( .A1(n19383), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13579) );
  OAI21_X1 U16922 ( .B1(n21309), .B2(n19350), .A(n13579), .ZN(P2_U2934) );
  AOI22_X1 U16923 ( .A1(n19383), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13580) );
  OAI21_X1 U16924 ( .B1(n15268), .B2(n19350), .A(n13580), .ZN(P2_U2926) );
  INV_X1 U16925 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14488) );
  AOI22_X1 U16926 ( .A1(n19383), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13581) );
  OAI21_X1 U16927 ( .B1(n14488), .B2(n19350), .A(n13581), .ZN(P2_U2930) );
  AOI22_X1 U16928 ( .A1(n19383), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13582) );
  OAI21_X1 U16929 ( .B1(n15256), .B2(n19350), .A(n13582), .ZN(P2_U2924) );
  AOI22_X1 U16930 ( .A1(n19383), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13583) );
  OAI21_X1 U16931 ( .B1(n13584), .B2(n19350), .A(n13583), .ZN(P2_U2923) );
  INV_X1 U16932 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13586) );
  AOI22_X1 U16933 ( .A1(n19383), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13585) );
  OAI21_X1 U16934 ( .B1(n13586), .B2(n19350), .A(n13585), .ZN(P2_U2933) );
  AOI22_X1 U16935 ( .A1(n19383), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13587) );
  OAI21_X1 U16936 ( .B1(n15245), .B2(n19350), .A(n13587), .ZN(P2_U2922) );
  NAND2_X1 U16937 ( .A1(n11284), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13588) );
  AND4_X1 U16938 ( .A1(n10187), .A2(n13588), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20033), .ZN(n13589) );
  MUX2_X1 U16939 ( .A(n10643), .B(n10348), .S(n15229), .Z(n13590) );
  OAI21_X1 U16940 ( .B1(n20035), .B2(n15242), .A(n13590), .ZN(P2_U2887) );
  AND2_X1 U16941 ( .A1(n13591), .A2(n20924), .ZN(n13592) );
  NAND2_X1 U16942 ( .A1(n13688), .A2(n20257), .ZN(n13712) );
  INV_X1 U16943 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13597) );
  NAND2_X1 U16944 ( .A1(n13688), .A2(n14026), .ZN(n13689) );
  INV_X1 U16945 ( .A(DATAI_15_), .ZN(n13595) );
  INV_X1 U16946 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13594) );
  MUX2_X1 U16947 ( .A(n13595), .B(n13594), .S(n20239), .Z(n14438) );
  INV_X1 U16948 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13596) );
  OAI222_X1 U16949 ( .A1(n13712), .A2(n13597), .B1(n13689), .B2(n14438), .C1(
        n13596), .C2(n13688), .ZN(P1_U2967) );
  MUX2_X1 U16950 ( .A(n19251), .B(n15835), .S(n15229), .Z(n13602) );
  OAI21_X1 U16951 ( .B1(n14061), .B2(n15242), .A(n13602), .ZN(P2_U2886) );
  NOR2_X1 U16952 ( .A1(n13605), .A2(n13604), .ZN(n13606) );
  NOR2_X1 U16953 ( .A1(n13607), .A2(n13606), .ZN(n19267) );
  NAND2_X1 U16954 ( .A1(n19277), .A2(n19267), .ZN(n19341) );
  OAI211_X1 U16955 ( .C1(n19277), .C2(n19267), .A(n19341), .B(n19343), .ZN(
        n13609) );
  AOI22_X1 U16956 ( .A1(n19339), .A2(n19267), .B1(n19338), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13608) );
  OAI211_X1 U16957 ( .C1(n19347), .C2(n14075), .A(n13609), .B(n13608), .ZN(
        P2_U2919) );
  INV_X1 U16958 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19951) );
  AOI21_X1 U16959 ( .B1(n15833), .B2(n13611), .A(n13610), .ZN(n15838) );
  AOI21_X1 U16960 ( .B1(n13613), .B2(n19254), .A(n13612), .ZN(n13614) );
  XOR2_X1 U16961 ( .A(n13614), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n15837) );
  AOI22_X1 U16962 ( .A1(n19404), .A2(n15838), .B1(n19400), .B2(n15837), .ZN(
        n13615) );
  OAI21_X1 U16963 ( .B1(n19951), .B2(n19214), .A(n13615), .ZN(n13616) );
  AOI21_X1 U16964 ( .B1(n16442), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13616), .ZN(n13618) );
  NAND2_X1 U16965 ( .A1(n19398), .A2(n12933), .ZN(n13617) );
  OAI211_X1 U16966 ( .C1(n15835), .C2(n15509), .A(n13618), .B(n13617), .ZN(
        P2_U3013) );
  XNOR2_X1 U16967 ( .A(n19271), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16470) );
  INV_X1 U16968 ( .A(n16470), .ZN(n13626) );
  OAI21_X1 U16969 ( .B1(n13620), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13619), .ZN(n16475) );
  OAI21_X1 U16970 ( .B1(n16442), .B2(n13621), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13623) );
  INV_X1 U16971 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19073) );
  NOR2_X1 U16972 ( .A1(n19214), .A2(n19073), .ZN(n16478) );
  INV_X1 U16973 ( .A(n16478), .ZN(n13622) );
  OAI211_X1 U16974 ( .C1(n16436), .C2(n16475), .A(n13623), .B(n13622), .ZN(
        n13624) );
  AOI21_X1 U16975 ( .B1(n11289), .B2(n19403), .A(n13624), .ZN(n13625) );
  OAI21_X1 U16976 ( .B1(n16435), .B2(n13626), .A(n13625), .ZN(P2_U3014) );
  INV_X1 U16977 ( .A(n15667), .ZN(n13641) );
  OAI21_X1 U16978 ( .B1(n13627), .B2(n15831), .A(n16469), .ZN(n13628) );
  AOI21_X1 U16979 ( .B1(n13641), .B2(n15831), .A(n13628), .ZN(n13648) );
  NAND2_X1 U16980 ( .A1(n13630), .A2(n13629), .ZN(n13633) );
  INV_X1 U16981 ( .A(n13631), .ZN(n13632) );
  AND2_X1 U16982 ( .A1(n13633), .A2(n13632), .ZN(n14153) );
  AOI21_X1 U16983 ( .B1(n13636), .B2(n13635), .A(n13634), .ZN(n13656) );
  INV_X1 U16984 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19953) );
  NOR2_X1 U16985 ( .A1(n19214), .A2(n19953), .ZN(n13658) );
  AOI21_X1 U16986 ( .B1(n16461), .B2(n13656), .A(n13658), .ZN(n13637) );
  OAI21_X1 U16987 ( .B1(n14153), .B2(n16474), .A(n13637), .ZN(n13646) );
  XNOR2_X1 U16988 ( .A(n13639), .B(n13638), .ZN(n13663) );
  OAI22_X1 U16989 ( .A1(n13663), .A2(n15800), .B1(n13668), .B2(n15834), .ZN(
        n13645) );
  NAND3_X1 U16990 ( .A1(n13641), .A2(n13640), .A3(n9747), .ZN(n13642) );
  NAND2_X1 U16991 ( .A1(n13643), .A2(n13642), .ZN(n13644) );
  NOR3_X1 U16992 ( .A1(n13646), .A2(n13645), .A3(n13644), .ZN(n13647) );
  OAI21_X1 U16993 ( .B1(n9747), .B2(n13648), .A(n13647), .ZN(P2_U3044) );
  INV_X1 U16994 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13652) );
  NAND2_X1 U16995 ( .A1(n13868), .A2(n16051), .ZN(n13650) );
  NOR2_X1 U16996 ( .A1(n20057), .A2(n16073), .ZN(n13649) );
  NAND2_X1 U16997 ( .A1(n20154), .A2(n20243), .ZN(n13852) );
  NAND2_X1 U16998 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16383) );
  NOR2_X1 U16999 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16383), .ZN(n13850) );
  AOI22_X1 U17000 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20163), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n13850), .ZN(n13651) );
  OAI21_X1 U17001 ( .B1(n13652), .B2(n13852), .A(n13651), .ZN(P1_U2916) );
  INV_X1 U17002 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13654) );
  AOI22_X1 U17003 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20163), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n13850), .ZN(n13653) );
  OAI21_X1 U17004 ( .B1(n13654), .B2(n13852), .A(n13653), .ZN(P1_U2911) );
  AOI22_X1 U17005 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20163), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n13850), .ZN(n13655) );
  OAI21_X1 U17006 ( .B1(n14747), .B2(n13852), .A(n13655), .ZN(P1_U2912) );
  INV_X1 U17007 ( .A(n13656), .ZN(n13660) );
  NOR2_X1 U17008 ( .A1(n19409), .A2(n12934), .ZN(n13657) );
  AOI211_X1 U17009 ( .C1(n19398), .C2(n14151), .A(n13658), .B(n13657), .ZN(
        n13659) );
  OAI21_X1 U17010 ( .B1(n13660), .B2(n16436), .A(n13659), .ZN(n13661) );
  AOI21_X1 U17011 ( .B1(n19403), .B2(n11277), .A(n13661), .ZN(n13662) );
  OAI21_X1 U17012 ( .B1(n13663), .B2(n16435), .A(n13662), .ZN(P2_U3012) );
  MUX2_X1 U17013 ( .A(n13668), .B(n14154), .S(n13900), .Z(n13669) );
  OAI21_X1 U17014 ( .B1(n20020), .B2(n15242), .A(n13669), .ZN(P2_U2885) );
  INV_X1 U17015 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13671) );
  AOI22_X1 U17016 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n13850), .B1(n20163), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13670) );
  OAI21_X1 U17017 ( .B1(n13671), .B2(n13852), .A(n13670), .ZN(P1_U2908) );
  INV_X1 U17018 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13673) );
  AOI22_X1 U17019 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n13850), .B1(n20163), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13672) );
  OAI21_X1 U17020 ( .B1(n13673), .B2(n13852), .A(n13672), .ZN(P1_U2914) );
  INV_X1 U17021 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13675) );
  AOI22_X1 U17022 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n13850), .B1(n20163), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13674) );
  OAI21_X1 U17023 ( .B1(n13675), .B2(n13852), .A(n13674), .ZN(P1_U2909) );
  INV_X1 U17024 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U17025 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21019), .B1(n20163), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13676) );
  OAI21_X1 U17026 ( .B1(n13677), .B2(n13852), .A(n13676), .ZN(P1_U2906) );
  INV_X1 U17027 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13679) );
  AOI22_X1 U17028 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n13850), .B1(n20163), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13678) );
  OAI21_X1 U17029 ( .B1(n13679), .B2(n13852), .A(n13678), .ZN(P1_U2913) );
  OAI21_X1 U17030 ( .B1(n13681), .B2(n13680), .A(n13823), .ZN(n20225) );
  OAI21_X1 U17031 ( .B1(n13684), .B2(n13683), .A(n13682), .ZN(n13917) );
  INV_X1 U17032 ( .A(n13917), .ZN(n14105) );
  OAI22_X1 U17033 ( .A1(n14727), .A2(n14105), .B1(n13685), .B2(n20153), .ZN(
        n13686) );
  INV_X1 U17034 ( .A(n13686), .ZN(n13687) );
  OAI21_X1 U17035 ( .B1(n20225), .B2(n14728), .A(n13687), .ZN(P1_U2871) );
  INV_X1 U17036 ( .A(n13712), .ZN(n20187) );
  INV_X2 U17037 ( .A(n13688), .ZN(n20215) );
  AOI22_X1 U17038 ( .A1(n20187), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20215), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13693) );
  NAND2_X1 U17039 ( .A1(n20237), .A2(DATAI_7_), .ZN(n13691) );
  NAND2_X1 U17040 ( .A1(n20239), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13690) );
  AND2_X1 U17041 ( .A1(n13691), .A2(n13690), .ZN(n20291) );
  INV_X1 U17042 ( .A(n20291), .ZN(n13692) );
  NAND2_X1 U17043 ( .A1(n20201), .A2(n13692), .ZN(n13727) );
  NAND2_X1 U17044 ( .A1(n13693), .A2(n13727), .ZN(P1_U2959) );
  AOI22_X1 U17045 ( .A1(n20187), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20215), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13696) );
  NAND2_X1 U17046 ( .A1(n20237), .A2(DATAI_6_), .ZN(n13695) );
  NAND2_X1 U17047 ( .A1(n20239), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13694) );
  AND2_X1 U17048 ( .A1(n13695), .A2(n13694), .ZN(n20283) );
  INV_X1 U17049 ( .A(n20283), .ZN(n14758) );
  NAND2_X1 U17050 ( .A1(n20201), .A2(n14758), .ZN(n13733) );
  NAND2_X1 U17051 ( .A1(n13696), .A2(n13733), .ZN(P1_U2958) );
  AOI22_X1 U17052 ( .A1(n20187), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20215), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13700) );
  NAND2_X1 U17053 ( .A1(n20237), .A2(DATAI_5_), .ZN(n13698) );
  NAND2_X1 U17054 ( .A1(n20239), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13697) );
  AND2_X1 U17055 ( .A1(n13698), .A2(n13697), .ZN(n20277) );
  INV_X1 U17056 ( .A(n20277), .ZN(n13699) );
  NAND2_X1 U17057 ( .A1(n20201), .A2(n13699), .ZN(n13719) );
  NAND2_X1 U17058 ( .A1(n13700), .A2(n13719), .ZN(P1_U2957) );
  AOI22_X1 U17059 ( .A1(n20187), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20215), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13704) );
  NAND2_X1 U17060 ( .A1(n20237), .A2(DATAI_2_), .ZN(n13702) );
  NAND2_X1 U17061 ( .A1(n20239), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13701) );
  AND2_X1 U17062 ( .A1(n13702), .A2(n13701), .ZN(n20263) );
  INV_X1 U17063 ( .A(n20263), .ZN(n13703) );
  NAND2_X1 U17064 ( .A1(n20201), .A2(n13703), .ZN(n13731) );
  NAND2_X1 U17065 ( .A1(n13704), .A2(n13731), .ZN(P1_U2954) );
  AOI22_X1 U17066 ( .A1(n20187), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20215), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13707) );
  NAND2_X1 U17067 ( .A1(n20237), .A2(DATAI_4_), .ZN(n13706) );
  NAND2_X1 U17068 ( .A1(n20239), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13705) );
  AND2_X1 U17069 ( .A1(n13706), .A2(n13705), .ZN(n20272) );
  INV_X1 U17070 ( .A(n20272), .ZN(n14768) );
  NAND2_X1 U17071 ( .A1(n20201), .A2(n14768), .ZN(n13735) );
  NAND2_X1 U17072 ( .A1(n13707), .A2(n13735), .ZN(P1_U2956) );
  AOI22_X1 U17073 ( .A1(n20187), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20215), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13711) );
  NAND2_X1 U17074 ( .A1(n20237), .A2(DATAI_3_), .ZN(n13709) );
  NAND2_X1 U17075 ( .A1(n20239), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13708) );
  AND2_X1 U17076 ( .A1(n13709), .A2(n13708), .ZN(n20267) );
  INV_X1 U17077 ( .A(n20267), .ZN(n13710) );
  NAND2_X1 U17078 ( .A1(n20201), .A2(n13710), .ZN(n13713) );
  NAND2_X1 U17079 ( .A1(n13711), .A2(n13713), .ZN(P1_U2955) );
  AOI22_X1 U17080 ( .A1(n20216), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13714) );
  NAND2_X1 U17081 ( .A1(n13714), .A2(n13713), .ZN(P1_U2940) );
  AOI22_X1 U17082 ( .A1(n20216), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13718) );
  NAND2_X1 U17083 ( .A1(n20237), .A2(DATAI_0_), .ZN(n13716) );
  NAND2_X1 U17084 ( .A1(n20239), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13715) );
  AND2_X1 U17085 ( .A1(n13716), .A2(n13715), .ZN(n20250) );
  INV_X1 U17086 ( .A(n20250), .ZN(n13717) );
  NAND2_X1 U17087 ( .A1(n20201), .A2(n13717), .ZN(n13725) );
  NAND2_X1 U17088 ( .A1(n13718), .A2(n13725), .ZN(P1_U2937) );
  AOI22_X1 U17089 ( .A1(n20216), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U17090 ( .A1(n13720), .A2(n13719), .ZN(P1_U2942) );
  AOI22_X1 U17091 ( .A1(n20216), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20215), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13724) );
  NAND2_X1 U17092 ( .A1(n20237), .A2(DATAI_1_), .ZN(n13722) );
  NAND2_X1 U17093 ( .A1(n20239), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13721) );
  AND2_X1 U17094 ( .A1(n13722), .A2(n13721), .ZN(n20258) );
  INV_X1 U17095 ( .A(n20258), .ZN(n13723) );
  NAND2_X1 U17096 ( .A1(n20201), .A2(n13723), .ZN(n13729) );
  NAND2_X1 U17097 ( .A1(n13724), .A2(n13729), .ZN(P1_U2953) );
  AOI22_X1 U17098 ( .A1(n20216), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20215), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13726) );
  NAND2_X1 U17099 ( .A1(n13726), .A2(n13725), .ZN(P1_U2952) );
  AOI22_X1 U17100 ( .A1(n20216), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13728) );
  NAND2_X1 U17101 ( .A1(n13728), .A2(n13727), .ZN(P1_U2944) );
  AOI22_X1 U17102 ( .A1(n20216), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13730) );
  NAND2_X1 U17103 ( .A1(n13730), .A2(n13729), .ZN(P1_U2938) );
  AOI22_X1 U17104 ( .A1(n20216), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13732) );
  NAND2_X1 U17105 ( .A1(n13732), .A2(n13731), .ZN(P1_U2939) );
  AOI22_X1 U17106 ( .A1(n20216), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13734) );
  NAND2_X1 U17107 ( .A1(n13734), .A2(n13733), .ZN(P1_U2943) );
  AOI22_X1 U17108 ( .A1(n20216), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13736) );
  NAND2_X1 U17109 ( .A1(n13736), .A2(n13735), .ZN(P1_U2941) );
  INV_X1 U17110 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n14141) );
  NOR2_X1 U17111 ( .A1(n15229), .A2(n14141), .ZN(n13740) );
  AOI21_X1 U17112 ( .B1(n10334), .B2(n15229), .A(n13740), .ZN(n13741) );
  OAI21_X1 U17113 ( .B1(n19503), .B2(n15242), .A(n13741), .ZN(P2_U2884) );
  INV_X1 U17114 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20726) );
  AOI21_X1 U17115 ( .B1(n15044), .B2(n21244), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13742) );
  NOR2_X1 U17116 ( .A1(n12986), .A2(n13742), .ZN(n13763) );
  OR2_X1 U17117 ( .A1(n13744), .A2(n12143), .ZN(n13747) );
  NAND2_X1 U17118 ( .A1(n13768), .A2(n13745), .ZN(n13746) );
  AOI21_X1 U17119 ( .B1(n13747), .B2(n14023), .A(n13746), .ZN(n13750) );
  INV_X1 U17120 ( .A(n13748), .ZN(n13749) );
  AND3_X1 U17121 ( .A1(n12204), .A2(n13750), .A3(n13749), .ZN(n15050) );
  INV_X1 U17122 ( .A(n15050), .ZN(n13866) );
  NAND2_X1 U17123 ( .A1(n20563), .A2(n13866), .ZN(n13762) );
  AND2_X1 U17124 ( .A1(n13769), .A2(n13751), .ZN(n13864) );
  MUX2_X1 U17125 ( .A(n13755), .B(n13752), .S(n15044), .Z(n13754) );
  NOR2_X1 U17126 ( .A1(n13754), .A2(n13753), .ZN(n13757) );
  AOI21_X1 U17127 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13753), .A(
        n13755), .ZN(n13756) );
  OAI22_X1 U17128 ( .A1(n13864), .A2(n13757), .B1(n13756), .B2(n13868), .ZN(
        n13758) );
  INV_X1 U17129 ( .A(n13758), .ZN(n13761) );
  NAND3_X1 U17130 ( .A1(n15050), .A2(n13863), .A3(n13763), .ZN(n13760) );
  NOR2_X1 U17131 ( .A1(n13868), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15046) );
  NAND2_X1 U17132 ( .A1(n15046), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13759) );
  NAND4_X1 U17133 ( .A1(n13762), .A2(n13761), .A3(n13760), .A4(n13759), .ZN(
        n13859) );
  AOI22_X1 U17134 ( .A1(n16058), .A2(n13763), .B1(n15060), .B2(n13859), .ZN(
        n13776) );
  NAND2_X1 U17135 ( .A1(n14025), .A2(n14026), .ZN(n14039) );
  OR2_X1 U17136 ( .A1(n14039), .A2(n20261), .ZN(n13764) );
  AND4_X1 U17137 ( .A1(n13767), .A2(n13766), .A3(n13765), .A4(n13764), .ZN(
        n13774) );
  NOR2_X1 U17138 ( .A1(n16073), .A2(n20924), .ZN(n13771) );
  NAND3_X1 U17139 ( .A1(n13769), .A2(n13768), .A3(n13868), .ZN(n13770) );
  OAI211_X1 U17140 ( .C1(n13772), .C2(n13771), .A(n14565), .B(n13770), .ZN(
        n13773) );
  INV_X1 U17141 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20063) );
  INV_X1 U17142 ( .A(n16383), .ZN(n16379) );
  NAND2_X1 U17143 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16379), .ZN(n13885) );
  OAI22_X1 U17144 ( .A1(n13879), .A2(n20057), .B1(n20063), .B2(n13885), .ZN(
        n13779) );
  AOI21_X1 U17145 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n11887), .A(n13779), 
        .ZN(n15065) );
  NAND2_X1 U17146 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n15065), .ZN(
        n13775) );
  OAI21_X1 U17147 ( .B1(n13776), .B2(n15065), .A(n13775), .ZN(P1_U3469) );
  INV_X1 U17148 ( .A(n20406), .ZN(n20724) );
  OR2_X1 U17149 ( .A1(n11969), .A2(n20724), .ZN(n13777) );
  XNOR2_X1 U17150 ( .A(n13777), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14056) );
  NAND2_X1 U17151 ( .A1(n14056), .A2(n13778), .ZN(n13877) );
  NAND2_X1 U17152 ( .A1(n15060), .A2(n13779), .ZN(n13781) );
  INV_X1 U17153 ( .A(n15065), .ZN(n13780) );
  OAI22_X1 U17154 ( .A1(n13877), .A2(n13781), .B1(n13878), .B2(n13780), .ZN(
        P1_U3468) );
  INV_X1 U17155 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13782) );
  NOR2_X1 U17156 ( .A1(n13783), .A2(n13782), .ZN(n13786) );
  INV_X1 U17157 ( .A(n13786), .ZN(n13784) );
  NAND2_X1 U17158 ( .A1(n13785), .A2(n13784), .ZN(n13788) );
  NAND2_X1 U17159 ( .A1(n13787), .A2(n13786), .ZN(n13902) );
  OAI21_X1 U17160 ( .B1(n13789), .B2(n13788), .A(n13902), .ZN(n19325) );
  OR2_X1 U17161 ( .A1(n13791), .A2(n13790), .ZN(n13792) );
  AND2_X1 U17162 ( .A1(n13792), .A2(n13809), .ZN(n19402) );
  NOR2_X1 U17163 ( .A1(n15229), .A2(n13793), .ZN(n13794) );
  AOI21_X1 U17164 ( .B1(n19402), .B2(n15229), .A(n13794), .ZN(n13795) );
  OAI21_X1 U17165 ( .B1(n19325), .B2(n15242), .A(n13795), .ZN(P2_U2883) );
  AOI22_X1 U17166 ( .A1(n20372), .A2(n13866), .B1(n15048), .B2(n12426), .ZN(
        n16022) );
  INV_X1 U17167 ( .A(n15060), .ZN(n13796) );
  OAI22_X1 U17168 ( .A1(n16022), .A2(n13796), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14021), .ZN(n13797) );
  AOI21_X1 U17169 ( .B1(n16058), .B2(n12426), .A(n13797), .ZN(n13799) );
  NOR2_X1 U17170 ( .A1(n13868), .A2(n12426), .ZN(n16029) );
  AOI22_X1 U17171 ( .A1(n16029), .A2(n15060), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15065), .ZN(n13798) );
  OAI21_X1 U17172 ( .B1(n13799), .B2(n15065), .A(n13798), .ZN(P1_U3474) );
  INV_X1 U17173 ( .A(n13800), .ZN(n13803) );
  OAI21_X1 U17174 ( .B1(n13803), .B2(n13802), .A(n13801), .ZN(n20235) );
  OR2_X1 U17175 ( .A1(n13804), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13806) );
  AND2_X1 U17176 ( .A1(n13806), .A2(n13805), .ZN(n14036) );
  INV_X1 U17177 ( .A(n14036), .ZN(n13807) );
  OAI222_X1 U17178 ( .A1(n20235), .A2(n14728), .B1(n14034), .B2(n20153), .C1(
        n13807), .C2(n14727), .ZN(P1_U2872) );
  INV_X1 U17179 ( .A(n13902), .ZN(n13904) );
  XNOR2_X1 U17180 ( .A(n13904), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13813) );
  AOI21_X1 U17181 ( .B1(n13810), .B2(n13809), .A(n13808), .ZN(n19245) );
  INV_X1 U17182 ( .A(n19245), .ZN(n14346) );
  NOR2_X1 U17183 ( .A1(n14346), .A2(n13900), .ZN(n13811) );
  AOI21_X1 U17184 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n13900), .A(n13811), .ZN(
        n13812) );
  OAI21_X1 U17185 ( .B1(n13813), .B2(n15242), .A(n13812), .ZN(P2_U2882) );
  OAI21_X1 U17186 ( .B1(n13815), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13814), .ZN(n20226) );
  AOI21_X1 U17187 ( .B1(n13958), .B2(n15051), .A(n15012), .ZN(n13816) );
  INV_X1 U17188 ( .A(n13816), .ZN(n13914) );
  OAI22_X1 U17189 ( .A1(n13914), .A2(n13818), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13817), .ZN(n13820) );
  AOI22_X1 U17190 ( .A1(n16367), .A2(n14036), .B1(n20232), .B2(
        P1_REIP_REG_0__SCAN_IN), .ZN(n13819) );
  OAI211_X1 U17191 ( .C1(n16370), .C2(n20226), .A(n13820), .B(n13819), .ZN(
        P1_U3031) );
  NAND2_X1 U17192 ( .A1(n12189), .A2(n20286), .ZN(n13821) );
  NAND2_X2 U17193 ( .A1(n14748), .A2(n13821), .ZN(n14785) );
  INV_X1 U17194 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20176) );
  OAI222_X1 U17195 ( .A1(n14785), .A2(n20225), .B1(n14748), .B2(n20176), .C1(
        n14439), .C2(n20258), .ZN(P1_U2903) );
  INV_X1 U17196 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20180) );
  OAI222_X1 U17197 ( .A1(n14785), .A2(n20235), .B1(n14748), .B2(n20180), .C1(
        n14439), .C2(n20250), .ZN(P1_U2904) );
  NAND2_X1 U17198 ( .A1(n13822), .A2(n13823), .ZN(n13824) );
  AND2_X1 U17199 ( .A1(n13825), .A2(n13824), .ZN(n20137) );
  INV_X1 U17200 ( .A(n20137), .ZN(n13826) );
  INV_X1 U17201 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20174) );
  OAI222_X1 U17202 ( .A1(n14785), .A2(n13826), .B1(n14748), .B2(n20174), .C1(
        n14439), .C2(n20263), .ZN(P1_U2902) );
  XNOR2_X1 U17203 ( .A(n14275), .B(n14153), .ZN(n13832) );
  XNOR2_X1 U17204 ( .A(n13828), .B(n13827), .ZN(n20030) );
  NOR2_X1 U17205 ( .A1(n20026), .A2(n20030), .ZN(n13829) );
  AOI21_X1 U17206 ( .B1(n20030), .B2(n20026), .A(n13829), .ZN(n19342) );
  NAND2_X1 U17207 ( .A1(n19342), .A2(n19341), .ZN(n19340) );
  INV_X1 U17208 ( .A(n13829), .ZN(n13830) );
  NAND2_X1 U17209 ( .A1(n19340), .A2(n13830), .ZN(n13831) );
  NAND2_X1 U17210 ( .A1(n13831), .A2(n13832), .ZN(n14114) );
  OAI21_X1 U17211 ( .B1(n13832), .B2(n13831), .A(n14114), .ZN(n13833) );
  NAND2_X1 U17212 ( .A1(n13833), .A2(n19343), .ZN(n13835) );
  INV_X1 U17213 ( .A(n19422), .ZN(n16417) );
  AOI22_X1 U17214 ( .A1(n19314), .A2(n16417), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19338), .ZN(n13834) );
  OAI211_X1 U17215 ( .C1(n14153), .C2(n19297), .A(n13835), .B(n13834), .ZN(
        P2_U2917) );
  OAI21_X1 U17216 ( .B1(n13838), .B2(n13837), .A(n13836), .ZN(n14517) );
  INV_X1 U17217 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20172) );
  OAI222_X1 U17218 ( .A1(n14785), .A2(n14517), .B1(n14748), .B2(n20172), .C1(
        n14439), .C2(n20267), .ZN(P1_U2901) );
  INV_X1 U17219 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13840) );
  AOI22_X1 U17220 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n13850), .B1(n20177), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13839) );
  OAI21_X1 U17221 ( .B1(n13840), .B2(n13852), .A(n13839), .ZN(P1_U2917) );
  INV_X1 U17222 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13842) );
  AOI22_X1 U17223 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13841) );
  OAI21_X1 U17224 ( .B1(n13842), .B2(n13852), .A(n13841), .ZN(P1_U2919) );
  INV_X1 U17225 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17226 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n13850), .B1(n20177), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13843) );
  OAI21_X1 U17227 ( .B1(n13844), .B2(n13852), .A(n13843), .ZN(P1_U2907) );
  INV_X1 U17228 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U17229 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13845) );
  OAI21_X1 U17230 ( .B1(n13846), .B2(n13852), .A(n13845), .ZN(P1_U2920) );
  INV_X1 U17231 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13848) );
  AOI22_X1 U17232 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n13850), .B1(n20177), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13847) );
  OAI21_X1 U17233 ( .B1(n13848), .B2(n13852), .A(n13847), .ZN(P1_U2915) );
  INV_X1 U17234 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14779) );
  AOI22_X1 U17235 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13849) );
  OAI21_X1 U17236 ( .B1(n14779), .B2(n13852), .A(n13849), .ZN(P1_U2918) );
  INV_X1 U17237 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U17238 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n13850), .B1(n20177), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13851) );
  OAI21_X1 U17239 ( .B1(n13853), .B2(n13852), .A(n13851), .ZN(P1_U2910) );
  OAI211_X1 U17240 ( .C1(n11318), .C2(n11317), .A(n15235), .B(n13978), .ZN(
        n13858) );
  NAND2_X1 U17241 ( .A1(n9834), .A2(n13920), .ZN(n13856) );
  AND2_X1 U17242 ( .A1(n13856), .A2(n13976), .ZN(n16439) );
  NAND2_X1 U17243 ( .A1(n16439), .A2(n15229), .ZN(n13857) );
  OAI211_X1 U17244 ( .C1(n15229), .C2(n10685), .A(n13858), .B(n13857), .ZN(
        P2_U2878) );
  NOR2_X1 U17245 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n14021), .ZN(n13882) );
  MUX2_X1 U17246 ( .A(n13859), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13879), .Z(n16035) );
  AOI22_X1 U17247 ( .A1(n13882), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n14021), .B2(n16035), .ZN(n13875) );
  OR2_X1 U17248 ( .A1(n13861), .A2(n15050), .ZN(n13873) );
  XNOR2_X1 U17249 ( .A(n15044), .B(n13862), .ZN(n15056) );
  NAND2_X1 U17250 ( .A1(n13863), .A2(n15056), .ZN(n13865) );
  OAI22_X1 U17251 ( .A1(n13866), .A2(n13865), .B1(n13864), .B2(n15056), .ZN(
        n13871) );
  NOR2_X1 U17252 ( .A1(n13868), .A2(n13867), .ZN(n13869) );
  MUX2_X1 U17253 ( .A(n13869), .B(n15046), .S(n21244), .Z(n13870) );
  NOR2_X1 U17254 ( .A1(n13871), .A2(n13870), .ZN(n13872) );
  NAND2_X1 U17255 ( .A1(n13873), .A2(n13872), .ZN(n15061) );
  INV_X1 U17256 ( .A(n13879), .ZN(n16023) );
  MUX2_X1 U17257 ( .A(n21244), .B(n15061), .S(n16023), .Z(n16030) );
  AOI22_X1 U17258 ( .A1(n16030), .A2(n14021), .B1(n21244), .B2(n13882), .ZN(
        n13874) );
  NOR2_X1 U17259 ( .A1(n13875), .A2(n13874), .ZN(n16041) );
  INV_X1 U17260 ( .A(n15045), .ZN(n13876) );
  NAND2_X1 U17261 ( .A1(n16041), .A2(n13876), .ZN(n13908) );
  NAND2_X1 U17262 ( .A1(n13877), .A2(n16023), .ZN(n13881) );
  AOI21_X1 U17263 ( .B1(n13879), .B2(n13878), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13880) );
  NAND2_X1 U17264 ( .A1(n13881), .A2(n13880), .ZN(n13884) );
  NAND2_X1 U17265 ( .A1(n13882), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13883) );
  AND2_X1 U17266 ( .A1(n16043), .A2(n20063), .ZN(n13886) );
  AOI21_X1 U17267 ( .B1(n13908), .B2(n13886), .A(n13885), .ZN(n13888) );
  NAND2_X1 U17268 ( .A1(n21011), .A2(n14021), .ZN(n21014) );
  INV_X1 U17269 ( .A(n21014), .ZN(n16059) );
  INV_X1 U17270 ( .A(n20412), .ZN(n13887) );
  NOR2_X1 U17271 ( .A1(n14021), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20994) );
  NOR2_X1 U17272 ( .A1(n13861), .A2(n20994), .ZN(n13892) );
  AOI21_X1 U17273 ( .B1(n13889), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20760), 
        .ZN(n20685) );
  NAND2_X1 U17274 ( .A1(n13889), .A2(n20689), .ZN(n20991) );
  NOR2_X1 U17275 ( .A1(n20991), .A2(n21012), .ZN(n13890) );
  MUX2_X1 U17276 ( .A(n20685), .B(n13890), .S(n12414), .Z(n13891) );
  OAI21_X1 U17277 ( .B1(n13892), .B2(n13891), .A(n20996), .ZN(n13893) );
  OAI21_X1 U17278 ( .B1(n20996), .B2(n20562), .A(n13893), .ZN(P1_U3476) );
  INV_X1 U17279 ( .A(n13894), .ZN(n13899) );
  INV_X1 U17280 ( .A(n13895), .ZN(n13897) );
  INV_X1 U17281 ( .A(n13808), .ZN(n13896) );
  NAND2_X1 U17282 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  NAND2_X1 U17283 ( .A1(n13899), .A2(n13898), .ZN(n19229) );
  NOR2_X1 U17284 ( .A1(n13902), .A2(n13901), .ZN(n13905) );
  NAND2_X1 U17285 ( .A1(n13904), .A2(n13903), .ZN(n13927) );
  OAI211_X1 U17286 ( .C1(n13905), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15235), .B(n13927), .ZN(n13907) );
  NAND2_X1 U17287 ( .A1(n13900), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13906) );
  OAI211_X1 U17288 ( .C1(n19229), .C2(n13900), .A(n13907), .B(n13906), .ZN(
        P2_U2881) );
  AND3_X1 U17289 ( .A1(n13908), .A2(n16043), .A3(n16379), .ZN(n16052) );
  INV_X1 U17290 ( .A(n20372), .ZN(n13909) );
  OAI22_X1 U17291 ( .A1(n12423), .A2(n20760), .B1(n13909), .B2(n20994), .ZN(
        n13910) );
  OAI21_X1 U17292 ( .B1(n16052), .B2(n13910), .A(n20996), .ZN(n13911) );
  OAI21_X1 U17293 ( .B1(n20996), .B2(n20759), .A(n13911), .ZN(P1_U3478) );
  XNOR2_X1 U17294 ( .A(n13912), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20221) );
  NOR2_X1 U17295 ( .A1(n14979), .A2(n13913), .ZN(n13915) );
  MUX2_X1 U17296 ( .A(n13915), .B(n13914), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n13916) );
  INV_X1 U17297 ( .A(n13916), .ZN(n13919) );
  INV_X1 U17298 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21000) );
  NOR2_X1 U17299 ( .A1(n20100), .A2(n21000), .ZN(n20223) );
  AOI21_X1 U17300 ( .B1(n16367), .B2(n13917), .A(n20223), .ZN(n13918) );
  OAI211_X1 U17301 ( .C1(n20221), .C2(n16370), .A(n13919), .B(n13918), .ZN(
        P1_U3030) );
  OAI21_X1 U17302 ( .B1(n13928), .B2(n13921), .A(n13920), .ZN(n14268) );
  INV_X1 U17303 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13923) );
  OAI21_X1 U17304 ( .B1(n13927), .B2(n13923), .A(n13922), .ZN(n13924) );
  NAND3_X1 U17305 ( .A1(n13924), .A2(n15235), .A3(n13854), .ZN(n13926) );
  NAND2_X1 U17306 ( .A1(n13900), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13925) );
  OAI211_X1 U17307 ( .C1(n14268), .C2(n13900), .A(n13926), .B(n13925), .ZN(
        P2_U2879) );
  XOR2_X1 U17308 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13927), .Z(n13932)
         );
  INV_X1 U17309 ( .A(n13928), .ZN(n13929) );
  OAI21_X1 U17310 ( .B1(n13894), .B2(n13930), .A(n13929), .ZN(n19217) );
  INV_X1 U17311 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n19216) );
  MUX2_X1 U17312 ( .A(n19217), .B(n19216), .S(n13900), .Z(n13931) );
  OAI21_X1 U17313 ( .B1(n13932), .B2(n15242), .A(n13931), .ZN(P2_U2880) );
  OAI21_X1 U17314 ( .B1(n13934), .B2(n13936), .A(n13935), .ZN(n16251) );
  NAND2_X1 U17315 ( .A1(n13964), .A2(n13937), .ZN(n13938) );
  AND2_X1 U17316 ( .A1(n14090), .A2(n13938), .ZN(n20104) );
  AOI22_X1 U17317 ( .A1(n20104), .A2(n20148), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14707), .ZN(n13939) );
  OAI21_X1 U17318 ( .B1(n16251), .B2(n14728), .A(n13939), .ZN(P1_U2867) );
  XNOR2_X1 U17319 ( .A(n13940), .B(n13941), .ZN(n13993) );
  INV_X1 U17320 ( .A(n14517), .ZN(n20120) );
  INV_X1 U17321 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13943) );
  NOR2_X1 U17322 ( .A1(n20100), .A2(n13943), .ZN(n13990) );
  AOI21_X1 U17323 ( .B1(n20228), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13990), .ZN(n13944) );
  OAI21_X1 U17324 ( .B1(n20219), .B2(n20114), .A(n13944), .ZN(n13945) );
  AOI21_X1 U17325 ( .B1(n20120), .B2(n13942), .A(n13945), .ZN(n13946) );
  OAI21_X1 U17326 ( .B1(n13993), .B2(n20220), .A(n13946), .ZN(P1_U2996) );
  XNOR2_X1 U17327 ( .A(n13948), .B(n13947), .ZN(n14521) );
  INV_X1 U17328 ( .A(n15016), .ZN(n16339) );
  NOR2_X1 U17329 ( .A1(n12212), .A2(n16339), .ZN(n13949) );
  AOI21_X1 U17330 ( .B1(n16338), .B2(n13984), .A(n15012), .ZN(n15026) );
  INV_X1 U17331 ( .A(n15026), .ZN(n16335) );
  MUX2_X1 U17332 ( .A(n13949), .B(n16335), .S(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n13950) );
  INV_X1 U17333 ( .A(n13950), .ZN(n13960) );
  NAND2_X1 U17334 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13952) );
  OAI21_X1 U17335 ( .B1(n13952), .B2(n13951), .A(n13985), .ZN(n13957) );
  NAND2_X1 U17336 ( .A1(n13954), .A2(n13953), .ZN(n13955) );
  NAND2_X1 U17337 ( .A1(n13988), .A2(n13955), .ZN(n20125) );
  INV_X1 U17338 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20138) );
  OAI22_X1 U17339 ( .A1(n16341), .A2(n20125), .B1(n20138), .B2(n20100), .ZN(
        n13956) );
  AOI21_X1 U17340 ( .B1(n13958), .B2(n13957), .A(n13956), .ZN(n13959) );
  OAI211_X1 U17341 ( .C1(n16370), .C2(n14521), .A(n13960), .B(n13959), .ZN(
        P1_U3029) );
  AOI21_X1 U17342 ( .B1(n13961), .B2(n13836), .A(n13934), .ZN(n13983) );
  INV_X1 U17343 ( .A(n14728), .ZN(n20149) );
  OR2_X1 U17344 ( .A1(n13987), .A2(n13962), .ZN(n13963) );
  NAND2_X1 U17345 ( .A1(n13964), .A2(n13963), .ZN(n14186) );
  OAI22_X1 U17346 ( .A1(n14186), .A2(n14727), .B1(n14054), .B2(n20153), .ZN(
        n13965) );
  AOI21_X1 U17347 ( .B1(n13983), .B2(n20149), .A(n13965), .ZN(n13966) );
  INV_X1 U17348 ( .A(n13966), .ZN(P1_U2868) );
  INV_X1 U17349 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20168) );
  OAI222_X1 U17350 ( .A1(n14785), .A2(n16251), .B1(n14748), .B2(n20168), .C1(
        n14439), .C2(n20277), .ZN(P1_U2899) );
  NAND2_X1 U17351 ( .A1(n9805), .A2(n13967), .ZN(n14046) );
  OAI211_X1 U17352 ( .C1(n9805), .C2(n13967), .A(n14046), .B(n15235), .ZN(
        n13973) );
  OR2_X1 U17353 ( .A1(n13969), .A2(n13970), .ZN(n13971) );
  NAND2_X1 U17354 ( .A1(n13968), .A2(n13971), .ZN(n19179) );
  INV_X1 U17355 ( .A(n19179), .ZN(n15754) );
  NAND2_X1 U17356 ( .A1(n15754), .A2(n15229), .ZN(n13972) );
  OAI211_X1 U17357 ( .C1(n15229), .C2(n13974), .A(n13973), .B(n13972), .ZN(
        P2_U2876) );
  AND2_X1 U17358 ( .A1(n13976), .A2(n13975), .ZN(n13977) );
  OR2_X1 U17359 ( .A1(n13977), .A2(n13969), .ZN(n19193) );
  INV_X1 U17360 ( .A(n19193), .ZN(n16430) );
  NOR2_X1 U17361 ( .A1(n15229), .A2(n19192), .ZN(n13981) );
  AOI211_X1 U17362 ( .C1(n13979), .C2(n13978), .A(n15242), .B(n9805), .ZN(
        n13980) );
  AOI211_X1 U17363 ( .C1(n16430), .C2(n15229), .A(n13981), .B(n13980), .ZN(
        n13982) );
  INV_X1 U17364 ( .A(n13982), .ZN(P2_U2877) );
  INV_X1 U17365 ( .A(n13983), .ZN(n14086) );
  INV_X1 U17366 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20170) );
  OAI222_X1 U17367 ( .A1(n14086), .A2(n14785), .B1(n20170), .B2(n14748), .C1(
        n14439), .C2(n20272), .ZN(P1_U2900) );
  OAI21_X1 U17368 ( .B1(n16333), .B2(n13985), .A(n15026), .ZN(n14183) );
  OAI21_X1 U17369 ( .B1(n13984), .B2(n16339), .A(n16333), .ZN(n16316) );
  NAND2_X1 U17370 ( .A1(n13985), .A2(n16316), .ZN(n16374) );
  INV_X1 U17371 ( .A(n16374), .ZN(n13986) );
  AOI22_X1 U17372 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14183), .B1(
        n13986), .B2(n14187), .ZN(n13992) );
  AOI21_X1 U17373 ( .B1(n13989), .B2(n13988), .A(n13987), .ZN(n20113) );
  AOI21_X1 U17374 ( .B1(n20113), .B2(n16367), .A(n13990), .ZN(n13991) );
  OAI211_X1 U17375 ( .C1(n16370), .C2(n13993), .A(n13992), .B(n13991), .ZN(
        P1_U3028) );
  NAND3_X1 U17376 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20032), .ZN(n19760) );
  NOR2_X1 U17377 ( .A1(n20040), .A2(n19760), .ZN(n19805) );
  NAND2_X1 U17378 ( .A1(n19921), .A2(n19763), .ZN(n19055) );
  NAND2_X1 U17379 ( .A1(n19055), .A2(n13994), .ZN(n13995) );
  INV_X1 U17380 ( .A(n19503), .ZN(n20011) );
  NAND2_X1 U17381 ( .A1(n20011), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19847) );
  OAI21_X1 U17382 ( .B1(n19550), .B2(n19847), .A(n19760), .ZN(n13996) );
  OAI211_X1 U17383 ( .C1(n19805), .C2(n20033), .A(n19851), .B(n13996), .ZN(
        n13997) );
  INV_X1 U17384 ( .A(n13997), .ZN(n14000) );
  NOR2_X1 U17385 ( .A1(n13998), .A2(n19805), .ZN(n14003) );
  NAND2_X1 U17386 ( .A1(n14003), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13999) );
  NAND2_X1 U17387 ( .A1(n14000), .A2(n13999), .ZN(n19798) );
  INV_X1 U17388 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U17389 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19433), .ZN(n19758) );
  NOR2_X2 U17390 ( .A1(n19730), .A2(n19550), .ZN(n19832) );
  AOI22_X1 U17391 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19433), .ZN(n19920) );
  INV_X1 U17392 ( .A(n19920), .ZN(n19831) );
  AOI22_X1 U17393 ( .A1(n19807), .A2(n19914), .B1(n19832), .B2(n19831), .ZN(
        n14005) );
  OAI22_X1 U17394 ( .A1(n14003), .A2(n19763), .B1(n19760), .B2(n20013), .ZN(
        n19806) );
  NOR2_X2 U17395 ( .A1(n19318), .A2(n19765), .ZN(n19907) );
  NAND2_X1 U17396 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19851), .ZN(n14010) );
  AOI22_X1 U17397 ( .A1(n19806), .A2(n19907), .B1(n19805), .B2(n19908), .ZN(
        n14004) );
  OAI211_X1 U17398 ( .C1(n19810), .C2(n14006), .A(n14005), .B(n14004), .ZN(
        P2_U3159) );
  AOI22_X1 U17399 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19433), .ZN(n19736) );
  AOI22_X1 U17400 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19433), .ZN(n19866) );
  AOI22_X1 U17401 ( .A1(n19807), .A2(n19863), .B1(n19832), .B2(n19811), .ZN(
        n14008) );
  NOR2_X2 U17402 ( .A1(n19348), .A2(n19765), .ZN(n19858) );
  AOI22_X1 U17403 ( .A1(n19806), .A2(n19858), .B1(n19859), .B2(n19805), .ZN(
        n14007) );
  OAI211_X1 U17404 ( .C1(n19810), .C2(n14009), .A(n14008), .B(n14007), .ZN(
        P2_U3153) );
  INV_X1 U17405 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14013) );
  AOI22_X1 U17406 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19433), .ZN(n19906) );
  INV_X1 U17407 ( .A(n19906), .ZN(n19748) );
  AOI22_X1 U17408 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19433), .ZN(n19751) );
  AOI22_X1 U17409 ( .A1(n19832), .A2(n19748), .B1(n19807), .B2(n19903), .ZN(
        n14012) );
  NOR2_X2 U17410 ( .A1(n19320), .A2(n19765), .ZN(n19782) );
  AOI22_X1 U17411 ( .A1(n19806), .A2(n19782), .B1(n19805), .B2(n9707), .ZN(
        n14011) );
  OAI211_X1 U17412 ( .C1(n19810), .C2(n14013), .A(n14012), .B(n14011), .ZN(
        P2_U3158) );
  NAND2_X1 U17413 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16059), .ZN(n16055) );
  NAND2_X1 U17414 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n11887), .ZN(n14014) );
  OAI21_X1 U17415 ( .B1(n14014), .B2(n12409), .A(n20100), .ZN(n14015) );
  INV_X1 U17416 ( .A(n14015), .ZN(n14016) );
  OAI21_X1 U17417 ( .B1(n16055), .B2(n11887), .A(n14016), .ZN(n14017) );
  NAND2_X1 U17418 ( .A1(n14018), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14020) );
  INV_X1 U17419 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14019) );
  XNOR2_X1 U17420 ( .A(n14020), .B(n14019), .ZN(n14512) );
  NOR2_X1 U17421 ( .A1(n14512), .A2(n14021), .ZN(n14022) );
  NAND2_X1 U17422 ( .A1(n21016), .A2(n14023), .ZN(n14024) );
  NAND2_X1 U17423 ( .A1(n16182), .A2(n14024), .ZN(n20136) );
  INV_X1 U17424 ( .A(n20136), .ZN(n14109) );
  NAND2_X1 U17425 ( .A1(n14026), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14029) );
  AND2_X1 U17426 ( .A1(n21018), .A2(n21012), .ZN(n16045) );
  NOR2_X1 U17427 ( .A1(n14029), .A2(n16045), .ZN(n14027) );
  AND2_X1 U17428 ( .A1(n14028), .A2(n16045), .ZN(n14037) );
  INV_X1 U17429 ( .A(n14029), .ZN(n14030) );
  NOR2_X1 U17430 ( .A1(n14037), .A2(n14030), .ZN(n14031) );
  AND2_X1 U17431 ( .A1(n14512), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14032) );
  OAI21_X1 U17432 ( .B1(n20128), .B2(n20131), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14033) );
  OAI21_X1 U17433 ( .B1(n20095), .B2(n14034), .A(n14033), .ZN(n14035) );
  AOI21_X1 U17434 ( .B1(n20127), .B2(n14036), .A(n14035), .ZN(n14042) );
  NAND2_X1 U17435 ( .A1(n20118), .A2(n20116), .ZN(n16166) );
  NOR2_X1 U17436 ( .A1(n14040), .A2(n14039), .ZN(n20129) );
  AOI22_X1 U17437 ( .A1(n16166), .A2(P1_REIP_REG_0__SCAN_IN), .B1(n20372), 
        .B2(n20129), .ZN(n14041) );
  OAI211_X1 U17438 ( .C1(n20235), .C2(n14109), .A(n14042), .B(n14041), .ZN(
        P1_U2840) );
  AOI21_X1 U17439 ( .B1(n14044), .B2(n13968), .A(n14043), .ZN(n15740) );
  INV_X1 U17440 ( .A(n15740), .ZN(n19169) );
  INV_X1 U17441 ( .A(n14046), .ZN(n14220) );
  INV_X1 U17442 ( .A(n14045), .ZN(n14047) );
  OAI211_X1 U17443 ( .C1(n14220), .C2(n14047), .A(n15235), .B(n14248), .ZN(
        n14049) );
  NAND2_X1 U17444 ( .A1(n13900), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14048) );
  OAI211_X1 U17445 ( .C1(n19169), .C2(n13900), .A(n14049), .B(n14048), .ZN(
        P2_U2875) );
  NAND4_X1 U17446 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_4__SCAN_IN), .ZN(n14539)
         );
  INV_X1 U17447 ( .A(n20116), .ZN(n14102) );
  NOR2_X1 U17448 ( .A1(n14539), .A2(n14102), .ZN(n14660) );
  INV_X1 U17449 ( .A(n14660), .ZN(n14050) );
  NAND2_X1 U17450 ( .A1(n16166), .A2(n14050), .ZN(n14675) );
  INV_X1 U17451 ( .A(n14675), .ZN(n20107) );
  NAND2_X1 U17452 ( .A1(n20107), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n14053) );
  OAI22_X1 U17453 ( .A1(n21293), .A2(n20094), .B1(n16168), .B2(n14186), .ZN(
        n14051) );
  AOI211_X1 U17454 ( .C1(n20131), .C2(n14083), .A(n14051), .B(n20232), .ZN(
        n14052) );
  OAI211_X1 U17455 ( .C1(n14054), .C2(n20095), .A(n14053), .B(n14052), .ZN(
        n14055) );
  AOI21_X1 U17456 ( .B1(n14056), .B2(n20129), .A(n14055), .ZN(n14060) );
  NAND3_X1 U17457 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n14057) );
  NOR2_X1 U17458 ( .A1(n20118), .A2(n14057), .ZN(n14058) );
  INV_X1 U17459 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20944) );
  NAND2_X1 U17460 ( .A1(n14058), .A2(n20944), .ZN(n14059) );
  OAI211_X1 U17461 ( .C1(n14086), .C2(n14109), .A(n14060), .B(n14059), .ZN(
        P1_U2836) );
  INV_X1 U17462 ( .A(n19455), .ZN(n14062) );
  NAND2_X1 U17463 ( .A1(n14062), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19449) );
  OR2_X1 U17464 ( .A1(n19449), .A2(n19503), .ZN(n14063) );
  NAND3_X1 U17465 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20024), .A3(
        n20032), .ZN(n19639) );
  NAND2_X1 U17466 ( .A1(n14063), .A2(n19639), .ZN(n14066) );
  NOR2_X1 U17467 ( .A1(n20040), .A2(n19639), .ZN(n19684) );
  INV_X1 U17468 ( .A(n19684), .ZN(n14064) );
  MUX2_X1 U17469 ( .A(n14066), .B(n14065), .S(n20013), .Z(n14067) );
  NAND2_X1 U17470 ( .A1(n14067), .A2(n19851), .ZN(n19687) );
  INV_X1 U17471 ( .A(n19639), .ZN(n14068) );
  NAND2_X1 U17472 ( .A1(n14068), .A2(n20004), .ZN(n14071) );
  OAI21_X1 U17473 ( .B1(n14069), .B2(n19684), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14070) );
  NAND2_X1 U17474 ( .A1(n14071), .A2(n14070), .ZN(n19686) );
  AOI22_X1 U17475 ( .A1(n19811), .A2(n19714), .B1(n19858), .B2(n19686), .ZN(
        n14073) );
  AOI22_X1 U17476 ( .A1(n19863), .A2(n19685), .B1(n19859), .B2(n19684), .ZN(
        n14072) );
  OAI211_X1 U17477 ( .C1(n19678), .C2(n14074), .A(n14073), .B(n14072), .ZN(
        P2_U3121) );
  INV_X1 U17478 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14079) );
  AOI22_X1 U17479 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19433), .ZN(n19857) );
  INV_X1 U17480 ( .A(n19857), .ZN(n19792) );
  NOR2_X2 U17481 ( .A1(n14075), .A2(n19765), .ZN(n19791) );
  AOI22_X1 U17482 ( .A1(n19792), .A2(n19714), .B1(n19791), .B2(n19686), .ZN(
        n14078) );
  AOI22_X1 U17483 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19433), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19432), .ZN(n19733) );
  AND2_X1 U17484 ( .A1(n9736), .A2(n19434), .ZN(n19842) );
  AOI22_X1 U17485 ( .A1(n19854), .A2(n19685), .B1(n19842), .B2(n19684), .ZN(
        n14077) );
  OAI211_X1 U17486 ( .C1(n19678), .C2(n14079), .A(n14078), .B(n14077), .ZN(
        P2_U3120) );
  XOR2_X1 U17487 ( .A(n14080), .B(n14081), .Z(n14190) );
  NAND2_X1 U17488 ( .A1(n14190), .A2(n20230), .ZN(n14085) );
  NAND2_X1 U17489 ( .A1(n20232), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n14184) );
  OAI21_X1 U17490 ( .B1(n16256), .B2(n21293), .A(n14184), .ZN(n14082) );
  AOI21_X1 U17491 ( .B1(n14083), .B2(n16252), .A(n14082), .ZN(n14084) );
  OAI211_X1 U17492 ( .C1(n20238), .C2(n14086), .A(n14085), .B(n14084), .ZN(
        P1_U2995) );
  INV_X1 U17493 ( .A(n14088), .ZN(n14210) );
  AOI21_X1 U17494 ( .B1(n14089), .B2(n13935), .A(n14210), .ZN(n16245) );
  INV_X1 U17495 ( .A(n16245), .ZN(n14099) );
  AOI21_X1 U17496 ( .B1(n14091), .B2(n14090), .A(n16350), .ZN(n16358) );
  AOI22_X1 U17497 ( .A1(n16358), .A2(n20148), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14707), .ZN(n14092) );
  OAI21_X1 U17498 ( .B1(n14099), .B2(n14728), .A(n14092), .ZN(P1_U2866) );
  OAI222_X1 U17499 ( .A1(n14785), .A2(n14099), .B1(n14748), .B2(n12454), .C1(
        n14439), .C2(n20283), .ZN(P1_U2898) );
  INV_X1 U17500 ( .A(n16166), .ZN(n16099) );
  INV_X1 U17501 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20948) );
  INV_X1 U17502 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20946) );
  NOR2_X1 U17503 ( .A1(n20948), .A2(n20946), .ZN(n20091) );
  OAI21_X1 U17504 ( .B1(n16099), .B2(n20091), .A(n14675), .ZN(n20098) );
  OAI22_X1 U17505 ( .A1(n20095), .A2(n14093), .B1(n16178), .B2(n16248), .ZN(
        n14097) );
  NAND2_X1 U17506 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20106), .ZN(n14095) );
  AOI22_X1 U17507 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20128), .B1(
        n20127), .B2(n16358), .ZN(n14094) );
  OAI211_X1 U17508 ( .C1(P1_REIP_REG_6__SCAN_IN), .C2(n14095), .A(n14094), .B(
        n20100), .ZN(n14096) );
  AOI211_X1 U17509 ( .C1(P1_REIP_REG_6__SCAN_IN), .C2(n20098), .A(n14097), .B(
        n14096), .ZN(n14098) );
  OAI21_X1 U17510 ( .B1(n16182), .B2(n14099), .A(n14098), .ZN(P1_U2834) );
  INV_X1 U17511 ( .A(n14101), .ZN(n20804) );
  NAND2_X1 U17512 ( .A1(n20133), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U17513 ( .A1(n20128), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14102), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14103) );
  OAI211_X1 U17514 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n16178), .A(
        n14104), .B(n14103), .ZN(n14107) );
  OAI22_X1 U17515 ( .A1(n16168), .A2(n14105), .B1(n20118), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14106) );
  AOI211_X1 U17516 ( .C1(n20804), .C2(n20129), .A(n14107), .B(n14106), .ZN(
        n14108) );
  OAI21_X1 U17517 ( .B1(n20225), .B2(n14109), .A(n14108), .ZN(P1_U2839) );
  OR2_X1 U17518 ( .A1(n14111), .A2(n14110), .ZN(n14113) );
  NAND2_X1 U17519 ( .A1(n14113), .A2(n14112), .ZN(n19331) );
  XOR2_X1 U17520 ( .A(n19331), .B(n19503), .Z(n19334) );
  INV_X1 U17521 ( .A(n14153), .ZN(n20022) );
  OAI21_X1 U17522 ( .B1(n14275), .B2(n20022), .A(n14114), .ZN(n19333) );
  NAND2_X1 U17523 ( .A1(n19334), .A2(n19333), .ZN(n19332) );
  NAND2_X1 U17524 ( .A1(n19503), .A2(n19331), .ZN(n14117) );
  INV_X1 U17525 ( .A(n14112), .ZN(n14115) );
  XNOR2_X1 U17526 ( .A(n14116), .B(n14115), .ZN(n15824) );
  AOI21_X1 U17527 ( .B1(n19332), .B2(n14117), .A(n15824), .ZN(n19326) );
  XNOR2_X1 U17528 ( .A(n19326), .B(n19325), .ZN(n14120) );
  AOI22_X1 U17529 ( .A1(n19339), .A2(n15824), .B1(n19338), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n14119) );
  INV_X1 U17530 ( .A(n19429), .ZN(n16410) );
  NAND2_X1 U17531 ( .A1(n19314), .A2(n16410), .ZN(n14118) );
  OAI211_X1 U17532 ( .C1(n14120), .C2(n19324), .A(n14119), .B(n14118), .ZN(
        P2_U2915) );
  OR2_X1 U17533 ( .A1(n14088), .A2(n14121), .ZN(n14212) );
  NAND2_X1 U17534 ( .A1(n14088), .A2(n14121), .ZN(n14122) );
  INV_X1 U17535 ( .A(n20150), .ZN(n14124) );
  OAI222_X1 U17536 ( .A1(n14124), .A2(n14785), .B1(n14123), .B2(n14748), .C1(
        n14439), .C2(n20291), .ZN(P1_U2897) );
  AND2_X1 U17537 ( .A1(n14126), .A2(n14127), .ZN(n14128) );
  OR2_X1 U17538 ( .A1(n14231), .A2(n14129), .ZN(n14130) );
  NAND2_X1 U17539 ( .A1(n14125), .A2(n14130), .ZN(n16183) );
  AND2_X1 U17540 ( .A1(n14399), .A2(n14131), .ZN(n14132) );
  NOR2_X1 U17541 ( .A1(n14446), .A2(n14132), .ZN(n16180) );
  AOI22_X1 U17542 ( .A1(n16180), .A2(n20148), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14707), .ZN(n14133) );
  OAI21_X1 U17543 ( .B1(n16183), .B2(n14728), .A(n14133), .ZN(P1_U2862) );
  INV_X1 U17544 ( .A(n14439), .ZN(n14136) );
  INV_X1 U17545 ( .A(DATAI_10_), .ZN(n14135) );
  NAND2_X1 U17546 ( .A1(n20239), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14134) );
  OAI21_X1 U17547 ( .B1(n20239), .B2(n14135), .A(n14134), .ZN(n20188) );
  AOI22_X1 U17548 ( .A1(n14136), .A2(n20188), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14767), .ZN(n14137) );
  OAI21_X1 U17549 ( .B1(n16183), .B2(n14785), .A(n14137), .ZN(P1_U2894) );
  NOR2_X1 U17550 ( .A1(n19242), .A2(n14138), .ZN(n14139) );
  XNOR2_X1 U17551 ( .A(n14139), .B(n14175), .ZN(n14140) );
  NAND2_X1 U17552 ( .A1(n14140), .A2(n19246), .ZN(n14148) );
  INV_X1 U17553 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14176) );
  OAI22_X1 U17554 ( .A1(n14141), .A2(n19252), .B1(n14174), .B2(n19222), .ZN(
        n14142) );
  AOI21_X1 U17555 ( .B1(n19279), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n14142), .ZN(n14143) );
  OAI21_X1 U17556 ( .B1(n14144), .B2(n19270), .A(n14143), .ZN(n14146) );
  NOR2_X1 U17557 ( .A1(n19331), .A2(n19258), .ZN(n14145) );
  AOI211_X1 U17558 ( .C1(n19273), .C2(n13739), .A(n14146), .B(n14145), .ZN(
        n14147) );
  OAI211_X1 U17559 ( .C1(n19503), .C2(n14201), .A(n14148), .B(n14147), .ZN(
        P2_U2852) );
  NAND2_X1 U17560 ( .A1(n19226), .A2(n14311), .ZN(n14150) );
  XNOR2_X1 U17561 ( .A(n14151), .B(n14150), .ZN(n14152) );
  NAND2_X1 U17562 ( .A1(n14152), .A2(n19246), .ZN(n14161) );
  OAI22_X1 U17563 ( .A1(n14153), .A2(n19258), .B1(n12934), .B2(n19250), .ZN(
        n14156) );
  NOR2_X1 U17564 ( .A1(n19252), .A2(n14154), .ZN(n14155) );
  AOI211_X1 U17565 ( .C1(n19265), .C2(P2_REIP_REG_2__SCAN_IN), .A(n14156), .B(
        n14155), .ZN(n14157) );
  OAI21_X1 U17566 ( .B1(n14158), .B2(n19270), .A(n14157), .ZN(n14159) );
  AOI21_X1 U17567 ( .B1(n11277), .B2(n19273), .A(n14159), .ZN(n14160) );
  OAI211_X1 U17568 ( .C1(n20020), .C2(n14201), .A(n14161), .B(n14160), .ZN(
        P2_U2853) );
  XNOR2_X1 U17569 ( .A(n15815), .B(n14164), .ZN(n15817) );
  XNOR2_X1 U17570 ( .A(n15817), .B(n15816), .ZN(n14182) );
  INV_X1 U17571 ( .A(n14162), .ZN(n14166) );
  NOR2_X1 U17572 ( .A1(n14163), .A2(n16482), .ZN(n14165) );
  MUX2_X1 U17573 ( .A(n14166), .B(n14165), .S(n14164), .Z(n14168) );
  OAI22_X1 U17574 ( .A1(n19331), .A2(n16474), .B1(n14174), .B2(n19214), .ZN(
        n14167) );
  AOI211_X1 U17575 ( .C1(n16479), .C2(n13739), .A(n14168), .B(n14167), .ZN(
        n14173) );
  NAND2_X1 U17576 ( .A1(n14171), .A2(n14170), .ZN(n14179) );
  NAND3_X1 U17577 ( .A1(n14169), .A2(n14179), .A3(n16461), .ZN(n14172) );
  OAI211_X1 U17578 ( .C1(n14182), .C2(n15800), .A(n14173), .B(n14172), .ZN(
        P2_U3043) );
  NOR2_X1 U17579 ( .A1(n19214), .A2(n14174), .ZN(n14178) );
  OAI22_X1 U17580 ( .A1(n14176), .A2(n19409), .B1(n16455), .B2(n14175), .ZN(
        n14177) );
  AOI211_X1 U17581 ( .C1(n19403), .C2(n10334), .A(n14178), .B(n14177), .ZN(
        n14181) );
  NAND3_X1 U17582 ( .A1(n14169), .A2(n14179), .A3(n19404), .ZN(n14180) );
  OAI211_X1 U17583 ( .C1(n14182), .C2(n16435), .A(n14181), .B(n14180), .ZN(
        P2_U3011) );
  NAND2_X1 U17584 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14183), .ZN(
        n14185) );
  OAI211_X1 U17585 ( .C1(n16341), .C2(n14186), .A(n14185), .B(n14184), .ZN(
        n14189) );
  AOI211_X1 U17586 ( .C1(n12228), .C2(n14187), .A(n16332), .B(n16374), .ZN(
        n14188) );
  AOI211_X1 U17587 ( .C1(n14190), .C2(n16360), .A(n14189), .B(n14188), .ZN(
        n14191) );
  INV_X1 U17588 ( .A(n14191), .ZN(P1_U3027) );
  AND2_X1 U17589 ( .A1(n19226), .A2(n14192), .ZN(n14194) );
  AOI21_X1 U17590 ( .B1(n19397), .B2(n14194), .A(n19928), .ZN(n14193) );
  OAI21_X1 U17591 ( .B1(n19397), .B2(n14194), .A(n14193), .ZN(n14200) );
  AOI22_X1 U17592 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19264), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19265), .ZN(n14195) );
  OAI211_X1 U17593 ( .C1(n19250), .C2(n19408), .A(n19214), .B(n14195), .ZN(
        n14196) );
  AOI21_X1 U17594 ( .B1(n19266), .B2(n15824), .A(n14196), .ZN(n14197) );
  OAI21_X1 U17595 ( .B1(n15818), .B2(n19270), .A(n14197), .ZN(n14198) );
  AOI21_X1 U17596 ( .B1(n19402), .B2(n19273), .A(n14198), .ZN(n14199) );
  OAI211_X1 U17597 ( .C1(n14201), .C2(n19325), .A(n14200), .B(n14199), .ZN(
        P2_U2851) );
  AND2_X1 U17598 ( .A1(n14247), .A2(n14238), .ZN(n14236) );
  NAND2_X1 U17599 ( .A1(n14247), .A2(n14202), .ZN(n14255) );
  OAI211_X1 U17600 ( .C1(n14236), .C2(n14203), .A(n14255), .B(n15235), .ZN(
        n14209) );
  OAI21_X1 U17601 ( .B1(n14204), .B2(n14206), .A(n14205), .ZN(n14207) );
  INV_X1 U17602 ( .A(n14207), .ZN(n19136) );
  NAND2_X1 U17603 ( .A1(n19136), .A2(n15229), .ZN(n14208) );
  OAI211_X1 U17604 ( .C1(n15229), .C2(n10707), .A(n14209), .B(n14208), .ZN(
        P2_U2872) );
  NAND2_X1 U17605 ( .A1(n14210), .A2(n14126), .ZN(n14229) );
  INV_X1 U17606 ( .A(n14229), .ZN(n14211) );
  AOI21_X1 U17607 ( .B1(n14213), .B2(n14212), .A(n14211), .ZN(n14297) );
  INV_X1 U17608 ( .A(n14297), .ZN(n14683) );
  INV_X1 U17609 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14215) );
  INV_X1 U17610 ( .A(DATAI_8_), .ZN(n14214) );
  INV_X1 U17611 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16618) );
  MUX2_X1 U17612 ( .A(n14214), .B(n16618), .S(n20239), .Z(n20181) );
  OAI222_X1 U17613 ( .A1(n14683), .A2(n14785), .B1(n14215), .B2(n14748), .C1(
        n14439), .C2(n20181), .ZN(P1_U2896) );
  INV_X1 U17614 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14217) );
  OAI21_X1 U17615 ( .B1(n16352), .B2(n14216), .A(n14397), .ZN(n16342) );
  OAI222_X1 U17616 ( .A1(n14683), .A2(n14728), .B1(n20153), .B2(n14217), .C1(
        n16342), .C2(n14727), .ZN(P1_U2864) );
  AND2_X1 U17617 ( .A1(n14247), .A2(n14218), .ZN(n14254) );
  NAND2_X1 U17618 ( .A1(n14220), .A2(n14219), .ZN(n14389) );
  OAI21_X1 U17619 ( .B1(n14254), .B2(n14221), .A(n14389), .ZN(n14444) );
  XNOR2_X1 U17620 ( .A(n14222), .B(n14223), .ZN(n15670) );
  INV_X1 U17621 ( .A(n15670), .ZN(n19113) );
  OAI22_X1 U17622 ( .A1(n15284), .A2(n19348), .B1(n19322), .B2(n21309), .ZN(
        n14226) );
  INV_X1 U17623 ( .A(n19291), .ZN(n15287) );
  INV_X1 U17624 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14224) );
  OAI22_X1 U17625 ( .A1(n15287), .A2(n16603), .B1(n19284), .B2(n14224), .ZN(
        n14225) );
  AOI211_X1 U17626 ( .C1(n19339), .C2(n19113), .A(n14226), .B(n14225), .ZN(
        n14227) );
  OAI21_X1 U17627 ( .B1(n14444), .B2(n19324), .A(n14227), .ZN(P2_U2902) );
  AND2_X1 U17628 ( .A1(n14229), .A2(n14228), .ZN(n14230) );
  INV_X1 U17629 ( .A(n20145), .ZN(n14235) );
  INV_X1 U17630 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14234) );
  INV_X1 U17631 ( .A(DATAI_9_), .ZN(n14233) );
  MUX2_X1 U17632 ( .A(n14233), .B(n14232), .S(n20239), .Z(n20184) );
  OAI222_X1 U17633 ( .A1(n14235), .A2(n14785), .B1(n14234), .B2(n14748), .C1(
        n14439), .C2(n20184), .ZN(P1_U2895) );
  INV_X1 U17634 ( .A(n14236), .ZN(n14237) );
  OAI211_X1 U17635 ( .C1(n14247), .C2(n14238), .A(n14237), .B(n15235), .ZN(
        n14241) );
  AOI21_X1 U17636 ( .B1(n14239), .B2(n14245), .A(n14204), .ZN(n19147) );
  NAND2_X1 U17637 ( .A1(n19147), .A2(n15229), .ZN(n14240) );
  OAI211_X1 U17638 ( .C1(n15229), .C2(n14242), .A(n14241), .B(n14240), .ZN(
        P2_U2873) );
  NAND2_X1 U17639 ( .A1(n10006), .A2(n14243), .ZN(n14244) );
  NAND2_X1 U17640 ( .A1(n14245), .A2(n14244), .ZN(n19156) );
  INV_X1 U17641 ( .A(n19156), .ZN(n14252) );
  INV_X1 U17642 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n14246) );
  NOR2_X1 U17643 ( .A1(n15229), .A2(n14246), .ZN(n14251) );
  AOI211_X1 U17644 ( .C1(n14249), .C2(n14248), .A(n15242), .B(n14247), .ZN(
        n14250) );
  AOI211_X1 U17645 ( .C1(n14252), .C2(n15229), .A(n14251), .B(n14250), .ZN(
        n14253) );
  INV_X1 U17646 ( .A(n14253), .ZN(P2_U2874) );
  AOI21_X1 U17647 ( .B1(n14256), .B2(n14255), .A(n14254), .ZN(n19293) );
  NAND2_X1 U17648 ( .A1(n19293), .A2(n15235), .ZN(n14260) );
  INV_X1 U17649 ( .A(n14257), .ZN(n14440) );
  AOI21_X1 U17650 ( .B1(n14258), .B2(n14205), .A(n14257), .ZN(n19125) );
  NAND2_X1 U17651 ( .A1(n19125), .A2(n15229), .ZN(n14259) );
  OAI211_X1 U17652 ( .C1(n15229), .C2(n14261), .A(n14260), .B(n14259), .ZN(
        P2_U2871) );
  AOI21_X1 U17653 ( .B1(n14264), .B2(n14262), .A(n14263), .ZN(n19316) );
  NAND2_X1 U17654 ( .A1(n19226), .A2(n14265), .ZN(n14266) );
  XOR2_X1 U17655 ( .A(n16454), .B(n14266), .Z(n14267) );
  AOI22_X1 U17656 ( .A1(n19316), .A2(n19266), .B1(n19246), .B2(n14267), .ZN(
        n14273) );
  INV_X1 U17657 ( .A(n14268), .ZN(n16460) );
  INV_X1 U17658 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n14269) );
  INV_X1 U17659 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21109) );
  OAI22_X1 U17660 ( .A1(n19222), .A2(n14269), .B1(n19250), .B2(n21109), .ZN(
        n14271) );
  OAI21_X1 U17661 ( .B1(n10831), .B2(n19252), .A(n19214), .ZN(n14270) );
  AOI211_X1 U17662 ( .C1(n16460), .C2(n19273), .A(n14271), .B(n14270), .ZN(
        n14272) );
  OAI211_X1 U17663 ( .C1(n14274), .C2(n19270), .A(n14273), .B(n14272), .ZN(
        P2_U2847) );
  OAI21_X1 U17664 ( .B1(n19832), .B2(n19915), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14276) );
  NAND2_X1 U17665 ( .A1(n14276), .A2(n20004), .ZN(n14278) );
  NAND2_X1 U17666 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19579), .ZN(
        n19849) );
  NOR2_X1 U17667 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19849), .ZN(
        n19830) );
  NOR2_X1 U17668 ( .A1(n19830), .A2(n19805), .ZN(n14281) );
  INV_X1 U17669 ( .A(n10524), .ZN(n14279) );
  OAI21_X1 U17670 ( .B1(n14279), .B2(n19830), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14277) );
  INV_X1 U17671 ( .A(n19833), .ZN(n14291) );
  INV_X1 U17672 ( .A(n19791), .ZN(n19844) );
  INV_X1 U17673 ( .A(n14278), .ZN(n14282) );
  AOI211_X1 U17674 ( .C1(n14279), .C2(n20033), .A(n19830), .B(n20004), .ZN(
        n14280) );
  AOI211_X2 U17675 ( .C1(n14282), .C2(n14281), .A(n14280), .B(n19765), .ZN(
        n19837) );
  INV_X1 U17676 ( .A(n19837), .ZN(n14289) );
  INV_X1 U17677 ( .A(n19832), .ZN(n14287) );
  AOI22_X1 U17678 ( .A1(n19792), .A2(n19915), .B1(n19842), .B2(n19830), .ZN(
        n14283) );
  OAI21_X1 U17679 ( .B1(n19733), .B2(n14287), .A(n14283), .ZN(n14284) );
  AOI21_X1 U17680 ( .B1(n14289), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n14284), .ZN(n14285) );
  OAI21_X1 U17681 ( .B1(n14291), .B2(n19844), .A(n14285), .ZN(P2_U3160) );
  INV_X1 U17682 ( .A(n19782), .ZN(n19901) );
  AOI22_X1 U17683 ( .A1(n19748), .A2(n19915), .B1(n9707), .B2(n19830), .ZN(
        n14286) );
  OAI21_X1 U17684 ( .B1(n14287), .B2(n19751), .A(n14286), .ZN(n14288) );
  AOI21_X1 U17685 ( .B1(n14289), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n14288), .ZN(n14290) );
  OAI21_X1 U17686 ( .B1(n14291), .B2(n19901), .A(n14290), .ZN(P2_U3166) );
  XNOR2_X1 U17687 ( .A(n14292), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14293) );
  XNOR2_X1 U17688 ( .A(n14294), .B(n14293), .ZN(n16344) );
  INV_X1 U17689 ( .A(n16344), .ZN(n14299) );
  AOI22_X1 U17690 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14295) );
  OAI21_X1 U17691 ( .B1(n20219), .B2(n14676), .A(n14295), .ZN(n14296) );
  AOI21_X1 U17692 ( .B1(n14297), .B2(n13942), .A(n14296), .ZN(n14298) );
  OAI21_X1 U17693 ( .B1(n14299), .B2(n20220), .A(n14298), .ZN(P1_U2991) );
  XNOR2_X1 U17694 ( .A(n14301), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14302) );
  XNOR2_X1 U17695 ( .A(n9763), .B(n14302), .ZN(n14350) );
  NOR2_X1 U17696 ( .A1(n14305), .A2(n14304), .ZN(n14306) );
  XNOR2_X1 U17697 ( .A(n14303), .B(n14306), .ZN(n14353) );
  NAND2_X1 U17698 ( .A1(n14353), .A2(n19404), .ZN(n14310) );
  INV_X1 U17699 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n14307) );
  NOR2_X1 U17700 ( .A1(n19214), .A2(n14307), .ZN(n14344) );
  INV_X1 U17701 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19237) );
  OAI22_X1 U17702 ( .A1(n16428), .A2(n19237), .B1(n16455), .B2(n19243), .ZN(
        n14308) );
  AOI211_X1 U17703 ( .C1(n19403), .C2(n19245), .A(n14344), .B(n14308), .ZN(
        n14309) );
  OAI211_X1 U17704 ( .C1(n16435), .C2(n14350), .A(n14310), .B(n14309), .ZN(
        P2_U3009) );
  OAI211_X1 U17705 ( .C1(n14313), .C2(n14312), .A(n19226), .B(n14311), .ZN(
        n19263) );
  OAI21_X1 U17706 ( .B1(n19226), .B2(n15833), .A(n19263), .ZN(n15861) );
  INV_X1 U17707 ( .A(n14313), .ZN(n19274) );
  AOI22_X1 U17708 ( .A1(n19242), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19274), .B2(n19226), .ZN(n15846) );
  NOR2_X1 U17709 ( .A1(n15846), .A2(n19921), .ZN(n15851) );
  NAND2_X1 U17710 ( .A1(n14315), .A2(n14314), .ZN(n15874) );
  INV_X1 U17711 ( .A(n10370), .ZN(n14316) );
  NAND2_X1 U17712 ( .A1(n14316), .A2(n16484), .ZN(n14319) );
  NAND2_X1 U17713 ( .A1(n15874), .A2(n14319), .ZN(n14318) );
  INV_X1 U17714 ( .A(n16505), .ZN(n14317) );
  NOR2_X1 U17715 ( .A1(n14317), .A2(n16503), .ZN(n15865) );
  MUX2_X1 U17716 ( .A(n14318), .B(n15865), .S(n10193), .Z(n14325) );
  INV_X1 U17717 ( .A(n15865), .ZN(n14320) );
  INV_X1 U17718 ( .A(n14319), .ZN(n15864) );
  NAND2_X1 U17719 ( .A1(n14320), .A2(n15864), .ZN(n15866) );
  OAI21_X1 U17720 ( .B1(n14323), .B2(n14321), .A(n14322), .ZN(n14324) );
  NAND3_X1 U17721 ( .A1(n14325), .A2(n15866), .A3(n14324), .ZN(n14326) );
  AOI21_X1 U17722 ( .B1(n11277), .B2(n15863), .A(n14326), .ZN(n16483) );
  OAI22_X1 U17723 ( .A1(n20020), .A2(n15882), .B1(n20006), .B2(n16483), .ZN(
        n14327) );
  AOI21_X1 U17724 ( .B1(n15861), .B2(n15851), .A(n14327), .ZN(n14328) );
  MUX2_X1 U17725 ( .A(n14328), .B(n16484), .S(n15883), .Z(n14329) );
  INV_X1 U17726 ( .A(n14329), .ZN(P2_U3599) );
  OAI21_X1 U17727 ( .B1(n9823), .B2(n10115), .A(n15233), .ZN(n15243) );
  NAND2_X1 U17728 ( .A1(n14331), .A2(n14332), .ZN(n14333) );
  AND2_X1 U17729 ( .A1(n15165), .A2(n14333), .ZN(n19089) );
  OAI22_X1 U17730 ( .A1(n15284), .A2(n19426), .B1(n19322), .B2(n14334), .ZN(
        n14338) );
  INV_X1 U17731 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14336) );
  INV_X1 U17732 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14335) );
  OAI22_X1 U17733 ( .A1(n15287), .A2(n14336), .B1(n19284), .B2(n14335), .ZN(
        n14337) );
  AOI211_X1 U17734 ( .C1(n19339), .C2(n19089), .A(n14338), .B(n14337), .ZN(
        n14339) );
  OAI21_X1 U17735 ( .B1(n15243), .B2(n19324), .A(n14339), .ZN(P2_U2900) );
  OAI21_X1 U17736 ( .B1(n14340), .B2(n14342), .A(n14341), .ZN(n19329) );
  OAI211_X1 U17737 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n15823), .B(n14343), .ZN(n14349) );
  INV_X1 U17738 ( .A(n14344), .ZN(n14345) );
  OAI21_X1 U17739 ( .B1(n15834), .B2(n14346), .A(n14345), .ZN(n14347) );
  AOI21_X1 U17740 ( .B1(n15822), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n14347), .ZN(n14348) );
  OAI211_X1 U17741 ( .C1(n19329), .C2(n16474), .A(n14349), .B(n14348), .ZN(
        n14352) );
  NOR2_X1 U17742 ( .A1(n14350), .A2(n15800), .ZN(n14351) );
  AOI211_X1 U17743 ( .C1(n14353), .C2(n16461), .A(n14352), .B(n14351), .ZN(
        n14354) );
  INV_X1 U17744 ( .A(n14354), .ZN(P2_U3041) );
  INV_X1 U17745 ( .A(n14125), .ZN(n14357) );
  INV_X1 U17746 ( .A(n14355), .ZN(n14356) );
  OAI21_X1 U17747 ( .B1(n14357), .B2(n14356), .A(n14358), .ZN(n14422) );
  OAI21_X1 U17748 ( .B1(n14422), .B2(n14423), .A(n14358), .ZN(n14360) );
  NAND2_X1 U17749 ( .A1(n14360), .A2(n14359), .ZN(n14406) );
  OAI21_X1 U17750 ( .B1(n14360), .B2(n14359), .A(n14406), .ZN(n16157) );
  INV_X1 U17751 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14364) );
  OR2_X1 U17752 ( .A1(n14361), .A2(n14362), .ZN(n14363) );
  NAND2_X1 U17753 ( .A1(n14408), .A2(n14363), .ZN(n16158) );
  OAI222_X1 U17754 ( .A1(n16157), .A2(n14728), .B1(n14364), .B2(n20153), .C1(
        n16158), .C2(n14727), .ZN(P1_U2860) );
  INV_X1 U17755 ( .A(DATAI_12_), .ZN(n14365) );
  MUX2_X1 U17756 ( .A(n14365), .B(n16611), .S(n20239), .Z(n20193) );
  OAI222_X1 U17757 ( .A1(n16157), .A2(n14785), .B1(n14366), .B2(n14748), .C1(
        n14439), .C2(n20193), .ZN(P1_U2892) );
  OAI21_X1 U17758 ( .B1(n14368), .B2(n14370), .A(n14369), .ZN(n16148) );
  INV_X1 U17759 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14373) );
  INV_X1 U17760 ( .A(DATAI_14_), .ZN(n14372) );
  MUX2_X1 U17761 ( .A(n14372), .B(n14371), .S(n20239), .Z(n20199) );
  OAI222_X1 U17762 ( .A1(n16148), .A2(n14785), .B1(n14373), .B2(n14748), .C1(
        n14439), .C2(n20199), .ZN(P1_U2890) );
  NAND2_X1 U17763 ( .A1(n14410), .A2(n14374), .ZN(n14375) );
  NAND2_X1 U17764 ( .A1(n14436), .A2(n14375), .ZN(n16313) );
  INV_X1 U17765 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14376) );
  OAI222_X1 U17766 ( .A1(n16313), .A2(n14727), .B1(n14376), .B2(n20153), .C1(
        n16148), .C2(n14728), .ZN(P1_U2858) );
  XNOR2_X1 U17767 ( .A(n12088), .B(n15030), .ZN(n14377) );
  XNOR2_X1 U17768 ( .A(n14378), .B(n14377), .ZN(n14403) );
  INV_X1 U17769 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14379) );
  NOR2_X1 U17770 ( .A1(n20100), .A2(n14379), .ZN(n14400) );
  AOI21_X1 U17771 ( .B1(n20228), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n14400), .ZN(n14381) );
  NAND2_X1 U17772 ( .A1(n16252), .A2(n20081), .ZN(n14380) );
  NAND2_X1 U17773 ( .A1(n14381), .A2(n14380), .ZN(n14382) );
  AOI21_X1 U17774 ( .B1(n20145), .B2(n13942), .A(n14382), .ZN(n14383) );
  OAI21_X1 U17775 ( .B1(n14403), .B2(n20220), .A(n14383), .ZN(P1_U2990) );
  NOR2_X1 U17776 ( .A1(n14385), .A2(n14386), .ZN(n14387) );
  OR2_X1 U17777 ( .A1(n14384), .A2(n14387), .ZN(n19102) );
  INV_X1 U17778 ( .A(n14388), .ZN(n14390) );
  AOI21_X1 U17779 ( .B1(n14390), .B2(n14389), .A(n9823), .ZN(n16418) );
  NAND2_X1 U17780 ( .A1(n16418), .A2(n15235), .ZN(n14392) );
  NAND2_X1 U17781 ( .A1(n13900), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14391) );
  OAI211_X1 U17782 ( .C1(n19102), .C2(n13900), .A(n14392), .B(n14391), .ZN(
        P2_U2869) );
  NAND3_X1 U17783 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14393) );
  NOR2_X1 U17784 ( .A1(n14393), .A2(n15007), .ZN(n15027) );
  AOI21_X1 U17785 ( .B1(n15027), .B2(n15026), .A(n15025), .ZN(n14395) );
  NAND2_X1 U17786 ( .A1(n15027), .A2(n16316), .ZN(n16331) );
  INV_X1 U17787 ( .A(n16331), .ZN(n14394) );
  AOI22_X1 U17788 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n14395), .B1(
        n14394), .B2(n15030), .ZN(n14402) );
  NAND2_X1 U17789 ( .A1(n14397), .A2(n14396), .ZN(n14398) );
  AND2_X1 U17790 ( .A1(n14399), .A2(n14398), .ZN(n20144) );
  AOI21_X1 U17791 ( .B1(n20144), .B2(n16367), .A(n14400), .ZN(n14401) );
  OAI211_X1 U17792 ( .C1(n14403), .C2(n16370), .A(n14402), .B(n14401), .ZN(
        P1_U3022) );
  INV_X1 U17793 ( .A(n14404), .ZN(n14405) );
  AOI21_X1 U17794 ( .B1(n14406), .B2(n14405), .A(n14368), .ZN(n14899) );
  INV_X1 U17795 ( .A(n14899), .ZN(n14431) );
  INV_X1 U17796 ( .A(n14897), .ZN(n14420) );
  NAND2_X1 U17797 ( .A1(n14408), .A2(n14407), .ZN(n14409) );
  NAND2_X1 U17798 ( .A1(n14410), .A2(n14409), .ZN(n14996) );
  INV_X1 U17799 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14430) );
  OAI22_X1 U17800 ( .A1(n14996), .A2(n16168), .B1(n14430), .B2(n20095), .ZN(
        n14411) );
  INV_X1 U17801 ( .A(n14411), .ZN(n14412) );
  OAI211_X1 U17802 ( .C1(n20094), .C2(n14413), .A(n14412), .B(n20100), .ZN(
        n14419) );
  NAND2_X1 U17803 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14415) );
  INV_X1 U17804 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20951) );
  NAND3_X1 U17805 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n14679) );
  NOR2_X1 U17806 ( .A1(n20951), .A2(n14679), .ZN(n20080) );
  NAND3_X1 U17807 ( .A1(n20080), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .ZN(n14537) );
  INV_X1 U17808 ( .A(n20106), .ZN(n14414) );
  NOR2_X1 U17809 ( .A1(n14415), .A2(n16174), .ZN(n14417) );
  NAND4_X1 U17810 ( .A1(n20080), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .A4(n14660), .ZN(n16165) );
  OAI21_X1 U17811 ( .B1(n14415), .B2(n16165), .A(n16166), .ZN(n16163) );
  INV_X1 U17812 ( .A(n16163), .ZN(n14416) );
  MUX2_X1 U17813 ( .A(n14417), .B(n14416), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14418) );
  AOI211_X1 U17814 ( .C1(n20131), .C2(n14420), .A(n14419), .B(n14418), .ZN(
        n14421) );
  OAI21_X1 U17815 ( .B1(n14431), .B2(n16182), .A(n14421), .ZN(P1_U2827) );
  XOR2_X1 U17816 ( .A(n14423), .B(n14422), .Z(n16231) );
  INV_X1 U17817 ( .A(n16231), .ZN(n14448) );
  INV_X1 U17818 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14426) );
  INV_X1 U17819 ( .A(DATAI_11_), .ZN(n14425) );
  MUX2_X1 U17820 ( .A(n14425), .B(n14424), .S(n20239), .Z(n20190) );
  OAI222_X1 U17821 ( .A1(n14448), .A2(n14785), .B1(n14426), .B2(n14748), .C1(
        n14439), .C2(n20190), .ZN(P1_U2893) );
  INV_X1 U17822 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14429) );
  INV_X1 U17823 ( .A(DATAI_13_), .ZN(n14428) );
  MUX2_X1 U17824 ( .A(n14428), .B(n14427), .S(n20239), .Z(n20196) );
  OAI222_X1 U17825 ( .A1(n14431), .A2(n14785), .B1(n14429), .B2(n14748), .C1(
        n14439), .C2(n20196), .ZN(P1_U2891) );
  OAI222_X1 U17826 ( .A1(n14431), .A2(n14728), .B1(n20153), .B2(n14430), .C1(
        n14996), .C2(n14727), .ZN(P1_U2859) );
  INV_X1 U17827 ( .A(n14432), .ZN(n14472) );
  NAND2_X1 U17828 ( .A1(n14369), .A2(n14433), .ZN(n14434) );
  NAND2_X1 U17829 ( .A1(n14472), .A2(n14434), .ZN(n14888) );
  INV_X1 U17830 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14437) );
  XNOR2_X1 U17831 ( .A(n14436), .B(n14435), .ZN(n14987) );
  OAI222_X1 U17832 ( .A1(n14888), .A2(n14728), .B1(n20153), .B2(n14437), .C1(
        n14987), .C2(n14727), .ZN(P1_U2857) );
  OAI222_X1 U17833 ( .A1(n14888), .A2(n14785), .B1(n14748), .B2(n13597), .C1(
        n14439), .C2(n14438), .ZN(P1_U2889) );
  AOI21_X1 U17834 ( .B1(n14441), .B2(n14440), .A(n14385), .ZN(n19114) );
  INV_X1 U17835 ( .A(n19114), .ZN(n15440) );
  NOR2_X1 U17836 ( .A1(n15440), .A2(n13900), .ZN(n14442) );
  AOI21_X1 U17837 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n13900), .A(n14442), .ZN(
        n14443) );
  OAI21_X1 U17838 ( .B1(n14444), .B2(n15242), .A(n14443), .ZN(P2_U2870) );
  NOR2_X1 U17839 ( .A1(n14446), .A2(n14445), .ZN(n14447) );
  OR2_X1 U17840 ( .A1(n14361), .A2(n14447), .ZN(n16324) );
  INV_X1 U17841 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n16167) );
  OAI222_X1 U17842 ( .A1(n16324), .A2(n14727), .B1(n16167), .B2(n20153), .C1(
        n14448), .C2(n14728), .ZN(P1_U2861) );
  XNOR2_X1 U17843 ( .A(n14449), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14469) );
  NAND2_X1 U17844 ( .A1(n9753), .A2(n14452), .ZN(n14453) );
  XOR2_X1 U17845 ( .A(n14450), .B(n14453), .Z(n14467) );
  INV_X1 U17846 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19958) );
  OAI22_X1 U17847 ( .A1(n16428), .A2(n19235), .B1(n19958), .B2(n19214), .ZN(
        n14456) );
  INV_X1 U17848 ( .A(n19228), .ZN(n14454) );
  OAI22_X1 U17849 ( .A1(n15509), .A2(n19229), .B1(n16455), .B2(n14454), .ZN(
        n14455) );
  AOI211_X1 U17850 ( .C1(n14467), .C2(n19400), .A(n14456), .B(n14455), .ZN(
        n14457) );
  OAI21_X1 U17851 ( .B1(n14469), .B2(n16436), .A(n14457), .ZN(P2_U3008) );
  NOR2_X1 U17852 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16463), .ZN(
        n14466) );
  XNOR2_X1 U17853 ( .A(n14458), .B(n14459), .ZN(n19321) );
  INV_X1 U17854 ( .A(n19229), .ZN(n14461) );
  NOR2_X1 U17855 ( .A1(n19958), .A2(n19214), .ZN(n14460) );
  AOI21_X1 U17856 ( .B1(n16479), .B2(n14461), .A(n14460), .ZN(n14464) );
  INV_X1 U17857 ( .A(n16456), .ZN(n14462) );
  NAND2_X1 U17858 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14463) );
  OAI211_X1 U17859 ( .C1(n19321), .C2(n16474), .A(n14464), .B(n14463), .ZN(
        n14465) );
  AOI211_X1 U17860 ( .C1(n14467), .C2(n16471), .A(n14466), .B(n14465), .ZN(
        n14468) );
  OAI21_X1 U17861 ( .B1(n14469), .B2(n16476), .A(n14468), .ZN(P2_U3040) );
  AOI21_X1 U17862 ( .B1(n14473), .B2(n14472), .A(n14471), .ZN(n16207) );
  INV_X1 U17863 ( .A(n16207), .ZN(n14481) );
  OAI21_X1 U17864 ( .B1(n14475), .B2(n14474), .A(n14725), .ZN(n16138) );
  INV_X1 U17865 ( .A(n16138), .ZN(n14476) );
  AOI22_X1 U17866 ( .A1(n14476), .A2(n20148), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14707), .ZN(n14477) );
  OAI21_X1 U17867 ( .B1(n14481), .B2(n14728), .A(n14477), .ZN(P1_U2856) );
  NAND3_X1 U17868 ( .A1(n14748), .A2(n12143), .A3(n20286), .ZN(n14780) );
  OAI22_X1 U17869 ( .A1(n14780), .A2(n20250), .B1(n14748), .B2(n13846), .ZN(
        n14478) );
  AOI21_X1 U17870 ( .B1(n14782), .B2(BUF1_REG_16__SCAN_IN), .A(n14478), .ZN(
        n14480) );
  NAND2_X1 U17871 ( .A1(n13035), .A2(DATAI_16_), .ZN(n14479) );
  OAI211_X1 U17872 ( .C1(n14481), .C2(n14785), .A(n14480), .B(n14479), .ZN(
        P1_U2888) );
  OAI21_X1 U17873 ( .B1(n14482), .B2(n14484), .A(n14483), .ZN(n15232) );
  AND2_X1 U17874 ( .A1(n15166), .A2(n14485), .ZN(n14487) );
  OR2_X1 U17875 ( .A1(n14487), .A2(n14486), .ZN(n15617) );
  INV_X1 U17876 ( .A(n15617), .ZN(n14493) );
  OAI22_X1 U17877 ( .A1(n15284), .A2(n19436), .B1(n19322), .B2(n14488), .ZN(
        n14492) );
  INV_X1 U17878 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14490) );
  INV_X1 U17879 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n14489) );
  OAI22_X1 U17880 ( .A1(n15287), .A2(n14490), .B1(n19284), .B2(n14489), .ZN(
        n14491) );
  AOI211_X1 U17881 ( .C1(n19339), .C2(n14493), .A(n14492), .B(n14491), .ZN(
        n14494) );
  OAI21_X1 U17882 ( .B1(n15232), .B2(n19324), .A(n14494), .ZN(P2_U2898) );
  NOR2_X1 U17883 ( .A1(n14471), .A2(n14496), .ZN(n14497) );
  OR2_X1 U17884 ( .A1(n14495), .A2(n14497), .ZN(n16130) );
  OAI22_X1 U17885 ( .A1(n14780), .A2(n20258), .B1(n14748), .B2(n13842), .ZN(
        n14498) );
  AOI21_X1 U17886 ( .B1(n14782), .B2(BUF1_REG_17__SCAN_IN), .A(n14498), .ZN(
        n14500) );
  NAND2_X1 U17887 ( .A1(n13035), .A2(DATAI_17_), .ZN(n14499) );
  OAI211_X1 U17888 ( .C1(n16130), .C2(n14785), .A(n14500), .B(n14499), .ZN(
        P1_U2887) );
  AOI21_X1 U17889 ( .B1(n14501), .B2(n14483), .A(n11471), .ZN(n14502) );
  INV_X1 U17890 ( .A(n14502), .ZN(n15228) );
  INV_X1 U17891 ( .A(n15143), .ZN(n14508) );
  OAI22_X1 U17892 ( .A1(n15284), .A2(n19320), .B1(n19322), .B2(n14503), .ZN(
        n14507) );
  INV_X1 U17893 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14505) );
  INV_X1 U17894 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n14504) );
  OAI22_X1 U17895 ( .A1(n15287), .A2(n14505), .B1(n19284), .B2(n14504), .ZN(
        n14506) );
  AOI211_X1 U17896 ( .C1(n19339), .C2(n14508), .A(n14507), .B(n14506), .ZN(
        n14509) );
  OAI21_X1 U17897 ( .B1(n15228), .B2(n19324), .A(n14509), .ZN(P2_U2897) );
  NAND2_X1 U17898 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14510) );
  OAI211_X1 U17899 ( .C1(n20219), .C2(n14512), .A(n14511), .B(n14510), .ZN(
        n14513) );
  AOI21_X1 U17900 ( .B1(n14576), .B2(n13942), .A(n14513), .ZN(n14514) );
  OAI21_X1 U17901 ( .B1(n14515), .B2(n20220), .A(n14514), .ZN(P1_U2968) );
  AOI22_X1 U17902 ( .A1(n20113), .A2(n20148), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14707), .ZN(n14516) );
  OAI21_X1 U17903 ( .B1(n14517), .B2(n14728), .A(n14516), .ZN(P1_U2869) );
  AOI22_X1 U17904 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14518) );
  OAI21_X1 U17905 ( .B1(n20219), .B2(n20130), .A(n14518), .ZN(n14519) );
  AOI21_X1 U17906 ( .B1(n20137), .B2(n13942), .A(n14519), .ZN(n14520) );
  OAI21_X1 U17907 ( .B1(n14521), .B2(n20220), .A(n14520), .ZN(P1_U2997) );
  OAI22_X1 U17908 ( .A1(n20125), .A2(n14727), .B1(n14522), .B2(n20153), .ZN(
        n14523) );
  AOI21_X1 U17909 ( .B1(n20137), .B2(n20149), .A(n14523), .ZN(n14524) );
  INV_X1 U17910 ( .A(n14524), .ZN(P1_U2870) );
  NAND2_X1 U17911 ( .A1(n13900), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14526) );
  OAI21_X1 U17912 ( .B1(n14525), .B2(n13900), .A(n14526), .ZN(P2_U2856) );
  NOR2_X1 U17913 ( .A1(n19242), .A2(n19928), .ZN(n19275) );
  NAND2_X1 U17914 ( .A1(n14527), .A2(n19275), .ZN(n14534) );
  INV_X1 U17915 ( .A(n19270), .ZN(n19255) );
  AOI22_X1 U17916 ( .A1(n19264), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19279), .ZN(n14530) );
  NAND2_X1 U17917 ( .A1(n19265), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14529) );
  OAI211_X1 U17918 ( .C1(n14528), .C2(n19258), .A(n14530), .B(n14529), .ZN(
        n14531) );
  AOI21_X1 U17919 ( .B1(n14532), .B2(n19255), .A(n14531), .ZN(n14533) );
  AOI22_X1 U17920 ( .A1(n14556), .A2(n20148), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14707), .ZN(n14536) );
  OAI21_X1 U17921 ( .B1(n14535), .B2(n14728), .A(n14536), .ZN(P1_U2843) );
  INV_X1 U17922 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n16312) );
  NAND3_X1 U17923 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n16146) );
  NOR2_X1 U17924 ( .A1(n16312), .A2(n16146), .ZN(n14669) );
  NAND4_X1 U17925 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14669), .A3(
        P1_REIP_REG_15__SCAN_IN), .A4(P1_REIP_REG_16__SCAN_IN), .ZN(n14663) );
  NOR2_X1 U17926 ( .A1(n14537), .A2(n14663), .ZN(n14661) );
  NAND3_X1 U17927 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .ZN(n14538) );
  NOR2_X1 U17928 ( .A1(n14539), .A2(n14538), .ZN(n14540) );
  AND3_X1 U17929 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n16098) );
  AND2_X1 U17930 ( .A1(n14540), .A2(n16098), .ZN(n14541) );
  AND2_X1 U17931 ( .A1(n14661), .A2(n14541), .ZN(n14645) );
  OR2_X1 U17932 ( .A1(n20118), .A2(n14645), .ZN(n14542) );
  NAND2_X1 U17933 ( .A1(n14542), .A2(n20116), .ZN(n16083) );
  NOR2_X1 U17934 ( .A1(n20118), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14543) );
  OR2_X1 U17935 ( .A1(n16083), .A2(n14543), .ZN(n14638) );
  AND2_X1 U17936 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14547) );
  NOR2_X1 U17937 ( .A1(n20118), .A2(n14547), .ZN(n14544) );
  NOR2_X1 U17938 ( .A1(n14638), .A2(n14544), .ZN(n14623) );
  NAND2_X1 U17939 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14549) );
  NAND2_X1 U17940 ( .A1(n16166), .A2(n14549), .ZN(n14545) );
  AND2_X1 U17941 ( .A1(n14623), .A2(n14545), .ZN(n14603) );
  NOR2_X1 U17942 ( .A1(n14603), .A2(n14546), .ZN(n14555) );
  INV_X1 U17943 ( .A(n14547), .ZN(n14548) );
  NAND2_X1 U17944 ( .A1(n14645), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14634) );
  OR3_X1 U17945 ( .A1(n20118), .A2(n14548), .A3(n14634), .ZN(n14614) );
  NOR2_X1 U17946 ( .A1(n14614), .A2(n14549), .ZN(n14586) );
  INV_X1 U17947 ( .A(n14586), .ZN(n14553) );
  AOI22_X1 U17948 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20128), .B1(
        n20131), .B2(n14550), .ZN(n14552) );
  NAND2_X1 U17949 ( .A1(n20133), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14551) );
  OAI211_X1 U17950 ( .C1(n14553), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14552), 
        .B(n14551), .ZN(n14554) );
  AOI211_X1 U17951 ( .C1(n14556), .C2(n20127), .A(n14555), .B(n14554), .ZN(
        n14557) );
  OAI21_X1 U17952 ( .B1(n14535), .B2(n16182), .A(n14557), .ZN(P1_U2811) );
  OAI22_X1 U17953 ( .A1(n14780), .A2(n20196), .B1(n14748), .B2(n13844), .ZN(
        n14558) );
  AOI21_X1 U17954 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14782), .A(n14558), .ZN(
        n14560) );
  NAND2_X1 U17955 ( .A1(n13035), .A2(DATAI_29_), .ZN(n14559) );
  OAI211_X1 U17956 ( .C1(n14535), .C2(n14785), .A(n14560), .B(n14559), .ZN(
        P1_U2875) );
  AOI22_X1 U17957 ( .A1(n12196), .A2(n14561), .B1(n14569), .B2(n14567), .ZN(
        n14564) );
  NAND2_X1 U17958 ( .A1(n14565), .A2(n14562), .ZN(n14563) );
  OAI211_X1 U17959 ( .C1(n14566), .C2(n14565), .A(n14564), .B(n14563), .ZN(
        n16038) );
  OR2_X1 U17960 ( .A1(n14568), .A2(n14567), .ZN(n14571) );
  NAND2_X1 U17961 ( .A1(n14569), .A2(n14573), .ZN(n14570) );
  AND2_X1 U17962 ( .A1(n14571), .A2(n14570), .ZN(n20056) );
  NAND3_X1 U17963 ( .A1(n14573), .A2(n16073), .A3(n14572), .ZN(n14574) );
  NAND2_X1 U17964 ( .A1(n14574), .A2(n21018), .ZN(n21010) );
  NAND2_X1 U17965 ( .A1(n20056), .A2(n21010), .ZN(n16036) );
  AND2_X1 U17966 ( .A1(n16036), .A2(n14575), .ZN(n20064) );
  MUX2_X1 U17967 ( .A(P1_MORE_REG_SCAN_IN), .B(n16038), .S(n20064), .Z(
        P1_U3484) );
  AND2_X1 U17968 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14577) );
  OAI21_X1 U17969 ( .B1(n14577), .B2(n16099), .A(n14603), .ZN(n14585) );
  INV_X1 U17970 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14578) );
  NAND4_X1 U17971 ( .A1(n14586), .A2(P1_REIP_REG_30__SCAN_IN), .A3(
        P1_REIP_REG_29__SCAN_IN), .A4(n14578), .ZN(n14580) );
  AOI22_X1 U17972 ( .A1(n20133), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20128), .ZN(n14579) );
  NAND2_X1 U17973 ( .A1(n14580), .A2(n14579), .ZN(n14581) );
  AOI21_X1 U17974 ( .B1(n14585), .B2(P1_REIP_REG_31__SCAN_IN), .A(n14581), 
        .ZN(n14582) );
  OAI211_X1 U17975 ( .C1(n14685), .C2(n16168), .A(n14583), .B(n14582), .ZN(
        P1_U2809) );
  NAND2_X1 U17976 ( .A1(n14794), .A2(n20099), .ZN(n14592) );
  INV_X1 U17977 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14584) );
  OAI22_X1 U17978 ( .A1(n14584), .A2(n20094), .B1(n16178), .B2(n14792), .ZN(
        n14590) );
  INV_X1 U17979 ( .A(n14585), .ZN(n14588) );
  AOI21_X1 U17980 ( .B1(n14586), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14587) );
  NOR2_X1 U17981 ( .A1(n14588), .A2(n14587), .ZN(n14589) );
  AOI211_X1 U17982 ( .C1(n20133), .C2(P1_EBX_REG_30__SCAN_IN), .A(n14590), .B(
        n14589), .ZN(n14591) );
  OAI211_X1 U17983 ( .C1(n16168), .C2(n14913), .A(n14592), .B(n14591), .ZN(
        P1_U2810) );
  BUF_X1 U17984 ( .A(n14593), .Z(n14607) );
  AOI21_X1 U17985 ( .B1(n14594), .B2(n14607), .A(n12875), .ZN(n14805) );
  INV_X1 U17986 ( .A(n14805), .ZN(n14736) );
  AND2_X1 U17987 ( .A1(n14609), .A2(n14595), .ZN(n14596) );
  NOR2_X1 U17988 ( .A1(n14597), .A2(n14596), .ZN(n14925) );
  INV_X1 U17989 ( .A(n14614), .ZN(n14598) );
  AOI21_X1 U17990 ( .B1(n14598), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14602) );
  INV_X1 U17991 ( .A(n14803), .ZN(n14599) );
  AOI22_X1 U17992 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20128), .B1(
        n20131), .B2(n14599), .ZN(n14601) );
  NAND2_X1 U17993 ( .A1(n20133), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14600) );
  OAI211_X1 U17994 ( .C1(n14603), .C2(n14602), .A(n14601), .B(n14600), .ZN(
        n14604) );
  AOI21_X1 U17995 ( .B1(n14925), .B2(n20127), .A(n14604), .ZN(n14605) );
  OAI21_X1 U17996 ( .B1(n14736), .B2(n16182), .A(n14605), .ZN(P1_U2812) );
  OAI21_X2 U17997 ( .B1(n14606), .B2(n14608), .A(n14607), .ZN(n14811) );
  INV_X1 U17998 ( .A(n14609), .ZN(n14610) );
  AOI21_X1 U17999 ( .B1(n14611), .B2(n14627), .A(n14610), .ZN(n16259) );
  INV_X1 U18000 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n16262) );
  NOR2_X1 U18001 ( .A1(n14623), .A2(n16262), .ZN(n14616) );
  AOI22_X1 U18002 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20128), .B1(
        n20131), .B2(n14814), .ZN(n14613) );
  NAND2_X1 U18003 ( .A1(n20133), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n14612) );
  OAI211_X1 U18004 ( .C1(n14614), .C2(P1_REIP_REG_27__SCAN_IN), .A(n14613), 
        .B(n14612), .ZN(n14615) );
  AOI211_X1 U18005 ( .C1(n16259), .C2(n20127), .A(n14616), .B(n14615), .ZN(
        n14617) );
  OAI21_X1 U18006 ( .B1(n14811), .B2(n16182), .A(n14617), .ZN(P1_U2813) );
  INV_X1 U18007 ( .A(n14606), .ZN(n14619) );
  OAI21_X1 U18008 ( .B1(n14620), .B2(n14618), .A(n14619), .ZN(n14824) );
  OAI22_X1 U18009 ( .A1(n14621), .A2(n20094), .B1(n16178), .B2(n14817), .ZN(
        n14626) );
  INV_X1 U18010 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14816) );
  INV_X1 U18011 ( .A(n20118), .ZN(n20139) );
  INV_X1 U18012 ( .A(n14634), .ZN(n14622) );
  NAND3_X1 U18013 ( .A1(n20139), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14622), 
        .ZN(n14624) );
  AOI21_X1 U18014 ( .B1(n14816), .B2(n14624), .A(n14623), .ZN(n14625) );
  AOI211_X1 U18015 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n20133), .A(n14626), .B(
        n14625), .ZN(n14631) );
  AOI21_X1 U18016 ( .B1(n14629), .B2(n14628), .A(n10068), .ZN(n14937) );
  NAND2_X1 U18017 ( .A1(n14937), .A2(n20127), .ZN(n14630) );
  OAI211_X1 U18018 ( .C1(n14824), .C2(n16182), .A(n14631), .B(n14630), .ZN(
        P1_U2814) );
  INV_X1 U18019 ( .A(n14632), .ZN(n14642) );
  AOI21_X1 U18020 ( .B1(n14633), .B2(n14642), .A(n14618), .ZN(n14825) );
  NAND2_X1 U18021 ( .A1(n14825), .A2(n20099), .ZN(n14640) );
  NOR3_X1 U18022 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n20118), .A3(n14634), 
        .ZN(n14637) );
  AOI22_X1 U18023 ( .A1(P1_EBX_REG_25__SCAN_IN), .A2(n20133), .B1(n20131), 
        .B2(n14828), .ZN(n14635) );
  OAI21_X1 U18024 ( .B1(n14826), .B2(n20094), .A(n14635), .ZN(n14636) );
  AOI211_X1 U18025 ( .C1(n14638), .C2(P1_REIP_REG_25__SCAN_IN), .A(n14637), 
        .B(n14636), .ZN(n14639) );
  OAI211_X1 U18026 ( .C1(n16168), .C2(n14689), .A(n14640), .B(n14639), .ZN(
        P1_U2815) );
  AOI21_X1 U18027 ( .B1(n14643), .B2(n14693), .A(n14632), .ZN(n14838) );
  INV_X1 U18028 ( .A(n14838), .ZN(n14752) );
  INV_X1 U18029 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14644) );
  NAND3_X1 U18030 ( .A1(n20139), .A2(n14645), .A3(n14644), .ZN(n14648) );
  INV_X1 U18031 ( .A(n14836), .ZN(n14646) );
  AOI22_X1 U18032 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20128), .B1(
        n20131), .B2(n14646), .ZN(n14647) );
  OAI211_X1 U18033 ( .C1(n20095), .C2(n14691), .A(n14648), .B(n14647), .ZN(
        n14653) );
  INV_X1 U18034 ( .A(n14649), .ZN(n14650) );
  OAI21_X1 U18035 ( .B1(n14696), .B2(n14651), .A(n14650), .ZN(n14944) );
  NOR2_X1 U18036 ( .A1(n14944), .A2(n16168), .ZN(n14652) );
  AOI211_X1 U18037 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n16083), .A(n14653), 
        .B(n14652), .ZN(n14654) );
  OAI21_X1 U18038 ( .B1(n14752), .B2(n16182), .A(n14654), .ZN(P1_U2816) );
  INV_X1 U18039 ( .A(n14656), .ZN(n14712) );
  AOI21_X1 U18040 ( .B1(n14657), .B2(n14655), .A(n14656), .ZN(n14854) );
  INV_X1 U18041 ( .A(n14854), .ZN(n14778) );
  NOR2_X1 U18042 ( .A1(n14720), .A2(n14658), .ZN(n14659) );
  OR2_X1 U18043 ( .A1(n14710), .A2(n14659), .ZN(n14715) );
  INV_X1 U18044 ( .A(n14715), .ZN(n16287) );
  AOI21_X1 U18045 ( .B1(n14661), .B2(n14660), .A(n16099), .ZN(n14662) );
  INV_X1 U18046 ( .A(n14662), .ZN(n16135) );
  NOR2_X1 U18047 ( .A1(n14663), .A2(n16174), .ZN(n16084) );
  INV_X1 U18048 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20963) );
  NAND2_X1 U18049 ( .A1(n16084), .A2(n20963), .ZN(n16121) );
  INV_X1 U18050 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20966) );
  AOI21_X1 U18051 ( .B1(n16135), .B2(n16121), .A(n20966), .ZN(n14667) );
  NAND2_X1 U18052 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n16084), .ZN(n16112) );
  AOI21_X1 U18053 ( .B1(n20128), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20232), .ZN(n14665) );
  AOI22_X1 U18054 ( .A1(n20133), .A2(P1_EBX_REG_19__SCAN_IN), .B1(n20131), 
        .B2(n14857), .ZN(n14664) );
  OAI211_X1 U18055 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(n16112), .A(n14665), 
        .B(n14664), .ZN(n14666) );
  AOI211_X1 U18056 ( .C1(n16287), .C2(n20127), .A(n14667), .B(n14666), .ZN(
        n14668) );
  OAI21_X1 U18057 ( .B1(n14778), .B2(n16182), .A(n14668), .ZN(P1_U2821) );
  NOR3_X1 U18058 ( .A1(n16312), .A2(n16146), .A3(n16174), .ZN(n16136) );
  INV_X1 U18059 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21267) );
  OAI22_X1 U18060 ( .A1(n14884), .A2(n16178), .B1(n16168), .B2(n14987), .ZN(
        n14673) );
  INV_X1 U18061 ( .A(n14669), .ZN(n14670) );
  OAI21_X1 U18062 ( .B1(n14670), .B2(n16165), .A(n16166), .ZN(n16154) );
  AOI22_X1 U18063 ( .A1(n20133), .A2(P1_EBX_REG_15__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20128), .ZN(n14671) );
  OAI211_X1 U18064 ( .C1(n21267), .C2(n16154), .A(n14671), .B(n20100), .ZN(
        n14672) );
  AOI211_X1 U18065 ( .C1(n16136), .C2(n21267), .A(n14673), .B(n14672), .ZN(
        n14674) );
  OAI21_X1 U18066 ( .B1(n14888), .B2(n16182), .A(n14674), .ZN(P1_U2825) );
  OAI21_X1 U18067 ( .B1(n16099), .B2(n20080), .A(n14675), .ZN(n20085) );
  OAI22_X1 U18068 ( .A1(n14676), .A2(n16178), .B1(n16168), .B2(n16342), .ZN(
        n14681) );
  NAND2_X1 U18069 ( .A1(n20106), .A2(n20951), .ZN(n14678) );
  AOI22_X1 U18070 ( .A1(n20133), .A2(P1_EBX_REG_8__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20128), .ZN(n14677) );
  OAI211_X1 U18071 ( .C1(n14679), .C2(n14678), .A(n14677), .B(n20100), .ZN(
        n14680) );
  AOI211_X1 U18072 ( .C1(P1_REIP_REG_8__SCAN_IN), .C2(n20085), .A(n14681), .B(
        n14680), .ZN(n14682) );
  OAI21_X1 U18073 ( .B1(n14683), .B2(n16182), .A(n14682), .ZN(P1_U2832) );
  INV_X1 U18074 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14684) );
  OAI22_X1 U18075 ( .A1(n14685), .A2(n14727), .B1(n20153), .B2(n14684), .ZN(
        P1_U2841) );
  AOI22_X1 U18076 ( .A1(n14925), .A2(n20148), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14707), .ZN(n14686) );
  OAI21_X1 U18077 ( .B1(n14736), .B2(n14728), .A(n14686), .ZN(P1_U2844) );
  AOI22_X1 U18078 ( .A1(n16259), .A2(n20148), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14707), .ZN(n14687) );
  OAI21_X1 U18079 ( .B1(n14811), .B2(n14728), .A(n14687), .ZN(P1_U2845) );
  AOI22_X1 U18080 ( .A1(n14937), .A2(n20148), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14707), .ZN(n14688) );
  OAI21_X1 U18081 ( .B1(n14824), .B2(n14728), .A(n14688), .ZN(P1_U2846) );
  INV_X1 U18082 ( .A(n14825), .ZN(n14746) );
  INV_X1 U18083 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14690) );
  OAI222_X1 U18084 ( .A1(n14728), .A2(n14746), .B1(n14690), .B2(n20153), .C1(
        n14689), .C2(n14727), .ZN(P1_U2847) );
  OAI222_X1 U18085 ( .A1(n14728), .A2(n14752), .B1(n14691), .B2(n20153), .C1(
        n14944), .C2(n14727), .ZN(P1_U2848) );
  OAI21_X1 U18086 ( .B1(n12743), .B2(n9828), .A(n14693), .ZN(n16088) );
  INV_X1 U18087 ( .A(n16096), .ZN(n14695) );
  AOI21_X1 U18088 ( .B1(n14695), .B2(n16095), .A(n14694), .ZN(n14697) );
  NOR2_X1 U18089 ( .A1(n14697), .A2(n14696), .ZN(n16272) );
  AOI22_X1 U18090 ( .A1(n16272), .A2(n20148), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14707), .ZN(n14698) );
  OAI21_X1 U18091 ( .B1(n16088), .B2(n14728), .A(n14698), .ZN(P1_U2849) );
  INV_X1 U18092 ( .A(n14699), .ZN(n14703) );
  INV_X1 U18093 ( .A(n14700), .ZN(n14702) );
  AOI21_X1 U18094 ( .B1(n14703), .B2(n14702), .A(n14701), .ZN(n16198) );
  INV_X1 U18095 ( .A(n16198), .ZN(n14766) );
  NAND2_X1 U18096 ( .A1(n14704), .A2(n14705), .ZN(n14706) );
  AND2_X1 U18097 ( .A1(n16096), .A2(n14706), .ZN(n16104) );
  AOI22_X1 U18098 ( .A1(n16104), .A2(n20148), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14707), .ZN(n14708) );
  OAI21_X1 U18099 ( .B1(n14766), .B2(n14728), .A(n14708), .ZN(P1_U2851) );
  OR2_X1 U18100 ( .A1(n14710), .A2(n14709), .ZN(n14711) );
  NAND2_X1 U18101 ( .A1(n14704), .A2(n14711), .ZN(n16117) );
  INV_X1 U18102 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14714) );
  AOI21_X1 U18103 ( .B1(n14713), .B2(n14712), .A(n14700), .ZN(n16203) );
  INV_X1 U18104 ( .A(n16203), .ZN(n14774) );
  OAI222_X1 U18105 ( .A1(n14727), .A2(n16117), .B1(n14714), .B2(n20153), .C1(
        n14774), .C2(n14728), .ZN(P1_U2852) );
  INV_X1 U18106 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14716) );
  OAI222_X1 U18107 ( .A1(n14728), .A2(n14778), .B1(n14716), .B2(n20153), .C1(
        n14715), .C2(n14727), .ZN(P1_U2853) );
  OR2_X1 U18108 ( .A1(n14495), .A2(n14717), .ZN(n14718) );
  AND2_X1 U18109 ( .A1(n14655), .A2(n14718), .ZN(n16124) );
  AND2_X1 U18110 ( .A1(n9786), .A2(n14719), .ZN(n14721) );
  OR2_X1 U18111 ( .A1(n14721), .A2(n14720), .ZN(n16298) );
  OAI22_X1 U18112 ( .A1(n16298), .A2(n14727), .B1(n16119), .B2(n20153), .ZN(
        n14722) );
  AOI21_X1 U18113 ( .B1(n16124), .B2(n20149), .A(n14722), .ZN(n14723) );
  INV_X1 U18114 ( .A(n14723), .ZN(P1_U2854) );
  INV_X1 U18115 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n16126) );
  NAND2_X1 U18116 ( .A1(n14725), .A2(n14724), .ZN(n14726) );
  AND2_X1 U18117 ( .A1(n9786), .A2(n14726), .ZN(n16306) );
  INV_X1 U18118 ( .A(n16306), .ZN(n16129) );
  OAI222_X1 U18119 ( .A1(n14728), .A2(n16130), .B1(n20153), .B2(n16126), .C1(
        n16129), .C2(n14727), .ZN(P1_U2855) );
  OAI22_X1 U18120 ( .A1(n14780), .A2(n20199), .B1(n14748), .B2(n13677), .ZN(
        n14729) );
  AOI21_X1 U18121 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14782), .A(n14729), .ZN(
        n14731) );
  NAND2_X1 U18122 ( .A1(n13035), .A2(DATAI_30_), .ZN(n14730) );
  OAI211_X1 U18123 ( .C1(n14732), .C2(n14785), .A(n14731), .B(n14730), .ZN(
        P1_U2874) );
  OAI22_X1 U18124 ( .A1(n14780), .A2(n20193), .B1(n14748), .B2(n13671), .ZN(
        n14733) );
  AOI21_X1 U18125 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14782), .A(n14733), .ZN(
        n14735) );
  NAND2_X1 U18126 ( .A1(n13035), .A2(DATAI_28_), .ZN(n14734) );
  OAI211_X1 U18127 ( .C1(n14736), .C2(n14785), .A(n14735), .B(n14734), .ZN(
        P1_U2876) );
  OAI22_X1 U18128 ( .A1(n14780), .A2(n20190), .B1(n14748), .B2(n13675), .ZN(
        n14737) );
  AOI21_X1 U18129 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14782), .A(n14737), .ZN(
        n14739) );
  NAND2_X1 U18130 ( .A1(n13035), .A2(DATAI_27_), .ZN(n14738) );
  OAI211_X1 U18131 ( .C1(n14811), .C2(n14785), .A(n14739), .B(n14738), .ZN(
        P1_U2877) );
  INV_X1 U18132 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16590) );
  INV_X1 U18133 ( .A(n14780), .ZN(n14769) );
  AOI22_X1 U18134 ( .A1(n14769), .A2(n20188), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n14767), .ZN(n14740) );
  OAI21_X1 U18135 ( .B1(n16590), .B2(n14771), .A(n14740), .ZN(n14741) );
  AOI21_X1 U18136 ( .B1(n13035), .B2(DATAI_26_), .A(n14741), .ZN(n14742) );
  OAI21_X1 U18137 ( .B1(n14824), .B2(n14785), .A(n14742), .ZN(P1_U2878) );
  OAI22_X1 U18138 ( .A1(n14780), .A2(n20184), .B1(n14748), .B2(n13654), .ZN(
        n14743) );
  AOI21_X1 U18139 ( .B1(BUF1_REG_25__SCAN_IN), .B2(n14782), .A(n14743), .ZN(
        n14745) );
  NAND2_X1 U18140 ( .A1(n13035), .A2(DATAI_25_), .ZN(n14744) );
  OAI211_X1 U18141 ( .C1(n14746), .C2(n14785), .A(n14745), .B(n14744), .ZN(
        P1_U2879) );
  OAI22_X1 U18142 ( .A1(n14780), .A2(n20181), .B1(n14748), .B2(n14747), .ZN(
        n14749) );
  AOI21_X1 U18143 ( .B1(n14782), .B2(BUF1_REG_24__SCAN_IN), .A(n14749), .ZN(
        n14751) );
  NAND2_X1 U18144 ( .A1(n13035), .A2(DATAI_24_), .ZN(n14750) );
  OAI211_X1 U18145 ( .C1(n14752), .C2(n14785), .A(n14751), .B(n14750), .ZN(
        P1_U2880) );
  OAI22_X1 U18146 ( .A1(n14780), .A2(n20291), .B1(n14748), .B2(n13679), .ZN(
        n14753) );
  AOI21_X1 U18147 ( .B1(n14782), .B2(BUF1_REG_23__SCAN_IN), .A(n14753), .ZN(
        n14755) );
  NAND2_X1 U18148 ( .A1(n13035), .A2(DATAI_23_), .ZN(n14754) );
  OAI211_X1 U18149 ( .C1(n16088), .C2(n14785), .A(n14755), .B(n14754), .ZN(
        P1_U2881) );
  OR2_X1 U18150 ( .A1(n14701), .A2(n14756), .ZN(n14757) );
  AND2_X1 U18151 ( .A1(n14692), .A2(n14757), .ZN(n16193) );
  INV_X1 U18152 ( .A(n16193), .ZN(n14762) );
  AOI22_X1 U18153 ( .A1(n14769), .A2(n14758), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n14767), .ZN(n14759) );
  OAI21_X1 U18154 ( .B1(n14505), .B2(n14771), .A(n14759), .ZN(n14760) );
  AOI21_X1 U18155 ( .B1(n13035), .B2(DATAI_22_), .A(n14760), .ZN(n14761) );
  OAI21_X1 U18156 ( .B1(n14762), .B2(n14785), .A(n14761), .ZN(P1_U2882) );
  OAI22_X1 U18157 ( .A1(n14780), .A2(n20277), .B1(n14748), .B2(n13848), .ZN(
        n14763) );
  AOI21_X1 U18158 ( .B1(n14782), .B2(BUF1_REG_21__SCAN_IN), .A(n14763), .ZN(
        n14765) );
  NAND2_X1 U18159 ( .A1(n13035), .A2(DATAI_21_), .ZN(n14764) );
  OAI211_X1 U18160 ( .C1(n14766), .C2(n14785), .A(n14765), .B(n14764), .ZN(
        P1_U2883) );
  INV_X1 U18161 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16598) );
  AOI22_X1 U18162 ( .A1(n14769), .A2(n14768), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n14767), .ZN(n14770) );
  OAI21_X1 U18163 ( .B1(n16598), .B2(n14771), .A(n14770), .ZN(n14772) );
  AOI21_X1 U18164 ( .B1(n13035), .B2(DATAI_20_), .A(n14772), .ZN(n14773) );
  OAI21_X1 U18165 ( .B1(n14774), .B2(n14785), .A(n14773), .ZN(P1_U2884) );
  OAI22_X1 U18166 ( .A1(n14780), .A2(n20267), .B1(n14748), .B2(n13840), .ZN(
        n14775) );
  AOI21_X1 U18167 ( .B1(n14782), .B2(BUF1_REG_19__SCAN_IN), .A(n14775), .ZN(
        n14777) );
  NAND2_X1 U18168 ( .A1(n13035), .A2(DATAI_19_), .ZN(n14776) );
  OAI211_X1 U18169 ( .C1(n14778), .C2(n14785), .A(n14777), .B(n14776), .ZN(
        P1_U2885) );
  INV_X1 U18170 ( .A(n16124), .ZN(n14786) );
  OAI22_X1 U18171 ( .A1(n14780), .A2(n20263), .B1(n14748), .B2(n14779), .ZN(
        n14781) );
  AOI21_X1 U18172 ( .B1(n14782), .B2(BUF1_REG_18__SCAN_IN), .A(n14781), .ZN(
        n14784) );
  NAND2_X1 U18173 ( .A1(n13035), .A2(DATAI_18_), .ZN(n14783) );
  OAI211_X1 U18174 ( .C1(n14786), .C2(n14785), .A(n14784), .B(n14783), .ZN(
        P1_U2886) );
  NAND2_X1 U18175 ( .A1(n14788), .A2(n14787), .ZN(n14789) );
  XNOR2_X1 U18176 ( .A(n14789), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14921) );
  INV_X1 U18177 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14790) );
  NOR2_X1 U18178 ( .A1(n20100), .A2(n14790), .ZN(n14914) );
  AOI21_X1 U18179 ( .B1(n20228), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14914), .ZN(n14791) );
  OAI21_X1 U18180 ( .B1(n20219), .B2(n14792), .A(n14791), .ZN(n14793) );
  AOI21_X1 U18181 ( .B1(n14794), .B2(n13942), .A(n14793), .ZN(n14795) );
  OAI21_X1 U18182 ( .B1(n14921), .B2(n20220), .A(n14795), .ZN(P1_U2969) );
  NAND2_X1 U18183 ( .A1(n12088), .A2(n14796), .ZN(n14819) );
  NAND2_X1 U18184 ( .A1(n14841), .A2(n14819), .ZN(n14800) );
  OAI21_X1 U18185 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14797), .A(
        n14800), .ZN(n14799) );
  INV_X1 U18186 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16264) );
  MUX2_X1 U18187 ( .A(n16264), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n12088), .Z(n14798) );
  OAI211_X1 U18188 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14800), .A(
        n14799), .B(n14798), .ZN(n14801) );
  XOR2_X1 U18189 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14801), .Z(
        n14931) );
  NAND2_X1 U18190 ( .A1(n20232), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14926) );
  NAND2_X1 U18191 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14802) );
  OAI211_X1 U18192 ( .C1(n20219), .C2(n14803), .A(n14926), .B(n14802), .ZN(
        n14804) );
  AOI21_X1 U18193 ( .B1(n14805), .B2(n13942), .A(n14804), .ZN(n14806) );
  OAI21_X1 U18194 ( .B1(n20220), .B2(n14931), .A(n14806), .ZN(P1_U2971) );
  MUX2_X1 U18195 ( .A(n14808), .B(n14807), .S(n9721), .Z(n14809) );
  OAI22_X1 U18196 ( .A1(n16256), .A2(n14810), .B1(n20100), .B2(n16262), .ZN(
        n14813) );
  NOR2_X1 U18197 ( .A1(n14811), .A2(n20238), .ZN(n14812) );
  OAI21_X1 U18198 ( .B1(n20220), .B2(n16258), .A(n14815), .ZN(P1_U2972) );
  NOR2_X1 U18199 ( .A1(n20100), .A2(n14816), .ZN(n14936) );
  NOR2_X1 U18200 ( .A1(n20219), .A2(n14817), .ZN(n14818) );
  AOI211_X1 U18201 ( .C1(n20228), .C2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14936), .B(n14818), .ZN(n14823) );
  OAI211_X1 U18202 ( .C1(n9721), .C2(n14841), .A(n14820), .B(n14819), .ZN(
        n14821) );
  XNOR2_X1 U18203 ( .A(n14821), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14932) );
  NAND2_X1 U18204 ( .A1(n14932), .A2(n20230), .ZN(n14822) );
  OAI211_X1 U18205 ( .C1(n14824), .C2(n20238), .A(n14823), .B(n14822), .ZN(
        P1_U2973) );
  NAND2_X1 U18206 ( .A1(n14825), .A2(n13942), .ZN(n14830) );
  INV_X1 U18207 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20973) );
  OAI22_X1 U18208 ( .A1(n16256), .A2(n14826), .B1(n20100), .B2(n20973), .ZN(
        n14827) );
  AOI21_X1 U18209 ( .B1(n16252), .B2(n14828), .A(n14827), .ZN(n14829) );
  OAI211_X1 U18210 ( .C1(n14831), .C2(n20220), .A(n14830), .B(n14829), .ZN(
        P1_U2974) );
  MUX2_X1 U18211 ( .A(n9721), .B(n14840), .S(n14832), .Z(n14834) );
  XNOR2_X1 U18212 ( .A(n14834), .B(n14833), .ZN(n14950) );
  AOI22_X1 U18213 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n14835) );
  OAI21_X1 U18214 ( .B1(n20219), .B2(n14836), .A(n14835), .ZN(n14837) );
  AOI21_X1 U18215 ( .B1(n14838), .B2(n13942), .A(n14837), .ZN(n14839) );
  OAI21_X1 U18216 ( .B1(n14950), .B2(n20220), .A(n14839), .ZN(P1_U2975) );
  INV_X1 U18217 ( .A(n14840), .ZN(n14846) );
  NOR2_X1 U18218 ( .A1(n9721), .A2(n14845), .ZN(n14843) );
  MUX2_X1 U18219 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n14845), .S(
        n12088), .Z(n14842) );
  MUX2_X1 U18220 ( .A(n14843), .B(n14842), .S(n14841), .Z(n14844) );
  AOI21_X1 U18221 ( .B1(n14846), .B2(n14845), .A(n14844), .ZN(n16271) );
  INV_X1 U18222 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14847) );
  OAI22_X1 U18223 ( .A1(n16256), .A2(n16092), .B1(n20100), .B2(n14847), .ZN(
        n14849) );
  NOR2_X1 U18224 ( .A1(n16088), .A2(n20238), .ZN(n14848) );
  AOI211_X1 U18225 ( .C1(n16252), .C2(n16082), .A(n14849), .B(n14848), .ZN(
        n14850) );
  OAI21_X1 U18226 ( .B1(n16271), .B2(n20220), .A(n14850), .ZN(P1_U2976) );
  NOR2_X1 U18227 ( .A1(n12088), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14852) );
  MUX2_X1 U18228 ( .A(n12088), .B(n14852), .S(n14851), .Z(n14853) );
  XNOR2_X1 U18229 ( .A(n14853), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16286) );
  NAND2_X1 U18230 ( .A1(n14854), .A2(n13942), .ZN(n14859) );
  OAI22_X1 U18231 ( .A1(n16256), .A2(n14855), .B1(n20100), .B2(n20966), .ZN(
        n14856) );
  AOI21_X1 U18232 ( .B1(n16252), .B2(n14857), .A(n14856), .ZN(n14858) );
  OAI211_X1 U18233 ( .C1(n16286), .C2(n20220), .A(n14859), .B(n14858), .ZN(
        P1_U2980) );
  OAI21_X1 U18234 ( .B1(n14861), .B2(n14860), .A(n14851), .ZN(n16299) );
  AOI22_X1 U18235 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14862) );
  OAI21_X1 U18236 ( .B1(n20219), .B2(n16118), .A(n14862), .ZN(n14863) );
  AOI21_X1 U18237 ( .B1(n16124), .B2(n13942), .A(n14863), .ZN(n14864) );
  OAI21_X1 U18238 ( .B1(n20220), .B2(n16299), .A(n14864), .ZN(P1_U2981) );
  NOR2_X1 U18239 ( .A1(n12088), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14870) );
  INV_X1 U18240 ( .A(n14866), .ZN(n14867) );
  NAND2_X1 U18241 ( .A1(n14903), .A2(n14867), .ZN(n16215) );
  OAI21_X1 U18242 ( .B1(n16215), .B2(n14965), .A(n14868), .ZN(n14869) );
  MUX2_X1 U18243 ( .A(n12088), .B(n14870), .S(n14869), .Z(n14872) );
  INV_X1 U18244 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14871) );
  XNOR2_X1 U18245 ( .A(n14872), .B(n14871), .ZN(n16307) );
  NAND2_X1 U18246 ( .A1(n16307), .A2(n20230), .ZN(n14876) );
  INV_X1 U18247 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14873) );
  OAI22_X1 U18248 ( .A1(n16256), .A2(n21087), .B1(n20100), .B2(n14873), .ZN(
        n14874) );
  AOI21_X1 U18249 ( .B1(n16128), .B2(n16252), .A(n14874), .ZN(n14875) );
  OAI211_X1 U18250 ( .C1(n20238), .C2(n16130), .A(n14876), .B(n14875), .ZN(
        P1_U2982) );
  INV_X1 U18251 ( .A(n16215), .ZN(n14878) );
  NOR2_X1 U18252 ( .A1(n14878), .A2(n14877), .ZN(n14966) );
  INV_X1 U18253 ( .A(n14966), .ZN(n14880) );
  NAND2_X1 U18254 ( .A1(n14880), .A2(n14879), .ZN(n14883) );
  NAND2_X1 U18255 ( .A1(n14881), .A2(n14964), .ZN(n14882) );
  XNOR2_X1 U18256 ( .A(n14883), .B(n14882), .ZN(n14986) );
  NAND2_X1 U18257 ( .A1(n14986), .A2(n20230), .ZN(n14887) );
  NOR2_X1 U18258 ( .A1(n20100), .A2(n21267), .ZN(n14991) );
  NOR2_X1 U18259 ( .A1(n20219), .A2(n14884), .ZN(n14885) );
  AOI211_X1 U18260 ( .C1(n20228), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n14991), .B(n14885), .ZN(n14886) );
  OAI211_X1 U18261 ( .C1(n20238), .C2(n14888), .A(n14887), .B(n14886), .ZN(
        P1_U2984) );
  INV_X1 U18262 ( .A(n14903), .ZN(n16227) );
  INV_X1 U18263 ( .A(n14889), .ZN(n14890) );
  AOI21_X1 U18264 ( .B1(n16227), .B2(n14891), .A(n14890), .ZN(n15010) );
  AND2_X1 U18265 ( .A1(n14892), .A2(n14893), .ZN(n15009) );
  NAND2_X1 U18266 ( .A1(n15010), .A2(n15009), .ZN(n15008) );
  NAND2_X1 U18267 ( .A1(n15008), .A2(n14893), .ZN(n14894) );
  XOR2_X1 U18268 ( .A(n14895), .B(n14894), .Z(n15005) );
  INV_X1 U18269 ( .A(n15005), .ZN(n14901) );
  AOI22_X1 U18270 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14896) );
  OAI21_X1 U18271 ( .B1(n20219), .B2(n14897), .A(n14896), .ZN(n14898) );
  AOI21_X1 U18272 ( .B1(n14899), .B2(n13942), .A(n14898), .ZN(n14900) );
  OAI21_X1 U18273 ( .B1(n14901), .B2(n20220), .A(n14900), .ZN(P1_U2986) );
  NAND2_X1 U18274 ( .A1(n14902), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14905) );
  XNOR2_X1 U18275 ( .A(n14903), .B(n14906), .ZN(n14904) );
  MUX2_X1 U18276 ( .A(n14905), .B(n14904), .S(n12088), .Z(n14908) );
  INV_X1 U18277 ( .A(n14902), .ZN(n14907) );
  NAND3_X1 U18278 ( .A1(n14907), .A2(n9721), .A3(n14906), .ZN(n16228) );
  NAND2_X1 U18279 ( .A1(n14908), .A2(n16228), .ZN(n15024) );
  NAND2_X1 U18280 ( .A1(n15024), .A2(n20230), .ZN(n14912) );
  INV_X1 U18281 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14909) );
  NOR2_X1 U18282 ( .A1(n20100), .A2(n14909), .ZN(n15029) );
  NOR2_X1 U18283 ( .A1(n20219), .A2(n16177), .ZN(n14910) );
  AOI211_X1 U18284 ( .C1(n20228), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15029), .B(n14910), .ZN(n14911) );
  OAI211_X1 U18285 ( .C1(n20238), .C2(n16183), .A(n14912), .B(n14911), .ZN(
        P1_U2989) );
  INV_X1 U18286 ( .A(n14913), .ZN(n14915) );
  AOI21_X1 U18287 ( .B1(n14915), .B2(n16367), .A(n14914), .ZN(n14920) );
  NAND2_X1 U18288 ( .A1(n14916), .A2(n12380), .ZN(n14917) );
  NAND2_X1 U18289 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  OAI211_X1 U18290 ( .C1(n14921), .C2(n16370), .A(n14920), .B(n14919), .ZN(
        P1_U3001) );
  INV_X1 U18291 ( .A(n14922), .ZN(n16266) );
  NOR3_X1 U18292 ( .A1(n14924), .A2(n14923), .A3(n16261), .ZN(n14929) );
  INV_X1 U18293 ( .A(n14925), .ZN(n14927) );
  OAI21_X1 U18294 ( .B1(n14927), .B2(n16341), .A(n14926), .ZN(n14928) );
  AOI211_X1 U18295 ( .C1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16266), .A(
        n14929), .B(n14928), .ZN(n14930) );
  OAI21_X1 U18296 ( .B1(n14931), .B2(n16370), .A(n14930), .ZN(P1_U3003) );
  INV_X1 U18297 ( .A(n14932), .ZN(n14940) );
  OAI22_X1 U18298 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n14935), .B1(
        n14934), .B2(n14933), .ZN(n14939) );
  AOI21_X1 U18299 ( .B1(n14937), .B2(n16367), .A(n14936), .ZN(n14938) );
  OAI211_X1 U18300 ( .C1(n14940), .C2(n16370), .A(n14939), .B(n14938), .ZN(
        P1_U3005) );
  NOR2_X1 U18301 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n14941), .ZN(
        n14943) );
  OAI21_X1 U18302 ( .B1(n14943), .B2(n14942), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14949) );
  INV_X1 U18303 ( .A(n14944), .ZN(n14947) );
  NOR2_X1 U18304 ( .A1(n20100), .A2(n14644), .ZN(n14946) );
  NOR3_X1 U18305 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14845), .A3(
        n16269), .ZN(n14945) );
  AOI211_X1 U18306 ( .C1(n14947), .C2(n16367), .A(n14946), .B(n14945), .ZN(
        n14948) );
  OAI211_X1 U18307 ( .C1(n14950), .C2(n16370), .A(n14949), .B(n14948), .ZN(
        P1_U3007) );
  NAND2_X1 U18308 ( .A1(n14951), .A2(n9721), .ZN(n16066) );
  NAND2_X1 U18309 ( .A1(n12088), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14952) );
  OR2_X1 U18310 ( .A1(n14851), .A2(n14952), .ZN(n16064) );
  NAND2_X1 U18311 ( .A1(n16066), .A2(n16064), .ZN(n14953) );
  XNOR2_X1 U18312 ( .A(n14953), .B(n16063), .ZN(n16202) );
  INV_X1 U18313 ( .A(n16202), .ZN(n14963) );
  NOR2_X1 U18314 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16292), .ZN(
        n14958) );
  NAND2_X1 U18315 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14998), .ZN(
        n14972) );
  OAI21_X1 U18316 ( .B1(n14974), .B2(n14972), .A(n14954), .ZN(n14978) );
  NAND2_X1 U18317 ( .A1(n14955), .A2(n14978), .ZN(n14959) );
  OAI21_X1 U18318 ( .B1(n14956), .B2(n14969), .A(n14959), .ZN(n16291) );
  INV_X1 U18319 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20965) );
  OAI22_X1 U18320 ( .A1(n16117), .A2(n16341), .B1(n20100), .B2(n20965), .ZN(
        n14957) );
  AOI21_X1 U18321 ( .B1(n14958), .B2(n16291), .A(n14957), .ZN(n14962) );
  OAI221_X1 U18322 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14969), 
        .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n14959), .A(n16289), .ZN(
        n14960) );
  NAND2_X1 U18323 ( .A1(n14960), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14961) );
  OAI211_X1 U18324 ( .C1(n14963), .C2(n16370), .A(n14962), .B(n14961), .ZN(
        P1_U3011) );
  OAI21_X1 U18325 ( .B1(n14966), .B2(n14965), .A(n14964), .ZN(n14968) );
  XNOR2_X1 U18326 ( .A(n14968), .B(n14967), .ZN(n16208) );
  NAND2_X1 U18327 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16304), .ZN(
        n14989) );
  NOR2_X1 U18328 ( .A1(n12102), .A2(n14989), .ZN(n14982) );
  NOR2_X1 U18329 ( .A1(n14970), .A2(n14969), .ZN(n14999) );
  OAI21_X1 U18330 ( .B1(n16318), .B2(n16333), .A(n14971), .ZN(n14976) );
  INV_X1 U18331 ( .A(n14972), .ZN(n14973) );
  NOR2_X1 U18332 ( .A1(n14974), .A2(n14973), .ZN(n14975) );
  OR2_X1 U18333 ( .A1(n14976), .A2(n14975), .ZN(n14977) );
  NOR2_X1 U18334 ( .A1(n14999), .A2(n14977), .ZN(n15003) );
  NAND2_X1 U18335 ( .A1(n15002), .A2(n14978), .ZN(n15001) );
  NAND2_X1 U18336 ( .A1(n15003), .A2(n15001), .ZN(n16315) );
  OAI22_X1 U18337 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n14989), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14979), .ZN(n14980) );
  NOR2_X1 U18338 ( .A1(n16315), .A2(n14980), .ZN(n14988) );
  INV_X1 U18339 ( .A(n14988), .ZN(n14981) );
  MUX2_X1 U18340 ( .A(n14982), .B(n14981), .S(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(n14984) );
  OAI22_X1 U18341 ( .A1(n16138), .A2(n16341), .B1(n20100), .B2(n21097), .ZN(
        n14983) );
  AOI211_X1 U18342 ( .C1(n16208), .C2(n16360), .A(n14984), .B(n14983), .ZN(
        n14985) );
  INV_X1 U18343 ( .A(n14985), .ZN(P1_U3015) );
  INV_X1 U18344 ( .A(n14986), .ZN(n14994) );
  INV_X1 U18345 ( .A(n14987), .ZN(n14992) );
  AOI21_X1 U18346 ( .B1(n12102), .B2(n14989), .A(n14988), .ZN(n14990) );
  AOI211_X1 U18347 ( .C1(n16367), .C2(n14992), .A(n14991), .B(n14990), .ZN(
        n14993) );
  OAI21_X1 U18348 ( .B1(n14994), .B2(n16370), .A(n14993), .ZN(P1_U3016) );
  INV_X1 U18349 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20957) );
  OR2_X1 U18350 ( .A1(n20100), .A2(n20957), .ZN(n14995) );
  OAI21_X1 U18351 ( .B1(n14996), .B2(n16341), .A(n14995), .ZN(n14997) );
  AOI21_X1 U18352 ( .B1(n14999), .B2(n14998), .A(n14997), .ZN(n15000) );
  OAI211_X1 U18353 ( .C1(n15003), .C2(n15002), .A(n15001), .B(n15000), .ZN(
        n15004) );
  AOI21_X1 U18354 ( .B1(n15005), .B2(n16360), .A(n15004), .ZN(n15006) );
  INV_X1 U18355 ( .A(n15006), .ZN(P1_U3018) );
  INV_X1 U18356 ( .A(n15007), .ZN(n16334) );
  NAND2_X1 U18357 ( .A1(n16334), .A2(n16316), .ZN(n16364) );
  NOR2_X1 U18358 ( .A1(n16364), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15021) );
  OAI21_X1 U18359 ( .B1(n15010), .B2(n15009), .A(n15008), .ZN(n15011) );
  INV_X1 U18360 ( .A(n15011), .ZN(n16226) );
  AOI221_X1 U18361 ( .B1(n15014), .B2(n16338), .C1(n15013), .C2(n16338), .A(
        n15012), .ZN(n15015) );
  OAI221_X1 U18362 ( .B1(n16333), .B2(n15020), .C1(n16333), .C2(n16334), .A(
        n15015), .ZN(n16327) );
  AOI21_X1 U18363 ( .B1(n15016), .B2(n16322), .A(n16327), .ZN(n15018) );
  OAI22_X1 U18364 ( .A1(n16226), .A2(n16370), .B1(n15018), .B2(n15017), .ZN(
        n15019) );
  AOI21_X1 U18365 ( .B1(n15021), .B2(n15020), .A(n15019), .ZN(n15023) );
  NAND2_X1 U18366 ( .A1(n20232), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15022) );
  OAI211_X1 U18367 ( .C1(n16341), .C2(n16158), .A(n15023), .B(n15022), .ZN(
        P1_U3019) );
  INV_X1 U18368 ( .A(n15024), .ZN(n15034) );
  AOI211_X1 U18369 ( .C1(n15027), .C2(n15026), .A(n15025), .B(n14906), .ZN(
        n15028) );
  AOI211_X1 U18370 ( .C1(n16367), .C2(n16180), .A(n15029), .B(n15028), .ZN(
        n15033) );
  AOI211_X1 U18371 ( .C1(n14906), .C2(n15030), .A(n16323), .B(n16331), .ZN(
        n15031) );
  INV_X1 U18372 ( .A(n15031), .ZN(n15032) );
  OAI211_X1 U18373 ( .C1(n15034), .C2(n16370), .A(n15033), .B(n15032), .ZN(
        P1_U3021) );
  INV_X1 U18374 ( .A(n13889), .ZN(n20721) );
  NOR2_X1 U18375 ( .A1(n20532), .A2(n20721), .ZN(n20480) );
  OAI21_X1 U18376 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20241), .A(n20637), 
        .ZN(n15037) );
  AOI21_X1 U18377 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20480), .A(n15037), 
        .ZN(n15042) );
  OR3_X1 U18378 ( .A1(n13889), .A2(n20760), .A3(n21012), .ZN(n20992) );
  INV_X1 U18379 ( .A(n20992), .ZN(n15039) );
  NAND2_X1 U18380 ( .A1(n20857), .A2(n15039), .ZN(n20766) );
  INV_X1 U18381 ( .A(n20994), .ZN(n15040) );
  NAND2_X1 U18382 ( .A1(n20563), .A2(n15040), .ZN(n15041) );
  OAI211_X1 U18383 ( .C1(n15042), .C2(n20760), .A(n20766), .B(n15041), .ZN(
        n15043) );
  MUX2_X1 U18384 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15043), .S(
        n20996), .Z(P1_U3475) );
  NOR2_X1 U18385 ( .A1(n15045), .A2(n15044), .ZN(n15047) );
  INV_X1 U18386 ( .A(n15047), .ZN(n15054) );
  AOI21_X1 U18387 ( .B1(n15048), .B2(n15047), .A(n15046), .ZN(n15049) );
  OAI21_X1 U18388 ( .B1(n14101), .B2(n15050), .A(n15049), .ZN(n16024) );
  NOR2_X1 U18389 ( .A1(n14021), .A2(n15051), .ZN(n15059) );
  OAI22_X1 U18390 ( .A1(n15052), .A2(n12212), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15057) );
  AOI22_X1 U18391 ( .A1(n16024), .A2(n15060), .B1(n15059), .B2(n15057), .ZN(
        n15053) );
  OAI21_X1 U18392 ( .B1(n15064), .B2(n15054), .A(n15053), .ZN(n15055) );
  MUX2_X1 U18393 ( .A(n15055), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15065), .Z(P1_U3473) );
  INV_X1 U18394 ( .A(n15056), .ZN(n15063) );
  INV_X1 U18395 ( .A(n15057), .ZN(n15058) );
  AOI22_X1 U18396 ( .A1(n15061), .A2(n15060), .B1(n15059), .B2(n15058), .ZN(
        n15062) );
  OAI21_X1 U18397 ( .B1(n15064), .B2(n15063), .A(n15062), .ZN(n15066) );
  MUX2_X1 U18398 ( .A(n15066), .B(n21244), .S(n15065), .Z(P1_U3472) );
  OAI21_X1 U18399 ( .B1(n15068), .B2(n19691), .A(n15067), .ZN(n15070) );
  NAND3_X1 U18400 ( .A1(n9722), .A2(n15068), .A3(n11284), .ZN(n15069) );
  AND2_X1 U18401 ( .A1(n15070), .A2(n15069), .ZN(n15072) );
  INV_X1 U18402 ( .A(n19055), .ZN(n16518) );
  OAI22_X1 U18403 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16518), .B1(n19942), 
        .B2(n19763), .ZN(n15071) );
  OAI21_X1 U18404 ( .B1(n15072), .B2(n12955), .A(n15071), .ZN(n15077) );
  OAI21_X1 U18405 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_0__SCAN_IN), .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n16516)
         );
  OAI21_X1 U18406 ( .B1(n19942), .B2(n15074), .A(n15073), .ZN(n15075) );
  AOI21_X1 U18407 ( .B1(n16516), .B2(n20033), .A(n15075), .ZN(n15076) );
  MUX2_X1 U18408 ( .A(n15077), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n15076), 
        .Z(P2_U3610) );
  NAND2_X1 U18409 ( .A1(n15093), .A2(n15078), .ZN(n15079) );
  NAND2_X1 U18410 ( .A1(n15080), .A2(n15079), .ZN(n15529) );
  OR2_X1 U18411 ( .A1(n15099), .A2(n15081), .ZN(n15082) );
  NAND2_X1 U18412 ( .A1(n9795), .A2(n15082), .ZN(n15532) );
  AOI22_X1 U18413 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19264), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19265), .ZN(n15085) );
  AOI22_X1 U18414 ( .A1(n15083), .A2(n19255), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19279), .ZN(n15084) );
  OAI211_X1 U18415 ( .C1(n15532), .C2(n19258), .A(n15085), .B(n15084), .ZN(
        n15089) );
  AOI211_X1 U18416 ( .C1(n15299), .C2(n15086), .A(n19928), .B(n15087), .ZN(
        n15088) );
  NOR2_X1 U18417 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  OAI21_X1 U18418 ( .B1(n15529), .B2(n19230), .A(n15090), .ZN(P2_U2826) );
  NAND2_X1 U18419 ( .A1(n13446), .A2(n15091), .ZN(n15092) );
  NAND2_X1 U18420 ( .A1(n15093), .A2(n15092), .ZN(n15544) );
  AOI211_X1 U18421 ( .C1(n15316), .C2(n15094), .A(n15095), .B(n19928), .ZN(
        n15096) );
  INV_X1 U18422 ( .A(n15096), .ZN(n15108) );
  AND2_X1 U18423 ( .A1(n15098), .A2(n15097), .ZN(n15100) );
  OR2_X1 U18424 ( .A1(n15100), .A2(n15099), .ZN(n15548) );
  NAND2_X1 U18425 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19279), .ZN(
        n15101) );
  OAI21_X1 U18426 ( .B1(n19252), .B2(n15102), .A(n15101), .ZN(n15103) );
  AOI21_X1 U18427 ( .B1(n19265), .B2(P2_REIP_REG_28__SCAN_IN), .A(n15103), 
        .ZN(n15104) );
  OAI21_X1 U18428 ( .B1(n15548), .B2(n19258), .A(n15104), .ZN(n15105) );
  AOI21_X1 U18429 ( .B1(n15106), .B2(n19255), .A(n15105), .ZN(n15107) );
  OAI211_X1 U18430 ( .C1(n19230), .C2(n15544), .A(n15108), .B(n15107), .ZN(
        P2_U2827) );
  AND2_X1 U18431 ( .A1(n15213), .A2(n15109), .ZN(n15111) );
  OR2_X1 U18432 ( .A1(n15111), .A2(n15110), .ZN(n15580) );
  AOI21_X1 U18433 ( .B1(n15113), .B2(n15275), .A(n15112), .ZN(n15577) );
  AOI22_X1 U18434 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19264), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19265), .ZN(n15114) );
  OAI21_X1 U18435 ( .B1(n15343), .B2(n19250), .A(n15114), .ZN(n15115) );
  AOI21_X1 U18436 ( .B1(n15577), .B2(n19266), .A(n15115), .ZN(n15116) );
  OAI21_X1 U18437 ( .B1(n15580), .B2(n19230), .A(n15116), .ZN(n15119) );
  AOI211_X1 U18438 ( .C1(n15117), .C2(n15346), .A(n9913), .B(n19928), .ZN(
        n15118) );
  AOI211_X1 U18439 ( .C1(n19255), .C2(n15120), .A(n15119), .B(n15118), .ZN(
        n15121) );
  INV_X1 U18440 ( .A(n15121), .ZN(P2_U2830) );
  OAI21_X1 U18441 ( .B1(n11230), .B2(n15123), .A(n15122), .ZN(n15605) );
  NAND2_X1 U18442 ( .A1(n15127), .A2(n15126), .ZN(n15128) );
  AND2_X1 U18443 ( .A1(n15125), .A2(n15128), .ZN(n15602) );
  AOI22_X1 U18444 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19264), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19265), .ZN(n15129) );
  OAI21_X1 U18445 ( .B1(n15371), .B2(n19250), .A(n15129), .ZN(n15130) );
  AOI21_X1 U18446 ( .B1(n15602), .B2(n19266), .A(n15130), .ZN(n15131) );
  OAI21_X1 U18447 ( .B1(n15605), .B2(n19230), .A(n15131), .ZN(n15135) );
  AOI211_X1 U18448 ( .C1(n15133), .C2(n15374), .A(n19928), .B(n15132), .ZN(
        n15134) );
  AOI211_X1 U18449 ( .C1(n19255), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        n15137) );
  INV_X1 U18450 ( .A(n15137), .ZN(P2_U2832) );
  AOI22_X1 U18451 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19264), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19265), .ZN(n15142) );
  OAI22_X1 U18452 ( .A1(n15139), .A2(n19270), .B1(n19250), .B2(n15138), .ZN(
        n15140) );
  INV_X1 U18453 ( .A(n15140), .ZN(n15141) );
  OAI211_X1 U18454 ( .C1(n15143), .C2(n19258), .A(n15142), .B(n15141), .ZN(
        n15147) );
  AOI211_X1 U18455 ( .C1(n15145), .C2(n9826), .A(n15144), .B(n19928), .ZN(
        n15146) );
  NOR2_X1 U18456 ( .A1(n15147), .A2(n15146), .ZN(n15148) );
  OAI21_X1 U18457 ( .B1(n19230), .B2(n15225), .A(n15148), .ZN(P2_U2833) );
  AND2_X1 U18458 ( .A1(n15164), .A2(n15149), .ZN(n15150) );
  NOR2_X1 U18459 ( .A1(n15151), .A2(n15150), .ZN(n15614) );
  NAND2_X1 U18460 ( .A1(n15614), .A2(n19273), .ZN(n15154) );
  OAI22_X1 U18461 ( .A1(n15396), .A2(n19250), .B1(n19979), .B2(n19222), .ZN(
        n15152) );
  AOI21_X1 U18462 ( .B1(n19264), .B2(P2_EBX_REG_21__SCAN_IN), .A(n15152), .ZN(
        n15153) );
  OAI211_X1 U18463 ( .C1(n19258), .C2(n15617), .A(n15154), .B(n15153), .ZN(
        n15158) );
  AOI211_X1 U18464 ( .C1(n15394), .C2(n15156), .A(n15155), .B(n19928), .ZN(
        n15157) );
  AOI211_X1 U18465 ( .C1(n19255), .C2(n15159), .A(n15158), .B(n15157), .ZN(
        n15160) );
  INV_X1 U18466 ( .A(n15160), .ZN(P2_U2834) );
  NAND2_X1 U18467 ( .A1(n15161), .A2(n15162), .ZN(n15163) );
  AND2_X1 U18468 ( .A1(n15164), .A2(n15163), .ZN(n15628) );
  INV_X1 U18469 ( .A(n15628), .ZN(n15238) );
  NOR2_X1 U18470 ( .A1(n19226), .A2(n19928), .ZN(n19278) );
  OAI21_X1 U18471 ( .B1(n14330), .B2(n10102), .A(n15166), .ZN(n16411) );
  OAI22_X1 U18472 ( .A1(n16411), .A2(n19258), .B1(n19250), .B2(n9904), .ZN(
        n15169) );
  INV_X1 U18473 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19978) );
  OAI22_X1 U18474 ( .A1(n15167), .A2(n19252), .B1(n19978), .B2(n19222), .ZN(
        n15168) );
  AOI211_X1 U18475 ( .C1(n15172), .C2(n19278), .A(n15169), .B(n15168), .ZN(
        n15175) );
  AOI21_X1 U18476 ( .B1(n15172), .B2(n15171), .A(n15170), .ZN(n15173) );
  NAND2_X1 U18477 ( .A1(n15173), .A2(n19275), .ZN(n15174) );
  OAI211_X1 U18478 ( .C1(n15238), .C2(n19230), .A(n15175), .B(n15174), .ZN(
        n15176) );
  AOI21_X1 U18479 ( .B1(n19255), .B2(n15177), .A(n15176), .ZN(n15178) );
  INV_X1 U18480 ( .A(n15178), .ZN(P2_U2835) );
  OR2_X1 U18481 ( .A1(n15180), .A2(n15179), .ZN(n15244) );
  NAND3_X1 U18482 ( .A1(n15244), .A2(n15181), .A3(n15235), .ZN(n15183) );
  NAND2_X1 U18483 ( .A1(n13900), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15182) );
  OAI211_X1 U18484 ( .C1(n13900), .C2(n15529), .A(n15183), .B(n15182), .ZN(
        P2_U2858) );
  INV_X1 U18485 ( .A(n15184), .ZN(n15185) );
  NAND2_X1 U18486 ( .A1(n15186), .A2(n15185), .ZN(n15188) );
  XNOR2_X1 U18487 ( .A(n15188), .B(n15187), .ZN(n15255) );
  NOR2_X1 U18488 ( .A1(n15544), .A2(n13900), .ZN(n15189) );
  AOI21_X1 U18489 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n13900), .A(n15189), .ZN(
        n15190) );
  OAI21_X1 U18490 ( .B1(n15255), .B2(n15242), .A(n15190), .ZN(P2_U2859) );
  OAI21_X1 U18491 ( .B1(n15193), .B2(n15192), .A(n15191), .ZN(n15260) );
  NOR2_X1 U18492 ( .A1(n15558), .A2(n13900), .ZN(n15194) );
  AOI21_X1 U18493 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n13900), .A(n15194), .ZN(
        n15195) );
  OAI21_X1 U18494 ( .B1(n15260), .B2(n15242), .A(n15195), .ZN(P2_U2860) );
  OAI21_X1 U18495 ( .B1(n15198), .B2(n15197), .A(n15196), .ZN(n15267) );
  NOR2_X1 U18496 ( .A1(n15110), .A2(n15199), .ZN(n15200) );
  OR2_X1 U18497 ( .A1(n15201), .A2(n15200), .ZN(n16388) );
  NOR2_X1 U18498 ( .A1(n16388), .A2(n13900), .ZN(n15202) );
  AOI21_X1 U18499 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n13900), .A(n15202), .ZN(
        n15203) );
  OAI21_X1 U18500 ( .B1(n15267), .B2(n15242), .A(n15203), .ZN(P2_U2861) );
  OAI21_X1 U18501 ( .B1(n15206), .B2(n15205), .A(n15204), .ZN(n15272) );
  MUX2_X1 U18502 ( .A(n15580), .B(n15207), .S(n13900), .Z(n15208) );
  OAI21_X1 U18503 ( .B1(n15272), .B2(n15242), .A(n15208), .ZN(P2_U2862) );
  AOI21_X1 U18504 ( .B1(n15210), .B2(n15209), .A(n9810), .ZN(n15211) );
  XOR2_X1 U18505 ( .A(n15212), .B(n15211), .Z(n15282) );
  INV_X1 U18506 ( .A(n15213), .ZN(n15214) );
  AOI21_X1 U18507 ( .B1(n15215), .B2(n15122), .A(n15214), .ZN(n16400) );
  NOR2_X1 U18508 ( .A1(n15229), .A2(n15216), .ZN(n15217) );
  AOI21_X1 U18509 ( .B1(n16400), .B2(n15229), .A(n15217), .ZN(n15218) );
  OAI21_X1 U18510 ( .B1(n15282), .B2(n15242), .A(n15218), .ZN(P2_U2863) );
  AOI21_X1 U18511 ( .B1(n15221), .B2(n15220), .A(n15219), .ZN(n15222) );
  INV_X1 U18512 ( .A(n15222), .ZN(n15291) );
  INV_X1 U18513 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n15223) );
  MUX2_X1 U18514 ( .A(n15223), .B(n15605), .S(n15229), .Z(n15224) );
  OAI21_X1 U18515 ( .B1(n15291), .B2(n15242), .A(n15224), .ZN(P2_U2864) );
  NOR2_X1 U18516 ( .A1(n15225), .A2(n13900), .ZN(n15226) );
  AOI21_X1 U18517 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n13900), .A(n15226), .ZN(
        n15227) );
  OAI21_X1 U18518 ( .B1(n15228), .B2(n15242), .A(n15227), .ZN(P2_U2865) );
  NAND2_X1 U18519 ( .A1(n13900), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15231) );
  NAND2_X1 U18520 ( .A1(n15614), .A2(n15229), .ZN(n15230) );
  OAI211_X1 U18521 ( .C1(n15232), .C2(n15242), .A(n15231), .B(n15230), .ZN(
        P2_U2866) );
  AOI21_X1 U18522 ( .B1(n15234), .B2(n15233), .A(n14482), .ZN(n16413) );
  NAND2_X1 U18523 ( .A1(n16413), .A2(n15235), .ZN(n15237) );
  NAND2_X1 U18524 ( .A1(n13900), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15236) );
  OAI211_X1 U18525 ( .C1(n15238), .C2(n13900), .A(n15237), .B(n15236), .ZN(
        P2_U2867) );
  OAI21_X1 U18526 ( .B1(n14384), .B2(n15239), .A(n15161), .ZN(n19088) );
  NOR2_X1 U18527 ( .A1(n19088), .A2(n13900), .ZN(n15240) );
  AOI21_X1 U18528 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n13900), .A(n15240), .ZN(
        n15241) );
  OAI21_X1 U18529 ( .B1(n15243), .B2(n15242), .A(n15241), .ZN(P2_U2868) );
  NAND3_X1 U18530 ( .A1(n15244), .A2(n15181), .A3(n19343), .ZN(n15250) );
  INV_X1 U18531 ( .A(n15532), .ZN(n15247) );
  OAI22_X1 U18532 ( .A1(n15284), .A2(n19302), .B1(n19322), .B2(n15245), .ZN(
        n15246) );
  AOI21_X1 U18533 ( .B1(n15247), .B2(n19339), .A(n15246), .ZN(n15249) );
  AOI22_X1 U18534 ( .A1(n19291), .A2(BUF1_REG_29__SCAN_IN), .B1(n19290), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15248) );
  NAND3_X1 U18535 ( .A1(n15250), .A2(n15249), .A3(n15248), .ZN(P2_U2890) );
  AOI22_X1 U18536 ( .A1(n19289), .A2(n19304), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n19338), .ZN(n15252) );
  AOI22_X1 U18537 ( .A1(n19291), .A2(BUF1_REG_28__SCAN_IN), .B1(n19290), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15251) );
  OAI211_X1 U18538 ( .C1(n15548), .C2(n19297), .A(n15252), .B(n15251), .ZN(
        n15253) );
  INV_X1 U18539 ( .A(n15253), .ZN(n15254) );
  OAI21_X1 U18540 ( .B1(n15255), .B2(n19324), .A(n15254), .ZN(P2_U2891) );
  OAI22_X1 U18541 ( .A1(n15284), .A2(n19307), .B1(n19322), .B2(n15256), .ZN(
        n15257) );
  AOI21_X1 U18542 ( .B1(n15555), .B2(n19339), .A(n15257), .ZN(n15259) );
  AOI22_X1 U18543 ( .A1(n19291), .A2(BUF1_REG_27__SCAN_IN), .B1(n19290), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15258) );
  OAI211_X1 U18544 ( .C1(n15260), .C2(n19324), .A(n15259), .B(n15258), .ZN(
        P2_U2892) );
  OR2_X1 U18545 ( .A1(n15112), .A2(n15261), .ZN(n15262) );
  AND2_X1 U18546 ( .A1(n15262), .A2(n13448), .ZN(n16398) );
  INV_X1 U18547 ( .A(n19309), .ZN(n15263) );
  OAI22_X1 U18548 ( .A1(n15284), .A2(n15263), .B1(n19322), .B2(n13573), .ZN(
        n15264) );
  AOI21_X1 U18549 ( .B1(n16398), .B2(n19339), .A(n15264), .ZN(n15266) );
  AOI22_X1 U18550 ( .A1(n19291), .A2(BUF1_REG_26__SCAN_IN), .B1(n19290), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15265) );
  OAI211_X1 U18551 ( .C1(n15267), .C2(n19324), .A(n15266), .B(n15265), .ZN(
        P2_U2893) );
  OAI22_X1 U18552 ( .A1(n15284), .A2(n19312), .B1(n19322), .B2(n15268), .ZN(
        n15269) );
  AOI21_X1 U18553 ( .B1(n15577), .B2(n19339), .A(n15269), .ZN(n15271) );
  AOI22_X1 U18554 ( .A1(n19291), .A2(BUF1_REG_25__SCAN_IN), .B1(n19290), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15270) );
  OAI211_X1 U18555 ( .C1(n15272), .C2(n19324), .A(n15271), .B(n15270), .ZN(
        P2_U2894) );
  NAND2_X1 U18556 ( .A1(n15125), .A2(n15273), .ZN(n15274) );
  MUX2_X1 U18557 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n15276), .Z(n19386) );
  INV_X1 U18558 ( .A(n19386), .ZN(n15278) );
  INV_X1 U18559 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15277) );
  OAI22_X1 U18560 ( .A1(n15284), .A2(n15278), .B1(n19322), .B2(n15277), .ZN(
        n15279) );
  AOI21_X1 U18561 ( .B1(n19339), .B2(n10118), .A(n15279), .ZN(n15281) );
  AOI22_X1 U18562 ( .A1(n19291), .A2(BUF1_REG_24__SCAN_IN), .B1(n19290), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15280) );
  OAI211_X1 U18563 ( .C1(n15282), .C2(n19324), .A(n15281), .B(n15280), .ZN(
        P2_U2895) );
  OAI22_X1 U18564 ( .A1(n15284), .A2(n19318), .B1(n19322), .B2(n15283), .ZN(
        n15289) );
  INV_X1 U18565 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n15286) );
  INV_X1 U18566 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15285) );
  OAI22_X1 U18567 ( .A1(n15287), .A2(n15286), .B1(n19284), .B2(n15285), .ZN(
        n15288) );
  AOI211_X1 U18568 ( .C1(n19339), .C2(n15602), .A(n15289), .B(n15288), .ZN(
        n15290) );
  OAI21_X1 U18569 ( .B1(n15291), .B2(n19324), .A(n15290), .ZN(P2_U2896) );
  NAND2_X1 U18570 ( .A1(n15293), .A2(n15292), .ZN(n15295) );
  XOR2_X1 U18571 ( .A(n15295), .B(n15294), .Z(n15539) );
  NAND2_X1 U18572 ( .A1(n19399), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15530) );
  OAI21_X1 U18573 ( .B1(n16428), .B2(n15296), .A(n15530), .ZN(n15298) );
  NOR2_X1 U18574 ( .A1(n15529), .A2(n15509), .ZN(n15297) );
  AOI211_X1 U18575 ( .C1(n19398), .C2(n15299), .A(n15298), .B(n15297), .ZN(
        n15303) );
  OAI211_X1 U18576 ( .C1(n15539), .C2(n16435), .A(n15303), .B(n15302), .ZN(
        P2_U2985) );
  OAI21_X1 U18577 ( .B1(n15304), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15305), .ZN(n15554) );
  OAI21_X1 U18578 ( .B1(n15307), .B2(n15340), .A(n15306), .ZN(n15309) );
  XNOR2_X1 U18579 ( .A(n15309), .B(n15308), .ZN(n15319) );
  INV_X1 U18580 ( .A(n15308), .ZN(n15310) );
  AOI22_X1 U18581 ( .A1(n15319), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n15310), .B2(n15309), .ZN(n15313) );
  XNOR2_X1 U18582 ( .A(n15311), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15312) );
  XNOR2_X1 U18583 ( .A(n15313), .B(n15312), .ZN(n15540) );
  NAND2_X1 U18584 ( .A1(n15540), .A2(n19400), .ZN(n15318) );
  NAND2_X1 U18585 ( .A1(n19399), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15546) );
  OAI21_X1 U18586 ( .B1(n16428), .B2(n9908), .A(n15546), .ZN(n15315) );
  NOR2_X1 U18587 ( .A1(n15544), .A2(n15509), .ZN(n15314) );
  AOI211_X1 U18588 ( .C1(n19398), .C2(n15316), .A(n15315), .B(n15314), .ZN(
        n15317) );
  OAI211_X1 U18589 ( .C1(n16436), .C2(n15554), .A(n15318), .B(n15317), .ZN(
        P2_U2986) );
  XNOR2_X1 U18590 ( .A(n15319), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15565) );
  NOR2_X1 U18591 ( .A1(n15320), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15321) );
  NOR2_X1 U18592 ( .A1(n15304), .A2(n15321), .ZN(n15562) );
  NAND2_X1 U18593 ( .A1(n19399), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15557) );
  OAI21_X1 U18594 ( .B1(n16428), .B2(n15322), .A(n15557), .ZN(n15323) );
  AOI21_X1 U18595 ( .B1(n19398), .B2(n15324), .A(n15323), .ZN(n15325) );
  OAI21_X1 U18596 ( .B1(n15558), .B2(n15509), .A(n15325), .ZN(n15326) );
  AOI21_X1 U18597 ( .B1(n15562), .B2(n19404), .A(n15326), .ZN(n15327) );
  OAI21_X1 U18598 ( .B1(n15565), .B2(n16435), .A(n15327), .ZN(P2_U2987) );
  INV_X1 U18599 ( .A(n15320), .ZN(n15329) );
  OAI21_X1 U18600 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15328), .A(
        n15329), .ZN(n15574) );
  INV_X1 U18601 ( .A(n15340), .ZN(n15330) );
  AOI21_X1 U18602 ( .B1(n15342), .B2(n15330), .A(n15339), .ZN(n15331) );
  XNOR2_X1 U18603 ( .A(n15332), .B(n15331), .ZN(n15572) );
  NOR2_X1 U18604 ( .A1(n19214), .A2(n15333), .ZN(n15568) );
  NOR2_X1 U18605 ( .A1(n16455), .A2(n15334), .ZN(n15335) );
  AOI211_X1 U18606 ( .C1(n16442), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15568), .B(n15335), .ZN(n15336) );
  OAI21_X1 U18607 ( .B1(n16388), .B2(n15509), .A(n15336), .ZN(n15337) );
  AOI21_X1 U18608 ( .B1(n15572), .B2(n19400), .A(n15337), .ZN(n15338) );
  OAI21_X1 U18609 ( .B1(n16436), .B2(n15574), .A(n15338), .ZN(P2_U2988) );
  NOR2_X1 U18610 ( .A1(n15340), .A2(n15339), .ZN(n15341) );
  XNOR2_X1 U18611 ( .A(n15342), .B(n15341), .ZN(n15588) );
  INV_X1 U18612 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19986) );
  OR2_X1 U18613 ( .A1(n19214), .A2(n19986), .ZN(n15579) );
  OAI21_X1 U18614 ( .B1(n19409), .B2(n15343), .A(n15579), .ZN(n15345) );
  NOR2_X1 U18615 ( .A1(n15580), .A2(n15509), .ZN(n15344) );
  AOI211_X1 U18616 ( .C1(n19398), .C2(n15346), .A(n15345), .B(n15344), .ZN(
        n15349) );
  INV_X1 U18617 ( .A(n15328), .ZN(n15585) );
  NAND2_X1 U18618 ( .A1(n15347), .A2(n21297), .ZN(n15584) );
  NAND3_X1 U18619 ( .A1(n15585), .A2(n19404), .A3(n15584), .ZN(n15348) );
  OAI211_X1 U18620 ( .C1(n15588), .C2(n16435), .A(n15349), .B(n15348), .ZN(
        P2_U2989) );
  INV_X1 U18621 ( .A(n15350), .ZN(n15351) );
  OAI21_X1 U18622 ( .B1(n15351), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15347), .ZN(n15599) );
  NOR2_X1 U18623 ( .A1(n15353), .A2(n15352), .ZN(n15362) );
  NOR2_X1 U18624 ( .A1(n15355), .A2(n15354), .ZN(n15370) );
  INV_X1 U18625 ( .A(n15370), .ZN(n15358) );
  XNOR2_X1 U18626 ( .A(n15356), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15369) );
  INV_X1 U18627 ( .A(n15369), .ZN(n15357) );
  NAND2_X1 U18628 ( .A1(n15358), .A2(n15357), .ZN(n15600) );
  OAI21_X1 U18629 ( .B1(n15360), .B2(n15359), .A(n15600), .ZN(n15361) );
  XOR2_X1 U18630 ( .A(n15362), .B(n15361), .Z(n15597) );
  NAND2_X1 U18631 ( .A1(n16400), .A2(n19403), .ZN(n15364) );
  NOR2_X1 U18632 ( .A1(n19214), .A2(n19984), .ZN(n15592) );
  AOI21_X1 U18633 ( .B1(n16442), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15592), .ZN(n15363) );
  OAI211_X1 U18634 ( .C1(n16455), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        n15366) );
  AOI21_X1 U18635 ( .B1(n15597), .B2(n19400), .A(n15366), .ZN(n15367) );
  OAI21_X1 U18636 ( .B1(n16436), .B2(n15599), .A(n15367), .ZN(P2_U2990) );
  OAI21_X1 U18637 ( .B1(n15368), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15350), .ZN(n15612) );
  NAND2_X1 U18638 ( .A1(n15370), .A2(n15369), .ZN(n15601) );
  NAND3_X1 U18639 ( .A1(n15601), .A2(n15600), .A3(n19400), .ZN(n15376) );
  OR2_X1 U18640 ( .A1(n19214), .A2(n19982), .ZN(n15604) );
  OAI21_X1 U18641 ( .B1(n16428), .B2(n15371), .A(n15604), .ZN(n15373) );
  NOR2_X1 U18642 ( .A1(n15605), .A2(n15509), .ZN(n15372) );
  AOI211_X1 U18643 ( .C1(n19398), .C2(n15374), .A(n15373), .B(n15372), .ZN(
        n15375) );
  OAI211_X1 U18644 ( .C1(n15612), .C2(n16436), .A(n15376), .B(n15375), .ZN(
        P2_U2991) );
  OAI21_X1 U18645 ( .B1(n15378), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15377), .ZN(n15624) );
  NAND2_X1 U18646 ( .A1(n15383), .A2(n15382), .ZN(n15434) );
  INV_X1 U18647 ( .A(n15383), .ZN(n15384) );
  NOR2_X1 U18648 ( .A1(n15388), .A2(n15389), .ZN(n15401) );
  NAND2_X1 U18649 ( .A1(n15402), .A2(n15401), .ZN(n15400) );
  INV_X1 U18650 ( .A(n15389), .ZN(n15390) );
  NAND2_X1 U18651 ( .A1(n15400), .A2(n15390), .ZN(n15393) );
  XNOR2_X1 U18652 ( .A(n15393), .B(n10100), .ZN(n15613) );
  NAND2_X1 U18653 ( .A1(n15613), .A2(n19400), .ZN(n15399) );
  NAND2_X1 U18654 ( .A1(n19398), .A2(n15394), .ZN(n15395) );
  NAND2_X1 U18655 ( .A1(n19399), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15615) );
  OAI211_X1 U18656 ( .C1(n19409), .C2(n15396), .A(n15395), .B(n15615), .ZN(
        n15397) );
  AOI21_X1 U18657 ( .B1(n15614), .B2(n19403), .A(n15397), .ZN(n15398) );
  OAI211_X1 U18658 ( .C1(n16436), .C2(n15624), .A(n15399), .B(n15398), .ZN(
        P2_U2993) );
  OAI21_X1 U18659 ( .B1(n15402), .B2(n15401), .A(n15400), .ZN(n15625) );
  NAND2_X1 U18660 ( .A1(n19399), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15629) );
  NAND2_X1 U18661 ( .A1(n16442), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15403) );
  OAI211_X1 U18662 ( .C1(n15404), .C2(n16455), .A(n15629), .B(n15403), .ZN(
        n15407) );
  NAND2_X1 U18663 ( .A1(n15409), .A2(n15408), .ZN(n15412) );
  NOR2_X1 U18664 ( .A1(n15410), .A2(n15420), .ZN(n15411) );
  XOR2_X1 U18665 ( .A(n15412), .B(n15411), .Z(n15646) );
  NAND2_X1 U18666 ( .A1(n19399), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15638) );
  OAI21_X1 U18667 ( .B1(n16428), .B2(n15413), .A(n15638), .ZN(n15415) );
  NOR2_X1 U18668 ( .A1(n19088), .A2(n15509), .ZN(n15414) );
  AOI211_X1 U18669 ( .C1(n19398), .C2(n15416), .A(n15415), .B(n15414), .ZN(
        n15419) );
  INV_X1 U18670 ( .A(n15417), .ZN(n15643) );
  NAND2_X1 U18671 ( .A1(n15424), .A2(n21279), .ZN(n15642) );
  NAND3_X1 U18672 ( .A1(n15643), .A2(n19404), .A3(n15642), .ZN(n15418) );
  OAI211_X1 U18673 ( .C1(n15646), .C2(n16435), .A(n15419), .B(n15418), .ZN(
        P2_U2995) );
  NOR2_X1 U18674 ( .A1(n15421), .A2(n15420), .ZN(n15422) );
  XNOR2_X1 U18675 ( .A(n15423), .B(n15422), .ZN(n15660) );
  OR2_X2 U18676 ( .A1(n15689), .A2(n15704), .ZN(n15690) );
  AOI21_X1 U18677 ( .B1(n15661), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15426) );
  INV_X1 U18678 ( .A(n15424), .ZN(n15425) );
  NOR2_X1 U18679 ( .A1(n15426), .A2(n15425), .ZN(n15658) );
  NOR2_X1 U18680 ( .A1(n19214), .A2(n19974), .ZN(n15653) );
  NOR2_X1 U18681 ( .A1(n15427), .A2(n16455), .ZN(n15428) );
  AOI211_X1 U18682 ( .C1(n16442), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15653), .B(n15428), .ZN(n15429) );
  OAI21_X1 U18683 ( .B1(n19102), .B2(n15509), .A(n15429), .ZN(n15430) );
  AOI21_X1 U18684 ( .B1(n15658), .B2(n19404), .A(n15430), .ZN(n15431) );
  OAI21_X1 U18685 ( .B1(n15660), .B2(n16435), .A(n15431), .ZN(P2_U2996) );
  XNOR2_X1 U18686 ( .A(n15661), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15443) );
  AOI21_X1 U18687 ( .B1(n15434), .B2(n15433), .A(n15432), .ZN(n15435) );
  INV_X1 U18688 ( .A(n15435), .ZN(n15672) );
  NOR2_X1 U18689 ( .A1(n19214), .A2(n15436), .ZN(n15668) );
  NOR2_X1 U18690 ( .A1(n19409), .A2(n21218), .ZN(n15437) );
  AOI211_X1 U18691 ( .C1(n15438), .C2(n19398), .A(n15668), .B(n15437), .ZN(
        n15439) );
  OAI21_X1 U18692 ( .B1(n15440), .B2(n15509), .A(n15439), .ZN(n15441) );
  AOI21_X1 U18693 ( .B1(n15672), .B2(n19400), .A(n15441), .ZN(n15442) );
  OAI21_X1 U18694 ( .B1(n16436), .B2(n15443), .A(n15442), .ZN(P2_U2997) );
  XNOR2_X1 U18695 ( .A(n15690), .B(n15687), .ZN(n15451) );
  XOR2_X1 U18696 ( .A(n15445), .B(n15444), .Z(n15681) );
  NOR2_X1 U18697 ( .A1(n10855), .A2(n19214), .ZN(n15446) );
  AOI21_X1 U18698 ( .B1(n19125), .B2(n19403), .A(n15446), .ZN(n15448) );
  AOI22_X1 U18699 ( .A1(n16442), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n19398), .B2(n19120), .ZN(n15447) );
  NAND2_X1 U18700 ( .A1(n15448), .A2(n15447), .ZN(n15449) );
  AOI21_X1 U18701 ( .B1(n15681), .B2(n19400), .A(n15449), .ZN(n15450) );
  OAI21_X1 U18702 ( .B1(n16436), .B2(n15451), .A(n15450), .ZN(P2_U2998) );
  NAND2_X1 U18703 ( .A1(n15761), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15483) );
  NOR2_X1 U18704 ( .A1(n15483), .A2(n15715), .ZN(n15466) );
  OAI21_X1 U18705 ( .B1(n15466), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15689), .ZN(n15721) );
  INV_X1 U18706 ( .A(n15452), .ZN(n15454) );
  NOR2_X1 U18707 ( .A1(n15454), .A2(n15453), .ZN(n15455) );
  XNOR2_X1 U18708 ( .A(n15456), .B(n15455), .ZN(n15718) );
  NAND2_X1 U18709 ( .A1(n19147), .A2(n19403), .ZN(n15458) );
  AOI22_X1 U18710 ( .A1(n16442), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19399), .ZN(n15457) );
  OAI211_X1 U18711 ( .C1(n16455), .C2(n15459), .A(n15458), .B(n15457), .ZN(
        n15460) );
  AOI21_X1 U18712 ( .B1(n15718), .B2(n19400), .A(n15460), .ZN(n15461) );
  OAI21_X1 U18713 ( .B1(n15721), .B2(n16436), .A(n15461), .ZN(P2_U3000) );
  NAND2_X1 U18714 ( .A1(n15463), .A2(n15462), .ZN(n15465) );
  XOR2_X1 U18715 ( .A(n15465), .B(n15464), .Z(n15734) );
  INV_X1 U18716 ( .A(n15483), .ZN(n15473) );
  AOI21_X1 U18717 ( .B1(n15473), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15467) );
  NOR2_X1 U18718 ( .A1(n15467), .A2(n15466), .ZN(n15722) );
  NAND2_X1 U18719 ( .A1(n15722), .A2(n19404), .ZN(n15472) );
  INV_X1 U18720 ( .A(n15468), .ZN(n19155) );
  NAND2_X1 U18721 ( .A1(n19399), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15727) );
  OAI21_X1 U18722 ( .B1(n19409), .B2(n19161), .A(n15727), .ZN(n15470) );
  NOR2_X1 U18723 ( .A1(n19156), .A2(n15509), .ZN(n15469) );
  AOI211_X1 U18724 ( .C1(n19398), .C2(n19155), .A(n15470), .B(n15469), .ZN(
        n15471) );
  OAI211_X1 U18725 ( .C1(n16435), .C2(n15734), .A(n15472), .B(n15471), .ZN(
        P2_U3001) );
  XNOR2_X1 U18726 ( .A(n15473), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15748) );
  OAI21_X1 U18727 ( .B1(n15475), .B2(n15477), .A(n15474), .ZN(n15476) );
  OAI21_X1 U18728 ( .B1(n15478), .B2(n15477), .A(n15476), .ZN(n15746) );
  NAND2_X1 U18729 ( .A1(n15740), .A2(n19403), .ZN(n15480) );
  NOR2_X1 U18730 ( .A1(n19214), .A2(n19967), .ZN(n15739) );
  AOI21_X1 U18731 ( .B1(n16442), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15739), .ZN(n15479) );
  OAI211_X1 U18732 ( .C1(n16455), .C2(n19163), .A(n15480), .B(n15479), .ZN(
        n15481) );
  AOI21_X1 U18733 ( .B1(n15746), .B2(n19400), .A(n15481), .ZN(n15482) );
  OAI21_X1 U18734 ( .B1(n15748), .B2(n16436), .A(n15482), .ZN(P2_U3002) );
  OAI21_X1 U18735 ( .B1(n15761), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15483), .ZN(n15760) );
  NAND2_X1 U18736 ( .A1(n16447), .A2(n16445), .ZN(n15485) );
  INV_X1 U18737 ( .A(n15790), .ZN(n15487) );
  INV_X1 U18738 ( .A(n15788), .ZN(n15486) );
  NAND2_X1 U18739 ( .A1(n15487), .A2(n15486), .ZN(n15772) );
  INV_X1 U18740 ( .A(n15772), .ZN(n15489) );
  AOI21_X1 U18741 ( .B1(n15489), .B2(n15774), .A(n15488), .ZN(n15494) );
  INV_X1 U18742 ( .A(n15490), .ZN(n15492) );
  NOR2_X1 U18743 ( .A1(n15492), .A2(n15491), .ZN(n15493) );
  XNOR2_X1 U18744 ( .A(n15494), .B(n15493), .ZN(n15758) );
  NOR2_X1 U18745 ( .A1(n19214), .A2(n19965), .ZN(n15753) );
  NOR2_X1 U18746 ( .A1(n16428), .A2(n19184), .ZN(n15495) );
  AOI211_X1 U18747 ( .C1(n19178), .C2(n19398), .A(n15753), .B(n15495), .ZN(
        n15496) );
  OAI21_X1 U18748 ( .B1(n15509), .B2(n19179), .A(n15496), .ZN(n15497) );
  AOI21_X1 U18749 ( .B1(n15758), .B2(n19400), .A(n15497), .ZN(n15498) );
  OAI21_X1 U18750 ( .B1(n15760), .B2(n16436), .A(n15498), .ZN(P2_U3003) );
  XNOR2_X1 U18751 ( .A(n9729), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15814) );
  AND2_X1 U18752 ( .A1(n15503), .A2(n15502), .ZN(n15501) );
  NAND2_X1 U18753 ( .A1(n15500), .A2(n15501), .ZN(n16446) );
  INV_X1 U18754 ( .A(n16445), .ZN(n15506) );
  AND2_X1 U18755 ( .A1(n15500), .A2(n15502), .ZN(n15505) );
  AND2_X1 U18756 ( .A1(n16445), .A2(n15503), .ZN(n15504) );
  OAI22_X1 U18757 ( .A1(n16446), .A2(n15506), .B1(n15505), .B2(n15504), .ZN(
        n15812) );
  INV_X1 U18758 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15507) );
  OAI22_X1 U18759 ( .A1(n19409), .A2(n15507), .B1(n16455), .B2(n19212), .ZN(
        n15511) );
  INV_X1 U18760 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n15508) );
  OAI22_X1 U18761 ( .A1(n19217), .A2(n15509), .B1(n19214), .B2(n15508), .ZN(
        n15510) );
  AOI211_X1 U18762 ( .C1(n15812), .C2(n19400), .A(n15511), .B(n15510), .ZN(
        n15512) );
  OAI21_X1 U18763 ( .B1(n15814), .B2(n16436), .A(n15512), .ZN(P2_U3007) );
  INV_X1 U18764 ( .A(n15513), .ZN(n15514) );
  NAND2_X1 U18765 ( .A1(n15514), .A2(n16471), .ZN(n15527) );
  INV_X1 U18766 ( .A(n15515), .ZN(n15524) );
  NAND2_X1 U18767 ( .A1(n15516), .A2(n16457), .ZN(n15517) );
  OAI211_X1 U18768 ( .C1(n15520), .C2(n15519), .A(n15518), .B(n15517), .ZN(
        n15521) );
  INV_X1 U18769 ( .A(n15521), .ZN(n15523) );
  INV_X1 U18770 ( .A(n15525), .ZN(n15526) );
  OAI211_X1 U18771 ( .C1(n15528), .C2(n16476), .A(n15527), .B(n15526), .ZN(
        P2_U3016) );
  NOR2_X1 U18772 ( .A1(n15543), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15559) );
  NOR2_X1 U18773 ( .A1(n15559), .A2(n15561), .ZN(n15541) );
  OAI21_X1 U18774 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15543), .A(
        n15541), .ZN(n15535) );
  NOR2_X1 U18775 ( .A1(n15529), .A2(n15834), .ZN(n15534) );
  OR4_X1 U18776 ( .A1(n10781), .A2(n15542), .A3(n15543), .A4(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15531) );
  OAI211_X1 U18777 ( .C1(n15532), .C2(n16474), .A(n15531), .B(n15530), .ZN(
        n15533) );
  NAND2_X1 U18778 ( .A1(n15536), .A2(n16461), .ZN(n15537) );
  OAI211_X1 U18779 ( .C1(n15539), .C2(n15800), .A(n15538), .B(n15537), .ZN(
        P2_U3017) );
  NAND2_X1 U18780 ( .A1(n15540), .A2(n16471), .ZN(n15553) );
  INV_X1 U18781 ( .A(n15541), .ZN(n15551) );
  NOR3_X1 U18782 ( .A1(n15543), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15542), .ZN(n15550) );
  INV_X1 U18783 ( .A(n15544), .ZN(n15545) );
  NAND2_X1 U18784 ( .A1(n15545), .A2(n16479), .ZN(n15547) );
  OAI211_X1 U18785 ( .C1(n16474), .C2(n15548), .A(n15547), .B(n15546), .ZN(
        n15549) );
  OAI211_X1 U18786 ( .C1(n15554), .C2(n16476), .A(n15553), .B(n15552), .ZN(
        P2_U3018) );
  NAND2_X1 U18787 ( .A1(n15555), .A2(n16457), .ZN(n15556) );
  OAI211_X1 U18788 ( .C1(n15558), .C2(n15834), .A(n15557), .B(n15556), .ZN(
        n15560) );
  AOI211_X1 U18789 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15561), .A(
        n15560), .B(n15559), .ZN(n15564) );
  NAND2_X1 U18790 ( .A1(n15562), .A2(n16461), .ZN(n15563) );
  OAI211_X1 U18791 ( .C1(n15565), .C2(n15800), .A(n15564), .B(n15563), .ZN(
        P2_U3019) );
  XNOR2_X1 U18792 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15566) );
  NOR2_X1 U18793 ( .A1(n15575), .A2(n15566), .ZN(n15571) );
  NOR2_X1 U18794 ( .A1(n16388), .A2(n15834), .ZN(n15567) );
  OAI21_X1 U18795 ( .B1(n21158), .B2(n15576), .A(n15569), .ZN(n15570) );
  AOI211_X1 U18796 ( .C1(n15572), .C2(n16471), .A(n15571), .B(n15570), .ZN(
        n15573) );
  OAI21_X1 U18797 ( .B1(n16476), .B2(n15574), .A(n15573), .ZN(P2_U3020) );
  INV_X1 U18798 ( .A(n15575), .ZN(n15583) );
  NOR2_X1 U18799 ( .A1(n15576), .A2(n21297), .ZN(n15582) );
  NAND2_X1 U18800 ( .A1(n15577), .A2(n16457), .ZN(n15578) );
  OAI211_X1 U18801 ( .C1(n15580), .C2(n15834), .A(n15579), .B(n15578), .ZN(
        n15581) );
  AOI211_X1 U18802 ( .C1(n15583), .C2(n21297), .A(n15582), .B(n15581), .ZN(
        n15587) );
  NAND3_X1 U18803 ( .A1(n15585), .A2(n16461), .A3(n15584), .ZN(n15586) );
  OAI211_X1 U18804 ( .C1(n15588), .C2(n15800), .A(n15587), .B(n15586), .ZN(
        P2_U3021) );
  INV_X1 U18805 ( .A(n16400), .ZN(n15595) );
  NOR2_X1 U18806 ( .A1(n15607), .A2(n15589), .ZN(n15591) );
  OAI21_X1 U18807 ( .B1(n15591), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15590), .ZN(n15594) );
  AOI21_X1 U18808 ( .B1(n16457), .B2(n10118), .A(n15592), .ZN(n15593) );
  OAI211_X1 U18809 ( .C1(n15595), .C2(n15834), .A(n15594), .B(n15593), .ZN(
        n15596) );
  AOI21_X1 U18810 ( .B1(n15597), .B2(n16471), .A(n15596), .ZN(n15598) );
  OAI21_X1 U18811 ( .B1(n16476), .B2(n15599), .A(n15598), .ZN(P2_U3022) );
  NAND3_X1 U18812 ( .A1(n15601), .A2(n15600), .A3(n16471), .ZN(n15611) );
  NAND2_X1 U18813 ( .A1(n16457), .A2(n15602), .ZN(n15603) );
  OAI211_X1 U18814 ( .C1(n15605), .C2(n15834), .A(n15604), .B(n15603), .ZN(
        n15609) );
  XNOR2_X1 U18815 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15606) );
  NOR2_X1 U18816 ( .A1(n15607), .A2(n15606), .ZN(n15608) );
  AOI211_X1 U18817 ( .C1(n15621), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15609), .B(n15608), .ZN(n15610) );
  OAI211_X1 U18818 ( .C1(n15612), .C2(n16476), .A(n15611), .B(n15610), .ZN(
        P2_U3023) );
  NAND2_X1 U18819 ( .A1(n15613), .A2(n16471), .ZN(n15623) );
  NAND2_X1 U18820 ( .A1(n15614), .A2(n16479), .ZN(n15616) );
  OAI211_X1 U18821 ( .C1(n16474), .C2(n15617), .A(n15616), .B(n15615), .ZN(
        n15620) );
  NOR3_X1 U18822 ( .A1(n15639), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15618), .ZN(n15619) );
  AOI211_X1 U18823 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15621), .A(
        n15620), .B(n15619), .ZN(n15622) );
  OAI211_X1 U18824 ( .C1(n15624), .C2(n16476), .A(n15623), .B(n15622), .ZN(
        P2_U3025) );
  INV_X1 U18825 ( .A(n15625), .ZN(n15626) );
  NAND2_X1 U18826 ( .A1(n15626), .A2(n16471), .ZN(n15635) );
  INV_X1 U18827 ( .A(n15708), .ZN(n15778) );
  AOI21_X1 U18828 ( .B1(n15664), .B2(n15627), .A(n15778), .ZN(n15649) );
  NAND2_X1 U18829 ( .A1(n15628), .A2(n16479), .ZN(n15630) );
  OAI211_X1 U18830 ( .C1(n16474), .C2(n16411), .A(n15630), .B(n15629), .ZN(
        n15633) );
  XNOR2_X1 U18831 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15631) );
  NOR2_X1 U18832 ( .A1(n15639), .A2(n15631), .ZN(n15632) );
  AOI211_X1 U18833 ( .C1(n15649), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15633), .B(n15632), .ZN(n15634) );
  OAI211_X1 U18834 ( .C1(n15636), .C2(n16476), .A(n15635), .B(n15634), .ZN(
        P2_U3026) );
  NAND2_X1 U18835 ( .A1(n16457), .A2(n19089), .ZN(n15637) );
  OAI211_X1 U18836 ( .C1(n19088), .C2(n15834), .A(n15638), .B(n15637), .ZN(
        n15641) );
  NOR2_X1 U18837 ( .A1(n15639), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15640) );
  AOI211_X1 U18838 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15649), .A(
        n15641), .B(n15640), .ZN(n15645) );
  NAND3_X1 U18839 ( .A1(n15643), .A2(n16461), .A3(n15642), .ZN(n15644) );
  OAI211_X1 U18840 ( .C1(n15646), .C2(n15800), .A(n15645), .B(n15644), .ZN(
        P2_U3027) );
  INV_X1 U18841 ( .A(n15647), .ZN(n15648) );
  NOR3_X1 U18842 ( .A1(n15691), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15648), .ZN(n15657) );
  NAND2_X1 U18843 ( .A1(n15649), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15655) );
  OR2_X1 U18844 ( .A1(n15651), .A2(n15650), .ZN(n15652) );
  AND2_X1 U18845 ( .A1(n14331), .A2(n15652), .ZN(n19100) );
  AOI21_X1 U18846 ( .B1(n16457), .B2(n19100), .A(n15653), .ZN(n15654) );
  OAI211_X1 U18847 ( .C1(n19102), .C2(n15834), .A(n15655), .B(n15654), .ZN(
        n15656) );
  AOI211_X1 U18848 ( .C1(n15658), .C2(n16461), .A(n15657), .B(n15656), .ZN(
        n15659) );
  OAI21_X1 U18849 ( .B1(n15660), .B2(n15800), .A(n15659), .ZN(P2_U3028) );
  INV_X1 U18850 ( .A(n15661), .ZN(n15662) );
  OAI21_X1 U18851 ( .B1(n16461), .B2(n15663), .A(n15662), .ZN(n15666) );
  INV_X1 U18852 ( .A(n15664), .ZN(n15665) );
  NAND2_X1 U18853 ( .A1(n15665), .A2(n15708), .ZN(n15697) );
  OAI211_X1 U18854 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15667), .A(
        n15666), .B(n15697), .ZN(n15677) );
  AOI21_X1 U18855 ( .B1(n15687), .B2(n15832), .A(n15677), .ZN(n15676) );
  AOI21_X1 U18856 ( .B1(n19114), .B2(n16479), .A(n15668), .ZN(n15669) );
  OAI21_X1 U18857 ( .B1(n15670), .B2(n16474), .A(n15669), .ZN(n15671) );
  AOI21_X1 U18858 ( .B1(n15672), .B2(n16471), .A(n15671), .ZN(n15674) );
  OAI22_X1 U18859 ( .A1(n15690), .A2(n16476), .B1(n15704), .B2(n15691), .ZN(
        n15685) );
  NAND3_X1 U18860 ( .A1(n15685), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15675), .ZN(n15673) );
  OAI211_X1 U18861 ( .C1(n15676), .C2(n15675), .A(n15674), .B(n15673), .ZN(
        P2_U3029) );
  INV_X1 U18862 ( .A(n15677), .ZN(n15688) );
  OR2_X1 U18863 ( .A1(n15679), .A2(n15678), .ZN(n15680) );
  NAND2_X1 U18864 ( .A1(n14222), .A2(n15680), .ZN(n19124) );
  NAND2_X1 U18865 ( .A1(n15681), .A2(n16471), .ZN(n15683) );
  AOI22_X1 U18866 ( .A1(n19125), .A2(n16479), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19399), .ZN(n15682) );
  OAI211_X1 U18867 ( .C1(n16474), .C2(n19124), .A(n15683), .B(n15682), .ZN(
        n15684) );
  AOI21_X1 U18868 ( .B1(n15687), .B2(n15685), .A(n15684), .ZN(n15686) );
  OAI21_X1 U18869 ( .B1(n15688), .B2(n15687), .A(n15686), .ZN(P2_U3030) );
  OAI21_X1 U18870 ( .B1(n9852), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15690), .ZN(n16423) );
  INV_X1 U18871 ( .A(n15691), .ZN(n15705) );
  XNOR2_X1 U18872 ( .A(n15693), .B(n15692), .ZN(n19299) );
  NAND2_X1 U18873 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19399), .ZN(n15694) );
  OAI21_X1 U18874 ( .B1(n16474), .B2(n19299), .A(n15694), .ZN(n15695) );
  AOI21_X1 U18875 ( .B1(n19136), .B2(n16479), .A(n15695), .ZN(n15696) );
  OAI21_X1 U18876 ( .B1(n15697), .B2(n15704), .A(n15696), .ZN(n15703) );
  NAND2_X1 U18877 ( .A1(n15699), .A2(n15698), .ZN(n15701) );
  XOR2_X1 U18878 ( .A(n15701), .B(n15700), .Z(n16424) );
  NOR2_X1 U18879 ( .A1(n16424), .A2(n15800), .ZN(n15702) );
  AOI211_X1 U18880 ( .C1(n15705), .C2(n15704), .A(n15703), .B(n15702), .ZN(
        n15706) );
  OAI21_X1 U18881 ( .B1(n16476), .B2(n16423), .A(n15706), .ZN(P2_U3031) );
  NAND2_X1 U18882 ( .A1(n15794), .A2(n15707), .ZN(n15735) );
  INV_X1 U18883 ( .A(n15715), .ZN(n15710) );
  INV_X1 U18884 ( .A(n15707), .ZN(n15709) );
  OAI21_X1 U18885 ( .B1(n15792), .B2(n15709), .A(n15708), .ZN(n15743) );
  OAI21_X1 U18886 ( .B1(n15735), .B2(n15710), .A(n15743), .ZN(n15731) );
  INV_X1 U18887 ( .A(n19147), .ZN(n15714) );
  AOI21_X1 U18888 ( .B1(n15712), .B2(n15711), .A(n15692), .ZN(n19300) );
  AOI22_X1 U18889 ( .A1(n16457), .A2(n19300), .B1(n19399), .B2(
        P2_REIP_REG_14__SCAN_IN), .ZN(n15713) );
  OAI21_X1 U18890 ( .B1(n15714), .B2(n15834), .A(n15713), .ZN(n15717) );
  NOR3_X1 U18891 ( .A1(n15735), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15715), .ZN(n15716) );
  AOI211_X1 U18892 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15731), .A(
        n15717), .B(n15716), .ZN(n15720) );
  NAND2_X1 U18893 ( .A1(n15718), .A2(n16471), .ZN(n15719) );
  OAI211_X1 U18894 ( .C1(n15721), .C2(n16476), .A(n15720), .B(n15719), .ZN(
        P2_U3032) );
  NAND2_X1 U18895 ( .A1(n15722), .A2(n16461), .ZN(n15733) );
  OAI21_X1 U18896 ( .B1(n15735), .B2(n15742), .A(n15723), .ZN(n15730) );
  OR2_X1 U18897 ( .A1(n15725), .A2(n15724), .ZN(n15726) );
  NAND2_X1 U18898 ( .A1(n15726), .A2(n15711), .ZN(n19303) );
  NOR2_X1 U18899 ( .A1(n16474), .A2(n19303), .ZN(n15729) );
  OAI21_X1 U18900 ( .B1(n19156), .B2(n15834), .A(n15727), .ZN(n15728) );
  AOI211_X1 U18901 ( .C1(n15731), .C2(n15730), .A(n15729), .B(n15728), .ZN(
        n15732) );
  OAI211_X1 U18902 ( .C1(n15734), .C2(n15800), .A(n15733), .B(n15732), .ZN(
        P2_U3033) );
  NOR2_X1 U18903 ( .A1(n15735), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15745) );
  XNOR2_X1 U18904 ( .A(n15736), .B(n15737), .ZN(n19306) );
  NOR2_X1 U18905 ( .A1(n16474), .A2(n19306), .ZN(n15738) );
  AOI211_X1 U18906 ( .C1(n15740), .C2(n16479), .A(n15739), .B(n15738), .ZN(
        n15741) );
  OAI21_X1 U18907 ( .B1(n15743), .B2(n15742), .A(n15741), .ZN(n15744) );
  AOI211_X1 U18908 ( .C1(n15746), .C2(n16471), .A(n15745), .B(n15744), .ZN(
        n15747) );
  OAI21_X1 U18909 ( .B1(n15748), .B2(n16476), .A(n15747), .ZN(P2_U3034) );
  NOR2_X1 U18910 ( .A1(n15792), .A2(n15793), .ZN(n15779) );
  NOR3_X1 U18911 ( .A1(n15779), .A2(n15778), .A3(n15749), .ZN(n15757) );
  OAI21_X1 U18912 ( .B1(n15765), .B2(n15750), .A(n15736), .ZN(n19308) );
  XNOR2_X1 U18913 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15751) );
  NAND2_X1 U18914 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15794), .ZN(
        n15766) );
  NOR2_X1 U18915 ( .A1(n15751), .A2(n15766), .ZN(n15752) );
  AOI211_X1 U18916 ( .C1(n16479), .C2(n15754), .A(n15753), .B(n15752), .ZN(
        n15755) );
  OAI21_X1 U18917 ( .B1(n16474), .B2(n19308), .A(n15755), .ZN(n15756) );
  AOI211_X1 U18918 ( .C1(n15758), .C2(n16471), .A(n15757), .B(n15756), .ZN(
        n15759) );
  OAI21_X1 U18919 ( .B1(n15760), .B2(n16476), .A(n15759), .ZN(P2_U3035) );
  AOI21_X1 U18920 ( .B1(n15777), .B2(n15784), .A(n15761), .ZN(n16429) );
  NAND2_X1 U18921 ( .A1(n16429), .A2(n16461), .ZN(n15783) );
  NOR2_X1 U18922 ( .A1(n15762), .A2(n15763), .ZN(n15764) );
  OR2_X1 U18923 ( .A1(n15765), .A2(n15764), .ZN(n19311) );
  NOR2_X1 U18924 ( .A1(n19188), .A2(n19214), .ZN(n15768) );
  NOR2_X1 U18925 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15766), .ZN(
        n15767) );
  NOR2_X1 U18926 ( .A1(n15768), .A2(n15767), .ZN(n15769) );
  OAI21_X1 U18927 ( .B1(n16474), .B2(n19311), .A(n15769), .ZN(n15771) );
  NOR2_X1 U18928 ( .A1(n15834), .A2(n19193), .ZN(n15770) );
  NOR2_X1 U18929 ( .A1(n15771), .A2(n15770), .ZN(n15782) );
  NAND2_X1 U18930 ( .A1(n15772), .A2(n15786), .ZN(n15776) );
  NAND2_X1 U18931 ( .A1(n15774), .A2(n15773), .ZN(n15775) );
  XNOR2_X1 U18932 ( .A(n15776), .B(n15775), .ZN(n16431) );
  NAND2_X1 U18933 ( .A1(n16431), .A2(n16471), .ZN(n15781) );
  OR3_X1 U18934 ( .A1(n15779), .A2(n15778), .A3(n15777), .ZN(n15780) );
  NAND4_X1 U18935 ( .A1(n15783), .A2(n15782), .A3(n15781), .A4(n15780), .ZN(
        P2_U3036) );
  OAI21_X1 U18936 ( .B1(n15785), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15784), .ZN(n16437) );
  INV_X1 U18937 ( .A(n15786), .ZN(n15787) );
  OR2_X1 U18938 ( .A1(n15788), .A2(n15787), .ZN(n15789) );
  XNOR2_X1 U18939 ( .A(n15790), .B(n15789), .ZN(n16434) );
  INV_X1 U18940 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19962) );
  NOR2_X1 U18941 ( .A1(n19962), .A2(n19214), .ZN(n15791) );
  AOI221_X1 U18942 ( .B1(n15794), .B2(n15793), .C1(n15792), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15791), .ZN(n15799) );
  INV_X1 U18943 ( .A(n16439), .ZN(n19204) );
  NOR2_X1 U18944 ( .A1(n15795), .A2(n14263), .ZN(n15796) );
  OR2_X1 U18945 ( .A1(n15762), .A2(n15796), .ZN(n19313) );
  OAI22_X1 U18946 ( .A1(n15834), .A2(n19204), .B1(n16474), .B2(n19313), .ZN(
        n15797) );
  INV_X1 U18947 ( .A(n15797), .ZN(n15798) );
  OAI211_X1 U18948 ( .C1(n16434), .C2(n15800), .A(n15799), .B(n15798), .ZN(
        n15801) );
  INV_X1 U18949 ( .A(n15801), .ZN(n15802) );
  OAI21_X1 U18950 ( .B1(n16437), .B2(n16476), .A(n15802), .ZN(P2_U3037) );
  NOR3_X1 U18951 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n16464), .A3(
        n16463), .ZN(n15811) );
  OR2_X1 U18952 ( .A1(n15804), .A2(n15803), .ZN(n15805) );
  NAND2_X1 U18953 ( .A1(n15805), .A2(n14262), .ZN(n19319) );
  OAI21_X1 U18954 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16463), .A(
        n16456), .ZN(n15806) );
  NAND2_X1 U18955 ( .A1(n15806), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15809) );
  INV_X1 U18956 ( .A(n19217), .ZN(n15807) );
  AOI22_X1 U18957 ( .A1(n16479), .A2(n15807), .B1(n19399), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n15808) );
  OAI211_X1 U18958 ( .C1(n16474), .C2(n19319), .A(n15809), .B(n15808), .ZN(
        n15810) );
  AOI211_X1 U18959 ( .C1(n15812), .C2(n16471), .A(n15811), .B(n15810), .ZN(
        n15813) );
  OAI21_X1 U18960 ( .B1(n15814), .B2(n16476), .A(n15813), .ZN(P2_U3039) );
  AOI22_X1 U18961 ( .A1(n15817), .A2(n15816), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15815), .ZN(n15820) );
  XNOR2_X1 U18962 ( .A(n15818), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15819) );
  XNOR2_X1 U18963 ( .A(n15820), .B(n15819), .ZN(n19401) );
  NAND2_X1 U18964 ( .A1(n19401), .A2(n16471), .ZN(n15830) );
  INV_X1 U18965 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19955) );
  NOR2_X1 U18966 ( .A1(n19955), .A2(n19214), .ZN(n15821) );
  AOI221_X1 U18967 ( .B1(n15823), .B2(n15826), .C1(n15822), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n15821), .ZN(n15829) );
  AOI22_X1 U18968 ( .A1(n19402), .A2(n16479), .B1(n16457), .B2(n15824), .ZN(
        n15828) );
  XNOR2_X1 U18969 ( .A(n15825), .B(n15826), .ZN(n19405) );
  NAND2_X1 U18970 ( .A1(n19405), .A2(n16461), .ZN(n15827) );
  NAND4_X1 U18971 ( .A1(n15830), .A2(n15829), .A3(n15828), .A4(n15827), .ZN(
        P2_U3042) );
  OAI211_X1 U18972 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15832), .B(n15831), .ZN(n15842) );
  OAI22_X1 U18973 ( .A1(n15835), .A2(n15834), .B1(n16469), .B2(n15833), .ZN(
        n15836) );
  INV_X1 U18974 ( .A(n15836), .ZN(n15841) );
  AOI22_X1 U18975 ( .A1(n15837), .A2(n16471), .B1(P2_REIP_REG_1__SCAN_IN), 
        .B2(n19399), .ZN(n15840) );
  AOI22_X1 U18976 ( .A1(n16461), .A2(n15838), .B1(n16457), .B2(n20030), .ZN(
        n15839) );
  NAND4_X1 U18977 ( .A1(n15842), .A2(n15841), .A3(n15840), .A4(n15839), .ZN(
        P2_U3045) );
  INV_X1 U18978 ( .A(n10985), .ZN(n15844) );
  NAND2_X1 U18979 ( .A1(n15844), .A2(n15843), .ZN(n15853) );
  MUX2_X1 U18980 ( .A(n15853), .B(n14322), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15845) );
  AOI21_X1 U18981 ( .B1(n11289), .B2(n15863), .A(n15845), .ZN(n16487) );
  INV_X1 U18982 ( .A(n16487), .ZN(n15847) );
  AOI22_X1 U18983 ( .A1(n15847), .A2(n15858), .B1(P2_STATE2_REG_1__SCAN_IN), 
        .B2(n15846), .ZN(n15848) );
  OAI21_X1 U18984 ( .B1(n15849), .B2(n15882), .A(n15848), .ZN(n15850) );
  MUX2_X1 U18985 ( .A(n15850), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15883), .Z(P2_U3601) );
  INV_X1 U18986 ( .A(n15851), .ZN(n15860) );
  INV_X1 U18987 ( .A(n15882), .ZN(n16519) );
  NAND2_X1 U18988 ( .A1(n11288), .A2(n15863), .ZN(n15857) );
  NOR2_X1 U18989 ( .A1(n15852), .A2(n10370), .ZN(n15854) );
  AOI22_X1 U18990 ( .A1(n14322), .A2(n15855), .B1(n15854), .B2(n15853), .ZN(
        n15856) );
  NAND2_X1 U18991 ( .A1(n15857), .A2(n15856), .ZN(n16485) );
  AOI22_X1 U18992 ( .A1(n20026), .A2(n16519), .B1(n15858), .B2(n16485), .ZN(
        n15859) );
  OAI21_X1 U18993 ( .B1(n15861), .B2(n15860), .A(n15859), .ZN(n15862) );
  MUX2_X1 U18994 ( .A(n15862), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15883), .Z(P2_U3600) );
  NAND2_X1 U18995 ( .A1(n11300), .A2(n15863), .ZN(n15880) );
  NOR2_X1 U18996 ( .A1(n15865), .A2(n15864), .ZN(n15868) );
  INV_X1 U18997 ( .A(n15866), .ZN(n15867) );
  MUX2_X1 U18998 ( .A(n15868), .B(n15867), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15878) );
  OAI211_X1 U18999 ( .C1(n15870), .C2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14322), .B(n15869), .ZN(n15876) );
  OAI21_X1 U19000 ( .B1(n10193), .B2(n15872), .A(n15871), .ZN(n15873) );
  NAND2_X1 U19001 ( .A1(n15874), .A2(n15873), .ZN(n15875) );
  NAND2_X1 U19002 ( .A1(n15876), .A2(n15875), .ZN(n15877) );
  NOR2_X1 U19003 ( .A1(n15878), .A2(n15877), .ZN(n15879) );
  NAND2_X1 U19004 ( .A1(n15880), .A2(n15879), .ZN(n16491) );
  INV_X1 U19005 ( .A(n16491), .ZN(n15881) );
  OAI22_X1 U19006 ( .A1(n19503), .A2(n15882), .B1(n20006), .B2(n15881), .ZN(
        n15884) );
  MUX2_X1 U19007 ( .A(n15884), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15883), .Z(P2_U3596) );
  OAI21_X1 U19008 ( .B1(n19545), .B2(n21345), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15885) );
  NAND2_X1 U19009 ( .A1(n15885), .A2(n20004), .ZN(n15889) );
  NOR2_X1 U19010 ( .A1(n15886), .A2(n19694), .ZN(n19764) );
  NAND2_X1 U19011 ( .A1(n19764), .A2(n20017), .ZN(n15893) );
  INV_X1 U19012 ( .A(n15890), .ZN(n15887) );
  NAND2_X1 U19013 ( .A1(n20017), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19610) );
  NOR2_X1 U19014 ( .A1(n19410), .A2(n19610), .ZN(n19544) );
  OAI21_X1 U19015 ( .B1(n15887), .B2(n19544), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15888) );
  INV_X1 U19016 ( .A(n15889), .ZN(n15894) );
  AOI21_X1 U19017 ( .B1(n15890), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n15891) );
  OAI21_X1 U19018 ( .B1(n15891), .B2(n19544), .A(n19851), .ZN(n15892) );
  INV_X1 U19019 ( .A(n19549), .ZN(n15895) );
  NAND2_X1 U19020 ( .A1(n15895), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n15897) );
  AOI22_X1 U19021 ( .A1(n19792), .A2(n21345), .B1(n19842), .B2(n19544), .ZN(
        n15896) );
  OAI211_X1 U19022 ( .C1(n19527), .C2(n19733), .A(n15897), .B(n15896), .ZN(
        n15898) );
  AOI21_X1 U19023 ( .B1(n19791), .B2(n19546), .A(n15898), .ZN(n15899) );
  INV_X1 U19024 ( .A(n15899), .ZN(P2_U3080) );
  AOI22_X1 U19025 ( .A1(n19811), .A2(n21345), .B1(n19859), .B2(n19544), .ZN(
        n15901) );
  NAND2_X1 U19026 ( .A1(n19863), .A2(n19545), .ZN(n15900) );
  OAI211_X1 U19027 ( .C1(n19549), .C2(n15902), .A(n15901), .B(n15900), .ZN(
        n15903) );
  AOI21_X1 U19028 ( .B1(n19858), .B2(n19546), .A(n15903), .ZN(n15904) );
  INV_X1 U19029 ( .A(n15904), .ZN(P2_U3081) );
  AOI22_X1 U19030 ( .A1(n19831), .A2(n21345), .B1(n19908), .B2(n19544), .ZN(
        n15906) );
  NAND2_X1 U19031 ( .A1(n19914), .A2(n19545), .ZN(n15905) );
  OAI211_X1 U19032 ( .C1(n19549), .C2(n15907), .A(n15906), .B(n15905), .ZN(
        n15908) );
  AOI21_X1 U19033 ( .B1(n19907), .B2(n19546), .A(n15908), .ZN(n15909) );
  INV_X1 U19034 ( .A(n15909), .ZN(P2_U3087) );
  INV_X1 U19035 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n21312) );
  INV_X1 U19036 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17143) );
  INV_X1 U19037 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17243) );
  INV_X1 U19038 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16912) );
  INV_X1 U19039 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17350) );
  NOR3_X4 U19040 ( .A1(n16077), .A2(n15912), .A3(n18883), .ZN(n17424) );
  INV_X1 U19041 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17049) );
  NOR2_X1 U19042 ( .A1(n17034), .A2(n17049), .ZN(n17396) );
  INV_X1 U19043 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17425) );
  INV_X1 U19044 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17420) );
  NOR2_X1 U19045 ( .A1(n17425), .A2(n17420), .ZN(n17395) );
  INV_X1 U19046 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17008) );
  NOR2_X2 U19047 ( .A1(n17401), .A2(n17008), .ZN(n17397) );
  NOR2_X2 U19048 ( .A1(n17389), .A2(n17390), .ZN(n17393) );
  INV_X1 U19050 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16936) );
  NOR2_X2 U19051 ( .A1(n17347), .A2(n16936), .ZN(n17310) );
  INV_X1 U19052 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n21242) );
  NOR2_X2 U19053 ( .A1(n17240), .A2(n21242), .ZN(n17197) );
  NOR2_X2 U19054 ( .A1(n17478), .A2(n17183), .ZN(n17194) );
  NAND3_X1 U19055 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n17194), .ZN(n17170) );
  NOR3_X2 U19056 ( .A1(n21312), .A2(n17143), .A3(n17170), .ZN(n17157) );
  AND2_X2 U19057 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17157), .ZN(n17142) );
  AND2_X2 U19058 ( .A1(n17142), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n17137) );
  AND2_X2 U19059 ( .A1(n17137), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n17134) );
  INV_X1 U19060 ( .A(n17126), .ZN(n17129) );
  NAND2_X1 U19061 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17129), .ZN(n17117) );
  INV_X1 U19062 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17118) );
  INV_X1 U19063 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17125) );
  NOR2_X1 U19064 ( .A1(n17118), .A2(n17125), .ZN(n17078) );
  NAND2_X1 U19065 ( .A1(n18410), .A2(n17424), .ZN(n17426) );
  INV_X2 U19066 ( .A(n17422), .ZN(n17414) );
  NAND2_X1 U19067 ( .A1(n17414), .A2(n17126), .ZN(n17124) );
  OAI21_X1 U19068 ( .B1(n17078), .B2(n17426), .A(n17124), .ZN(n17120) );
  AOI22_X1 U19069 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15913) );
  OAI21_X1 U19070 ( .B1(n17322), .B2(n17313), .A(n15913), .ZN(n15924) );
  AOI22_X1 U19071 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15921) );
  INV_X1 U19072 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17321) );
  OAI22_X1 U19073 ( .A1(n17317), .A2(n17321), .B1(n13090), .B2(n21200), .ZN(
        n15919) );
  AOI22_X1 U19074 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17314), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15917) );
  AOI22_X1 U19075 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15916) );
  AOI22_X1 U19076 ( .A1(n17377), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15915) );
  NAND3_X1 U19077 ( .A1(n15917), .A2(n15916), .A3(n15915), .ZN(n15918) );
  AOI211_X1 U19078 ( .C1(n17086), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n15919), .B(n15918), .ZN(n15920) );
  OAI211_X1 U19079 ( .C1(n15914), .C2(n15922), .A(n15921), .B(n15920), .ZN(
        n15923) );
  AOI211_X1 U19080 ( .C1(n9720), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n15924), .B(n15923), .ZN(n17127) );
  AOI22_X1 U19081 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n9716), .ZN(n15925) );
  OAI21_X1 U19082 ( .B1(n17354), .B2(n17205), .A(n15925), .ZN(n15935) );
  AOI22_X1 U19083 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17215), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15933) );
  AOI22_X1 U19084 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n13113), .ZN(n15926) );
  OAI21_X1 U19085 ( .B1(n13090), .B2(n18601), .A(n15926), .ZN(n15931) );
  AOI22_X1 U19086 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15928) );
  AOI22_X1 U19087 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17367), .B1(
        n9720), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15927) );
  OAI211_X1 U19088 ( .C1(n15929), .C2(n17298), .A(n15928), .B(n15927), .ZN(
        n15930) );
  AOI211_X1 U19089 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n17375), .A(
        n15931), .B(n15930), .ZN(n15932) );
  OAI211_X1 U19090 ( .C1(n17210), .C2(n18421), .A(n15933), .B(n15932), .ZN(
        n15934) );
  AOI211_X1 U19091 ( .C1(n9765), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n15935), .B(n15934), .ZN(n17135) );
  AOI22_X1 U19092 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15945) );
  AOI22_X1 U19093 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9720), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15944) );
  AOI22_X1 U19094 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15943) );
  OAI22_X1 U19095 ( .A1(n17210), .A2(n18418), .B1(n15914), .B2(n21155), .ZN(
        n15941) );
  AOI22_X1 U19096 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15939) );
  AOI22_X1 U19097 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15938) );
  AOI22_X1 U19098 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15937) );
  NAND2_X1 U19099 ( .A1(n17377), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n15936) );
  NAND4_X1 U19100 ( .A1(n15939), .A2(n15938), .A3(n15937), .A4(n15936), .ZN(
        n15940) );
  AOI211_X1 U19101 ( .C1(n9767), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n15941), .B(n15940), .ZN(n15942) );
  NAND4_X1 U19102 ( .A1(n15945), .A2(n15944), .A3(n15943), .A4(n15942), .ZN(
        n17139) );
  AOI22_X1 U19103 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17332), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15955) );
  AOI22_X1 U19104 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15954) );
  OAI22_X1 U19105 ( .A1(n17371), .A2(n21093), .B1(n17210), .B2(n21122), .ZN(
        n15952) );
  INV_X1 U19106 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n21266) );
  AOI22_X1 U19107 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15950) );
  AOI22_X1 U19108 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15947) );
  AOI22_X1 U19109 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15946) );
  OAI211_X1 U19110 ( .C1(n17317), .C2(n18438), .A(n15947), .B(n15946), .ZN(
        n15948) );
  AOI21_X1 U19111 ( .B1(n13113), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n15948), .ZN(n15949) );
  OAI211_X1 U19112 ( .C1(n13090), .C2(n21266), .A(n15950), .B(n15949), .ZN(
        n15951) );
  AOI211_X1 U19113 ( .C1(n17377), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n15952), .B(n15951), .ZN(n15953) );
  NAND3_X1 U19114 ( .A1(n15955), .A2(n15954), .A3(n15953), .ZN(n17140) );
  NAND2_X1 U19115 ( .A1(n17139), .A2(n17140), .ZN(n17138) );
  NOR2_X1 U19116 ( .A1(n17135), .A2(n17138), .ZN(n17132) );
  INV_X1 U19117 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18424) );
  AOI22_X1 U19118 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15966) );
  AOI22_X1 U19119 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15957) );
  AOI22_X1 U19120 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15956) );
  OAI211_X1 U19121 ( .C1(n17298), .C2(n15958), .A(n15957), .B(n15956), .ZN(
        n15964) );
  AOI22_X1 U19122 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15962) );
  AOI22_X1 U19123 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15961) );
  AOI22_X1 U19124 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15960) );
  NAND2_X1 U19125 ( .A1(n13113), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n15959) );
  NAND4_X1 U19126 ( .A1(n15962), .A2(n15961), .A3(n15960), .A4(n15959), .ZN(
        n15963) );
  AOI211_X1 U19127 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n15964), .B(n15963), .ZN(n15965) );
  OAI211_X1 U19128 ( .C1(n17210), .C2(n18424), .A(n15966), .B(n15965), .ZN(
        n17131) );
  NAND2_X1 U19129 ( .A1(n17132), .A2(n17131), .ZN(n17130) );
  NOR2_X1 U19130 ( .A1(n17127), .A2(n17130), .ZN(n17452) );
  AOI22_X1 U19131 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9716), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15978) );
  AOI22_X1 U19132 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17332), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15977) );
  AOI22_X1 U19133 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15976) );
  OAI22_X1 U19134 ( .A1(n13148), .A2(n15968), .B1(n13090), .B2(n15967), .ZN(
        n15974) );
  AOI22_X1 U19135 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15972) );
  AOI22_X1 U19136 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15971) );
  AOI22_X1 U19137 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15970) );
  NAND2_X1 U19138 ( .A1(n17377), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n15969) );
  NAND4_X1 U19139 ( .A1(n15972), .A2(n15971), .A3(n15970), .A4(n15969), .ZN(
        n15973) );
  AOI211_X1 U19140 ( .C1(n17086), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n15974), .B(n15973), .ZN(n15975) );
  NAND4_X1 U19141 ( .A1(n15978), .A2(n15977), .A3(n15976), .A4(n15975), .ZN(
        n17451) );
  NAND2_X1 U19142 ( .A1(n17452), .A2(n17451), .ZN(n17450) );
  INV_X1 U19143 ( .A(n17450), .ZN(n17113) );
  AOI22_X1 U19144 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15988) );
  AOI22_X1 U19145 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15987) );
  AOI22_X1 U19146 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15986) );
  INV_X1 U19147 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n21226) );
  OAI22_X1 U19148 ( .A1(n17327), .A2(n21226), .B1(n13090), .B2(n17278), .ZN(
        n15984) );
  AOI22_X1 U19149 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15982) );
  AOI22_X1 U19150 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9716), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15981) );
  AOI22_X1 U19151 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15980) );
  NAND2_X1 U19152 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n15979) );
  NAND4_X1 U19153 ( .A1(n15982), .A2(n15981), .A3(n15980), .A4(n15979), .ZN(
        n15983) );
  AOI211_X1 U19154 ( .C1(n17377), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n15984), .B(n15983), .ZN(n15985) );
  NAND4_X1 U19155 ( .A1(n15988), .A2(n15987), .A3(n15986), .A4(n15985), .ZN(
        n17114) );
  XOR2_X1 U19156 ( .A(n17113), .B(n17114), .Z(n17445) );
  AOI22_X1 U19157 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17120), .B1(n17422), 
        .B2(n17445), .ZN(n15989) );
  OAI21_X1 U19158 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17117), .A(n15989), .ZN(
        P3_U2675) );
  NOR2_X1 U19159 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18983), .ZN(
        n18414) );
  INV_X1 U19160 ( .A(n18414), .ZN(n15991) );
  INV_X1 U19161 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18365) );
  NAND3_X1 U19162 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18982)
         );
  INV_X1 U19163 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21141) );
  NAND3_X1 U19164 ( .A1(n17210), .A2(n16008), .A3(n21141), .ZN(n18364) );
  INV_X1 U19165 ( .A(n18364), .ZN(n15990) );
  OAI221_X1 U19166 ( .B1(n18365), .B2(n18982), .C1(n15990), .C2(n18982), .A(
        n18620), .ZN(n18370) );
  NAND2_X1 U19167 ( .A1(n15991), .A2(n18370), .ZN(n15994) );
  INV_X1 U19168 ( .A(n15994), .ZN(n15993) );
  INV_X1 U19169 ( .A(n15997), .ZN(n18718) );
  OAI22_X1 U19170 ( .A1(n17851), .A2(n19028), .B1(n18834), .B2(n18983), .ZN(
        n15996) );
  NAND3_X1 U19171 ( .A1(n18833), .A2(n18370), .A3(n15996), .ZN(n15992) );
  OAI221_X1 U19172 ( .B1(n18833), .B2(n15993), .C1(n18833), .C2(n18718), .A(
        n15992), .ZN(P3_U2864) );
  NOR2_X1 U19173 ( .A1(n18833), .A2(n18855), .ZN(n18524) );
  INV_X1 U19174 ( .A(n18524), .ZN(n18372) );
  NOR2_X1 U19175 ( .A1(n17851), .A2(n19028), .ZN(n15995) );
  AOI221_X1 U19176 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18372), .C1(n15995), 
        .C2(n18372), .A(n15994), .ZN(n18369) );
  OAI221_X1 U19177 ( .B1(n15997), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n15997), .C2(n15996), .A(n18370), .ZN(n18367) );
  AOI22_X1 U19178 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18369), .B1(
        n18367), .B2(n18855), .ZN(P3_U2865) );
  INV_X1 U19179 ( .A(n19034), .ZN(n18894) );
  NOR2_X1 U19180 ( .A1(n18894), .A2(n16677), .ZN(n16004) );
  NAND2_X1 U19181 ( .A1(n19033), .A2(n17639), .ZN(n18869) );
  AOI21_X1 U19182 ( .B1(n16004), .B2(n17578), .A(n15999), .ZN(n16006) );
  NAND2_X1 U19183 ( .A1(n18809), .A2(n16000), .ZN(n16005) );
  NAND3_X1 U19184 ( .A1(n16006), .A2(n16005), .A3(n16078), .ZN(n18852) );
  NOR2_X1 U19185 ( .A1(n18365), .A2(n18982), .ZN(n16007) );
  NOR2_X1 U19186 ( .A1(n18983), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18378) );
  INV_X1 U19187 ( .A(n16697), .ZN(n18841) );
  AOI21_X1 U19188 ( .B1(n16008), .B2(n21141), .A(n18841), .ZN(n18865) );
  NAND3_X1 U19189 ( .A1(n19012), .A2(n19010), .A3(n18865), .ZN(n16009) );
  OAI21_X1 U19190 ( .B1(n19012), .B2(n21141), .A(n16009), .ZN(P3_U3284) );
  NAND2_X1 U19191 ( .A1(n18267), .A2(n18832), .ZN(n18252) );
  OAI21_X1 U19192 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18237), .A(
        n16010), .ZN(n16568) );
  OAI21_X1 U19193 ( .B1(n16011), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18338), .ZN(n16013) );
  AOI221_X1 U19194 ( .B1(n16568), .B2(n18358), .C1(n16013), .C2(n18358), .A(
        n16012), .ZN(n16020) );
  NAND2_X1 U19195 ( .A1(n16015), .A2(n16014), .ZN(n16016) );
  XOR2_X1 U19196 ( .A(n16016), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16540) );
  NOR3_X1 U19197 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16017), .A3(
        n16533), .ZN(n16018) );
  AOI21_X1 U19198 ( .B1(n18263), .B2(n16540), .A(n16018), .ZN(n16019) );
  INV_X2 U19199 ( .A(n18358), .ZN(n18348) );
  NAND2_X1 U19200 ( .A1(n18348), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16545) );
  OAI211_X1 U19201 ( .C1(n16020), .C2(n16537), .A(n16019), .B(n16545), .ZN(
        P3_U2833) );
  INV_X1 U19202 ( .A(n16022), .ZN(n16028) );
  INV_X1 U19203 ( .A(n20720), .ZN(n16027) );
  INV_X1 U19204 ( .A(n16029), .ZN(n16021) );
  AOI21_X1 U19205 ( .B1(n16022), .B2(n16021), .A(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16026) );
  AND2_X1 U19206 ( .A1(n16024), .A2(n16023), .ZN(n16025) );
  OAI33_X1 U19207 ( .A1(n20368), .A2(n16029), .A3(n16028), .B1(n16027), .B2(
        n16026), .B3(n16025), .ZN(n16033) );
  INV_X1 U19208 ( .A(n16033), .ZN(n16031) );
  OAI21_X1 U19209 ( .B1(n16031), .B2(n20562), .A(n16030), .ZN(n16032) );
  OAI21_X1 U19210 ( .B1(n16033), .B2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16032), .ZN(n16034) );
  AOI222_X1 U19211 ( .A1(n21136), .A2(n16035), .B1(n21136), .B2(n16034), .C1(
        n16035), .C2(n16034), .ZN(n16044) );
  INV_X1 U19212 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n16037) );
  AOI21_X1 U19213 ( .B1(n20063), .B2(n16037), .A(n16036), .ZN(n16039) );
  NOR4_X1 U19214 ( .A1(n16041), .A2(n16040), .A3(n16039), .A4(n16038), .ZN(
        n16042) );
  OAI211_X1 U19215 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n16044), .A(
        n16043), .B(n16042), .ZN(n16053) );
  INV_X1 U19216 ( .A(n16073), .ZN(n16046) );
  NAND2_X1 U19217 ( .A1(n16046), .A2(n16045), .ZN(n16050) );
  OAI21_X1 U19218 ( .B1(n16048), .B2(n21018), .A(n16047), .ZN(n16049) );
  OAI21_X1 U19219 ( .B1(n16051), .B2(n16050), .A(n16049), .ZN(n16378) );
  AOI221_X1 U19220 ( .B1(n11887), .B2(n14021), .C1(n16053), .C2(n14021), .A(
        n16378), .ZN(n16382) );
  AOI21_X1 U19221 ( .B1(n16054), .B2(n16053), .A(n16052), .ZN(n16056) );
  OAI211_X1 U19222 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21018), .A(n16056), 
        .B(n16055), .ZN(n16057) );
  NOR2_X1 U19223 ( .A1(n16382), .A2(n16057), .ZN(n16062) );
  NAND2_X1 U19224 ( .A1(n16059), .A2(n16058), .ZN(n16060) );
  NAND2_X1 U19225 ( .A1(n11887), .A2(n16060), .ZN(n16061) );
  OAI22_X1 U19226 ( .A1(n16062), .A2(n11887), .B1(n16382), .B2(n16061), .ZN(
        P1_U3161) );
  OR2_X1 U19227 ( .A1(n16064), .A2(n16063), .ZN(n16065) );
  OAI21_X1 U19228 ( .B1(n16066), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16065), .ZN(n16067) );
  XOR2_X1 U19229 ( .A(n16069), .B(n16067), .Z(n16201) );
  AND2_X1 U19230 ( .A1(n16068), .A2(n16291), .ZN(n16281) );
  AOI22_X1 U19231 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n20232), .B1(n16281), 
        .B2(n16069), .ZN(n16071) );
  AOI22_X1 U19232 ( .A1(n16278), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n16104), .B2(n16367), .ZN(n16070) );
  OAI211_X1 U19233 ( .C1(n16201), .C2(n16370), .A(n16071), .B(n16070), .ZN(
        P1_U3010) );
  INV_X1 U19234 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20940) );
  OAI221_X1 U19235 ( .B1(n20924), .B2(HOLD), .C1(n20924), .C2(n20940), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n16074) );
  INV_X1 U19236 ( .A(HOLD), .ZN(n20937) );
  OAI211_X1 U19237 ( .C1(n20940), .C2(n20937), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n16072) );
  NAND3_X1 U19238 ( .A1(n16074), .A2(n16073), .A3(n16072), .ZN(P1_U3195) );
  AND2_X1 U19239 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n20163), .ZN(P1_U2905)
         );
  NOR3_X1 U19240 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16075) );
  NOR2_X1 U19241 ( .A1(n19922), .A2(n19923), .ZN(n16513) );
  NOR4_X1 U19242 ( .A1(n16075), .A2(n16518), .A3(n16527), .A4(n16513), .ZN(
        P2_U3178) );
  AOI221_X1 U19243 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16527), .C1(n20045), .C2(
        n16527), .A(n19851), .ZN(n20041) );
  INV_X1 U19244 ( .A(n20041), .ZN(n20038) );
  NOR2_X1 U19245 ( .A1(n16493), .A2(n20038), .ZN(P2_U3047) );
  INV_X1 U19246 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17637) );
  NAND2_X1 U19247 ( .A1(n18410), .A2(n17427), .ZN(n17479) );
  NOR2_X1 U19248 ( .A1(n17637), .A2(n17479), .ZN(n17566) );
  INV_X1 U19249 ( .A(n17566), .ZN(n17577) );
  NAND2_X1 U19250 ( .A1(n17565), .A2(n17577), .ZN(n17576) );
  AOI22_X1 U19251 ( .A1(n17574), .A2(BUF2_REG_0__SCAN_IN), .B1(n17573), .B2(
        n16080), .ZN(n16081) );
  OAI221_X1 U19252 ( .B1(n17576), .B2(n17637), .C1(n17576), .C2(n17479), .A(
        n16081), .ZN(P3_U2735) );
  AOI22_X1 U19253 ( .A1(n20133), .A2(P1_EBX_REG_23__SCAN_IN), .B1(n20131), 
        .B2(n16082), .ZN(n16091) );
  INV_X1 U19254 ( .A(n16083), .ZN(n16087) );
  INV_X1 U19255 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n16085) );
  NAND2_X1 U19256 ( .A1(n16098), .A2(n16084), .ZN(n16097) );
  NOR2_X1 U19257 ( .A1(n16085), .A2(n16097), .ZN(n16093) );
  AOI21_X1 U19258 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n16093), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n16086) );
  OAI22_X1 U19259 ( .A1(n16088), .A2(n16182), .B1(n16087), .B2(n16086), .ZN(
        n16089) );
  AOI21_X1 U19260 ( .B1(n20127), .B2(n16272), .A(n16089), .ZN(n16090) );
  OAI211_X1 U19261 ( .C1(n16092), .C2(n20094), .A(n16091), .B(n16090), .ZN(
        P1_U2817) );
  AOI22_X1 U19262 ( .A1(n20133), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20128), .ZN(n16103) );
  INV_X1 U19263 ( .A(n16196), .ZN(n16094) );
  INV_X1 U19264 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20970) );
  AOI22_X1 U19265 ( .A1(n16094), .A2(n20131), .B1(n16093), .B2(n20970), .ZN(
        n16102) );
  XNOR2_X1 U19266 ( .A(n16096), .B(n16095), .ZN(n16279) );
  AOI22_X1 U19267 ( .A1(n16193), .A2(n20099), .B1(n20127), .B2(n16279), .ZN(
        n16101) );
  NOR2_X1 U19268 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n16097), .ZN(n16105) );
  OAI21_X1 U19269 ( .B1(n16099), .B2(n16098), .A(n16135), .ZN(n16113) );
  OAI21_X1 U19270 ( .B1(n16105), .B2(n16113), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n16100) );
  NAND4_X1 U19271 ( .A1(n16103), .A2(n16102), .A3(n16101), .A4(n16100), .ZN(
        P1_U2818) );
  AOI22_X1 U19272 ( .A1(n20133), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20128), .ZN(n16109) );
  AOI22_X1 U19273 ( .A1(n16197), .A2(n20131), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n16113), .ZN(n16108) );
  AOI22_X1 U19274 ( .A1(n16198), .A2(n20099), .B1(n20127), .B2(n16104), .ZN(
        n16107) );
  INV_X1 U19275 ( .A(n16105), .ZN(n16106) );
  NAND4_X1 U19276 ( .A1(n16109), .A2(n16108), .A3(n16107), .A4(n16106), .ZN(
        P1_U2819) );
  INV_X1 U19277 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16110) );
  OAI22_X1 U19278 ( .A1(n16110), .A2(n20094), .B1(n16178), .B2(n16206), .ZN(
        n16111) );
  AOI21_X1 U19279 ( .B1(n20133), .B2(P1_EBX_REG_20__SCAN_IN), .A(n16111), .ZN(
        n16116) );
  OAI21_X1 U19280 ( .B1(n20966), .B2(n16112), .A(n20965), .ZN(n16114) );
  AOI22_X1 U19281 ( .A1(n16203), .A2(n20099), .B1(n16114), .B2(n16113), .ZN(
        n16115) );
  OAI211_X1 U19282 ( .C1(n16168), .C2(n16117), .A(n16116), .B(n16115), .ZN(
        P1_U2820) );
  OAI22_X1 U19283 ( .A1(n20095), .A2(n16119), .B1(n16178), .B2(n16118), .ZN(
        n16120) );
  AOI211_X1 U19284 ( .C1(n20128), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20232), .B(n16120), .ZN(n16122) );
  OAI211_X1 U19285 ( .C1(n16135), .C2(n20963), .A(n16122), .B(n16121), .ZN(
        n16123) );
  AOI21_X1 U19286 ( .B1(n16124), .B2(n20099), .A(n16123), .ZN(n16125) );
  OAI21_X1 U19287 ( .B1(n16168), .B2(n16298), .A(n16125), .ZN(P1_U2822) );
  INV_X1 U19288 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21097) );
  NOR2_X1 U19289 ( .A1(n21267), .A2(n21097), .ZN(n16145) );
  AOI21_X1 U19290 ( .B1(n16145), .B2(n16136), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n16134) );
  OAI22_X1 U19291 ( .A1(n20095), .A2(n16126), .B1(n21087), .B2(n20094), .ZN(
        n16127) );
  AOI211_X1 U19292 ( .C1(n20131), .C2(n16128), .A(n20232), .B(n16127), .ZN(
        n16133) );
  OAI22_X1 U19293 ( .A1(n16130), .A2(n16182), .B1(n16168), .B2(n16129), .ZN(
        n16131) );
  INV_X1 U19294 ( .A(n16131), .ZN(n16132) );
  OAI211_X1 U19295 ( .C1(n16135), .C2(n16134), .A(n16133), .B(n16132), .ZN(
        P1_U2823) );
  OAI21_X1 U19296 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), 
        .A(n16136), .ZN(n16144) );
  NAND2_X1 U19297 ( .A1(n20128), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16137) );
  OAI211_X1 U19298 ( .C1(n16178), .C2(n16211), .A(n16137), .B(n20100), .ZN(
        n16140) );
  NOR2_X1 U19299 ( .A1(n16138), .A2(n16168), .ZN(n16139) );
  AOI211_X1 U19300 ( .C1(n20133), .C2(P1_EBX_REG_16__SCAN_IN), .A(n16140), .B(
        n16139), .ZN(n16141) );
  OAI21_X1 U19301 ( .B1(n16154), .B2(n21097), .A(n16141), .ZN(n16142) );
  AOI21_X1 U19302 ( .B1(n16207), .B2(n20099), .A(n16142), .ZN(n16143) );
  OAI21_X1 U19303 ( .B1(n16145), .B2(n16144), .A(n16143), .ZN(P1_U2824) );
  NOR2_X1 U19304 ( .A1(n16146), .A2(n16174), .ZN(n16147) );
  NOR2_X1 U19305 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16147), .ZN(n16155) );
  AOI22_X1 U19306 ( .A1(n20133), .A2(P1_EBX_REG_14__SCAN_IN), .B1(n20131), 
        .B2(n16218), .ZN(n16153) );
  INV_X1 U19307 ( .A(n16148), .ZN(n16219) );
  NOR2_X1 U19308 ( .A1(n16313), .A2(n16168), .ZN(n16151) );
  INV_X1 U19309 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16149) );
  OAI21_X1 U19310 ( .B1(n20094), .B2(n16149), .A(n20100), .ZN(n16150) );
  AOI211_X1 U19311 ( .C1(n16219), .C2(n20099), .A(n16151), .B(n16150), .ZN(
        n16152) );
  OAI211_X1 U19312 ( .C1(n16155), .C2(n16154), .A(n16153), .B(n16152), .ZN(
        P1_U2826) );
  AOI21_X1 U19313 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16156), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16164) );
  AOI22_X1 U19314 ( .A1(n20133), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n20131), 
        .B2(n16223), .ZN(n16162) );
  INV_X1 U19315 ( .A(n16157), .ZN(n16222) );
  OAI22_X1 U19316 ( .A1(n16159), .A2(n20094), .B1(n16168), .B2(n16158), .ZN(
        n16160) );
  AOI211_X1 U19317 ( .C1(n16222), .C2(n20099), .A(n20232), .B(n16160), .ZN(
        n16161) );
  OAI211_X1 U19318 ( .C1(n16164), .C2(n16163), .A(n16162), .B(n16161), .ZN(
        P1_U2828) );
  INV_X1 U19319 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20955) );
  NAND2_X1 U19320 ( .A1(n16166), .A2(n16165), .ZN(n16186) );
  AOI21_X1 U19321 ( .B1(n20128), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20232), .ZN(n16171) );
  OAI22_X1 U19322 ( .A1(n16324), .A2(n16168), .B1(n20095), .B2(n16167), .ZN(
        n16169) );
  INV_X1 U19323 ( .A(n16169), .ZN(n16170) );
  OAI211_X1 U19324 ( .C1(n16234), .C2(n16178), .A(n16171), .B(n16170), .ZN(
        n16172) );
  AOI21_X1 U19325 ( .B1(n20099), .B2(n16231), .A(n16172), .ZN(n16173) );
  OAI221_X1 U19326 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16174), .C1(n20955), 
        .C2(n16186), .A(n16173), .ZN(P1_U2829) );
  NAND3_X1 U19327 ( .A1(n20080), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n20106), 
        .ZN(n16187) );
  NAND2_X1 U19328 ( .A1(n20133), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n16176) );
  AOI21_X1 U19329 ( .B1(n20128), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20232), .ZN(n16175) );
  OAI211_X1 U19330 ( .C1(n16178), .C2(n16177), .A(n16176), .B(n16175), .ZN(
        n16179) );
  AOI21_X1 U19331 ( .B1(n16180), .B2(n20127), .A(n16179), .ZN(n16181) );
  OAI21_X1 U19332 ( .B1(n16183), .B2(n16182), .A(n16181), .ZN(n16184) );
  INV_X1 U19333 ( .A(n16184), .ZN(n16185) );
  OAI221_X1 U19334 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n16187), .C1(n14909), 
        .C2(n16186), .A(n16185), .ZN(P1_U2830) );
  AOI22_X1 U19335 ( .A1(n16193), .A2(n20149), .B1(n20148), .B2(n16279), .ZN(
        n16188) );
  OAI21_X1 U19336 ( .B1(n20153), .B2(n16189), .A(n16188), .ZN(P1_U2850) );
  AOI22_X1 U19337 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16195) );
  NAND2_X1 U19338 ( .A1(n16191), .A2(n16190), .ZN(n16192) );
  XNOR2_X1 U19339 ( .A(n16192), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16277) );
  AOI22_X1 U19340 ( .A1(n16193), .A2(n13942), .B1(n20230), .B2(n16277), .ZN(
        n16194) );
  OAI211_X1 U19341 ( .C1(n20219), .C2(n16196), .A(n16195), .B(n16194), .ZN(
        P1_U2977) );
  AOI22_X1 U19342 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n16200) );
  AOI22_X1 U19343 ( .A1(n16198), .A2(n13942), .B1(n16252), .B2(n16197), .ZN(
        n16199) );
  OAI211_X1 U19344 ( .C1(n16201), .C2(n20220), .A(n16200), .B(n16199), .ZN(
        P1_U2978) );
  AOI22_X1 U19345 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n16205) );
  AOI22_X1 U19346 ( .A1(n16203), .A2(n13942), .B1(n20230), .B2(n16202), .ZN(
        n16204) );
  OAI211_X1 U19347 ( .C1(n20219), .C2(n16206), .A(n16205), .B(n16204), .ZN(
        P1_U2979) );
  AOI22_X1 U19348 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16210) );
  AOI22_X1 U19349 ( .A1(n16208), .A2(n20230), .B1(n13942), .B2(n16207), .ZN(
        n16209) );
  OAI211_X1 U19350 ( .C1(n20219), .C2(n16211), .A(n16210), .B(n16209), .ZN(
        P1_U2983) );
  INV_X1 U19351 ( .A(n16212), .ZN(n16213) );
  AOI21_X1 U19352 ( .B1(n16215), .B2(n16214), .A(n16213), .ZN(n16217) );
  XNOR2_X1 U19353 ( .A(n12088), .B(n16317), .ZN(n16216) );
  XNOR2_X1 U19354 ( .A(n16217), .B(n16216), .ZN(n16321) );
  AOI22_X1 U19355 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16221) );
  AOI22_X1 U19356 ( .A1(n16219), .A2(n13942), .B1(n16252), .B2(n16218), .ZN(
        n16220) );
  OAI211_X1 U19357 ( .C1(n16321), .C2(n20220), .A(n16221), .B(n16220), .ZN(
        P1_U2985) );
  AOI22_X1 U19358 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16225) );
  AOI22_X1 U19359 ( .A1(n16252), .A2(n16223), .B1(n13942), .B2(n16222), .ZN(
        n16224) );
  OAI211_X1 U19360 ( .C1(n16226), .C2(n20220), .A(n16225), .B(n16224), .ZN(
        P1_U2987) );
  AOI22_X1 U19361 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16233) );
  NAND3_X1 U19362 ( .A1(n16227), .A2(n12088), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16229) );
  NAND2_X1 U19363 ( .A1(n16229), .A2(n16228), .ZN(n16230) );
  XOR2_X1 U19364 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16230), .Z(
        n16326) );
  AOI22_X1 U19365 ( .A1(n20230), .A2(n16326), .B1(n13942), .B2(n16231), .ZN(
        n16232) );
  OAI211_X1 U19366 ( .C1(n20219), .C2(n16234), .A(n16233), .B(n16232), .ZN(
        P1_U2988) );
  AOI22_X1 U19367 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16240) );
  XNOR2_X1 U19368 ( .A(n16236), .B(n16235), .ZN(n16237) );
  XNOR2_X1 U19369 ( .A(n16238), .B(n16237), .ZN(n16354) );
  AOI22_X1 U19370 ( .A1(n16354), .A2(n20230), .B1(n13942), .B2(n20150), .ZN(
        n16239) );
  OAI211_X1 U19371 ( .C1(n20219), .C2(n20089), .A(n16240), .B(n16239), .ZN(
        P1_U2992) );
  AOI22_X1 U19372 ( .A1(n20228), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20232), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16247) );
  NAND2_X1 U19373 ( .A1(n16242), .A2(n16241), .ZN(n16243) );
  XNOR2_X1 U19374 ( .A(n16244), .B(n16243), .ZN(n16359) );
  AOI22_X1 U19375 ( .A1(n16359), .A2(n20230), .B1(n13942), .B2(n16245), .ZN(
        n16246) );
  OAI211_X1 U19376 ( .C1(n20219), .C2(n16248), .A(n16247), .B(n16246), .ZN(
        P1_U2993) );
  XNOR2_X1 U19377 ( .A(n16250), .B(n16249), .ZN(n16371) );
  INV_X1 U19378 ( .A(n16371), .ZN(n16253) );
  INV_X1 U19379 ( .A(n16251), .ZN(n20108) );
  AOI222_X1 U19380 ( .A1(n16253), .A2(n20230), .B1(n13942), .B2(n20108), .C1(
        n20105), .C2(n16252), .ZN(n16255) );
  NOR2_X1 U19381 ( .A1(n20100), .A2(n20946), .ZN(n16366) );
  INV_X1 U19382 ( .A(n16366), .ZN(n16254) );
  OAI211_X1 U19383 ( .C1(n16257), .C2(n16256), .A(n16255), .B(n16254), .ZN(
        P1_U2994) );
  INV_X1 U19384 ( .A(n16258), .ZN(n16260) );
  INV_X1 U19385 ( .A(n16261), .ZN(n16265) );
  NOR2_X1 U19386 ( .A1(n20100), .A2(n16262), .ZN(n16263) );
  AOI221_X1 U19387 ( .B1(n16266), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n16265), .C2(n16264), .A(n16263), .ZN(n16267) );
  NAND2_X1 U19388 ( .A1(n16268), .A2(n16267), .ZN(P1_U3004) );
  INV_X1 U19389 ( .A(n16269), .ZN(n16270) );
  AOI22_X1 U19390 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n20232), .B1(n16270), 
        .B2(n14845), .ZN(n16275) );
  INV_X1 U19391 ( .A(n16271), .ZN(n16273) );
  AOI22_X1 U19392 ( .A1(n16273), .A2(n16360), .B1(n16367), .B2(n16272), .ZN(
        n16274) );
  OAI211_X1 U19393 ( .C1(n16276), .C2(n14845), .A(n16275), .B(n16274), .ZN(
        P1_U3008) );
  AOI22_X1 U19394 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16278), .B1(
        n16360), .B2(n16277), .ZN(n16285) );
  NAND2_X1 U19395 ( .A1(n20232), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n16284) );
  NAND2_X1 U19396 ( .A1(n16279), .A2(n16367), .ZN(n16283) );
  OAI211_X1 U19397 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16281), .B(n16280), .ZN(
        n16282) );
  NAND4_X1 U19398 ( .A1(n16285), .A2(n16284), .A3(n16283), .A4(n16282), .ZN(
        P1_U3009) );
  INV_X1 U19399 ( .A(n16286), .ZN(n16288) );
  AOI22_X1 U19400 ( .A1(n16288), .A2(n16360), .B1(n16367), .B2(n16287), .ZN(
        n16295) );
  INV_X1 U19401 ( .A(n16289), .ZN(n16293) );
  NOR2_X1 U19402 ( .A1(n20100), .A2(n20966), .ZN(n16290) );
  AOI221_X1 U19403 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16293), 
        .C1(n16292), .C2(n16291), .A(n16290), .ZN(n16294) );
  NAND2_X1 U19404 ( .A1(n16295), .A2(n16294), .ZN(P1_U3012) );
  AOI21_X1 U19405 ( .B1(n16340), .B2(n16296), .A(n16315), .ZN(n16311) );
  INV_X1 U19406 ( .A(n16304), .ZN(n16297) );
  NOR3_X1 U19407 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16297), .A3(
        n16296), .ZN(n16301) );
  OAI22_X1 U19408 ( .A1(n16299), .A2(n16370), .B1(n16341), .B2(n16298), .ZN(
        n16300) );
  AOI211_X1 U19409 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n20232), .A(n16301), 
        .B(n16300), .ZN(n16302) );
  OAI21_X1 U19410 ( .B1(n16311), .B2(n21294), .A(n16302), .ZN(P1_U3013) );
  NOR3_X1 U19411 ( .A1(n16317), .A2(n12102), .A3(n16303), .ZN(n16305) );
  AOI21_X1 U19412 ( .B1(n16305), .B2(n16304), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16310) );
  AOI22_X1 U19413 ( .A1(n16307), .A2(n16360), .B1(n16367), .B2(n16306), .ZN(
        n16309) );
  NAND2_X1 U19414 ( .A1(n20232), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16308) );
  OAI211_X1 U19415 ( .C1(n16311), .C2(n16310), .A(n16309), .B(n16308), .ZN(
        P1_U3014) );
  OAI22_X1 U19416 ( .A1(n16313), .A2(n16341), .B1(n16312), .B2(n20100), .ZN(
        n16314) );
  AOI21_X1 U19417 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16315), .A(
        n16314), .ZN(n16320) );
  NAND4_X1 U19418 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16318), .A3(
        n16317), .A4(n16316), .ZN(n16319) );
  OAI211_X1 U19419 ( .C1(n16321), .C2(n16370), .A(n16320), .B(n16319), .ZN(
        P1_U3017) );
  NAND2_X1 U19420 ( .A1(n16323), .A2(n16322), .ZN(n16330) );
  OAI22_X1 U19421 ( .A1(n16324), .A2(n16341), .B1(n20100), .B2(n20955), .ZN(
        n16325) );
  INV_X1 U19422 ( .A(n16325), .ZN(n16329) );
  AOI22_X1 U19423 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16327), .B1(
        n16360), .B2(n16326), .ZN(n16328) );
  OAI211_X1 U19424 ( .C1(n16331), .C2(n16330), .A(n16329), .B(n16328), .ZN(
        P1_U3020) );
  NAND2_X1 U19425 ( .A1(n16332), .A2(n12046), .ZN(n16375) );
  NOR2_X1 U19426 ( .A1(n16334), .A2(n16333), .ZN(n16336) );
  AOI211_X1 U19427 ( .C1(n16338), .C2(n16337), .A(n16336), .B(n16335), .ZN(
        n16365) );
  OAI21_X1 U19428 ( .B1(n16339), .B2(n16375), .A(n16365), .ZN(n16361) );
  AOI21_X1 U19429 ( .B1(n16345), .B2(n16340), .A(n16361), .ZN(n16357) );
  INV_X1 U19430 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16348) );
  OAI22_X1 U19431 ( .A1(n16342), .A2(n16341), .B1(n20951), .B2(n20100), .ZN(
        n16343) );
  AOI21_X1 U19432 ( .B1(n16344), .B2(n16360), .A(n16343), .ZN(n16347) );
  NOR2_X1 U19433 ( .A1(n16345), .A2(n16364), .ZN(n16353) );
  OAI221_X1 U19434 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16348), .C2(n16235), .A(
        n16353), .ZN(n16346) );
  OAI211_X1 U19435 ( .C1(n16357), .C2(n16348), .A(n16347), .B(n16346), .ZN(
        P1_U3023) );
  NOR2_X1 U19436 ( .A1(n16350), .A2(n16349), .ZN(n16351) );
  AOI22_X1 U19437 ( .A1(n9822), .A2(n16367), .B1(n20232), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16356) );
  AOI22_X1 U19438 ( .A1(n16360), .A2(n16354), .B1(n16353), .B2(n16235), .ZN(
        n16355) );
  OAI211_X1 U19439 ( .C1(n16357), .C2(n16235), .A(n16356), .B(n16355), .ZN(
        P1_U3024) );
  AOI22_X1 U19440 ( .A1(n16358), .A2(n16367), .B1(n20232), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16363) );
  AOI22_X1 U19441 ( .A1(n16361), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16360), .B2(n16359), .ZN(n16362) );
  OAI211_X1 U19442 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16364), .A(
        n16363), .B(n16362), .ZN(P1_U3025) );
  OR2_X1 U19443 ( .A1(n16365), .A2(n12046), .ZN(n16369) );
  AOI21_X1 U19444 ( .B1(n20104), .B2(n16367), .A(n16366), .ZN(n16368) );
  OAI211_X1 U19445 ( .C1(n16371), .C2(n16370), .A(n16369), .B(n16368), .ZN(
        n16372) );
  INV_X1 U19446 ( .A(n16372), .ZN(n16373) );
  OAI21_X1 U19447 ( .B1(n16375), .B2(n16374), .A(n16373), .ZN(P1_U3026) );
  NAND4_X1 U19448 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n21011), .A4(n21018), .ZN(n16376) );
  NAND2_X1 U19449 ( .A1(n16377), .A2(n16376), .ZN(n20920) );
  OAI21_X1 U19450 ( .B1(n16379), .B2(n20920), .A(n16378), .ZN(n16380) );
  OAI221_X1 U19451 ( .B1(n21014), .B2(n20726), .C1(n21014), .C2(n21018), .A(
        n16380), .ZN(n16381) );
  AOI221_X1 U19452 ( .B1(n16382), .B2(n14021), .C1(n11887), .C2(n14021), .A(
        n16381), .ZN(P1_U3162) );
  NOR2_X1 U19453 ( .A1(n16382), .A2(n11887), .ZN(n16384) );
  OAI22_X1 U19454 ( .A1(n20726), .A2(n16384), .B1(n16383), .B2(n11887), .ZN(
        P1_U3466) );
  AOI211_X1 U19455 ( .C1(n16387), .C2(n16386), .A(n16385), .B(n19928), .ZN(
        n16397) );
  INV_X1 U19456 ( .A(n16388), .ZN(n16389) );
  NAND2_X1 U19457 ( .A1(n16389), .A2(n19273), .ZN(n16394) );
  INV_X1 U19458 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16391) );
  OAI22_X1 U19459 ( .A1(n19252), .A2(n16391), .B1(n19250), .B2(n16390), .ZN(
        n16392) );
  AOI21_X1 U19460 ( .B1(n19265), .B2(P2_REIP_REG_26__SCAN_IN), .A(n16392), 
        .ZN(n16393) );
  OAI211_X1 U19461 ( .C1(n19270), .C2(n16395), .A(n16394), .B(n16393), .ZN(
        n16396) );
  AOI211_X1 U19462 ( .C1(n19266), .C2(n16398), .A(n16397), .B(n16396), .ZN(
        n16399) );
  INV_X1 U19463 ( .A(n16399), .ZN(P2_U2829) );
  AOI22_X1 U19464 ( .A1(n16400), .A2(n19273), .B1(n19266), .B2(n10118), .ZN(
        n16409) );
  AOI211_X1 U19465 ( .C1(n16403), .C2(n16402), .A(n16401), .B(n19928), .ZN(
        n16407) );
  AOI22_X1 U19466 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19279), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19265), .ZN(n16404) );
  OAI21_X1 U19467 ( .B1(n16405), .B2(n19270), .A(n16404), .ZN(n16406) );
  AOI211_X1 U19468 ( .C1(n19264), .C2(P2_EBX_REG_24__SCAN_IN), .A(n16407), .B(
        n16406), .ZN(n16408) );
  NAND2_X1 U19469 ( .A1(n16409), .A2(n16408), .ZN(P2_U2831) );
  AOI22_X1 U19470 ( .A1(n19289), .A2(n16410), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19338), .ZN(n16416) );
  AOI22_X1 U19471 ( .A1(n19291), .A2(BUF1_REG_20__SCAN_IN), .B1(n19290), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16415) );
  INV_X1 U19472 ( .A(n16411), .ZN(n16412) );
  AOI22_X1 U19473 ( .A1(n16413), .A2(n19343), .B1(n19339), .B2(n16412), .ZN(
        n16414) );
  NAND3_X1 U19474 ( .A1(n16416), .A2(n16415), .A3(n16414), .ZN(P2_U2899) );
  AOI22_X1 U19475 ( .A1(n19289), .A2(n16417), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19338), .ZN(n16421) );
  AOI22_X1 U19476 ( .A1(n19291), .A2(BUF1_REG_18__SCAN_IN), .B1(n19290), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16420) );
  AOI22_X1 U19477 ( .A1(n16418), .A2(n19343), .B1(n19339), .B2(n19100), .ZN(
        n16419) );
  NAND3_X1 U19478 ( .A1(n16421), .A2(n16420), .A3(n16419), .ZN(P2_U2901) );
  AOI22_X1 U19479 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19399), .B1(n19398), 
        .B2(n16422), .ZN(n16427) );
  OAI22_X1 U19480 ( .A1(n16424), .A2(n16435), .B1(n16436), .B2(n16423), .ZN(
        n16425) );
  AOI21_X1 U19481 ( .B1(n19403), .B2(n19136), .A(n16425), .ZN(n16426) );
  OAI211_X1 U19482 ( .C1(n16428), .C2(n21179), .A(n16427), .B(n16426), .ZN(
        P2_U2999) );
  AOI22_X1 U19483 ( .A1(n16442), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19399), .ZN(n16433) );
  AOI222_X1 U19484 ( .A1(n16431), .A2(n19400), .B1(n19403), .B2(n16430), .C1(
        n19404), .C2(n16429), .ZN(n16432) );
  OAI211_X1 U19485 ( .C1(n16455), .C2(n19186), .A(n16433), .B(n16432), .ZN(
        P2_U3004) );
  AOI22_X1 U19486 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19399), .B1(n19398), 
        .B2(n19203), .ZN(n16441) );
  OAI22_X1 U19487 ( .A1(n16437), .A2(n16436), .B1(n16435), .B2(n16434), .ZN(
        n16438) );
  AOI21_X1 U19488 ( .B1(n19403), .B2(n16439), .A(n16438), .ZN(n16440) );
  OAI211_X1 U19489 ( .C1(n19409), .C2(n19209), .A(n16441), .B(n16440), .ZN(
        P2_U3005) );
  AOI22_X1 U19490 ( .A1(n16442), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19399), .ZN(n16453) );
  XOR2_X1 U19491 ( .A(n16443), .B(n16444), .Z(n16462) );
  NAND2_X1 U19492 ( .A1(n16446), .A2(n16445), .ZN(n16451) );
  INV_X1 U19493 ( .A(n16447), .ZN(n16449) );
  NOR2_X1 U19494 ( .A1(n16449), .A2(n16448), .ZN(n16450) );
  XNOR2_X1 U19495 ( .A(n16451), .B(n16450), .ZN(n16459) );
  AOI222_X1 U19496 ( .A1(n16462), .A2(n19404), .B1(n19403), .B2(n16460), .C1(
        n19400), .C2(n16459), .ZN(n16452) );
  OAI211_X1 U19497 ( .C1(n16455), .C2(n16454), .A(n16453), .B(n16452), .ZN(
        P2_U3006) );
  OAI221_X1 U19498 ( .B1(n16463), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n16463), .C2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n16456), .ZN(
        n16458) );
  AOI22_X1 U19499 ( .A1(n16458), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16457), .B2(n19316), .ZN(n16468) );
  AOI222_X1 U19500 ( .A1(n16462), .A2(n16461), .B1(n16479), .B2(n16460), .C1(
        n16471), .C2(n16459), .ZN(n16467) );
  NAND2_X1 U19501 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19399), .ZN(n16466) );
  OR4_X1 U19502 ( .A1(n16464), .A2(n10677), .A3(n16463), .A4(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16465) );
  NAND4_X1 U19503 ( .A1(n16468), .A2(n16467), .A3(n16466), .A4(n16465), .ZN(
        P2_U3038) );
  INV_X1 U19504 ( .A(n16469), .ZN(n16472) );
  AOI22_X1 U19505 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16472), .B1(
        n16471), .B2(n16470), .ZN(n16481) );
  INV_X1 U19506 ( .A(n19267), .ZN(n16473) );
  OAI22_X1 U19507 ( .A1(n16476), .A2(n16475), .B1(n16474), .B2(n16473), .ZN(
        n16477) );
  AOI211_X1 U19508 ( .C1(n16479), .C2(n11289), .A(n16478), .B(n16477), .ZN(
        n16480) );
  OAI211_X1 U19509 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16482), .A(
        n16481), .B(n16480), .ZN(P2_U3046) );
  MUX2_X1 U19510 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16491), .S(
        n16486), .Z(n16494) );
  INV_X1 U19511 ( .A(n16494), .ZN(n16512) );
  MUX2_X1 U19512 ( .A(n16484), .B(n16483), .S(n16486), .Z(n16511) );
  INV_X1 U19513 ( .A(n16485), .ZN(n16488) );
  INV_X1 U19514 ( .A(n16486), .ZN(n16508) );
  AOI21_X1 U19515 ( .B1(n16488), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16508), .ZN(n16490) );
  OAI211_X1 U19516 ( .C1(n16488), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16487), .ZN(n16489) );
  OAI211_X1 U19517 ( .C1(n16491), .C2(n20017), .A(n16490), .B(n16489), .ZN(
        n16492) );
  NAND2_X1 U19518 ( .A1(n20017), .A2(n20024), .ZN(n19504) );
  AOI222_X1 U19519 ( .A1(n16511), .A2(n16492), .B1(n16511), .B2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C1(n16492), .C2(n19504), .ZN(
        n16495) );
  OAI221_X1 U19520 ( .B1(n16495), .B2(n16494), .C1(n16495), .C2(n20017), .A(
        n16493), .ZN(n16510) );
  OAI21_X1 U19521 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16496), .ZN(n16500) );
  INV_X1 U19522 ( .A(n16497), .ZN(n16499) );
  NAND3_X1 U19523 ( .A1(n16500), .A2(n16499), .A3(n16498), .ZN(n16507) );
  INV_X1 U19524 ( .A(n16501), .ZN(n16506) );
  AOI22_X1 U19525 ( .A1(n16506), .A2(n16503), .B1(n10997), .B2(n16502), .ZN(
        n16504) );
  OAI21_X1 U19526 ( .B1(n16506), .B2(n16505), .A(n16504), .ZN(n20043) );
  AOI211_X1 U19527 ( .C1(n16508), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16507), .B(n20043), .ZN(n16509) );
  OAI211_X1 U19528 ( .C1(n16512), .C2(n16511), .A(n16510), .B(n16509), .ZN(
        n16520) );
  AOI211_X1 U19529 ( .C1(n19927), .C2(n16520), .A(n16514), .B(n16513), .ZN(
        n16525) );
  AOI21_X1 U19530 ( .B1(n16515), .B2(n16517), .A(n16516), .ZN(n16521) );
  AOI22_X1 U19531 ( .A1(n16519), .A2(n16518), .B1(n19942), .B2(n16521), .ZN(
        n16523) );
  OAI21_X1 U19532 ( .B1(n16520), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16522) );
  NAND2_X1 U19533 ( .A1(n16522), .A2(n16521), .ZN(n19926) );
  NAND2_X1 U19534 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19926), .ZN(n16528) );
  OAI21_X1 U19535 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16523), .A(n16528), 
        .ZN(n16524) );
  OAI211_X1 U19536 ( .C1(n20045), .C2(n16526), .A(n16525), .B(n16524), .ZN(
        P2_U3176) );
  AOI21_X1 U19537 ( .B1(n16528), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16527), 
        .ZN(n16529) );
  INV_X1 U19538 ( .A(n16529), .ZN(P2_U3593) );
  INV_X1 U19539 ( .A(n16530), .ZN(n16531) );
  AOI22_X1 U19540 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16532), .B1(
        n9836), .B2(n16531), .ZN(n16547) );
  INV_X1 U19541 ( .A(n16533), .ZN(n16535) );
  INV_X1 U19542 ( .A(n18063), .ZN(n17699) );
  NAND2_X1 U19543 ( .A1(n16535), .A2(n17699), .ZN(n16567) );
  AOI211_X1 U19544 ( .C1(n16537), .C2(n16567), .A(n16534), .B(n17887), .ZN(
        n16539) );
  NAND2_X1 U19545 ( .A1(n17700), .A2(n16535), .ZN(n16569) );
  AOI211_X1 U19546 ( .C1(n16537), .C2(n16569), .A(n16536), .B(n18058), .ZN(
        n16538) );
  AOI211_X1 U19547 ( .C1(n17953), .C2(n16540), .A(n16539), .B(n16538), .ZN(
        n16546) );
  OAI21_X1 U19548 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16703), .A(
        n16541), .ZN(n16542) );
  INV_X1 U19549 ( .A(n16542), .ZN(n16736) );
  OAI21_X1 U19550 ( .B1(n16543), .B2(n17914), .A(n16736), .ZN(n16544) );
  NAND4_X1 U19551 ( .A1(n16547), .A2(n16546), .A3(n16545), .A4(n16544), .ZN(
        P3_U2801) );
  NAND2_X1 U19552 ( .A1(n18338), .A2(n18270), .ZN(n18344) );
  OAI21_X1 U19553 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18344), .A(
        n16548), .ZN(n16554) );
  NAND2_X1 U19554 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18993), .ZN(
        n16550) );
  NOR4_X1 U19555 ( .A1(n16551), .A2(n16550), .A3(n18359), .A4(n16549), .ZN(
        n16552) );
  AOI211_X1 U19556 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16554), .A(
        n16553), .B(n16552), .ZN(n16558) );
  INV_X1 U19557 ( .A(n18210), .ZN(n18275) );
  AOI22_X1 U19558 ( .A1(n16556), .A2(n18275), .B1(n16555), .B2(n18263), .ZN(
        n16557) );
  OAI211_X1 U19559 ( .C1(n16559), .C2(n18317), .A(n16558), .B(n16557), .ZN(
        P3_U2831) );
  AOI21_X1 U19560 ( .B1(n17958), .B2(n16560), .A(n16561), .ZN(n17704) );
  INV_X1 U19561 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17701) );
  AOI22_X1 U19562 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17847), .B1(
        n17958), .B2(n17701), .ZN(n17703) );
  NOR2_X1 U19563 ( .A1(n18814), .A2(n18359), .ZN(n18357) );
  NOR3_X1 U19564 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17847), .A3(
        n18351), .ZN(n16562) );
  AOI21_X1 U19565 ( .B1(n18263), .B2(n16561), .A(n16562), .ZN(n16576) );
  AOI22_X1 U19566 ( .A1(n18808), .A2(n17869), .B1(n16563), .B2(n18191), .ZN(
        n18164) );
  NAND2_X1 U19567 ( .A1(n18338), .A2(n18121), .ZN(n18130) );
  NOR2_X1 U19568 ( .A1(n16565), .A2(n18130), .ZN(n18066) );
  NOR2_X1 U19569 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18059), .ZN(
        n17708) );
  AOI22_X1 U19570 ( .A1(n18348), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n18066), 
        .B2(n17708), .ZN(n16575) );
  INV_X1 U19571 ( .A(n16567), .ZN(n16571) );
  AOI211_X1 U19572 ( .C1(n18808), .C2(n16569), .A(n18291), .B(n16568), .ZN(
        n16570) );
  OAI21_X1 U19573 ( .B1(n16571), .B2(n18239), .A(n16570), .ZN(n16572) );
  OAI211_X1 U19574 ( .C1(n16573), .C2(n16572), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18358), .ZN(n16574) );
  OAI211_X1 U19575 ( .C1(n16577), .C2(n16576), .A(n16574), .B(n16575), .ZN(
        P3_U2834) );
  NOR3_X1 U19576 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n16579) );
  NOR4_X1 U19577 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16578) );
  NAND4_X1 U19578 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16579), .A3(n16578), .A4(
        U215), .ZN(U213) );
  INV_X1 U19579 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19349) );
  INV_X2 U19580 ( .A(U214), .ZN(n16630) );
  NOR2_X2 U19581 ( .A1(n16630), .A2(n16580), .ZN(n16627) );
  INV_X1 U19582 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16666) );
  OAI222_X1 U19583 ( .A1(U212), .A2(n19349), .B1(n16632), .B2(n16581), .C1(
        U214), .C2(n16666), .ZN(U216) );
  AOI222_X1 U19584 ( .A1(n16629), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16627), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16630), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n16582) );
  INV_X1 U19585 ( .A(n16582), .ZN(U217) );
  INV_X1 U19586 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16584) );
  AOI22_X1 U19587 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16629), .ZN(n16583) );
  OAI21_X1 U19588 ( .B1(n16584), .B2(n16632), .A(n16583), .ZN(U218) );
  INV_X1 U19589 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16586) );
  AOI22_X1 U19590 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16629), .ZN(n16585) );
  OAI21_X1 U19591 ( .B1(n16586), .B2(n16632), .A(n16585), .ZN(U219) );
  INV_X1 U19592 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16588) );
  AOI22_X1 U19593 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16629), .ZN(n16587) );
  OAI21_X1 U19594 ( .B1(n16588), .B2(n16632), .A(n16587), .ZN(U220) );
  AOI22_X1 U19595 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16629), .ZN(n16589) );
  OAI21_X1 U19596 ( .B1(n16590), .B2(n16632), .A(n16589), .ZN(U221) );
  INV_X1 U19597 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16592) );
  AOI22_X1 U19598 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16629), .ZN(n16591) );
  OAI21_X1 U19599 ( .B1(n16592), .B2(n16632), .A(n16591), .ZN(U222) );
  AOI222_X1 U19600 ( .A1(n16629), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(n16627), 
        .B2(BUF1_REG_24__SCAN_IN), .C1(n16630), .C2(P1_DATAO_REG_24__SCAN_IN), 
        .ZN(n16593) );
  INV_X1 U19601 ( .A(n16593), .ZN(U223) );
  AOI22_X1 U19602 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16629), .ZN(n16594) );
  OAI21_X1 U19603 ( .B1(n15286), .B2(n16632), .A(n16594), .ZN(U224) );
  AOI22_X1 U19604 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16629), .ZN(n16595) );
  OAI21_X1 U19605 ( .B1(n14505), .B2(n16632), .A(n16595), .ZN(U225) );
  AOI22_X1 U19606 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16629), .ZN(n16596) );
  OAI21_X1 U19607 ( .B1(n14490), .B2(n16632), .A(n16596), .ZN(U226) );
  AOI22_X1 U19608 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16629), .ZN(n16597) );
  OAI21_X1 U19609 ( .B1(n16598), .B2(n16632), .A(n16597), .ZN(U227) );
  AOI22_X1 U19610 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16629), .ZN(n16599) );
  OAI21_X1 U19611 ( .B1(n14336), .B2(n16632), .A(n16599), .ZN(U228) );
  INV_X1 U19612 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16601) );
  AOI22_X1 U19613 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16629), .ZN(n16600) );
  OAI21_X1 U19614 ( .B1(n16601), .B2(n16632), .A(n16600), .ZN(U229) );
  INV_X1 U19615 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16603) );
  AOI22_X1 U19616 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16629), .ZN(n16602) );
  OAI21_X1 U19617 ( .B1(n16603), .B2(n16632), .A(n16602), .ZN(U230) );
  INV_X1 U19618 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n19358) );
  AOI22_X1 U19619 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16630), .ZN(n16604) );
  OAI21_X1 U19620 ( .B1(n19358), .B2(U212), .A(n16604), .ZN(U231) );
  INV_X1 U19621 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n16606) );
  AOI22_X1 U19622 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16630), .ZN(n16605) );
  OAI21_X1 U19623 ( .B1(n16606), .B2(U212), .A(n16605), .ZN(U232) );
  INV_X1 U19624 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16608) );
  AOI22_X1 U19625 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16630), .ZN(n16607) );
  OAI21_X1 U19626 ( .B1(n16608), .B2(U212), .A(n16607), .ZN(U233) );
  INV_X1 U19627 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16647) );
  AOI22_X1 U19628 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16630), .ZN(n16609) );
  OAI21_X1 U19629 ( .B1(n16647), .B2(U212), .A(n16609), .ZN(U234) );
  AOI22_X1 U19630 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16629), .ZN(n16610) );
  OAI21_X1 U19631 ( .B1(n16611), .B2(n16632), .A(n16610), .ZN(U235) );
  INV_X1 U19632 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16613) );
  AOI22_X1 U19633 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16630), .ZN(n16612) );
  OAI21_X1 U19634 ( .B1(n16613), .B2(U212), .A(n16612), .ZN(U236) );
  AOI22_X1 U19635 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16629), .ZN(n16614) );
  OAI21_X1 U19636 ( .B1(n16615), .B2(n16632), .A(n16614), .ZN(U237) );
  INV_X1 U19637 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16643) );
  AOI22_X1 U19638 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16630), .ZN(n16616) );
  OAI21_X1 U19639 ( .B1(n16643), .B2(U212), .A(n16616), .ZN(U238) );
  AOI22_X1 U19640 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16629), .ZN(n16617) );
  OAI21_X1 U19641 ( .B1(n16618), .B2(n16632), .A(n16617), .ZN(U239) );
  INV_X1 U19642 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16641) );
  AOI22_X1 U19643 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16630), .ZN(n16619) );
  OAI21_X1 U19644 ( .B1(n16641), .B2(U212), .A(n16619), .ZN(U240) );
  INV_X1 U19645 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16640) );
  AOI22_X1 U19646 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16630), .ZN(n16620) );
  OAI21_X1 U19647 ( .B1(n16640), .B2(U212), .A(n16620), .ZN(U241) );
  INV_X1 U19648 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16639) );
  AOI22_X1 U19649 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16630), .ZN(n16621) );
  OAI21_X1 U19650 ( .B1(n16639), .B2(U212), .A(n16621), .ZN(U242) );
  INV_X1 U19651 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16623) );
  AOI22_X1 U19652 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16629), .ZN(n16622) );
  OAI21_X1 U19653 ( .B1(n16623), .B2(n16632), .A(n16622), .ZN(U243) );
  INV_X1 U19654 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16637) );
  AOI22_X1 U19655 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16630), .ZN(n16624) );
  OAI21_X1 U19656 ( .B1(n16637), .B2(U212), .A(n16624), .ZN(U244) );
  INV_X1 U19657 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16626) );
  AOI22_X1 U19658 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16629), .ZN(n16625) );
  OAI21_X1 U19659 ( .B1(n16626), .B2(n16632), .A(n16625), .ZN(U245) );
  INV_X1 U19660 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16635) );
  AOI22_X1 U19661 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16627), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16630), .ZN(n16628) );
  OAI21_X1 U19662 ( .B1(n16635), .B2(U212), .A(n16628), .ZN(U246) );
  INV_X1 U19663 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16633) );
  AOI22_X1 U19664 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16630), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16629), .ZN(n16631) );
  OAI21_X1 U19665 ( .B1(n16633), .B2(n16632), .A(n16631), .ZN(U247) );
  OAI22_X1 U19666 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16664), .ZN(n16634) );
  INV_X1 U19667 ( .A(n16634), .ZN(U251) );
  INV_X1 U19668 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18382) );
  AOI22_X1 U19669 ( .A1(n16664), .A2(n16635), .B1(n18382), .B2(U215), .ZN(U252) );
  OAI22_X1 U19670 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16653), .ZN(n16636) );
  INV_X1 U19671 ( .A(n16636), .ZN(U253) );
  INV_X1 U19672 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18390) );
  AOI22_X1 U19673 ( .A1(n16664), .A2(n16637), .B1(n18390), .B2(U215), .ZN(U254) );
  OAI22_X1 U19674 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16653), .ZN(n16638) );
  INV_X1 U19675 ( .A(n16638), .ZN(U255) );
  INV_X1 U19676 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18400) );
  AOI22_X1 U19677 ( .A1(n16664), .A2(n16639), .B1(n18400), .B2(U215), .ZN(U256) );
  INV_X1 U19678 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18403) );
  AOI22_X1 U19679 ( .A1(n16664), .A2(n16640), .B1(n18403), .B2(U215), .ZN(U257) );
  INV_X1 U19680 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18407) );
  AOI22_X1 U19681 ( .A1(n16664), .A2(n16641), .B1(n18407), .B2(U215), .ZN(U258) );
  OAI22_X1 U19682 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16653), .ZN(n16642) );
  INV_X1 U19683 ( .A(n16642), .ZN(U259) );
  INV_X1 U19684 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17677) );
  AOI22_X1 U19685 ( .A1(n16664), .A2(n16643), .B1(n17677), .B2(U215), .ZN(U260) );
  OAI22_X1 U19686 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16653), .ZN(n16644) );
  INV_X1 U19687 ( .A(n16644), .ZN(U261) );
  OAI22_X1 U19688 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16653), .ZN(n16645) );
  INV_X1 U19689 ( .A(n16645), .ZN(U262) );
  OAI22_X1 U19690 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16653), .ZN(n16646) );
  INV_X1 U19691 ( .A(n16646), .ZN(U263) );
  INV_X1 U19692 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17687) );
  AOI22_X1 U19693 ( .A1(n16664), .A2(n16647), .B1(n17687), .B2(U215), .ZN(U264) );
  OAI22_X1 U19694 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16653), .ZN(n16648) );
  INV_X1 U19695 ( .A(n16648), .ZN(U265) );
  OAI22_X1 U19696 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16664), .ZN(n16649) );
  INV_X1 U19697 ( .A(n16649), .ZN(U266) );
  INV_X1 U19698 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18371) );
  AOI22_X1 U19699 ( .A1(n16664), .A2(n19358), .B1(n18371), .B2(U215), .ZN(U267) );
  OAI22_X1 U19700 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16653), .ZN(n16650) );
  INV_X1 U19701 ( .A(n16650), .ZN(U268) );
  OAI22_X1 U19702 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16664), .ZN(n16651) );
  INV_X1 U19703 ( .A(n16651), .ZN(U269) );
  OAI22_X1 U19704 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16653), .ZN(n16652) );
  INV_X1 U19705 ( .A(n16652), .ZN(U270) );
  OAI22_X1 U19706 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16653), .ZN(n16654) );
  INV_X1 U19707 ( .A(n16654), .ZN(U271) );
  OAI22_X1 U19708 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16664), .ZN(n16655) );
  INV_X1 U19709 ( .A(n16655), .ZN(U272) );
  OAI22_X1 U19710 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16664), .ZN(n16656) );
  INV_X1 U19711 ( .A(n16656), .ZN(U273) );
  OAI22_X1 U19712 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16664), .ZN(n16657) );
  INV_X1 U19713 ( .A(n16657), .ZN(U274) );
  OAI22_X1 U19714 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16664), .ZN(n16658) );
  INV_X1 U19715 ( .A(n16658), .ZN(U275) );
  OAI22_X1 U19716 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16664), .ZN(n16659) );
  INV_X1 U19717 ( .A(n16659), .ZN(U276) );
  OAI22_X1 U19718 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16664), .ZN(n16660) );
  INV_X1 U19719 ( .A(n16660), .ZN(U277) );
  OAI22_X1 U19720 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16664), .ZN(n16661) );
  INV_X1 U19721 ( .A(n16661), .ZN(U278) );
  OAI22_X1 U19722 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16664), .ZN(n16662) );
  INV_X1 U19723 ( .A(n16662), .ZN(U279) );
  OAI22_X1 U19724 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16664), .ZN(n16663) );
  INV_X1 U19725 ( .A(n16663), .ZN(U280) );
  INV_X1 U19726 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19352) );
  INV_X1 U19727 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n21126) );
  AOI22_X1 U19728 ( .A1(n16664), .A2(n19352), .B1(n21126), .B2(U215), .ZN(U281) );
  OAI22_X1 U19729 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n16664), .ZN(n16665) );
  INV_X1 U19730 ( .A(n16665), .ZN(U282) );
  INV_X1 U19731 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16667) );
  AOI222_X1 U19732 ( .A1(n19349), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16667), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .C1(n16666), .C2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n16668) );
  INV_X2 U19733 ( .A(n16670), .ZN(n16669) );
  INV_X1 U19734 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18930) );
  INV_X1 U19735 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19964) );
  AOI22_X1 U19736 ( .A1(n16669), .A2(n18930), .B1(n19964), .B2(n16670), .ZN(
        U347) );
  INV_X1 U19737 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18928) );
  INV_X1 U19738 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19963) );
  AOI22_X1 U19739 ( .A1(n16669), .A2(n18928), .B1(n19963), .B2(n16670), .ZN(
        U348) );
  INV_X1 U19740 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n21321) );
  INV_X1 U19741 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19961) );
  AOI22_X1 U19742 ( .A1(n16669), .A2(n21321), .B1(n19961), .B2(n16670), .ZN(
        U349) );
  INV_X1 U19743 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18926) );
  INV_X1 U19744 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19960) );
  AOI22_X1 U19745 ( .A1(n16669), .A2(n18926), .B1(n19960), .B2(n16670), .ZN(
        U350) );
  INV_X1 U19746 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18924) );
  INV_X1 U19747 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19959) );
  AOI22_X1 U19748 ( .A1(n16669), .A2(n18924), .B1(n19959), .B2(n16670), .ZN(
        U351) );
  INV_X1 U19749 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18921) );
  INV_X1 U19750 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19957) );
  AOI22_X1 U19751 ( .A1(n16669), .A2(n18921), .B1(n19957), .B2(n16670), .ZN(
        U352) );
  INV_X1 U19752 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18920) );
  INV_X1 U19753 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19956) );
  AOI22_X1 U19754 ( .A1(n16669), .A2(n18920), .B1(n19956), .B2(n16670), .ZN(
        U353) );
  INV_X1 U19755 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18918) );
  INV_X1 U19756 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19954) );
  AOI22_X1 U19757 ( .A1(n16669), .A2(n18918), .B1(n19954), .B2(n16670), .ZN(
        U354) );
  INV_X1 U19758 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18971) );
  INV_X1 U19759 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19994) );
  AOI22_X1 U19760 ( .A1(n16669), .A2(n18971), .B1(n19994), .B2(n16670), .ZN(
        U355) );
  INV_X1 U19761 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18969) );
  INV_X1 U19762 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19992) );
  AOI22_X1 U19763 ( .A1(n16669), .A2(n18969), .B1(n19992), .B2(n16670), .ZN(
        U356) );
  INV_X1 U19764 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18965) );
  INV_X1 U19765 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19990) );
  AOI22_X1 U19766 ( .A1(n16669), .A2(n18965), .B1(n19990), .B2(n16670), .ZN(
        U357) );
  INV_X1 U19767 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18963) );
  INV_X1 U19768 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n21152) );
  AOI22_X1 U19769 ( .A1(n16669), .A2(n18963), .B1(n21152), .B2(n16670), .ZN(
        U358) );
  INV_X1 U19770 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18961) );
  INV_X1 U19771 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19988) );
  AOI22_X1 U19772 ( .A1(n16669), .A2(n18961), .B1(n19988), .B2(n16670), .ZN(
        U359) );
  INV_X1 U19773 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18959) );
  INV_X1 U19774 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19987) );
  AOI22_X1 U19775 ( .A1(n16669), .A2(n18959), .B1(n19987), .B2(n16670), .ZN(
        U360) );
  INV_X1 U19776 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18957) );
  INV_X1 U19777 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19985) );
  AOI22_X1 U19778 ( .A1(n16669), .A2(n18957), .B1(n19985), .B2(n16670), .ZN(
        U361) );
  INV_X1 U19779 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18954) );
  INV_X1 U19780 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19983) );
  AOI22_X1 U19781 ( .A1(n16669), .A2(n18954), .B1(n19983), .B2(n16670), .ZN(
        U362) );
  INV_X1 U19782 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18953) );
  INV_X1 U19783 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U19784 ( .A1(n16669), .A2(n18953), .B1(n19981), .B2(n16670), .ZN(
        U363) );
  INV_X1 U19785 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18951) );
  INV_X1 U19786 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n21186) );
  AOI22_X1 U19787 ( .A1(n16669), .A2(n18951), .B1(n21186), .B2(n16670), .ZN(
        U364) );
  INV_X1 U19788 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18916) );
  INV_X1 U19789 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n21183) );
  AOI22_X1 U19790 ( .A1(n16669), .A2(n18916), .B1(n21183), .B2(n16670), .ZN(
        U365) );
  INV_X1 U19791 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18949) );
  INV_X1 U19792 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n21121) );
  AOI22_X1 U19793 ( .A1(n16669), .A2(n18949), .B1(n21121), .B2(n16670), .ZN(
        U366) );
  INV_X1 U19794 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18947) );
  INV_X1 U19795 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19977) );
  AOI22_X1 U19796 ( .A1(n16669), .A2(n18947), .B1(n19977), .B2(n16670), .ZN(
        U367) );
  INV_X1 U19797 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18945) );
  INV_X1 U19798 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19975) );
  AOI22_X1 U19799 ( .A1(n16669), .A2(n18945), .B1(n19975), .B2(n16670), .ZN(
        U368) );
  INV_X1 U19800 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18942) );
  INV_X1 U19801 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n21304) );
  AOI22_X1 U19802 ( .A1(n16669), .A2(n18942), .B1(n21304), .B2(n16670), .ZN(
        U369) );
  INV_X1 U19803 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18941) );
  INV_X1 U19804 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19973) );
  AOI22_X1 U19805 ( .A1(n16669), .A2(n18941), .B1(n19973), .B2(n16670), .ZN(
        U370) );
  INV_X1 U19806 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18939) );
  INV_X1 U19807 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19972) );
  AOI22_X1 U19808 ( .A1(n16669), .A2(n18939), .B1(n19972), .B2(n16670), .ZN(
        U371) );
  INV_X1 U19809 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18936) );
  INV_X1 U19810 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19970) );
  AOI22_X1 U19811 ( .A1(n16669), .A2(n18936), .B1(n19970), .B2(n16670), .ZN(
        U372) );
  INV_X1 U19812 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18935) );
  INV_X1 U19813 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n21157) );
  AOI22_X1 U19814 ( .A1(n16669), .A2(n18935), .B1(n21157), .B2(n16670), .ZN(
        U373) );
  INV_X1 U19815 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18933) );
  INV_X1 U19816 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19968) );
  AOI22_X1 U19817 ( .A1(n16669), .A2(n18933), .B1(n19968), .B2(n16670), .ZN(
        U374) );
  INV_X1 U19818 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18931) );
  INV_X1 U19819 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19966) );
  AOI22_X1 U19820 ( .A1(n16669), .A2(n18931), .B1(n19966), .B2(n16670), .ZN(
        U375) );
  INV_X1 U19821 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18914) );
  AOI22_X1 U19822 ( .A1(n16669), .A2(n18914), .B1(n19952), .B2(n16670), .ZN(
        U376) );
  INV_X1 U19823 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18913) );
  NAND2_X1 U19824 ( .A1(n18913), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18899) );
  INV_X1 U19825 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18903) );
  NAND2_X1 U19826 ( .A1(n18910), .A2(n18903), .ZN(n18895) );
  OAI21_X1 U19827 ( .B1(n18899), .B2(n18903), .A(n18895), .ZN(n18981) );
  AOI21_X1 U19828 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18981), .ZN(n16671) );
  INV_X1 U19829 ( .A(n16671), .ZN(P3_U2633) );
  NOR2_X1 U19830 ( .A1(n17639), .A2(n16672), .ZN(n16678) );
  OAI21_X1 U19831 ( .B1(n17640), .B2(n16678), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16673) );
  NAND2_X1 U19832 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19045), .ZN(n18882) );
  NAND2_X1 U19833 ( .A1(n16673), .A2(n18882), .ZN(P3_U2634) );
  NOR2_X1 U19834 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16675) );
  AOI22_X1 U19835 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n19042), .B1(n16675), .B2(
        n18910), .ZN(n16674) );
  OAI21_X1 U19836 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n19042), .A(n16674), 
        .ZN(P3_U2635) );
  OAI21_X1 U19837 ( .B1(n16675), .B2(BS16), .A(n18981), .ZN(n18979) );
  OAI21_X1 U19838 ( .B1(n18981), .B2(n19032), .A(n18979), .ZN(P3_U2636) );
  INV_X1 U19839 ( .A(n16676), .ZN(n16679) );
  NOR3_X1 U19840 ( .A1(n16679), .A2(n16678), .A3(n16677), .ZN(n18815) );
  NOR2_X1 U19841 ( .A1(n18815), .A2(n18883), .ZN(n19026) );
  OAI21_X1 U19842 ( .B1(n19026), .B2(n18365), .A(n16680), .ZN(P3_U2637) );
  NOR4_X1 U19843 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16684) );
  NOR4_X1 U19844 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16683) );
  NOR4_X1 U19845 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16682) );
  NOR4_X1 U19846 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16681) );
  NAND4_X1 U19847 ( .A1(n16684), .A2(n16683), .A3(n16682), .A4(n16681), .ZN(
        n16690) );
  NOR4_X1 U19848 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16688) );
  AOI211_X1 U19849 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16687) );
  NOR4_X1 U19850 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16686) );
  NOR4_X1 U19851 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16685) );
  NAND4_X1 U19852 ( .A1(n16688), .A2(n16687), .A3(n16686), .A4(n16685), .ZN(
        n16689) );
  NOR2_X1 U19853 ( .A1(n16690), .A2(n16689), .ZN(n19020) );
  INV_X1 U19854 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16692) );
  NOR3_X1 U19855 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16693) );
  OAI21_X1 U19856 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16693), .A(n19020), .ZN(
        n16691) );
  OAI21_X1 U19857 ( .B1(n19020), .B2(n16692), .A(n16691), .ZN(P3_U2638) );
  INV_X1 U19858 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19016) );
  INV_X1 U19859 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18980) );
  AOI21_X1 U19860 ( .B1(n19016), .B2(n18980), .A(n16693), .ZN(n16695) );
  INV_X1 U19861 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16694) );
  INV_X1 U19862 ( .A(n19020), .ZN(n19023) );
  AOI22_X1 U19863 ( .A1(n19020), .A2(n16695), .B1(n16694), .B2(n19023), .ZN(
        P3_U2639) );
  NOR2_X1 U19864 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19036) );
  NAND2_X1 U19865 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19036), .ZN(n18872) );
  NAND4_X1 U19866 ( .A1(n18866), .A2(n18871), .A3(n19032), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n17060) );
  NOR2_X1 U19867 ( .A1(n18348), .A2(n18885), .ZN(n16698) );
  AOI211_X1 U19868 ( .C1(n19033), .C2(n19031), .A(n18894), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16699) );
  AOI211_X4 U19869 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n17642), .A(n16699), .B(
        n16702), .ZN(n17069) );
  INV_X1 U19870 ( .A(n16699), .ZN(n18868) );
  INV_X1 U19871 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18958) );
  INV_X1 U19872 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18955) );
  INV_X1 U19873 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18950) );
  INV_X1 U19874 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18937) );
  INV_X1 U19875 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18934) );
  INV_X1 U19876 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n21241) );
  INV_X1 U19877 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18922) );
  INV_X1 U19878 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18919) );
  NAND3_X1 U19879 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17017) );
  NOR3_X1 U19880 ( .A1(n18922), .A2(n18919), .A3(n17017), .ZN(n16967) );
  NAND4_X1 U19881 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16967), .A3(
        P3_REIP_REG_7__SCAN_IN), .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n16940) );
  INV_X1 U19882 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21094) );
  INV_X1 U19883 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18929) );
  NOR2_X1 U19884 ( .A1(n21094), .A2(n18929), .ZN(n16928) );
  INV_X1 U19885 ( .A(n16928), .ZN(n16943) );
  NOR3_X1 U19886 ( .A1(n21241), .A2(n16940), .A3(n16943), .ZN(n16921) );
  NAND2_X1 U19887 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16921), .ZN(n16902) );
  NOR3_X1 U19888 ( .A1(n18937), .A2(n18934), .A3(n16902), .ZN(n16895) );
  NAND4_X1 U19889 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16895), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n16834) );
  NAND2_X1 U19890 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16843) );
  NOR2_X1 U19891 ( .A1(n16834), .A2(n16843), .ZN(n16831) );
  NAND2_X1 U19892 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16831), .ZN(n16806) );
  NOR2_X1 U19893 ( .A1(n18950), .A2(n16806), .ZN(n16805) );
  NAND2_X1 U19894 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16805), .ZN(n16796) );
  NOR2_X1 U19895 ( .A1(n18955), .A2(n16796), .ZN(n16794) );
  NAND2_X1 U19896 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16794), .ZN(n16776) );
  NOR2_X1 U19897 ( .A1(n18958), .A2(n16776), .ZN(n16764) );
  NAND2_X1 U19898 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16764), .ZN(n16715) );
  NAND4_X1 U19899 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16758), .ZN(n16717) );
  NOR3_X1 U19900 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18972), .A3(n16717), 
        .ZN(n16700) );
  AOI21_X1 U19901 ( .B1(n17069), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16700), .ZN(
        n16722) );
  NAND2_X1 U19902 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17642), .ZN(n16701) );
  AOI211_X4 U19903 ( .C1(n19032), .C2(n19034), .A(n16702), .B(n16701), .ZN(
        n17068) );
  NAND3_X1 U19904 ( .A1(n17425), .A2(n17420), .A3(n17049), .ZN(n17048) );
  INV_X1 U19905 ( .A(n17048), .ZN(n17035) );
  NAND2_X1 U19906 ( .A1(n17035), .A2(n17034), .ZN(n17033) );
  NOR2_X1 U19907 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17033), .ZN(n17012) );
  NAND2_X1 U19908 ( .A1(n17012), .A2(n17008), .ZN(n17007) );
  NOR2_X1 U19909 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17007), .ZN(n16991) );
  NAND2_X1 U19910 ( .A1(n16991), .A2(n17390), .ZN(n16988) );
  NOR2_X1 U19911 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16988), .ZN(n16961) );
  NAND2_X1 U19912 ( .A1(n16961), .A2(n17350), .ZN(n16942) );
  NAND2_X1 U19913 ( .A1(n16941), .A2(n16936), .ZN(n16935) );
  NAND2_X1 U19914 ( .A1(n16915), .A2(n16912), .ZN(n16911) );
  NAND2_X1 U19915 ( .A1(n16891), .A2(n17243), .ZN(n16884) );
  NAND2_X1 U19916 ( .A1(n16870), .A2(n21242), .ZN(n16861) );
  NOR2_X1 U19917 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16861), .ZN(n16846) );
  INV_X1 U19918 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17196) );
  NAND2_X1 U19919 ( .A1(n16846), .A2(n17196), .ZN(n16839) );
  NOR2_X1 U19920 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16839), .ZN(n16827) );
  NAND2_X1 U19921 ( .A1(n16827), .A2(n17143), .ZN(n16821) );
  NOR2_X1 U19922 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16821), .ZN(n16807) );
  INV_X1 U19923 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16800) );
  NAND2_X1 U19924 ( .A1(n16807), .A2(n16800), .ZN(n16799) );
  NOR2_X1 U19925 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16799), .ZN(n16785) );
  INV_X1 U19926 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16780) );
  NAND2_X1 U19927 ( .A1(n16785), .A2(n16780), .ZN(n16779) );
  NOR2_X1 U19928 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16779), .ZN(n16765) );
  NAND2_X1 U19929 ( .A1(n16765), .A2(n17125), .ZN(n16759) );
  NOR2_X1 U19930 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16759), .ZN(n16745) );
  INV_X1 U19931 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17121) );
  NAND2_X1 U19932 ( .A1(n16745), .A2(n17121), .ZN(n16724) );
  NOR2_X1 U19933 ( .A1(n17011), .A2(n16724), .ZN(n16731) );
  INV_X1 U19934 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17084) );
  AOI21_X1 U19935 ( .B1(n16705), .B2(n16704), .A(n16703), .ZN(n17698) );
  OAI21_X1 U19936 ( .B1(n16706), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16705), .ZN(n17717) );
  INV_X1 U19937 ( .A(n17717), .ZN(n16755) );
  AOI21_X1 U19938 ( .B1(n10020), .B2(n17695), .A(n16706), .ZN(n17730) );
  INV_X1 U19939 ( .A(n16710), .ZN(n16708) );
  INV_X1 U19940 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17751) );
  NOR2_X1 U19941 ( .A1(n16708), .A2(n17751), .ZN(n16707) );
  OAI21_X1 U19942 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16707), .A(
        n17695), .ZN(n17742) );
  INV_X1 U19943 ( .A(n17742), .ZN(n16774) );
  AOI21_X1 U19944 ( .B1(n16708), .B2(n17751), .A(n16707), .ZN(n17750) );
  INV_X1 U19945 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17767) );
  NOR2_X1 U19946 ( .A1(n21104), .A2(n17779), .ZN(n16714) );
  INV_X1 U19947 ( .A(n16714), .ZN(n16713) );
  NOR2_X1 U19948 ( .A1(n16709), .A2(n16713), .ZN(n16711) );
  INV_X1 U19949 ( .A(n16711), .ZN(n17738) );
  AOI21_X1 U19950 ( .B1(n17767), .B2(n17738), .A(n16710), .ZN(n17761) );
  NAND2_X1 U19951 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16714), .ZN(
        n16712) );
  AOI21_X1 U19952 ( .B1(n21288), .B2(n16712), .A(n16711), .ZN(n17778) );
  OAI22_X1 U19953 ( .A1(n17792), .A2(n16713), .B1(n16714), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17789) );
  INV_X1 U19954 ( .A(n17789), .ZN(n16818) );
  NOR2_X1 U19955 ( .A1(n21104), .A2(n17812), .ZN(n17811) );
  INV_X1 U19956 ( .A(n17811), .ZN(n16856) );
  NOR2_X1 U19957 ( .A1(n17814), .A2(n16856), .ZN(n17776) );
  INV_X1 U19958 ( .A(n17776), .ZN(n16835) );
  AOI21_X1 U19959 ( .B1(n10018), .B2(n16835), .A(n16714), .ZN(n17804) );
  NOR2_X1 U19960 ( .A1(n21104), .A2(n17850), .ZN(n17852) );
  NAND2_X1 U19961 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17852), .ZN(
        n16878) );
  OAI21_X1 U19962 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16878), .A(
        n17002), .ZN(n16881) );
  OAI21_X1 U19963 ( .B1(n17776), .B2(n17025), .A(n16881), .ZN(n16826) );
  NOR2_X1 U19964 ( .A1(n17804), .A2(n16826), .ZN(n16825) );
  NOR2_X1 U19965 ( .A1(n16825), .A2(n17025), .ZN(n16817) );
  NOR2_X1 U19966 ( .A1(n16818), .A2(n16817), .ZN(n16816) );
  NOR2_X1 U19967 ( .A1(n16816), .A2(n17025), .ZN(n16809) );
  NOR2_X1 U19968 ( .A1(n17750), .A2(n9774), .ZN(n16786) );
  NOR2_X1 U19969 ( .A1(n16786), .A2(n17025), .ZN(n16773) );
  NOR2_X1 U19970 ( .A1(n16755), .A2(n9776), .ZN(n16754) );
  NOR2_X1 U19971 ( .A1(n16734), .A2(n17025), .ZN(n16725) );
  NAND2_X1 U19972 ( .A1(n17002), .A2(n18885), .ZN(n17041) );
  NOR3_X1 U19973 ( .A1(n16726), .A2(n16725), .A3(n17041), .ZN(n16720) );
  NAND3_X1 U19974 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16716) );
  AND2_X1 U19975 ( .A1(n17051), .A2(n16715), .ZN(n16763) );
  NOR2_X1 U19976 ( .A1(n17058), .A2(n16763), .ZN(n16762) );
  INV_X1 U19977 ( .A(n16762), .ZN(n16769) );
  AOI21_X1 U19978 ( .B1(n17051), .B2(n16716), .A(n16769), .ZN(n16744) );
  NOR2_X1 U19979 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16717), .ZN(n16729) );
  INV_X1 U19980 ( .A(n16729), .ZN(n16718) );
  AOI21_X1 U19981 ( .B1(n16744), .B2(n16718), .A(n18970), .ZN(n16719) );
  AOI211_X1 U19982 ( .C1(n16731), .C2(n17084), .A(n16720), .B(n16719), .ZN(
        n16721) );
  OAI211_X1 U19983 ( .C1(n16723), .C2(n17059), .A(n16722), .B(n16721), .ZN(
        P3_U2640) );
  NAND2_X1 U19984 ( .A1(n17068), .A2(n16724), .ZN(n16740) );
  XOR2_X1 U19985 ( .A(n16726), .B(n16725), .Z(n16730) );
  OAI22_X1 U19986 ( .A1(n16744), .A2(n18972), .B1(n16727), .B2(n17059), .ZN(
        n16728) );
  AOI211_X1 U19987 ( .C1(n16730), .C2(n18885), .A(n16729), .B(n16728), .ZN(
        n16733) );
  OAI21_X1 U19988 ( .B1(n17069), .B2(n16731), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16732) );
  OAI211_X1 U19989 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16740), .A(n16733), .B(
        n16732), .ZN(P3_U2641) );
  INV_X1 U19990 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18968) );
  AOI211_X1 U19991 ( .C1(n16736), .C2(n16735), .A(n16734), .B(n17060), .ZN(
        n16739) );
  NAND3_X1 U19992 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16758), .ZN(n16737) );
  OAI22_X1 U19993 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16737), .B1(n10021), 
        .B2(n17059), .ZN(n16738) );
  AOI211_X1 U19994 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17069), .A(n16739), .B(
        n16738), .ZN(n16743) );
  INV_X1 U19995 ( .A(n16740), .ZN(n16741) );
  OAI21_X1 U19996 ( .B1(n16745), .B2(n17121), .A(n16741), .ZN(n16742) );
  OAI211_X1 U19997 ( .C1(n16744), .C2(n18968), .A(n16743), .B(n16742), .ZN(
        P3_U2642) );
  AOI22_X1 U19998 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17038), .B1(
        n17069), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16753) );
  AOI211_X1 U19999 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16759), .A(n16745), .B(
        n17011), .ZN(n16749) );
  AOI211_X1 U20000 ( .C1(n17698), .C2(n16747), .A(n16746), .B(n17060), .ZN(
        n16748) );
  AOI211_X1 U20001 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16769), .A(n16749), 
        .B(n16748), .ZN(n16752) );
  NAND2_X1 U20002 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16750) );
  OAI211_X1 U20003 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16758), .B(n16750), .ZN(n16751) );
  NAND3_X1 U20004 ( .A1(n16753), .A2(n16752), .A3(n16751), .ZN(P3_U2643) );
  INV_X1 U20005 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18962) );
  AOI211_X1 U20006 ( .C1(n16755), .C2(n9776), .A(n16754), .B(n17060), .ZN(
        n16757) );
  INV_X1 U20007 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17720) );
  OAI22_X1 U20008 ( .A1(n17720), .A2(n17059), .B1(n17062), .B2(n17125), .ZN(
        n16756) );
  AOI211_X1 U20009 ( .C1(n16758), .C2(n18962), .A(n16757), .B(n16756), .ZN(
        n16761) );
  OAI211_X1 U20010 ( .C1(n16765), .C2(n17125), .A(n17068), .B(n16759), .ZN(
        n16760) );
  OAI211_X1 U20011 ( .C1(n16762), .C2(n18962), .A(n16761), .B(n16760), .ZN(
        P3_U2644) );
  AOI22_X1 U20012 ( .A1(n17069), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16764), 
        .B2(n16763), .ZN(n16771) );
  AOI211_X1 U20013 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16779), .A(n16765), .B(
        n17011), .ZN(n16768) );
  AOI211_X1 U20014 ( .C1(n17730), .C2(n9820), .A(n16766), .B(n17060), .ZN(
        n16767) );
  AOI211_X1 U20015 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16769), .A(n16768), 
        .B(n16767), .ZN(n16770) );
  OAI211_X1 U20016 ( .C1(n10020), .C2(n17059), .A(n16771), .B(n16770), .ZN(
        P3_U2645) );
  INV_X1 U20017 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18956) );
  OAI21_X1 U20018 ( .B1(n16794), .B2(n17070), .A(n17073), .ZN(n16791) );
  AOI21_X1 U20019 ( .B1(n17051), .B2(n18956), .A(n16791), .ZN(n16783) );
  AOI211_X1 U20020 ( .C1(n16774), .C2(n16773), .A(n16772), .B(n17060), .ZN(
        n16778) );
  NAND2_X1 U20021 ( .A1(n17051), .A2(n18958), .ZN(n16775) );
  OAI22_X1 U20022 ( .A1(n17062), .A2(n16780), .B1(n16776), .B2(n16775), .ZN(
        n16777) );
  AOI211_X1 U20023 ( .C1(n17038), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16778), .B(n16777), .ZN(n16782) );
  OAI211_X1 U20024 ( .C1(n16785), .C2(n16780), .A(n17068), .B(n16779), .ZN(
        n16781) );
  OAI211_X1 U20025 ( .C1(n16783), .C2(n18958), .A(n16782), .B(n16781), .ZN(
        P3_U2646) );
  NOR2_X1 U20026 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17070), .ZN(n16784) );
  AOI22_X1 U20027 ( .A1(n17069), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16794), 
        .B2(n16784), .ZN(n16790) );
  AOI211_X1 U20028 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16799), .A(n16785), .B(
        n17011), .ZN(n16788) );
  AOI211_X1 U20029 ( .C1(n17750), .C2(n9774), .A(n16786), .B(n17060), .ZN(
        n16787) );
  AOI211_X1 U20030 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16791), .A(n16788), 
        .B(n16787), .ZN(n16789) );
  OAI211_X1 U20031 ( .C1(n17751), .C2(n17059), .A(n16790), .B(n16789), .ZN(
        P3_U2647) );
  INV_X1 U20032 ( .A(n16791), .ZN(n16803) );
  AOI211_X1 U20033 ( .C1(n17761), .C2(n16793), .A(n16792), .B(n17060), .ZN(
        n16798) );
  OR2_X1 U20034 ( .A1(n17070), .A2(n16794), .ZN(n16795) );
  OAI22_X1 U20035 ( .A1(n17062), .A2(n16800), .B1(n16796), .B2(n16795), .ZN(
        n16797) );
  AOI211_X1 U20036 ( .C1(n17038), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16798), .B(n16797), .ZN(n16802) );
  OAI211_X1 U20037 ( .C1(n16807), .C2(n16800), .A(n17068), .B(n16799), .ZN(
        n16801) );
  OAI211_X1 U20038 ( .C1(n16803), .C2(n18955), .A(n16802), .B(n16801), .ZN(
        P3_U2648) );
  NOR2_X1 U20039 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17070), .ZN(n16804) );
  AOI22_X1 U20040 ( .A1(n17069), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n16805), 
        .B2(n16804), .ZN(n16814) );
  AOI21_X1 U20041 ( .B1(n17051), .B2(n16806), .A(n17058), .ZN(n16815) );
  NAND4_X1 U20042 ( .A1(n17051), .A2(P3_REIP_REG_20__SCAN_IN), .A3(n16831), 
        .A4(n18950), .ZN(n16823) );
  NAND2_X1 U20043 ( .A1(n16815), .A2(n16823), .ZN(n16812) );
  AOI211_X1 U20044 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16821), .A(n16807), .B(
        n17011), .ZN(n16811) );
  AOI211_X1 U20045 ( .C1(n17778), .C2(n16809), .A(n16808), .B(n17060), .ZN(
        n16810) );
  AOI211_X1 U20046 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16812), .A(n16811), 
        .B(n16810), .ZN(n16813) );
  OAI211_X1 U20047 ( .C1(n21288), .C2(n17059), .A(n16814), .B(n16813), .ZN(
        P3_U2649) );
  INV_X1 U20048 ( .A(n16815), .ZN(n16830) );
  AOI211_X1 U20049 ( .C1(n16818), .C2(n16817), .A(n16816), .B(n17060), .ZN(
        n16820) );
  OAI22_X1 U20050 ( .A1(n17792), .A2(n17059), .B1(n17062), .B2(n17143), .ZN(
        n16819) );
  AOI211_X1 U20051 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16830), .A(n16820), 
        .B(n16819), .ZN(n16824) );
  OAI211_X1 U20052 ( .C1(n16827), .C2(n17143), .A(n17068), .B(n16821), .ZN(
        n16822) );
  NAND3_X1 U20053 ( .A1(n16824), .A2(n16823), .A3(n16822), .ZN(P3_U2650) );
  AOI211_X1 U20054 ( .C1(n17804), .C2(n16826), .A(n16825), .B(n17060), .ZN(
        n16829) );
  AOI211_X1 U20055 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16839), .A(n16827), .B(
        n17011), .ZN(n16828) );
  AOI211_X1 U20056 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17069), .A(n16829), .B(
        n16828), .ZN(n16833) );
  OAI221_X1 U20057 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n17051), .C1(
        P3_REIP_REG_20__SCAN_IN), .C2(n16831), .A(n16830), .ZN(n16832) );
  OAI211_X1 U20058 ( .C1(n17059), .C2(n10018), .A(n16833), .B(n16832), .ZN(
        P3_U2651) );
  AOI21_X1 U20059 ( .B1(n17051), .B2(n16834), .A(n17058), .ZN(n16859) );
  INV_X1 U20060 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18946) );
  NAND2_X1 U20061 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17811), .ZN(
        n16848) );
  INV_X1 U20062 ( .A(n16881), .ZN(n16868) );
  AOI21_X1 U20063 ( .B1(n17002), .B2(n16848), .A(n16868), .ZN(n16838) );
  INV_X1 U20064 ( .A(n16848), .ZN(n16836) );
  OAI21_X1 U20065 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16836), .A(
        n16835), .ZN(n17816) );
  OAI21_X1 U20066 ( .B1(n16838), .B2(n17816), .A(n18885), .ZN(n16837) );
  AOI21_X1 U20067 ( .B1(n16838), .B2(n17816), .A(n16837), .ZN(n16842) );
  OAI211_X1 U20068 ( .C1(n16846), .C2(n17196), .A(n17068), .B(n16839), .ZN(
        n16840) );
  OAI211_X1 U20069 ( .C1(n17062), .C2(n17196), .A(n18358), .B(n16840), .ZN(
        n16841) );
  AOI211_X1 U20070 ( .C1(n17038), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16842), .B(n16841), .ZN(n16845) );
  INV_X1 U20071 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18943) );
  NAND3_X1 U20072 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n16883), .ZN(n16860) );
  NOR2_X1 U20073 ( .A1(n18943), .A2(n16860), .ZN(n16852) );
  OAI211_X1 U20074 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16852), .B(n16843), .ZN(n16844) );
  OAI211_X1 U20075 ( .C1(n16859), .C2(n18946), .A(n16845), .B(n16844), .ZN(
        P3_U2652) );
  INV_X1 U20076 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17830) );
  AOI211_X1 U20077 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16861), .A(n16846), .B(
        n17011), .ZN(n16847) );
  AOI211_X1 U20078 ( .C1(n17069), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18348), .B(
        n16847), .ZN(n16855) );
  INV_X1 U20079 ( .A(n16859), .ZN(n16853) );
  INV_X1 U20080 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18944) );
  AOI21_X1 U20081 ( .B1(n17002), .B2(n16856), .A(n16868), .ZN(n16850) );
  OAI21_X1 U20082 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17811), .A(
        n16848), .ZN(n17827) );
  OAI21_X1 U20083 ( .B1(n16850), .B2(n17827), .A(n18885), .ZN(n16849) );
  AOI21_X1 U20084 ( .B1(n16850), .B2(n17827), .A(n16849), .ZN(n16851) );
  AOI221_X1 U20085 ( .B1(n16853), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n16852), 
        .C2(n18944), .A(n16851), .ZN(n16854) );
  OAI211_X1 U20086 ( .C1(n17830), .C2(n17059), .A(n16855), .B(n16854), .ZN(
        P3_U2653) );
  AND2_X1 U20087 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17836), .ZN(
        n16857) );
  INV_X1 U20088 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17040) );
  AOI21_X1 U20089 ( .B1(n16857), .B2(n17040), .A(n17025), .ZN(n16858) );
  OAI21_X1 U20090 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16857), .A(
        n16856), .ZN(n17840) );
  XNOR2_X1 U20091 ( .A(n16858), .B(n17840), .ZN(n16865) );
  AOI21_X1 U20092 ( .B1(n18943), .B2(n16860), .A(n16859), .ZN(n16864) );
  OAI211_X1 U20093 ( .C1(n16870), .C2(n21242), .A(n17068), .B(n16861), .ZN(
        n16862) );
  OAI21_X1 U20094 ( .B1(n17059), .B2(n10017), .A(n16862), .ZN(n16863) );
  AOI211_X1 U20095 ( .C1(n16865), .C2(n18885), .A(n16864), .B(n16863), .ZN(
        n16866) );
  OAI211_X1 U20096 ( .C1(n17062), .C2(n21242), .A(n16866), .B(n18358), .ZN(
        P3_U2654) );
  NAND2_X1 U20097 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16883), .ZN(n16877) );
  INV_X1 U20098 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18940) );
  INV_X1 U20099 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18938) );
  OAI21_X1 U20100 ( .B1(n16895), .B2(n17070), .A(n17073), .ZN(n16898) );
  AOI21_X1 U20101 ( .B1(n16883), .B2(n18938), .A(n16898), .ZN(n16876) );
  INV_X1 U20102 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16867) );
  AOI22_X1 U20103 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17836), .B1(
        n16867), .B2(n16878), .ZN(n17853) );
  INV_X1 U20104 ( .A(n17853), .ZN(n16869) );
  AOI221_X1 U20105 ( .B1(n16881), .B2(n16869), .C1(n16868), .C2(n17853), .A(
        n17060), .ZN(n16874) );
  AOI211_X1 U20106 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16884), .A(n16870), .B(
        n17011), .ZN(n16873) );
  AOI22_X1 U20107 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17038), .B1(
        n17069), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16871) );
  INV_X1 U20108 ( .A(n16871), .ZN(n16872) );
  NOR4_X1 U20109 ( .A1(n18348), .A2(n16874), .A3(n16873), .A4(n16872), .ZN(
        n16875) );
  OAI221_X1 U20110 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16877), .C1(n18940), 
        .C2(n16876), .A(n16875), .ZN(P3_U2655) );
  AOI22_X1 U20111 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17038), .B1(
        n17069), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n16887) );
  OAI21_X1 U20112 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17852), .A(
        n16878), .ZN(n17863) );
  NOR2_X1 U20113 ( .A1(n17060), .A2(n17002), .ZN(n17047) );
  INV_X1 U20114 ( .A(n17047), .ZN(n16880) );
  OAI221_X1 U20115 ( .B1(n17863), .B2(n17852), .C1(n17863), .C2(n17040), .A(
        n18885), .ZN(n16879) );
  AOI22_X1 U20116 ( .A1(n16881), .A2(n17863), .B1(n16880), .B2(n16879), .ZN(
        n16882) );
  AOI221_X1 U20117 ( .B1(n16898), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n16883), 
        .C2(n18938), .A(n16882), .ZN(n16886) );
  OAI211_X1 U20118 ( .C1(n16891), .C2(n17243), .A(n17068), .B(n16884), .ZN(
        n16885) );
  NAND4_X1 U20119 ( .A1(n16887), .A2(n16886), .A3(n18358), .A4(n16885), .ZN(
        P3_U2656) );
  INV_X1 U20120 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17994) );
  NAND2_X1 U20121 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9772), .ZN(
        n17001) );
  NOR2_X1 U20122 ( .A1(n17994), .A2(n17001), .ZN(n16992) );
  INV_X1 U20123 ( .A(n16992), .ZN(n16981) );
  NOR2_X1 U20124 ( .A1(n16888), .A2(n16981), .ZN(n16925) );
  AND2_X1 U20125 ( .A1(n17891), .A2(n16925), .ZN(n16903) );
  INV_X1 U20126 ( .A(n17852), .ZN(n16889) );
  OAI21_X1 U20127 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16903), .A(
        n16889), .ZN(n17883) );
  NAND2_X1 U20128 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16925), .ZN(
        n16904) );
  INV_X1 U20129 ( .A(n16904), .ZN(n16917) );
  NAND2_X1 U20130 ( .A1(n16917), .A2(n17040), .ZN(n16918) );
  INV_X1 U20131 ( .A(n16918), .ZN(n16890) );
  AOI21_X1 U20132 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16890), .A(
        n17025), .ZN(n16906) );
  XOR2_X1 U20133 ( .A(n17883), .B(n16906), .Z(n16901) );
  AOI211_X1 U20134 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16911), .A(n16891), .B(
        n17011), .ZN(n16894) );
  AOI21_X1 U20135 ( .B1(n17069), .B2(P3_EBX_REG_14__SCAN_IN), .A(n18348), .ZN(
        n16892) );
  INV_X1 U20136 ( .A(n16892), .ZN(n16893) );
  AOI211_X1 U20137 ( .C1(n17038), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16894), .B(n16893), .ZN(n16900) );
  NOR3_X1 U20138 ( .A1(n17070), .A2(n18934), .A3(n16902), .ZN(n16897) );
  INV_X1 U20139 ( .A(n16895), .ZN(n16896) );
  AOI22_X1 U20140 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16898), .B1(n16897), 
        .B2(n16896), .ZN(n16899) );
  OAI211_X1 U20141 ( .C1(n17060), .C2(n16901), .A(n16900), .B(n16899), .ZN(
        P3_U2657) );
  OR2_X1 U20142 ( .A1(n17070), .A2(n16902), .ZN(n16909) );
  INV_X1 U20143 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18932) );
  OAI21_X1 U20144 ( .B1(n16921), .B2(n17070), .A(n17073), .ZN(n16916) );
  AOI21_X1 U20145 ( .B1(n17051), .B2(n18932), .A(n16916), .ZN(n16908) );
  AOI21_X1 U20146 ( .B1(n17896), .B2(n16904), .A(n16903), .ZN(n17899) );
  AOI21_X1 U20147 ( .B1(n17899), .B2(n16918), .A(n17060), .ZN(n16905) );
  OAI22_X1 U20148 ( .A1(n17899), .A2(n16906), .B1(n17047), .B2(n16905), .ZN(
        n16907) );
  OAI221_X1 U20149 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n16909), .C1(n18934), 
        .C2(n16908), .A(n16907), .ZN(n16910) );
  AOI211_X1 U20150 ( .C1(n17069), .C2(P3_EBX_REG_13__SCAN_IN), .A(n18348), .B(
        n16910), .ZN(n16914) );
  OAI211_X1 U20151 ( .C1(n16915), .C2(n16912), .A(n17068), .B(n16911), .ZN(
        n16913) );
  OAI211_X1 U20152 ( .C1(n17059), .C2(n17896), .A(n16914), .B(n16913), .ZN(
        P3_U2658) );
  AOI211_X1 U20153 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16935), .A(n16915), .B(
        n17011), .ZN(n16924) );
  INV_X1 U20154 ( .A(n16916), .ZN(n16932) );
  NOR2_X1 U20155 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17070), .ZN(n16920) );
  INV_X1 U20156 ( .A(n16925), .ZN(n17894) );
  AOI21_X1 U20157 ( .B1(n17910), .B2(n17894), .A(n16917), .ZN(n17913) );
  NOR2_X1 U20158 ( .A1(n17913), .A2(n17041), .ZN(n16919) );
  AOI22_X1 U20159 ( .A1(n16921), .A2(n16920), .B1(n16919), .B2(n16918), .ZN(
        n16922) );
  OAI211_X1 U20160 ( .C1(n18932), .C2(n16932), .A(n16922), .B(n18358), .ZN(
        n16923) );
  AOI211_X1 U20161 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17069), .A(n16924), .B(
        n16923), .ZN(n16927) );
  NAND2_X1 U20162 ( .A1(n17002), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17061) );
  AND2_X1 U20163 ( .A1(n17061), .A2(n18885), .ZN(n17065) );
  OAI211_X1 U20164 ( .C1(n16925), .C2(n17025), .A(n17913), .B(n17065), .ZN(
        n16926) );
  OAI211_X1 U20165 ( .C1(n17059), .C2(n17910), .A(n16927), .B(n16926), .ZN(
        P3_U2659) );
  INV_X1 U20166 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16939) );
  NOR2_X1 U20167 ( .A1(n17070), .A2(n16940), .ZN(n16955) );
  AOI21_X1 U20168 ( .B1(n16928), .B2(n16955), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16933) );
  NAND2_X1 U20169 ( .A1(n17040), .A2(n16992), .ZN(n16982) );
  INV_X1 U20170 ( .A(n16982), .ZN(n16993) );
  AOI21_X1 U20171 ( .B1(n16929), .B2(n16993), .A(n17025), .ZN(n16930) );
  NOR2_X1 U20172 ( .A1(n17960), .A2(n16981), .ZN(n16957) );
  INV_X1 U20173 ( .A(n16957), .ZN(n16969) );
  NOR2_X1 U20174 ( .A1(n17922), .A2(n16969), .ZN(n16948) );
  OAI21_X1 U20175 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16948), .A(
        n17894), .ZN(n17923) );
  XOR2_X1 U20176 ( .A(n16930), .B(n17923), .Z(n16931) );
  OAI22_X1 U20177 ( .A1(n16933), .A2(n16932), .B1(n17060), .B2(n16931), .ZN(
        n16934) );
  AOI211_X1 U20178 ( .C1(n17069), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18348), .B(
        n16934), .ZN(n16938) );
  OAI211_X1 U20179 ( .C1(n16941), .C2(n16936), .A(n17068), .B(n16935), .ZN(
        n16937) );
  OAI211_X1 U20180 ( .C1(n17059), .C2(n16939), .A(n16938), .B(n16937), .ZN(
        P3_U2660) );
  AOI21_X1 U20181 ( .B1(n17051), .B2(n16940), .A(n17058), .ZN(n16977) );
  AOI211_X1 U20182 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16942), .A(n16941), .B(
        n17011), .ZN(n16947) );
  INV_X1 U20183 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n16945) );
  OAI211_X1 U20184 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(P3_REIP_REG_10__SCAN_IN), 
        .A(n16955), .B(n16943), .ZN(n16944) );
  OAI211_X1 U20185 ( .C1(n17062), .C2(n16945), .A(n18358), .B(n16944), .ZN(
        n16946) );
  AOI211_X1 U20186 ( .C1(n17038), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16947), .B(n16946), .ZN(n16954) );
  INV_X1 U20187 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16949) );
  NAND2_X1 U20188 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16957), .ZN(
        n16950) );
  AOI21_X1 U20189 ( .B1(n16949), .B2(n16950), .A(n16948), .ZN(n16952) );
  INV_X1 U20190 ( .A(n16950), .ZN(n16956) );
  AOI21_X1 U20191 ( .B1(n17040), .B2(n16956), .A(n17025), .ZN(n16951) );
  INV_X1 U20192 ( .A(n16952), .ZN(n17935) );
  INV_X1 U20193 ( .A(n16951), .ZN(n16959) );
  OAI221_X1 U20194 ( .B1(n16952), .B2(n16951), .C1(n17935), .C2(n16959), .A(
        n18885), .ZN(n16953) );
  OAI211_X1 U20195 ( .C1(n16977), .C2(n18929), .A(n16954), .B(n16953), .ZN(
        P3_U2661) );
  NOR2_X1 U20196 ( .A1(n16961), .A2(n17011), .ZN(n16970) );
  AOI22_X1 U20197 ( .A1(n16955), .A2(n21094), .B1(n16970), .B2(n17350), .ZN(
        n16966) );
  INV_X1 U20198 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17934) );
  AOI21_X1 U20199 ( .B1(n17934), .B2(n16969), .A(n16956), .ZN(n16960) );
  INV_X1 U20200 ( .A(n16960), .ZN(n17949) );
  NAND3_X1 U20201 ( .A1(n16957), .A2(n17934), .A3(n17040), .ZN(n16958) );
  OAI221_X1 U20202 ( .B1(n16960), .B2(n16959), .C1(n17949), .C2(n17002), .A(
        n16958), .ZN(n16964) );
  AOI21_X1 U20203 ( .B1(n17068), .B2(n16961), .A(n17069), .ZN(n16962) );
  OAI22_X1 U20204 ( .A1(n17934), .A2(n17059), .B1(n17350), .B2(n16962), .ZN(
        n16963) );
  AOI211_X1 U20205 ( .C1(n18885), .C2(n16964), .A(n18348), .B(n16963), .ZN(
        n16965) );
  OAI211_X1 U20206 ( .C1(n16977), .C2(n21094), .A(n16966), .B(n16965), .ZN(
        P3_U2662) );
  NAND2_X1 U20207 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16979) );
  INV_X1 U20208 ( .A(n16979), .ZN(n16968) );
  INV_X1 U20209 ( .A(n16967), .ZN(n16978) );
  NOR2_X1 U20210 ( .A1(n17070), .A2(n16978), .ZN(n16995) );
  AOI21_X1 U20211 ( .B1(n16968), .B2(n16995), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n16976) );
  AOI22_X1 U20212 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17038), .B1(
        n17069), .B2(P3_EBX_REG_8__SCAN_IN), .ZN(n16975) );
  INV_X1 U20213 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17976) );
  NOR2_X1 U20214 ( .A1(n17976), .A2(n16981), .ZN(n16980) );
  AOI21_X1 U20215 ( .B1(n16980), .B2(n17040), .A(n17025), .ZN(n16984) );
  OAI21_X1 U20216 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16980), .A(
        n16969), .ZN(n17962) );
  XNOR2_X1 U20217 ( .A(n16984), .B(n17962), .ZN(n16973) );
  INV_X1 U20218 ( .A(n16970), .ZN(n16971) );
  AOI21_X1 U20219 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n16988), .A(n16971), .ZN(
        n16972) );
  AOI211_X1 U20220 ( .C1(n18885), .C2(n16973), .A(n18348), .B(n16972), .ZN(
        n16974) );
  OAI211_X1 U20221 ( .C1(n16977), .C2(n16976), .A(n16975), .B(n16974), .ZN(
        P3_U2663) );
  AOI21_X1 U20222 ( .B1(n17051), .B2(n16978), .A(n17058), .ZN(n17004) );
  INV_X1 U20223 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18925) );
  OAI211_X1 U20224 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16995), .B(n16979), .ZN(n16986) );
  AOI21_X1 U20225 ( .B1(n17976), .B2(n16981), .A(n16980), .ZN(n17981) );
  AOI21_X1 U20226 ( .B1(n17981), .B2(n16982), .A(n17060), .ZN(n16983) );
  OAI22_X1 U20227 ( .A1(n17981), .A2(n16984), .B1(n17047), .B2(n16983), .ZN(
        n16985) );
  OAI211_X1 U20228 ( .C1(n17004), .C2(n18925), .A(n16986), .B(n16985), .ZN(
        n16987) );
  AOI211_X1 U20229 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n17038), .A(
        n18348), .B(n16987), .ZN(n16990) );
  OAI211_X1 U20230 ( .C1(n16991), .C2(n17390), .A(n17068), .B(n16988), .ZN(
        n16989) );
  OAI211_X1 U20231 ( .C1(n17390), .C2(n17062), .A(n16990), .B(n16989), .ZN(
        P3_U2664) );
  INV_X1 U20232 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18923) );
  AOI211_X1 U20233 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17007), .A(n16991), .B(
        n17011), .ZN(n16999) );
  INV_X1 U20234 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17398) );
  AOI21_X1 U20235 ( .B1(n17994), .B2(n17001), .A(n16992), .ZN(n17991) );
  NOR3_X1 U20236 ( .A1(n17991), .A2(n16993), .A3(n17041), .ZN(n16994) );
  AOI211_X1 U20237 ( .C1(n16995), .C2(n18923), .A(n18348), .B(n16994), .ZN(
        n16997) );
  OAI211_X1 U20238 ( .C1(n17994), .C2(n17025), .A(n17991), .B(n17065), .ZN(
        n16996) );
  OAI211_X1 U20239 ( .C1(n17398), .C2(n17062), .A(n16997), .B(n16996), .ZN(
        n16998) );
  AOI211_X1 U20240 ( .C1(n17038), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16999), .B(n16998), .ZN(n17000) );
  OAI21_X1 U20241 ( .B1(n18923), .B2(n17004), .A(n17000), .ZN(P3_U2665) );
  NOR2_X1 U20242 ( .A1(n17070), .A2(n17017), .ZN(n17014) );
  AOI21_X1 U20243 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17014), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17005) );
  NOR2_X1 U20244 ( .A1(n21104), .A2(n17996), .ZN(n17015) );
  OAI21_X1 U20245 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17015), .A(
        n17001), .ZN(n18004) );
  NAND2_X1 U20246 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17040), .ZN(
        n17043) );
  OAI21_X1 U20247 ( .B1(n17996), .B2(n17043), .A(n17002), .ZN(n17016) );
  XNOR2_X1 U20248 ( .A(n18004), .B(n17016), .ZN(n17003) );
  OAI22_X1 U20249 ( .A1(n17005), .A2(n17004), .B1(n17060), .B2(n17003), .ZN(
        n17006) );
  AOI211_X1 U20250 ( .C1(n17069), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18348), .B(
        n17006), .ZN(n17010) );
  OAI211_X1 U20251 ( .C1(n17012), .C2(n17008), .A(n17068), .B(n17007), .ZN(
        n17009) );
  OAI211_X1 U20252 ( .C1(n17059), .C2(n17995), .A(n17010), .B(n17009), .ZN(
        P3_U2666) );
  AOI211_X1 U20253 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17033), .A(n17012), .B(
        n17011), .ZN(n17013) );
  AOI21_X1 U20254 ( .B1(n17014), .B2(n18919), .A(n17013), .ZN(n17023) );
  NAND2_X1 U20255 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18018), .ZN(
        n17026) );
  AOI21_X1 U20256 ( .B1(n10015), .B2(n17026), .A(n17015), .ZN(n18019) );
  NAND2_X1 U20257 ( .A1(n18018), .A2(n10015), .ZN(n18015) );
  OAI22_X1 U20258 ( .A1(n18019), .A2(n17016), .B1(n17043), .B2(n18015), .ZN(
        n17021) );
  AOI21_X1 U20259 ( .B1(n17051), .B2(n17017), .A(n17058), .ZN(n17028) );
  AOI22_X1 U20260 ( .A1(n17069), .A2(P3_EBX_REG_4__SCAN_IN), .B1(n18019), .B2(
        n17047), .ZN(n17019) );
  NAND2_X1 U20261 ( .A1(n18379), .A2(n19044), .ZN(n19049) );
  INV_X1 U20262 ( .A(n19049), .ZN(n17071) );
  OAI21_X1 U20263 ( .B1(n17215), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n17071), .ZN(n17018) );
  OAI211_X1 U20264 ( .C1(n17028), .C2(n18919), .A(n17019), .B(n17018), .ZN(
        n17020) );
  AOI211_X1 U20265 ( .C1(n18885), .C2(n17021), .A(n18348), .B(n17020), .ZN(
        n17022) );
  OAI211_X1 U20266 ( .C1(n10015), .C2(n17059), .A(n17023), .B(n17022), .ZN(
        P3_U2667) );
  NOR2_X1 U20267 ( .A1(n13063), .A2(n9732), .ZN(n18840) );
  NAND2_X1 U20268 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18840), .ZN(
        n18825) );
  INV_X1 U20269 ( .A(n18825), .ZN(n17024) );
  OAI21_X1 U20270 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n17024), .A(
        n17373), .ZN(n18987) );
  NOR2_X1 U20271 ( .A1(n21104), .A2(n18039), .ZN(n17039) );
  AOI21_X1 U20272 ( .B1(n17039), .B2(n17040), .A(n17025), .ZN(n17027) );
  OAI21_X1 U20273 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17039), .A(
        n17026), .ZN(n18033) );
  XNOR2_X1 U20274 ( .A(n17027), .B(n18033), .ZN(n17032) );
  INV_X1 U20275 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18917) );
  NAND2_X1 U20276 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17050) );
  AOI221_X1 U20277 ( .B1(n17070), .B2(n18917), .C1(n17050), .C2(n18917), .A(
        n17028), .ZN(n17031) );
  OAI22_X1 U20278 ( .A1(n17029), .A2(n17059), .B1(n17062), .B2(n17034), .ZN(
        n17030) );
  AOI211_X1 U20279 ( .C1(n17032), .C2(n18885), .A(n17031), .B(n17030), .ZN(
        n17037) );
  OAI211_X1 U20280 ( .C1(n17035), .C2(n17034), .A(n17068), .B(n17033), .ZN(
        n17036) );
  OAI211_X1 U20281 ( .C1(n19049), .C2(n18987), .A(n17037), .B(n17036), .ZN(
        P3_U2668) );
  AOI22_X1 U20282 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17038), .B1(
        n17069), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n17055) );
  AOI21_X1 U20283 ( .B1(n21104), .B2(n18039), .A(n17039), .ZN(n18042) );
  AND2_X1 U20284 ( .A1(n17040), .A2(n17039), .ZN(n17042) );
  AOI211_X1 U20285 ( .C1(n18042), .C2(n17043), .A(n17042), .B(n17041), .ZN(
        n17046) );
  INV_X1 U20286 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18915) );
  INV_X1 U20287 ( .A(n17044), .ZN(n18839) );
  NAND2_X1 U20288 ( .A1(n13063), .A2(n18839), .ZN(n18823) );
  NAND2_X1 U20289 ( .A1(n18823), .A2(n18825), .ZN(n18995) );
  OAI22_X1 U20290 ( .A1(n17073), .A2(n18915), .B1(n18995), .B2(n19049), .ZN(
        n17045) );
  AOI211_X1 U20291 ( .C1(n17047), .C2(n18042), .A(n17046), .B(n17045), .ZN(
        n17054) );
  NOR2_X1 U20292 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17057) );
  OAI211_X1 U20293 ( .C1(n17057), .C2(n17049), .A(n17068), .B(n17048), .ZN(
        n17053) );
  OAI211_X1 U20294 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17051), .B(n17050), .ZN(n17052) );
  NAND4_X1 U20295 ( .A1(n17055), .A2(n17054), .A3(n17053), .A4(n17052), .ZN(
        P3_U2669) );
  NAND2_X1 U20296 ( .A1(n17056), .A2(n18839), .ZN(n19001) );
  NOR2_X1 U20297 ( .A1(n17057), .A2(n17395), .ZN(n17418) );
  AOI22_X1 U20298 ( .A1(n17068), .A2(n17418), .B1(n17058), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17067) );
  OAI21_X1 U20299 ( .B1(n17061), .B2(n17060), .A(n17059), .ZN(n17064) );
  OAI22_X1 U20300 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17070), .B1(n17062), 
        .B2(n17420), .ZN(n17063) );
  AOI221_X1 U20301 ( .B1(n17065), .B2(n21104), .C1(n17064), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17063), .ZN(n17066) );
  OAI211_X1 U20302 ( .C1(n19001), .C2(n19049), .A(n17067), .B(n17066), .ZN(
        P3_U2670) );
  NOR2_X1 U20303 ( .A1(n17069), .A2(n17068), .ZN(n17076) );
  NAND2_X1 U20304 ( .A1(n17073), .A2(n17070), .ZN(n17072) );
  AOI22_X1 U20305 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17072), .B1(n17071), 
        .B2(n19014), .ZN(n17075) );
  NAND3_X1 U20306 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18996), .A3(
        n17073), .ZN(n17074) );
  OAI211_X1 U20307 ( .C1(n17076), .C2(n17425), .A(n17075), .B(n17074), .ZN(
        P3_U2671) );
  INV_X1 U20308 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17077) );
  NOR3_X1 U20309 ( .A1(n17077), .A2(n17196), .A3(n17183), .ZN(n17158) );
  NAND4_X1 U20310 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n17078), .A4(n17158), .ZN(n17079) );
  NOR4_X1 U20311 ( .A1(n17121), .A2(n21312), .A3(n17143), .A4(n17079), .ZN(
        n17080) );
  NAND3_X1 U20312 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17080), .ZN(n17083) );
  NAND2_X1 U20313 ( .A1(n17414), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17082) );
  NAND2_X1 U20314 ( .A1(n17112), .A2(n18410), .ZN(n17081) );
  OAI22_X1 U20315 ( .A1(n17112), .A2(n17082), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17081), .ZN(P3_U2672) );
  NAND2_X1 U20316 ( .A1(n17084), .A2(n17083), .ZN(n17085) );
  NAND2_X1 U20317 ( .A1(n17085), .A2(n17414), .ZN(n17111) );
  AOI22_X1 U20318 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20319 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9765), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20320 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17087) );
  OAI211_X1 U20321 ( .C1(n17298), .C2(n21214), .A(n17088), .B(n17087), .ZN(
        n17094) );
  AOI22_X1 U20322 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17332), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20323 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17091) );
  AOI22_X1 U20324 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17090) );
  NAND2_X1 U20325 ( .A1(n13113), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n17089) );
  NAND4_X1 U20326 ( .A1(n17092), .A2(n17091), .A3(n17090), .A4(n17089), .ZN(
        n17093) );
  AOI211_X1 U20327 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17094), .B(n17093), .ZN(n17095) );
  OAI211_X1 U20328 ( .C1(n13090), .C2(n18614), .A(n17096), .B(n17095), .ZN(
        n17116) );
  NAND3_X1 U20329 ( .A1(n17114), .A2(n17113), .A3(n17116), .ZN(n17110) );
  AOI22_X1 U20330 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17097) );
  OAI21_X1 U20331 ( .B1(n9785), .B2(n21122), .A(n17097), .ZN(n17108) );
  AOI22_X1 U20332 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U20333 ( .A1(n13113), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17098) );
  OAI21_X1 U20334 ( .B1(n17210), .B2(n18438), .A(n17098), .ZN(n17103) );
  AOI22_X1 U20335 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17314), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20336 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17099) );
  OAI211_X1 U20337 ( .C1(n17298), .C2(n17101), .A(n17100), .B(n17099), .ZN(
        n17102) );
  AOI211_X1 U20338 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n17103), .B(n17102), .ZN(n17104) );
  OAI211_X1 U20339 ( .C1(n15914), .C2(n17106), .A(n17105), .B(n17104), .ZN(
        n17107) );
  AOI211_X1 U20340 ( .C1(n9765), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n17108), .B(n17107), .ZN(n17109) );
  XNOR2_X1 U20341 ( .A(n17110), .B(n17109), .ZN(n17440) );
  OAI22_X1 U20342 ( .A1(n17112), .A2(n17111), .B1(n17440), .B2(n17414), .ZN(
        P3_U2673) );
  NAND2_X1 U20343 ( .A1(n17114), .A2(n17113), .ZN(n17115) );
  XOR2_X1 U20344 ( .A(n17116), .B(n17115), .Z(n17444) );
  OAI21_X1 U20345 ( .B1(n17118), .B2(n17117), .A(n17121), .ZN(n17119) );
  OAI21_X1 U20346 ( .B1(n17121), .B2(n17120), .A(n17119), .ZN(n17122) );
  OAI21_X1 U20347 ( .B1(n17414), .B2(n17444), .A(n17122), .ZN(P3_U2674) );
  OAI211_X1 U20348 ( .C1(n17452), .C2(n17451), .A(n17422), .B(n17450), .ZN(
        n17123) );
  OAI221_X1 U20349 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17126), .C1(n17125), 
        .C2(n17124), .A(n17123), .ZN(P3_U2676) );
  AOI21_X1 U20350 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17414), .A(n17134), .ZN(
        n17128) );
  XNOR2_X1 U20351 ( .A(n17127), .B(n17130), .ZN(n17461) );
  OAI22_X1 U20352 ( .A1(n17129), .A2(n17128), .B1(n17414), .B2(n17461), .ZN(
        P3_U2677) );
  AOI21_X1 U20353 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17414), .A(n17137), .ZN(
        n17133) );
  OAI21_X1 U20354 ( .B1(n17132), .B2(n17131), .A(n17130), .ZN(n17465) );
  OAI22_X1 U20355 ( .A1(n17134), .A2(n17133), .B1(n17414), .B2(n17465), .ZN(
        P3_U2678) );
  AOI21_X1 U20356 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17414), .A(n17142), .ZN(
        n17136) );
  XNOR2_X1 U20357 ( .A(n17135), .B(n17138), .ZN(n17471) );
  OAI22_X1 U20358 ( .A1(n17137), .A2(n17136), .B1(n17414), .B2(n17471), .ZN(
        P3_U2679) );
  AOI21_X1 U20359 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17414), .A(n17157), .ZN(
        n17141) );
  OAI21_X1 U20360 ( .B1(n17140), .B2(n17139), .A(n17138), .ZN(n17476) );
  OAI22_X1 U20361 ( .A1(n17142), .A2(n17141), .B1(n17414), .B2(n17476), .ZN(
        P3_U2680) );
  OAI22_X1 U20362 ( .A1(n21312), .A2(n17422), .B1(n17143), .B2(n17170), .ZN(
        n17144) );
  INV_X1 U20363 ( .A(n17144), .ZN(n17156) );
  INV_X1 U20364 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17260) );
  AOI22_X1 U20365 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17145) );
  OAI21_X1 U20366 ( .B1(n17327), .B2(n17260), .A(n17145), .ZN(n17155) );
  AOI22_X1 U20367 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17153) );
  OAI22_X1 U20368 ( .A1(n17338), .A2(n17146), .B1(n15914), .B2(n18614), .ZN(
        n17151) );
  AOI22_X1 U20369 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20370 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20371 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17377), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17147) );
  NAND3_X1 U20372 ( .A1(n17149), .A2(n17148), .A3(n17147), .ZN(n17150) );
  AOI211_X1 U20373 ( .C1(n17368), .C2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n17151), .B(n17150), .ZN(n17152) );
  OAI211_X1 U20374 ( .C1(n17295), .C2(n21214), .A(n17153), .B(n17152), .ZN(
        n17154) );
  AOI211_X1 U20375 ( .C1(n9720), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n17155), .B(n17154), .ZN(n17481) );
  OAI22_X1 U20376 ( .A1(n17157), .A2(n17156), .B1(n17481), .B2(n17414), .ZN(
        P3_U2681) );
  NOR2_X1 U20377 ( .A1(n17422), .A2(n17158), .ZN(n17181) );
  AOI22_X1 U20378 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U20379 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17159) );
  OAI21_X1 U20380 ( .B1(n17327), .B2(n17286), .A(n17159), .ZN(n17166) );
  AOI22_X1 U20381 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17377), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17164) );
  INV_X1 U20382 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20383 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20384 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17160) );
  OAI211_X1 U20385 ( .C1(n17317), .C2(n17276), .A(n17161), .B(n17160), .ZN(
        n17162) );
  AOI21_X1 U20386 ( .B1(n13113), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n17162), .ZN(n17163) );
  OAI211_X1 U20387 ( .C1(n17210), .C2(n17405), .A(n17164), .B(n17163), .ZN(
        n17165) );
  AOI211_X1 U20388 ( .C1(n17086), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n17166), .B(n17165), .ZN(n17167) );
  OAI211_X1 U20389 ( .C1(n13089), .C2(n21226), .A(n17168), .B(n17167), .ZN(
        n17486) );
  AOI22_X1 U20390 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17181), .B1(n17422), 
        .B2(n17486), .ZN(n17169) );
  OAI21_X1 U20391 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17170), .A(n17169), .ZN(
        P3_U2682) );
  AOI22_X1 U20392 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17171) );
  OAI21_X1 U20393 ( .B1(n17327), .B2(n17306), .A(n17171), .ZN(n17180) );
  AOI22_X1 U20394 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20395 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17172) );
  OAI21_X1 U20396 ( .B1(n17298), .B2(n17294), .A(n17172), .ZN(n17176) );
  INV_X1 U20397 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21261) );
  AOI22_X1 U20398 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9720), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20399 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17173) );
  OAI211_X1 U20400 ( .C1(n17338), .C2(n21261), .A(n17174), .B(n17173), .ZN(
        n17175) );
  AOI211_X1 U20401 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17176), .B(n17175), .ZN(n17177) );
  OAI211_X1 U20402 ( .C1(n17210), .C2(n17407), .A(n17178), .B(n17177), .ZN(
        n17179) );
  AOI211_X1 U20403 ( .C1(n17314), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17180), .B(n17179), .ZN(n17494) );
  OAI221_X1 U20404 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(P3_EBX_REG_19__SCAN_IN), 
        .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17194), .A(n17181), .ZN(n17182) );
  OAI21_X1 U20405 ( .B1(n17494), .B2(n17414), .A(n17182), .ZN(P3_U2683) );
  NAND2_X1 U20406 ( .A1(n17414), .A2(n17183), .ZN(n17212) );
  INV_X1 U20407 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U20408 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20409 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9716), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20410 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17184) );
  OAI211_X1 U20411 ( .C1(n17338), .C2(n17313), .A(n17185), .B(n17184), .ZN(
        n17191) );
  AOI22_X1 U20412 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20413 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20414 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17187) );
  NAND2_X1 U20415 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n17186) );
  NAND4_X1 U20416 ( .A1(n17189), .A2(n17188), .A3(n17187), .A4(n17186), .ZN(
        n17190) );
  AOI211_X1 U20417 ( .C1(n17377), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n17191), .B(n17190), .ZN(n17192) );
  OAI211_X1 U20418 ( .C1(n17210), .C2(n17411), .A(n17193), .B(n17192), .ZN(
        n17495) );
  AOI22_X1 U20419 ( .A1(n17422), .A2(n17495), .B1(n17194), .B2(n17196), .ZN(
        n17195) );
  OAI21_X1 U20420 ( .B1(n17196), .B2(n17212), .A(n17195), .ZN(P3_U2684) );
  NAND2_X1 U20421 ( .A1(n18410), .A2(n17197), .ZN(n17226) );
  INV_X1 U20422 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20423 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20424 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17198) );
  OAI21_X1 U20425 ( .B1(n17327), .B2(n17346), .A(n17198), .ZN(n17207) );
  AOI22_X1 U20426 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U20427 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U20428 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17200) );
  OAI211_X1 U20429 ( .C1(n17317), .C2(n18424), .A(n17201), .B(n17200), .ZN(
        n17202) );
  AOI21_X1 U20430 ( .B1(n17377), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17202), .ZN(n17203) );
  OAI211_X1 U20431 ( .C1(n17205), .C2(n21323), .A(n17204), .B(n17203), .ZN(
        n17206) );
  AOI211_X1 U20432 ( .C1(n9720), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n17207), .B(n17206), .ZN(n17208) );
  OAI211_X1 U20433 ( .C1(n17210), .C2(n17416), .A(n17209), .B(n17208), .ZN(
        n17499) );
  NAND2_X1 U20434 ( .A1(n17422), .A2(n17499), .ZN(n17211) );
  OAI221_X1 U20435 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17226), .C1(n17213), 
        .C2(n17212), .A(n17211), .ZN(P3_U2685) );
  OAI22_X1 U20436 ( .A1(n17214), .A2(n17338), .B1(n17327), .B2(n17353), .ZN(
        n17225) );
  AOI22_X1 U20437 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17215), .ZN(n17223) );
  AOI22_X1 U20438 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17367), .B1(
        n17314), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20439 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17334), .ZN(n17216) );
  OAI21_X1 U20440 ( .B1(n9785), .B2(n17354), .A(n17216), .ZN(n17220) );
  AOI22_X1 U20441 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n9767), .ZN(n17218) );
  AOI22_X1 U20442 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n9717), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17199), .ZN(n17217) );
  OAI211_X1 U20443 ( .C1(n17317), .C2(n18421), .A(n17218), .B(n17217), .ZN(
        n17219) );
  AOI211_X1 U20444 ( .C1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .C2(n17377), .A(
        n17220), .B(n17219), .ZN(n17221) );
  NAND3_X1 U20445 ( .A1(n17223), .A2(n17222), .A3(n17221), .ZN(n17224) );
  AOI211_X1 U20446 ( .C1(n17368), .C2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n17225), .B(n17224), .ZN(n17509) );
  INV_X1 U20447 ( .A(n17240), .ZN(n17227) );
  OAI21_X1 U20448 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17227), .A(n17226), .ZN(
        n17228) );
  AOI22_X1 U20449 ( .A1(n17422), .A2(n17509), .B1(n17228), .B2(n17414), .ZN(
        P3_U2686) );
  OAI22_X1 U20450 ( .A1(n17229), .A2(n17372), .B1(n17327), .B2(n21155), .ZN(
        n17239) );
  AOI22_X1 U20451 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20452 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17236) );
  INV_X1 U20453 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17370) );
  AOI22_X1 U20454 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17230) );
  OAI21_X1 U20455 ( .B1(n17338), .B2(n17370), .A(n17230), .ZN(n17234) );
  AOI22_X1 U20456 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U20457 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17231) );
  OAI211_X1 U20458 ( .C1(n17317), .C2(n18418), .A(n17232), .B(n17231), .ZN(
        n17233) );
  AOI211_X1 U20459 ( .C1(n17377), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n17234), .B(n17233), .ZN(n17235) );
  NAND3_X1 U20460 ( .A1(n17237), .A2(n17236), .A3(n17235), .ZN(n17238) );
  AOI211_X1 U20461 ( .C1(n17368), .C2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n17239), .B(n17238), .ZN(n17515) );
  OAI21_X1 U20462 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17257), .A(n17240), .ZN(
        n17241) );
  AOI22_X1 U20463 ( .A1(n17422), .A2(n17515), .B1(n17241), .B2(n17414), .ZN(
        P3_U2687) );
  AOI21_X1 U20464 ( .B1(n17243), .B2(n17242), .A(n17422), .ZN(n17244) );
  INV_X1 U20465 ( .A(n17244), .ZN(n17256) );
  AOI22_X1 U20466 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9716), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17245) );
  OAI21_X1 U20467 ( .B1(n15914), .B2(n21266), .A(n17245), .ZN(n17255) );
  AOI22_X1 U20468 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17253) );
  INV_X1 U20469 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20470 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17246) );
  OAI21_X1 U20471 ( .B1(n17298), .B2(n17247), .A(n17246), .ZN(n17251) );
  AOI22_X1 U20472 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17249) );
  AOI22_X1 U20473 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17314), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17248) );
  OAI211_X1 U20474 ( .C1(n17317), .C2(n21122), .A(n17249), .B(n17248), .ZN(
        n17250) );
  AOI211_X1 U20475 ( .C1(n13113), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n17251), .B(n17250), .ZN(n17252) );
  OAI211_X1 U20476 ( .C1(n17373), .C2(n18438), .A(n17253), .B(n17252), .ZN(
        n17254) );
  AOI211_X1 U20477 ( .C1(n17086), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n17255), .B(n17254), .ZN(n17519) );
  OAI22_X1 U20478 ( .A1(n17257), .A2(n17256), .B1(n17519), .B2(n17414), .ZN(
        P3_U2688) );
  NAND2_X1 U20479 ( .A1(n18410), .A2(n17258), .ZN(n17273) );
  NOR2_X1 U20480 ( .A1(n17422), .A2(n17258), .ZN(n17290) );
  AOI22_X1 U20481 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20482 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17270) );
  OAI22_X1 U20483 ( .A1(n13089), .A2(n17260), .B1(n13090), .B2(n17259), .ZN(
        n17268) );
  AOI22_X1 U20484 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17375), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17266) );
  AOI22_X1 U20485 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9716), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17262) );
  AOI22_X1 U20486 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17261) );
  OAI211_X1 U20487 ( .C1(n17338), .C2(n17263), .A(n17262), .B(n17261), .ZN(
        n17264) );
  AOI21_X1 U20488 ( .B1(n17377), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17264), .ZN(n17265) );
  OAI211_X1 U20489 ( .C1(n17327), .C2(n18614), .A(n17266), .B(n17265), .ZN(
        n17267) );
  AOI211_X1 U20490 ( .C1(n17199), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n17268), .B(n17267), .ZN(n17269) );
  NAND3_X1 U20491 ( .A1(n17271), .A2(n17270), .A3(n17269), .ZN(n17522) );
  AOI22_X1 U20492 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17290), .B1(n17422), 
        .B2(n17522), .ZN(n17272) );
  OAI21_X1 U20493 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17273), .A(n17272), .ZN(
        P3_U2689) );
  AOI22_X1 U20494 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17275) );
  OAI21_X1 U20495 ( .B1(n17373), .B2(n17276), .A(n17275), .ZN(n17288) );
  AOI22_X1 U20496 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17285) );
  OAI22_X1 U20497 ( .A1(n17327), .A2(n17278), .B1(n17338), .B2(n17277), .ZN(
        n17283) );
  AOI22_X1 U20498 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20499 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U20500 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17377), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17279) );
  NAND3_X1 U20501 ( .A1(n17281), .A2(n17280), .A3(n17279), .ZN(n17282) );
  AOI211_X1 U20502 ( .C1(n17368), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n17283), .B(n17282), .ZN(n17284) );
  OAI211_X1 U20503 ( .C1(n13089), .C2(n17286), .A(n17285), .B(n17284), .ZN(
        n17287) );
  AOI211_X1 U20504 ( .C1(n9720), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n17288), .B(n17287), .ZN(n17526) );
  INV_X1 U20505 ( .A(n17289), .ZN(n17291) );
  OAI21_X1 U20506 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17291), .A(n17290), .ZN(
        n17292) );
  OAI21_X1 U20507 ( .B1(n17526), .B2(n17414), .A(n17292), .ZN(P3_U2690) );
  AOI22_X1 U20508 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17293) );
  OAI21_X1 U20509 ( .B1(n17295), .B2(n17294), .A(n17293), .ZN(n17308) );
  AOI22_X1 U20510 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17305) );
  INV_X1 U20511 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17297) );
  AOI22_X1 U20512 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17296) );
  OAI21_X1 U20513 ( .B1(n17298), .B2(n17297), .A(n17296), .ZN(n17303) );
  AOI22_X1 U20514 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20515 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17299) );
  OAI211_X1 U20516 ( .C1(n17338), .C2(n17301), .A(n17300), .B(n17299), .ZN(
        n17302) );
  AOI211_X1 U20517 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n17303), .B(n17302), .ZN(n17304) );
  OAI211_X1 U20518 ( .C1(n13089), .C2(n17306), .A(n17305), .B(n17304), .ZN(
        n17307) );
  AOI211_X1 U20519 ( .C1(n9767), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n17308), .B(n17307), .ZN(n17530) );
  NOR2_X1 U20520 ( .A1(n17422), .A2(n17310), .ZN(n17328) );
  NOR2_X1 U20521 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17478), .ZN(n17309) );
  AOI22_X1 U20522 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17328), .B1(n17310), 
        .B2(n17309), .ZN(n17311) );
  OAI21_X1 U20523 ( .B1(n17530), .B2(n17414), .A(n17311), .ZN(P3_U2691) );
  AOI22_X1 U20524 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17326) );
  AOI22_X1 U20525 ( .A1(n9767), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17312) );
  OAI21_X1 U20526 ( .B1(n17371), .B2(n17313), .A(n17312), .ZN(n17324) );
  AOI22_X1 U20527 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17377), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17320) );
  AOI22_X1 U20528 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17316) );
  AOI22_X1 U20529 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17315) );
  OAI211_X1 U20530 ( .C1(n17317), .C2(n17411), .A(n17316), .B(n17315), .ZN(
        n17318) );
  AOI21_X1 U20531 ( .B1(n13113), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17318), .ZN(n17319) );
  OAI211_X1 U20532 ( .C1(n17322), .C2(n17321), .A(n17320), .B(n17319), .ZN(
        n17323) );
  AOI211_X1 U20533 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17324), .B(n17323), .ZN(n17325) );
  OAI211_X1 U20534 ( .C1(n17327), .C2(n21200), .A(n17326), .B(n17325), .ZN(
        n17533) );
  INV_X1 U20535 ( .A(n17533), .ZN(n17331) );
  INV_X1 U20536 ( .A(n17347), .ZN(n17329) );
  OAI21_X1 U20537 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17329), .A(n17328), .ZN(
        n17330) );
  OAI21_X1 U20538 ( .B1(n17331), .B2(n17414), .A(n17330), .ZN(P3_U2692) );
  AOI22_X1 U20539 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17332), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17345) );
  AOI22_X1 U20540 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17333) );
  OAI21_X1 U20541 ( .B1(n9785), .B2(n21323), .A(n17333), .ZN(n17343) );
  AOI22_X1 U20542 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17334), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17341) );
  INV_X1 U20543 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17337) );
  AOI22_X1 U20544 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9767), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17336) );
  AOI22_X1 U20545 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17199), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17335) );
  OAI211_X1 U20546 ( .C1(n17338), .C2(n17337), .A(n17336), .B(n17335), .ZN(
        n17339) );
  AOI21_X1 U20547 ( .B1(n17377), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n17339), .ZN(n17340) );
  OAI211_X1 U20548 ( .C1(n17317), .C2(n17416), .A(n17341), .B(n17340), .ZN(
        n17342) );
  AOI211_X1 U20549 ( .C1(n9720), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n17343), .B(n17342), .ZN(n17344) );
  OAI211_X1 U20550 ( .C1(n13089), .C2(n17346), .A(n17345), .B(n17344), .ZN(
        n17536) );
  INV_X1 U20551 ( .A(n17536), .ZN(n17349) );
  OAI21_X1 U20552 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17366), .A(n17347), .ZN(
        n17348) );
  AOI22_X1 U20553 ( .A1(n17422), .A2(n17349), .B1(n17348), .B2(n17414), .ZN(
        P3_U2693) );
  AOI21_X1 U20554 ( .B1(n17350), .B2(n17386), .A(n17422), .ZN(n17351) );
  INV_X1 U20555 ( .A(n17351), .ZN(n17365) );
  AOI22_X1 U20556 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n9716), .ZN(n17352) );
  OAI21_X1 U20557 ( .B1(n13089), .B2(n17353), .A(n17352), .ZN(n17364) );
  INV_X1 U20558 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17362) );
  AOI22_X1 U20559 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17334), .B1(
        n17377), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17361) );
  OAI22_X1 U20560 ( .A1(n17210), .A2(n17354), .B1(n17373), .B2(n18421), .ZN(
        n17359) );
  AOI22_X1 U20561 ( .A1(n9765), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n9767), .ZN(n17357) );
  AOI22_X1 U20562 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17367), .B1(
        n9720), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17356) );
  AOI22_X1 U20563 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13113), .B1(
        n17375), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17355) );
  NAND3_X1 U20564 ( .A1(n17357), .A2(n17356), .A3(n17355), .ZN(n17358) );
  AOI211_X1 U20565 ( .C1(n17274), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n17359), .B(n17358), .ZN(n17360) );
  OAI211_X1 U20566 ( .C1(n17362), .C2(n15914), .A(n17361), .B(n17360), .ZN(
        n17363) );
  AOI211_X1 U20567 ( .C1(n17086), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n17364), .B(n17363), .ZN(n17540) );
  OAI22_X1 U20568 ( .A1(n17366), .A2(n17365), .B1(n17540), .B2(n17414), .ZN(
        P3_U2694) );
  AOI22_X1 U20569 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U20570 ( .A1(n17199), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17369) );
  OAI21_X1 U20571 ( .B1(n17371), .B2(n17370), .A(n17369), .ZN(n17383) );
  OAI22_X1 U20572 ( .A1(n17373), .A2(n18418), .B1(n13090), .B2(n17372), .ZN(
        n17374) );
  AOI21_X1 U20573 ( .B1(n17375), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n17374), .ZN(n17381) );
  AOI22_X1 U20574 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9767), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U20575 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17379) );
  AOI22_X1 U20576 ( .A1(n17377), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13113), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17378) );
  NAND4_X1 U20577 ( .A1(n17381), .A2(n17380), .A3(n17379), .A4(n17378), .ZN(
        n17382) );
  AOI211_X1 U20578 ( .C1(n9765), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n17383), .B(n17382), .ZN(n17384) );
  OAI211_X1 U20579 ( .C1(n13089), .C2(n21155), .A(n17385), .B(n17384), .ZN(
        n17546) );
  INV_X1 U20580 ( .A(n17546), .ZN(n17388) );
  OAI21_X1 U20581 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17393), .A(n17386), .ZN(
        n17387) );
  AOI22_X1 U20582 ( .A1(n17422), .A2(n17388), .B1(n17387), .B2(n17414), .ZN(
        P3_U2695) );
  AOI21_X1 U20583 ( .B1(n17390), .B2(n17389), .A(n17422), .ZN(n17391) );
  INV_X1 U20584 ( .A(n17391), .ZN(n17392) );
  OAI22_X1 U20585 ( .A1(n17393), .A2(n17392), .B1(n21122), .B2(n17414), .ZN(
        P3_U2696) );
  INV_X1 U20586 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n21138) );
  INV_X1 U20587 ( .A(n17426), .ZN(n17394) );
  NAND2_X1 U20588 ( .A1(n17395), .A2(n17394), .ZN(n17417) );
  INV_X1 U20589 ( .A(n17417), .ZN(n17410) );
  NAND2_X1 U20590 ( .A1(n17396), .A2(n17410), .ZN(n17406) );
  NOR2_X1 U20591 ( .A1(n21138), .A2(n17406), .ZN(n17409) );
  NOR2_X1 U20592 ( .A1(n17422), .A2(n17397), .ZN(n17402) );
  OAI222_X1 U20593 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17409), .C1(n17402), .C2(n17398), 
        .ZN(n17399) );
  OAI21_X1 U20594 ( .B1(n17400), .B2(n17414), .A(n17399), .ZN(P3_U2697) );
  INV_X1 U20595 ( .A(n17401), .ZN(n17403) );
  OAI21_X1 U20596 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17403), .A(n17402), .ZN(
        n17404) );
  OAI21_X1 U20597 ( .B1(n17414), .B2(n17405), .A(n17404), .ZN(P3_U2698) );
  INV_X1 U20598 ( .A(n17406), .ZN(n17413) );
  AOI21_X1 U20599 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17414), .A(n17413), .ZN(
        n17408) );
  OAI22_X1 U20600 ( .A1(n17409), .A2(n17408), .B1(n17407), .B2(n17414), .ZN(
        P3_U2699) );
  AOI22_X1 U20601 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17414), .B1(
        P3_EBX_REG_2__SCAN_IN), .B2(n17410), .ZN(n17412) );
  OAI22_X1 U20602 ( .A1(n17413), .A2(n17412), .B1(n17411), .B2(n17414), .ZN(
        P3_U2700) );
  NAND3_X1 U20603 ( .A1(n17417), .A2(P3_EBX_REG_2__SCAN_IN), .A3(n17414), .ZN(
        n17415) );
  OAI221_X1 U20604 ( .B1(n17417), .B2(P3_EBX_REG_2__SCAN_IN), .C1(n17414), 
        .C2(n17416), .A(n17415), .ZN(P3_U2701) );
  INV_X1 U20605 ( .A(n17418), .ZN(n17421) );
  INV_X1 U20606 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17419) );
  OAI222_X1 U20607 ( .A1(n17421), .A2(n17426), .B1(n17420), .B2(n17424), .C1(
        n17419), .C2(n17414), .ZN(P3_U2702) );
  NAND2_X1 U20608 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17422), .ZN(
        n17423) );
  OAI221_X1 U20609 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17426), .C1(n17425), 
        .C2(n17424), .A(n17423), .ZN(P3_U2703) );
  INV_X1 U20610 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17585) );
  INV_X1 U20611 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17588) );
  NAND4_X1 U20612 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_1__SCAN_IN), .ZN(n17428) );
  INV_X1 U20613 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17620) );
  NOR2_X2 U20614 ( .A1(n17549), .A2(n17620), .ZN(n17543) );
  INV_X1 U20615 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17611) );
  INV_X1 U20616 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17613) );
  INV_X1 U20617 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17681) );
  INV_X1 U20618 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17616) );
  NOR4_X1 U20619 ( .A1(n17611), .A2(n17613), .A3(n17681), .A4(n17616), .ZN(
        n17521) );
  AND2_X1 U20620 ( .A1(n17521), .A2(n10103), .ZN(n17430) );
  INV_X1 U20621 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17694) );
  INV_X1 U20622 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17603) );
  INV_X1 U20623 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17597) );
  NOR2_X1 U20624 ( .A1(n17603), .A2(n17597), .ZN(n17431) );
  NAND4_X1 U20625 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n17431), .ZN(n17477) );
  INV_X1 U20626 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17595) );
  NAND2_X1 U20627 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17473), .ZN(n17472) );
  NOR2_X2 U20628 ( .A1(n17472), .A2(n17478), .ZN(n17468) );
  NAND2_X1 U20629 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17446), .ZN(n17441) );
  NAND2_X1 U20630 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17437), .ZN(n17436) );
  NAND2_X1 U20631 ( .A1(n17432), .A2(n17544), .ZN(n17480) );
  OAI22_X1 U20632 ( .A1(n17544), .A2(n17437), .B1(P3_EAX_REG_30__SCAN_IN), 
        .B2(n17479), .ZN(n17433) );
  AOI22_X1 U20633 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17510), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17433), .ZN(n17434) );
  OAI21_X1 U20634 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17436), .A(n17434), .ZN(
        P3_U2704) );
  NAND2_X1 U20635 ( .A1(n17435), .A2(n17544), .ZN(n17504) );
  AOI22_X1 U20636 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17511), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17510), .ZN(n17439) );
  OAI211_X1 U20637 ( .C1(n17437), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17565), .B(
        n17436), .ZN(n17438) );
  OAI211_X1 U20638 ( .C1(n17440), .C2(n17568), .A(n17439), .B(n17438), .ZN(
        P3_U2705) );
  AOI22_X1 U20639 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17511), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17510), .ZN(n17443) );
  OAI211_X1 U20640 ( .C1(n17446), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17565), .B(
        n17441), .ZN(n17442) );
  OAI211_X1 U20641 ( .C1(n17568), .C2(n17444), .A(n17443), .B(n17442), .ZN(
        P3_U2706) );
  INV_X1 U20642 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18395) );
  AOI22_X1 U20643 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17511), .B1(n17445), .B2(
        n17573), .ZN(n17449) );
  AOI211_X1 U20644 ( .C1(n17585), .C2(n17453), .A(n17446), .B(n17544), .ZN(
        n17447) );
  INV_X1 U20645 ( .A(n17447), .ZN(n17448) );
  OAI211_X1 U20646 ( .C1(n17480), .C2(n18395), .A(n17449), .B(n17448), .ZN(
        P3_U2707) );
  OAI21_X1 U20647 ( .B1(n17452), .B2(n17451), .A(n17450), .ZN(n17456) );
  AOI22_X1 U20648 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17511), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17510), .ZN(n17455) );
  OAI211_X1 U20649 ( .C1(n17457), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17565), .B(
        n17453), .ZN(n17454) );
  OAI211_X1 U20650 ( .C1(n17568), .C2(n17456), .A(n17455), .B(n17454), .ZN(
        P3_U2708) );
  AOI22_X1 U20651 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17511), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17510), .ZN(n17460) );
  AOI211_X1 U20652 ( .C1(n17588), .C2(n17462), .A(n17457), .B(n17544), .ZN(
        n17458) );
  INV_X1 U20653 ( .A(n17458), .ZN(n17459) );
  OAI211_X1 U20654 ( .C1(n17568), .C2(n17461), .A(n17460), .B(n17459), .ZN(
        P3_U2709) );
  AOI22_X1 U20655 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17511), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17510), .ZN(n17464) );
  OAI211_X1 U20656 ( .C1(n17466), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17565), .B(
        n17462), .ZN(n17463) );
  OAI211_X1 U20657 ( .C1(n17568), .C2(n17465), .A(n17464), .B(n17463), .ZN(
        P3_U2710) );
  AOI22_X1 U20658 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17511), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17510), .ZN(n17470) );
  INV_X1 U20659 ( .A(n17466), .ZN(n17467) );
  OAI211_X1 U20660 ( .C1(n17468), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17565), .B(
        n17467), .ZN(n17469) );
  OAI211_X1 U20661 ( .C1(n17568), .C2(n17471), .A(n17470), .B(n17469), .ZN(
        P3_U2711) );
  AOI22_X1 U20662 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17511), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17510), .ZN(n17475) );
  OAI211_X1 U20663 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17473), .A(n17565), .B(
        n17472), .ZN(n17474) );
  OAI211_X1 U20664 ( .C1(n17476), .C2(n17568), .A(n17475), .B(n17474), .ZN(
        P3_U2712) );
  NOR3_X1 U20665 ( .A1(n17478), .A2(n17512), .A3(n17477), .ZN(n17484) );
  INV_X1 U20666 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17599) );
  INV_X1 U20667 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17645) );
  NAND2_X1 U20668 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17500), .ZN(n17496) );
  NOR2_X1 U20669 ( .A1(n17599), .A2(n17496), .ZN(n17490) );
  OR2_X1 U20670 ( .A1(n17544), .A2(n17490), .ZN(n17489) );
  OAI21_X1 U20671 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17479), .A(n17489), .ZN(
        n17483) );
  OAI22_X1 U20672 ( .A1(n17481), .A2(n17568), .B1(n14504), .B2(n17480), .ZN(
        n17482) );
  AOI221_X1 U20673 ( .B1(n17484), .B2(n17595), .C1(n17483), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n17482), .ZN(n17485) );
  OAI21_X1 U20674 ( .B1(n18403), .B2(n17504), .A(n17485), .ZN(P3_U2713) );
  AOI22_X1 U20675 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17510), .B1(n17573), .B2(
        n17486), .ZN(n17488) );
  AOI22_X1 U20676 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17511), .B1(n17490), .B2(
        n17597), .ZN(n17487) );
  OAI211_X1 U20677 ( .C1(n17597), .C2(n17489), .A(n17488), .B(n17487), .ZN(
        P3_U2714) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17511), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17510), .ZN(n17493) );
  AOI211_X1 U20679 ( .C1(n17599), .C2(n17496), .A(n17490), .B(n17544), .ZN(
        n17491) );
  INV_X1 U20680 ( .A(n17491), .ZN(n17492) );
  OAI211_X1 U20681 ( .C1(n17494), .C2(n17568), .A(n17493), .B(n17492), .ZN(
        P3_U2715) );
  AOI22_X1 U20682 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n17510), .B1(n17573), .B2(
        n17495), .ZN(n17498) );
  OAI211_X1 U20683 ( .C1(n17500), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17565), .B(
        n17496), .ZN(n17497) );
  OAI211_X1 U20684 ( .C1(n17504), .C2(n18390), .A(n17498), .B(n17497), .ZN(
        P3_U2716) );
  INV_X1 U20685 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18385) );
  AOI22_X1 U20686 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17510), .B1(n17573), .B2(
        n17499), .ZN(n17503) );
  AOI211_X1 U20687 ( .C1(n17603), .C2(n17505), .A(n17500), .B(n17544), .ZN(
        n17501) );
  INV_X1 U20688 ( .A(n17501), .ZN(n17502) );
  OAI211_X1 U20689 ( .C1(n17504), .C2(n18385), .A(n17503), .B(n17502), .ZN(
        P3_U2717) );
  AOI22_X1 U20690 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17511), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17510), .ZN(n17508) );
  INV_X1 U20691 ( .A(n17512), .ZN(n17506) );
  OAI211_X1 U20692 ( .C1(n17506), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17565), .B(
        n17505), .ZN(n17507) );
  OAI211_X1 U20693 ( .C1(n17509), .C2(n17568), .A(n17508), .B(n17507), .ZN(
        P3_U2718) );
  AOI22_X1 U20694 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17511), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17510), .ZN(n17514) );
  OAI211_X1 U20695 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17516), .A(n17565), .B(
        n17512), .ZN(n17513) );
  OAI211_X1 U20696 ( .C1(n17515), .C2(n17568), .A(n17514), .B(n17513), .ZN(
        P3_U2719) );
  AOI211_X1 U20697 ( .C1(n17694), .C2(n17520), .A(n17544), .B(n17516), .ZN(
        n17517) );
  AOI21_X1 U20698 ( .B1(n17574), .B2(BUF2_REG_15__SCAN_IN), .A(n17517), .ZN(
        n17518) );
  OAI21_X1 U20699 ( .B1(n17519), .B2(n17568), .A(n17518), .ZN(P3_U2720) );
  INV_X1 U20700 ( .A(n17520), .ZN(n17525) );
  NAND3_X1 U20701 ( .A1(n18410), .A2(P3_EAX_REG_9__SCAN_IN), .A3(n17543), .ZN(
        n17538) );
  AND2_X1 U20702 ( .A1(n17521), .A2(n17542), .ZN(n17527) );
  AOI21_X1 U20703 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17565), .A(n17527), .ZN(
        n17524) );
  AOI22_X1 U20704 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17574), .B1(n17573), .B2(
        n17522), .ZN(n17523) );
  OAI21_X1 U20705 ( .B1(n17525), .B2(n17524), .A(n17523), .ZN(P3_U2721) );
  NAND2_X1 U20706 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17542), .ZN(n17535) );
  NOR2_X1 U20707 ( .A1(n17681), .A2(n17535), .ZN(n17529) );
  AND2_X1 U20708 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17529), .ZN(n17532) );
  AOI21_X1 U20709 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17565), .A(n17532), .ZN(
        n17528) );
  OAI222_X1 U20710 ( .A1(n17571), .A2(n17687), .B1(n17528), .B2(n17527), .C1(
        n17568), .C2(n17526), .ZN(P3_U2722) );
  INV_X1 U20711 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17683) );
  AOI21_X1 U20712 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17565), .A(n17529), .ZN(
        n17531) );
  OAI222_X1 U20713 ( .A1(n17571), .A2(n17683), .B1(n17532), .B2(n17531), .C1(
        n17568), .C2(n17530), .ZN(P3_U2723) );
  NAND2_X1 U20714 ( .A1(n17565), .A2(n17535), .ZN(n17539) );
  AOI22_X1 U20715 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17574), .B1(n17573), .B2(
        n17533), .ZN(n17534) );
  OAI221_X1 U20716 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17535), .C1(n17681), 
        .C2(n17539), .A(n17534), .ZN(P3_U2724) );
  AOI22_X1 U20717 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17574), .B1(n17573), .B2(
        n17536), .ZN(n17537) );
  OAI221_X1 U20718 ( .B1(n17539), .B2(n17616), .C1(n17539), .C2(n17538), .A(
        n17537), .ZN(P3_U2725) );
  AOI22_X1 U20719 ( .A1(n18410), .A2(n17543), .B1(P3_EAX_REG_9__SCAN_IN), .B2(
        n17565), .ZN(n17541) );
  OAI222_X1 U20720 ( .A1(n17571), .A2(n17677), .B1(n17542), .B2(n17541), .C1(
        n17568), .C2(n17540), .ZN(P3_U2726) );
  INV_X1 U20721 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17675) );
  AOI211_X1 U20722 ( .C1(n17620), .C2(n17549), .A(n17544), .B(n17543), .ZN(
        n17545) );
  AOI21_X1 U20723 ( .B1(n17573), .B2(n17546), .A(n17545), .ZN(n17547) );
  OAI21_X1 U20724 ( .B1(n17675), .B2(n17571), .A(n17547), .ZN(P3_U2727) );
  AOI22_X1 U20725 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17574), .B1(n17573), .B2(
        n17548), .ZN(n17551) );
  OAI211_X1 U20726 ( .C1(P3_EAX_REG_7__SCAN_IN), .C2(n17554), .A(n17565), .B(
        n17549), .ZN(n17550) );
  NAND2_X1 U20727 ( .A1(n17551), .A2(n17550), .ZN(P3_U2728) );
  INV_X1 U20728 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17625) );
  INV_X1 U20729 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17632) );
  INV_X1 U20730 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17665) );
  NOR3_X1 U20731 ( .A1(n17632), .A2(n17665), .A3(n17577), .ZN(n17570) );
  AND2_X1 U20732 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17570), .ZN(n17564) );
  NAND2_X1 U20733 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17564), .ZN(n17555) );
  NOR2_X1 U20734 ( .A1(n17625), .A2(n17555), .ZN(n17558) );
  AOI21_X1 U20735 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17565), .A(n17558), .ZN(
        n17553) );
  OAI222_X1 U20736 ( .A1(n18403), .A2(n17571), .B1(n17554), .B2(n17553), .C1(
        n17568), .C2(n17552), .ZN(P3_U2729) );
  INV_X1 U20737 ( .A(n17555), .ZN(n17561) );
  AOI21_X1 U20738 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17565), .A(n17561), .ZN(
        n17557) );
  OAI222_X1 U20739 ( .A1(n18400), .A2(n17571), .B1(n17558), .B2(n17557), .C1(
        n17568), .C2(n17556), .ZN(P3_U2730) );
  INV_X1 U20740 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18394) );
  AOI21_X1 U20741 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17565), .A(n17564), .ZN(
        n17560) );
  OAI222_X1 U20742 ( .A1(n18394), .A2(n17571), .B1(n17561), .B2(n17560), .C1(
        n17568), .C2(n9718), .ZN(P3_U2731) );
  AOI21_X1 U20743 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17565), .A(n17570), .ZN(
        n17563) );
  OAI222_X1 U20744 ( .A1(n18390), .A2(n17571), .B1(n17564), .B2(n17563), .C1(
        n17568), .C2(n17562), .ZN(P3_U2732) );
  AOI22_X1 U20745 ( .A1(n17566), .A2(P3_EAX_REG_1__SCAN_IN), .B1(
        P3_EAX_REG_2__SCAN_IN), .B2(n17565), .ZN(n17569) );
  OAI222_X1 U20746 ( .A1(n18385), .A2(n17571), .B1(n17570), .B2(n17569), .C1(
        n17568), .C2(n17567), .ZN(P3_U2733) );
  AOI22_X1 U20747 ( .A1(n17574), .A2(BUF2_REG_1__SCAN_IN), .B1(n17573), .B2(
        n17572), .ZN(n17575) );
  OAI221_X1 U20748 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17577), .C1(n17665), 
        .C2(n17576), .A(n17575), .ZN(P3_U2734) );
  AND2_X1 U20749 ( .A1(P3_DATAO_REG_31__SCAN_IN), .A2(n17628), .ZN(P3_U2736)
         );
  INV_X1 U20750 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17662) );
  NAND2_X1 U20751 ( .A1(n17580), .A2(n17579), .ZN(n17606) );
  AOI22_X1 U20752 ( .A1(n19030), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17628), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17581) );
  OAI21_X1 U20753 ( .B1(n17662), .B2(n17606), .A(n17581), .ZN(P3_U2737) );
  INV_X1 U20754 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17583) );
  AOI22_X1 U20755 ( .A1(n18874), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17582) );
  OAI21_X1 U20756 ( .B1(n17583), .B2(n17606), .A(n17582), .ZN(P3_U2738) );
  AOI22_X1 U20757 ( .A1(n19030), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17628), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17584) );
  OAI21_X1 U20758 ( .B1(n17585), .B2(n17606), .A(n17584), .ZN(P3_U2739) );
  INV_X1 U20759 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17657) );
  AOI22_X1 U20760 ( .A1(n18874), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17628), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17586) );
  OAI21_X1 U20761 ( .B1(n17657), .B2(n17606), .A(n17586), .ZN(P3_U2740) );
  AOI22_X1 U20762 ( .A1(P3_DATAO_REG_26__SCAN_IN), .A2(n17634), .B1(n19030), 
        .B2(P3_UWORD_REG_10__SCAN_IN), .ZN(n17587) );
  OAI21_X1 U20763 ( .B1(n17588), .B2(n17606), .A(n17587), .ZN(P3_U2741) );
  INV_X1 U20764 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17590) );
  AOI22_X1 U20765 ( .A1(n18874), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17628), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17589) );
  OAI21_X1 U20766 ( .B1(n17590), .B2(n17606), .A(n17589), .ZN(P3_U2742) );
  INV_X1 U20767 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17592) );
  AOI22_X1 U20768 ( .A1(n18874), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17628), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17591) );
  OAI21_X1 U20769 ( .B1(n17592), .B2(n17606), .A(n17591), .ZN(P3_U2743) );
  INV_X1 U20770 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17652) );
  AOI22_X1 U20771 ( .A1(n18874), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17593) );
  OAI21_X1 U20772 ( .B1(n17652), .B2(n17606), .A(n17593), .ZN(P3_U2744) );
  AOI22_X1 U20773 ( .A1(n18874), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17628), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17594) );
  OAI21_X1 U20774 ( .B1(n17595), .B2(n17606), .A(n17594), .ZN(P3_U2745) );
  AOI22_X1 U20775 ( .A1(n18874), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17596) );
  OAI21_X1 U20776 ( .B1(n17597), .B2(n17606), .A(n17596), .ZN(P3_U2746) );
  AOI22_X1 U20777 ( .A1(n18874), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17598) );
  OAI21_X1 U20778 ( .B1(n17599), .B2(n17606), .A(n17598), .ZN(P3_U2747) );
  INV_X1 U20779 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17601) );
  AOI22_X1 U20780 ( .A1(n18874), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17600) );
  OAI21_X1 U20781 ( .B1(n17601), .B2(n17606), .A(n17600), .ZN(P3_U2748) );
  AOI22_X1 U20782 ( .A1(n18874), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17602) );
  OAI21_X1 U20783 ( .B1(n17603), .B2(n17606), .A(n17602), .ZN(P3_U2749) );
  AOI22_X1 U20784 ( .A1(n18874), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17604) );
  OAI21_X1 U20785 ( .B1(n17645), .B2(n17606), .A(n17604), .ZN(P3_U2750) );
  INV_X1 U20786 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17607) );
  AOI22_X1 U20787 ( .A1(P3_DATAO_REG_16__SCAN_IN), .A2(n17634), .B1(n19030), 
        .B2(P3_UWORD_REG_0__SCAN_IN), .ZN(n17605) );
  OAI21_X1 U20788 ( .B1(n17607), .B2(n17606), .A(n17605), .ZN(P3_U2751) );
  AOI22_X1 U20789 ( .A1(n18874), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17608) );
  OAI21_X1 U20790 ( .B1(n17694), .B2(n17636), .A(n17608), .ZN(P3_U2752) );
  INV_X1 U20791 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17689) );
  AOI22_X1 U20792 ( .A1(n18874), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17609) );
  OAI21_X1 U20793 ( .B1(n17689), .B2(n17636), .A(n17609), .ZN(P3_U2753) );
  AOI22_X1 U20794 ( .A1(n18874), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17610) );
  OAI21_X1 U20795 ( .B1(n17611), .B2(n17636), .A(n17610), .ZN(P3_U2754) );
  AOI22_X1 U20796 ( .A1(P3_LWORD_REG_12__SCAN_IN), .A2(n19030), .B1(n17634), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17612) );
  OAI21_X1 U20797 ( .B1(n17613), .B2(n17636), .A(n17612), .ZN(P3_U2755) );
  AOI22_X1 U20798 ( .A1(n18874), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17614) );
  OAI21_X1 U20799 ( .B1(n17681), .B2(n17636), .A(n17614), .ZN(P3_U2756) );
  AOI22_X1 U20800 ( .A1(n18874), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17615) );
  OAI21_X1 U20801 ( .B1(n17616), .B2(n17636), .A(n17615), .ZN(P3_U2757) );
  INV_X1 U20802 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17618) );
  AOI22_X1 U20803 ( .A1(P3_LWORD_REG_9__SCAN_IN), .A2(n19030), .B1(n17634), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17617) );
  OAI21_X1 U20804 ( .B1(n17618), .B2(n17636), .A(n17617), .ZN(P3_U2758) );
  AOI22_X1 U20805 ( .A1(n18874), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17628), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17619) );
  OAI21_X1 U20806 ( .B1(n17620), .B2(n17636), .A(n17619), .ZN(P3_U2759) );
  INV_X1 U20807 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17672) );
  AOI22_X1 U20808 ( .A1(n18874), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17621) );
  OAI21_X1 U20809 ( .B1(n17672), .B2(n17636), .A(n17621), .ZN(P3_U2760) );
  INV_X1 U20810 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17623) );
  AOI22_X1 U20811 ( .A1(n18874), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17628), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17622) );
  OAI21_X1 U20812 ( .B1(n17623), .B2(n17636), .A(n17622), .ZN(P3_U2761) );
  AOI22_X1 U20813 ( .A1(n18874), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17628), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17624) );
  OAI21_X1 U20814 ( .B1(n17625), .B2(n17636), .A(n17624), .ZN(P3_U2762) );
  INV_X1 U20815 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17627) );
  AOI22_X1 U20816 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(n17634), .B1(n19030), 
        .B2(P3_LWORD_REG_4__SCAN_IN), .ZN(n17626) );
  OAI21_X1 U20817 ( .B1(n17627), .B2(n17636), .A(n17626), .ZN(P3_U2763) );
  INV_X1 U20818 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17630) );
  AOI22_X1 U20819 ( .A1(n18874), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17628), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17629) );
  OAI21_X1 U20820 ( .B1(n17630), .B2(n17636), .A(n17629), .ZN(P3_U2764) );
  AOI22_X1 U20821 ( .A1(n18874), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17631) );
  OAI21_X1 U20822 ( .B1(n17632), .B2(n17636), .A(n17631), .ZN(P3_U2765) );
  AOI22_X1 U20823 ( .A1(n18874), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17633) );
  OAI21_X1 U20824 ( .B1(n17665), .B2(n17636), .A(n17633), .ZN(P3_U2766) );
  AOI22_X1 U20825 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(n17634), .B1(n19030), 
        .B2(P3_LWORD_REG_0__SCAN_IN), .ZN(n17635) );
  OAI21_X1 U20826 ( .B1(n17637), .B2(n17636), .A(n17635), .ZN(P3_U2767) );
  INV_X1 U20827 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U20828 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17684), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17690), .ZN(n17643) );
  OAI21_X1 U20829 ( .B1(n18373), .B2(n17686), .A(n17643), .ZN(P3_U2768) );
  INV_X1 U20830 ( .A(n17673), .ZN(n17693) );
  AOI22_X1 U20831 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17691), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17690), .ZN(n17644) );
  OAI21_X1 U20832 ( .B1(n17645), .B2(n17693), .A(n17644), .ZN(P3_U2769) );
  AOI22_X1 U20833 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17684), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17690), .ZN(n17646) );
  OAI21_X1 U20834 ( .B1(n18385), .B2(n17686), .A(n17646), .ZN(P3_U2770) );
  AOI22_X1 U20835 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17684), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17659), .ZN(n17647) );
  OAI21_X1 U20836 ( .B1(n18390), .B2(n17686), .A(n17647), .ZN(P3_U2771) );
  AOI22_X1 U20837 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17684), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17659), .ZN(n17648) );
  OAI21_X1 U20838 ( .B1(n18394), .B2(n17686), .A(n17648), .ZN(P3_U2772) );
  AOI22_X1 U20839 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17673), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17659), .ZN(n17649) );
  OAI21_X1 U20840 ( .B1(n18400), .B2(n17686), .A(n17649), .ZN(P3_U2773) );
  AOI22_X1 U20841 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17684), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17659), .ZN(n17650) );
  OAI21_X1 U20842 ( .B1(n18403), .B2(n17686), .A(n17650), .ZN(P3_U2774) );
  AOI22_X1 U20843 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17691), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17690), .ZN(n17651) );
  OAI21_X1 U20844 ( .B1(n17652), .B2(n17693), .A(n17651), .ZN(P3_U2775) );
  AOI22_X1 U20845 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17673), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17659), .ZN(n17653) );
  OAI21_X1 U20846 ( .B1(n17675), .B2(n17686), .A(n17653), .ZN(P3_U2776) );
  AOI22_X1 U20847 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17684), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17659), .ZN(n17654) );
  OAI21_X1 U20848 ( .B1(n17677), .B2(n17686), .A(n17654), .ZN(P3_U2777) );
  INV_X1 U20849 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17679) );
  AOI22_X1 U20850 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17684), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17659), .ZN(n17655) );
  OAI21_X1 U20851 ( .B1(n17679), .B2(n17686), .A(n17655), .ZN(P3_U2778) );
  AOI22_X1 U20852 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17691), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17659), .ZN(n17656) );
  OAI21_X1 U20853 ( .B1(n17657), .B2(n17693), .A(n17656), .ZN(P3_U2779) );
  AOI22_X1 U20854 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17684), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17659), .ZN(n17658) );
  OAI21_X1 U20855 ( .B1(n17683), .B2(n17686), .A(n17658), .ZN(P3_U2780) );
  AOI22_X1 U20856 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17684), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17659), .ZN(n17660) );
  OAI21_X1 U20857 ( .B1(n17687), .B2(n17686), .A(n17660), .ZN(P3_U2781) );
  AOI22_X1 U20858 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17691), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17690), .ZN(n17661) );
  OAI21_X1 U20859 ( .B1(n17662), .B2(n17693), .A(n17661), .ZN(P3_U2782) );
  AOI22_X1 U20860 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17684), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17690), .ZN(n17663) );
  OAI21_X1 U20861 ( .B1(n18373), .B2(n17686), .A(n17663), .ZN(P3_U2783) );
  AOI22_X1 U20862 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17691), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17690), .ZN(n17664) );
  OAI21_X1 U20863 ( .B1(n17665), .B2(n17693), .A(n17664), .ZN(P3_U2784) );
  AOI22_X1 U20864 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17684), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17690), .ZN(n17666) );
  OAI21_X1 U20865 ( .B1(n18385), .B2(n17686), .A(n17666), .ZN(P3_U2785) );
  AOI22_X1 U20866 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17673), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17690), .ZN(n17667) );
  OAI21_X1 U20867 ( .B1(n18390), .B2(n17686), .A(n17667), .ZN(P3_U2786) );
  AOI22_X1 U20868 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17684), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17690), .ZN(n17668) );
  OAI21_X1 U20869 ( .B1(n18394), .B2(n17686), .A(n17668), .ZN(P3_U2787) );
  AOI22_X1 U20870 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17673), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17690), .ZN(n17669) );
  OAI21_X1 U20871 ( .B1(n18400), .B2(n17686), .A(n17669), .ZN(P3_U2788) );
  AOI22_X1 U20872 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17684), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17690), .ZN(n17670) );
  OAI21_X1 U20873 ( .B1(n18403), .B2(n17686), .A(n17670), .ZN(P3_U2789) );
  AOI22_X1 U20874 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17691), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17690), .ZN(n17671) );
  OAI21_X1 U20875 ( .B1(n17672), .B2(n17693), .A(n17671), .ZN(P3_U2790) );
  AOI22_X1 U20876 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17673), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17690), .ZN(n17674) );
  OAI21_X1 U20877 ( .B1(n17675), .B2(n17686), .A(n17674), .ZN(P3_U2791) );
  AOI22_X1 U20878 ( .A1(P3_LWORD_REG_9__SCAN_IN), .A2(n17690), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17684), .ZN(n17676) );
  OAI21_X1 U20879 ( .B1(n17677), .B2(n17686), .A(n17676), .ZN(P3_U2792) );
  AOI22_X1 U20880 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17684), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17690), .ZN(n17678) );
  OAI21_X1 U20881 ( .B1(n17679), .B2(n17686), .A(n17678), .ZN(P3_U2793) );
  AOI22_X1 U20882 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17691), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17690), .ZN(n17680) );
  OAI21_X1 U20883 ( .B1(n17681), .B2(n17693), .A(n17680), .ZN(P3_U2794) );
  AOI22_X1 U20884 ( .A1(P3_LWORD_REG_12__SCAN_IN), .A2(n17690), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n17684), .ZN(n17682) );
  OAI21_X1 U20885 ( .B1(n17683), .B2(n17686), .A(n17682), .ZN(P3_U2795) );
  AOI22_X1 U20886 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17684), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17690), .ZN(n17685) );
  OAI21_X1 U20887 ( .B1(n17687), .B2(n17686), .A(n17685), .ZN(P3_U2796) );
  AOI22_X1 U20888 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17691), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17690), .ZN(n17688) );
  OAI21_X1 U20889 ( .B1(n17689), .B2(n17693), .A(n17688), .ZN(P3_U2797) );
  AOI22_X1 U20890 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17691), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17690), .ZN(n17692) );
  OAI21_X1 U20891 ( .B1(n17694), .B2(n17693), .A(n17692), .ZN(P3_U2798) );
  INV_X1 U20892 ( .A(n18054), .ZN(n18029) );
  AOI21_X1 U20893 ( .B1(n17695), .B2(n17895), .A(n18029), .ZN(n17696) );
  INV_X1 U20894 ( .A(n17696), .ZN(n17697) );
  AOI21_X1 U20895 ( .B1(n17851), .B2(n17709), .A(n17697), .ZN(n17727) );
  OAI21_X1 U20896 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17837), .A(
        n17727), .ZN(n17719) );
  AOI22_X1 U20897 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17719), .B1(
        n17914), .B2(n17698), .ZN(n17714) );
  NOR2_X1 U20898 ( .A1(n18047), .A2(n17968), .ZN(n17805) );
  OAI22_X1 U20899 ( .A1(n17700), .A2(n18058), .B1(n17699), .B2(n17887), .ZN(
        n17734) );
  NOR2_X1 U20900 ( .A1(n18059), .A2(n17734), .ZN(n17702) );
  NOR3_X1 U20901 ( .A1(n17805), .A2(n17702), .A3(n17701), .ZN(n17707) );
  AOI211_X1 U20902 ( .C1(n9792), .C2(n17708), .A(n17707), .B(n10105), .ZN(
        n17713) );
  NAND2_X1 U20903 ( .A1(n18348), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17712) );
  NOR2_X1 U20904 ( .A1(n17813), .A2(n17709), .ZN(n17721) );
  OAI211_X1 U20905 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17721), .B(n17710), .ZN(n17711) );
  NAND4_X1 U20906 ( .A1(n17714), .A2(n17713), .A3(n17712), .A4(n17711), .ZN(
        P3_U2802) );
  NOR2_X1 U20907 ( .A1(n16561), .A2(n17715), .ZN(n17716) );
  XOR2_X1 U20908 ( .A(n17716), .B(n17958), .Z(n18071) );
  OAI22_X1 U20909 ( .A1(n18358), .A2(n18962), .B1(n17864), .B2(n17717), .ZN(
        n17718) );
  AOI221_X1 U20910 ( .B1(n17721), .B2(n17720), .C1(n17719), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17718), .ZN(n17723) );
  AOI22_X1 U20911 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17734), .B1(
        n9792), .B2(n18059), .ZN(n17722) );
  OAI211_X1 U20912 ( .C1(n18071), .C2(n17971), .A(n17723), .B(n17722), .ZN(
        P3_U2803) );
  INV_X1 U20913 ( .A(n17724), .ZN(n17758) );
  INV_X1 U20914 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21254) );
  NAND3_X1 U20915 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n21254), .ZN(n18072) );
  INV_X1 U20916 ( .A(n17837), .ZN(n17729) );
  AOI21_X1 U20917 ( .B1(n18753), .B2(n17725), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17726) );
  NAND2_X1 U20918 ( .A1(n18348), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18079) );
  OAI21_X1 U20919 ( .B1(n17727), .B2(n17726), .A(n18079), .ZN(n17728) );
  AOI221_X1 U20920 ( .B1(n17914), .B2(n17730), .C1(n17729), .C2(n17730), .A(
        n17728), .ZN(n17736) );
  AOI21_X1 U20921 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17732), .A(
        n17731), .ZN(n18075) );
  INV_X1 U20922 ( .A(n18075), .ZN(n17733) );
  AOI22_X1 U20923 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17734), .B1(
        n17953), .B2(n17733), .ZN(n17735) );
  OAI211_X1 U20924 ( .C1(n17758), .C2(n18072), .A(n17736), .B(n17735), .ZN(
        P3_U2804) );
  XOR2_X1 U20925 ( .A(n21220), .B(n17737), .Z(n18091) );
  AND2_X1 U20926 ( .A1(n17739), .A2(n18753), .ZN(n17764) );
  AOI211_X1 U20927 ( .C1(n17895), .C2(n17738), .A(n17764), .B(n18029), .ZN(
        n17768) );
  OAI21_X1 U20928 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17837), .A(
        n17768), .ZN(n17753) );
  NOR2_X1 U20929 ( .A1(n17813), .A2(n17739), .ZN(n17752) );
  OAI211_X1 U20930 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17752), .B(n17740), .ZN(n17741) );
  NAND2_X1 U20931 ( .A1(n18348), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18088) );
  OAI211_X1 U20932 ( .C1(n17864), .C2(n17742), .A(n17741), .B(n18088), .ZN(
        n17747) );
  XOR2_X1 U20933 ( .A(n17743), .B(n21220), .Z(n18095) );
  OAI21_X1 U20934 ( .B1(n17847), .B2(n9775), .A(n17744), .ZN(n17745) );
  XOR2_X1 U20935 ( .A(n17745), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18090) );
  OAI22_X1 U20936 ( .A1(n18058), .A2(n18095), .B1(n17971), .B2(n18090), .ZN(
        n17746) );
  AOI211_X1 U20937 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17753), .A(
        n17747), .B(n17746), .ZN(n17748) );
  OAI21_X1 U20938 ( .B1(n17887), .B2(n18091), .A(n17748), .ZN(P3_U2805) );
  AOI22_X1 U20939 ( .A1(n18047), .A2(n18097), .B1(n17968), .B2(n18096), .ZN(
        n17775) );
  OAI21_X1 U20940 ( .B1(n9818), .B2(n18082), .A(n17749), .ZN(n18105) );
  INV_X1 U20941 ( .A(n17750), .ZN(n17755) );
  AOI22_X1 U20942 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17753), .B1(
        n17752), .B2(n17751), .ZN(n17754) );
  NAND2_X1 U20943 ( .A1(n18348), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18106) );
  OAI211_X1 U20944 ( .C1(n17755), .C2(n17864), .A(n17754), .B(n18106), .ZN(
        n17756) );
  AOI21_X1 U20945 ( .B1(n17953), .B2(n18105), .A(n17756), .ZN(n17757) );
  OAI221_X1 U20946 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17758), 
        .C1(n18082), .C2(n17775), .A(n17757), .ZN(P3_U2806) );
  INV_X1 U20947 ( .A(n13192), .ZN(n17806) );
  AOI21_X1 U20948 ( .B1(n18109), .B2(n17825), .A(n17783), .ZN(n17759) );
  AOI211_X1 U20949 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17847), .A(
        n17806), .B(n17759), .ZN(n17760) );
  XOR2_X1 U20950 ( .A(n17760), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n18110) );
  AOI22_X1 U20951 ( .A1(n18348), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17914), 
        .B2(n17761), .ZN(n17766) );
  NOR2_X1 U20952 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17837), .ZN(
        n17763) );
  OAI221_X1 U20953 ( .B1(n17764), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C1(
        n17764), .C2(n17763), .A(n17762), .ZN(n17765) );
  OAI211_X1 U20954 ( .C1(n17768), .C2(n17767), .A(n17766), .B(n17765), .ZN(
        n17769) );
  AOI21_X1 U20955 ( .B1(n17953), .B2(n18110), .A(n17769), .ZN(n17774) );
  INV_X1 U20956 ( .A(n17869), .ZN(n18115) );
  NAND2_X1 U20957 ( .A1(n18047), .A2(n18097), .ZN(n17771) );
  NAND2_X1 U20958 ( .A1(n17968), .A2(n18096), .ZN(n17770) );
  OAI22_X1 U20959 ( .A1(n18115), .A2(n17771), .B1(n18190), .B2(n17770), .ZN(
        n17772) );
  NAND3_X1 U20960 ( .A1(n18109), .A2(n18158), .A3(n17772), .ZN(n17773) );
  OAI211_X1 U20961 ( .C1(n17775), .C2(n18113), .A(n17774), .B(n17773), .ZN(
        P3_U2807) );
  OAI21_X1 U20962 ( .B1(n17776), .B2(n18891), .A(n18054), .ZN(n17777) );
  AOI21_X1 U20963 ( .B1(n17851), .B2(n17779), .A(n17777), .ZN(n17802) );
  OAI21_X1 U20964 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17837), .A(
        n17802), .ZN(n17791) );
  AOI22_X1 U20965 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17791), .B1(
        n17914), .B2(n17778), .ZN(n17788) );
  NOR2_X1 U20966 ( .A1(n17813), .A2(n17779), .ZN(n17793) );
  AOI21_X1 U20967 ( .B1(n21288), .B2(n17792), .A(n17780), .ZN(n17781) );
  AOI22_X1 U20968 ( .A1(n18348), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17793), 
        .B2(n17781), .ZN(n17787) );
  NOR2_X1 U20969 ( .A1(n17832), .A2(n17782), .ZN(n18118) );
  AOI22_X1 U20970 ( .A1(n18047), .A2(n18115), .B1(n17968), .B2(n18190), .ZN(
        n17861) );
  OAI21_X1 U20971 ( .B1(n17805), .B2(n18118), .A(n17861), .ZN(n17798) );
  OAI221_X1 U20972 ( .B1(n17783), .B2(n18122), .C1(n17783), .C2(n17794), .A(
        n13192), .ZN(n17784) );
  XOR2_X1 U20973 ( .A(n18129), .B(n17784), .Z(n18126) );
  AOI22_X1 U20974 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17798), .B1(
        n17953), .B2(n18126), .ZN(n17786) );
  NAND3_X1 U20975 ( .A1(n17833), .A2(n18118), .A3(n18129), .ZN(n17785) );
  NAND4_X1 U20976 ( .A1(n17788), .A2(n17787), .A3(n17786), .A4(n17785), .ZN(
        P3_U2808) );
  OR2_X1 U20977 ( .A1(n17796), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18142) );
  NOR2_X1 U20978 ( .A1(n17832), .A2(n18131), .ZN(n18133) );
  NAND2_X1 U20979 ( .A1(n17833), .A2(n18133), .ZN(n17823) );
  OAI22_X1 U20980 ( .A1(n18358), .A2(n18950), .B1(n17864), .B2(n17789), .ZN(
        n17790) );
  AOI221_X1 U20981 ( .B1(n17793), .B2(n17792), .C1(n17791), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17790), .ZN(n17800) );
  NAND3_X1 U20982 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17958), .A3(
        n17794), .ZN(n17818) );
  OAI22_X1 U20983 ( .A1(n17796), .A2(n17818), .B1(n17795), .B2(n17825), .ZN(
        n17797) );
  XOR2_X1 U20984 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17797), .Z(
        n18132) );
  AOI22_X1 U20985 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17798), .B1(
        n17953), .B2(n18132), .ZN(n17799) );
  OAI211_X1 U20986 ( .C1(n18142), .C2(n17823), .A(n17800), .B(n17799), .ZN(
        P3_U2809) );
  NAND2_X1 U20987 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21224), .ZN(
        n18149) );
  AOI21_X1 U20988 ( .B1(n9835), .B2(n18753), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17801) );
  INV_X1 U20989 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18948) );
  OAI22_X1 U20990 ( .A1(n17802), .A2(n17801), .B1(n18358), .B2(n18948), .ZN(
        n17803) );
  AOI221_X1 U20991 ( .B1(n17914), .B2(n17804), .C1(n17729), .C2(n17804), .A(
        n17803), .ZN(n17810) );
  AND2_X1 U20992 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18133), .ZN(
        n18145) );
  OAI21_X1 U20993 ( .B1(n17805), .B2(n18145), .A(n17861), .ZN(n17820) );
  INV_X1 U20994 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17807) );
  AOI221_X1 U20995 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17818), 
        .C1(n17807), .C2(n17824), .A(n17806), .ZN(n17808) );
  XOR2_X1 U20996 ( .A(n17808), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n18143) );
  AOI22_X1 U20997 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17820), .B1(
        n17953), .B2(n18143), .ZN(n17809) );
  OAI211_X1 U20998 ( .C1(n17823), .C2(n18149), .A(n17810), .B(n17809), .ZN(
        P3_U2810) );
  AOI21_X1 U20999 ( .B1(n17851), .B2(n17812), .A(n18029), .ZN(n17846) );
  OAI21_X1 U21000 ( .B1(n17811), .B2(n18891), .A(n17846), .ZN(n17829) );
  NOR2_X1 U21001 ( .A1(n17813), .A2(n17812), .ZN(n17831) );
  OAI211_X1 U21002 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17831), .B(n17814), .ZN(n17815) );
  NAND2_X1 U21003 ( .A1(n18348), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18152) );
  OAI211_X1 U21004 ( .C1(n17864), .C2(n17816), .A(n17815), .B(n18152), .ZN(
        n17817) );
  AOI21_X1 U21005 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17829), .A(
        n17817), .ZN(n17822) );
  OAI21_X1 U21006 ( .B1(n17824), .B2(n17825), .A(n17818), .ZN(n17819) );
  XOR2_X1 U21007 ( .A(n17819), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n18150) );
  AOI22_X1 U21008 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17820), .B1(
        n17953), .B2(n18150), .ZN(n17821) );
  OAI211_X1 U21009 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17823), .A(
        n17822), .B(n17821), .ZN(P3_U2811) );
  OAI21_X1 U21010 ( .B1(n17847), .B2(n18131), .A(n17824), .ZN(n17826) );
  XNOR2_X1 U21011 ( .A(n17826), .B(n17825), .ZN(n18169) );
  OAI22_X1 U21012 ( .A1(n18358), .A2(n18944), .B1(n17864), .B2(n17827), .ZN(
        n17828) );
  AOI221_X1 U21013 ( .B1(n17831), .B2(n17830), .C1(n17829), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17828), .ZN(n17835) );
  OAI21_X1 U21014 ( .B1(n18158), .B2(n17862), .A(n17861), .ZN(n17843) );
  NOR2_X1 U21015 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17832), .ZN(
        n18165) );
  AOI22_X1 U21016 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17843), .B1(
        n17833), .B2(n18165), .ZN(n17834) );
  OAI211_X1 U21017 ( .C1(n17971), .C2(n18169), .A(n17835), .B(n17834), .ZN(
        P3_U2812) );
  AOI21_X1 U21018 ( .B1(n17836), .B2(n18753), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17845) );
  OAI21_X1 U21019 ( .B1(n18182), .B2(n17862), .A(n18171), .ZN(n17842) );
  AOI21_X1 U21020 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17839), .A(
        n17838), .ZN(n18175) );
  OAI22_X1 U21021 ( .A1(n18034), .A2(n17840), .B1(n18175), .B2(n17971), .ZN(
        n17841) );
  AOI21_X1 U21022 ( .B1(n17843), .B2(n17842), .A(n17841), .ZN(n17844) );
  NAND2_X1 U21023 ( .A1(n18348), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18173) );
  OAI211_X1 U21024 ( .C1(n17846), .C2(n17845), .A(n17844), .B(n18173), .ZN(
        P3_U2813) );
  NOR2_X1 U21025 ( .A1(n17847), .A2(n17927), .ZN(n17932) );
  INV_X1 U21026 ( .A(n17932), .ZN(n17945) );
  OAI22_X1 U21027 ( .A1(n17958), .A2(n17848), .B1(n18163), .B2(n17945), .ZN(
        n17849) );
  XOR2_X1 U21028 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17849), .Z(
        n18184) );
  AOI21_X1 U21029 ( .B1(n17851), .B2(n17850), .A(n18029), .ZN(n17881) );
  OAI21_X1 U21030 ( .B1(n17852), .B2(n18891), .A(n17881), .ZN(n17866) );
  AOI22_X1 U21031 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17866), .B1(
        n17914), .B2(n17853), .ZN(n17858) );
  NAND2_X1 U21032 ( .A1(n17891), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17855) );
  NAND2_X1 U21033 ( .A1(n17892), .A2(n17854), .ZN(n17911) );
  NOR2_X1 U21034 ( .A1(n17855), .A2(n17911), .ZN(n17868) );
  OAI211_X1 U21035 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17868), .B(n17856), .ZN(n17857) );
  OAI211_X1 U21036 ( .C1(n18940), .C2(n18358), .A(n17858), .B(n17857), .ZN(
        n17859) );
  AOI21_X1 U21037 ( .B1(n17953), .B2(n18184), .A(n17859), .ZN(n17860) );
  OAI221_X1 U21038 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17862), 
        .C1(n18182), .C2(n17861), .A(n17860), .ZN(P3_U2814) );
  AOI21_X1 U21039 ( .B1(n18180), .B2(n18240), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18193) );
  NAND2_X1 U21040 ( .A1(n17968), .A2(n18190), .ZN(n17877) );
  INV_X1 U21041 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17867) );
  OAI22_X1 U21042 ( .A1(n18358), .A2(n18938), .B1(n17864), .B2(n17863), .ZN(
        n17865) );
  AOI221_X1 U21043 ( .B1(n17868), .B2(n17867), .C1(n17866), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17865), .ZN(n17876) );
  INV_X1 U21044 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17874) );
  NOR2_X1 U21045 ( .A1(n18245), .A2(n18204), .ZN(n17885) );
  NAND2_X1 U21046 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17885), .ZN(
        n17884) );
  AOI21_X1 U21047 ( .B1(n17874), .B2(n17884), .A(n17869), .ZN(n18187) );
  NAND3_X1 U21048 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n18240), .ZN(n17871) );
  OAI21_X1 U21049 ( .B1(n18228), .B2(n17871), .A(n17870), .ZN(n17872) );
  OAI221_X1 U21050 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18203), 
        .C1(n18227), .C2(n17958), .A(n17872), .ZN(n17873) );
  XOR2_X1 U21051 ( .A(n17874), .B(n17873), .Z(n18196) );
  AOI22_X1 U21052 ( .A1(n18047), .A2(n18187), .B1(n17953), .B2(n18196), .ZN(
        n17875) );
  OAI211_X1 U21053 ( .C1(n18193), .C2(n17877), .A(n17876), .B(n17875), .ZN(
        P3_U2815) );
  INV_X1 U21054 ( .A(n18204), .ZN(n17879) );
  AOI21_X1 U21055 ( .B1(n17932), .B2(n17879), .A(n17878), .ZN(n17880) );
  XOR2_X1 U21056 ( .A(n17880), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18215) );
  AND2_X1 U21057 ( .A1(n17892), .A2(n18753), .ZN(n17925) );
  AOI21_X1 U21058 ( .B1(n17891), .B2(n17925), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17882) );
  OAI22_X1 U21059 ( .A1(n18034), .A2(n17883), .B1(n17882), .B2(n17881), .ZN(
        n17889) );
  OAI21_X1 U21060 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17885), .A(
        n17884), .ZN(n18211) );
  NAND2_X1 U21061 ( .A1(n18202), .A2(n18240), .ZN(n17902) );
  INV_X1 U21062 ( .A(n17902), .ZN(n18219) );
  NAND2_X1 U21063 ( .A1(n18180), .A2(n18240), .ZN(n17886) );
  OAI221_X1 U21064 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18219), .A(n17886), .ZN(
        n18209) );
  OAI22_X1 U21065 ( .A1(n18058), .A2(n18211), .B1(n17887), .B2(n18209), .ZN(
        n17888) );
  AOI211_X1 U21066 ( .C1(n18348), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17889), 
        .B(n17888), .ZN(n17890) );
  OAI21_X1 U21067 ( .B1(n18215), .B2(n17971), .A(n17890), .ZN(P3_U2816) );
  NAND2_X1 U21068 ( .A1(n18202), .A2(n17904), .ZN(n18226) );
  AOI211_X1 U21069 ( .C1(n17910), .C2(n17896), .A(n17891), .B(n17911), .ZN(
        n17898) );
  OAI21_X1 U21070 ( .B1(n17892), .B2(n18017), .A(n18054), .ZN(n17893) );
  AOI21_X1 U21071 ( .B1(n17895), .B2(n17894), .A(n17893), .ZN(n17909) );
  OAI22_X1 U21072 ( .A1(n17909), .A2(n17896), .B1(n18358), .B2(n18934), .ZN(
        n17897) );
  AOI211_X1 U21073 ( .C1(n17914), .C2(n17899), .A(n17898), .B(n17897), .ZN(
        n17907) );
  NAND2_X1 U21074 ( .A1(n18202), .A2(n9878), .ZN(n18222) );
  AOI22_X1 U21075 ( .A1(n17902), .A2(n17968), .B1(n18222), .B2(n18047), .ZN(
        n17900) );
  INV_X1 U21076 ( .A(n17900), .ZN(n17915) );
  OAI21_X1 U21077 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17958), .A(
        n17902), .ZN(n17903) );
  OAI21_X1 U21078 ( .B1(n17958), .B2(n17901), .A(n17903), .ZN(n17905) );
  XOR2_X1 U21079 ( .A(n17905), .B(n17904), .Z(n18218) );
  AOI22_X1 U21080 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17915), .B1(
        n17953), .B2(n18218), .ZN(n17906) );
  OAI211_X1 U21081 ( .C1(n17956), .C2(n18226), .A(n17907), .B(n17906), .ZN(
        P3_U2817) );
  INV_X1 U21082 ( .A(n18228), .ZN(n18238) );
  AOI21_X1 U21083 ( .B1(n17932), .B2(n18238), .A(n17901), .ZN(n17908) );
  XOR2_X1 U21084 ( .A(n17908), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18234) );
  NAND2_X1 U21085 ( .A1(n18348), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18232) );
  OAI221_X1 U21086 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17911), .C1(
        n17910), .C2(n17909), .A(n18232), .ZN(n17912) );
  AOI21_X1 U21087 ( .B1(n17914), .B2(n17913), .A(n17912), .ZN(n17918) );
  OAI21_X1 U21088 ( .B1(n18228), .B2(n17956), .A(n18227), .ZN(n17916) );
  NAND2_X1 U21089 ( .A1(n17916), .A2(n17915), .ZN(n17917) );
  OAI211_X1 U21090 ( .C1(n18234), .C2(n17971), .A(n17918), .B(n17917), .ZN(
        P3_U2818) );
  OR2_X1 U21091 ( .A1(n17920), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18251) );
  OAI21_X1 U21092 ( .B1(n17920), .B2(n17945), .A(n17919), .ZN(n17921) );
  XOR2_X1 U21093 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17921), .Z(
        n18236) );
  NOR2_X1 U21094 ( .A1(n18358), .A2(n21241), .ZN(n18235) );
  NOR3_X1 U21095 ( .A1(n17974), .A2(n17976), .A3(n18693), .ZN(n17964) );
  NAND2_X1 U21096 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17964), .ZN(
        n17947) );
  NOR2_X1 U21097 ( .A1(n17922), .A2(n17947), .ZN(n17937) );
  AOI21_X1 U21098 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18049), .A(
        n17937), .ZN(n17924) );
  OAI22_X1 U21099 ( .A1(n17925), .A2(n17924), .B1(n18034), .B2(n17923), .ZN(
        n17926) );
  AOI211_X1 U21100 ( .C1(n17953), .C2(n18236), .A(n18235), .B(n17926), .ZN(
        n17930) );
  NOR2_X1 U21101 ( .A1(n18247), .A2(n17956), .ZN(n17940) );
  AOI22_X1 U21102 ( .A1(n17927), .A2(n17968), .B1(n18047), .B2(n18245), .ZN(
        n17955) );
  INV_X1 U21103 ( .A(n17955), .ZN(n17928) );
  OAI21_X1 U21104 ( .B1(n17940), .B2(n17928), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17929) );
  OAI211_X1 U21105 ( .C1(n17956), .C2(n18251), .A(n17930), .B(n17929), .ZN(
        P3_U2819) );
  AOI21_X1 U21106 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17932), .A(
        n17931), .ZN(n17933) );
  XOR2_X1 U21107 ( .A(n17943), .B(n17933), .Z(n18255) );
  NOR2_X1 U21108 ( .A1(n18358), .A2(n18929), .ZN(n17939) );
  NOR2_X1 U21109 ( .A1(n17934), .A2(n17947), .ZN(n17951) );
  AOI21_X1 U21110 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18049), .A(
        n17951), .ZN(n17936) );
  OAI22_X1 U21111 ( .A1(n17937), .A2(n17936), .B1(n18034), .B2(n17935), .ZN(
        n17938) );
  AOI211_X1 U21112 ( .C1(n17953), .C2(n18255), .A(n17939), .B(n17938), .ZN(
        n17942) );
  OAI21_X1 U21113 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17940), .ZN(n17941) );
  OAI211_X1 U21114 ( .C1(n17955), .C2(n17943), .A(n17942), .B(n17941), .ZN(
        P3_U2820) );
  INV_X1 U21115 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18258) );
  NAND2_X1 U21116 ( .A1(n17945), .A2(n17944), .ZN(n17946) );
  XOR2_X1 U21117 ( .A(n17946), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18262) );
  NOR2_X1 U21118 ( .A1(n18358), .A2(n21094), .ZN(n18261) );
  INV_X1 U21119 ( .A(n17947), .ZN(n17948) );
  AOI21_X1 U21120 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18049), .A(
        n17948), .ZN(n17950) );
  OAI22_X1 U21121 ( .A1(n17951), .A2(n17950), .B1(n18034), .B2(n17949), .ZN(
        n17952) );
  AOI211_X1 U21122 ( .C1(n17953), .C2(n18262), .A(n18261), .B(n17952), .ZN(
        n17954) );
  OAI221_X1 U21123 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17956), .C1(
        n18258), .C2(n17955), .A(n17954), .ZN(P3_U2821) );
  NOR2_X1 U21124 ( .A1(n18240), .A2(n17957), .ZN(n18274) );
  XOR2_X1 U21125 ( .A(n18274), .B(n17958), .Z(n18280) );
  INV_X1 U21126 ( .A(n17974), .ZN(n17959) );
  OAI21_X1 U21127 ( .B1(n18017), .B2(n17959), .A(n18054), .ZN(n17975) );
  AOI21_X1 U21128 ( .B1(n17960), .B2(n18753), .A(n17975), .ZN(n17961) );
  INV_X1 U21129 ( .A(n17961), .ZN(n17965) );
  INV_X1 U21130 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18927) );
  OAI22_X1 U21131 ( .A1(n18034), .A2(n17962), .B1(n18358), .B2(n18927), .ZN(
        n17963) );
  AOI221_X1 U21132 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17965), .C1(
        n17964), .C2(n17965), .A(n17963), .ZN(n17970) );
  AOI21_X1 U21133 ( .B1(n17967), .B2(n9918), .A(n17966), .ZN(n18276) );
  AOI22_X1 U21134 ( .A1(n18047), .A2(n18276), .B1(n17968), .B2(n18274), .ZN(
        n17969) );
  OAI211_X1 U21135 ( .C1(n18280), .C2(n17971), .A(n17970), .B(n17969), .ZN(
        P3_U2822) );
  OAI21_X1 U21136 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17973), .A(
        n17972), .ZN(n18290) );
  NOR2_X1 U21137 ( .A1(n17974), .A2(n18693), .ZN(n17977) );
  NOR2_X1 U21138 ( .A1(n18358), .A2(n18925), .ZN(n18281) );
  AOI221_X1 U21139 ( .B1(n17977), .B2(n17976), .C1(n17975), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18281), .ZN(n17983) );
  NAND2_X1 U21140 ( .A1(n17979), .A2(n17978), .ZN(n17980) );
  XOR2_X1 U21141 ( .A(n17980), .B(n18285), .Z(n18286) );
  AOI22_X1 U21142 ( .A1(n18047), .A2(n18286), .B1(n17981), .B2(n18048), .ZN(
        n17982) );
  OAI211_X1 U21143 ( .C1(n18057), .C2(n18290), .A(n17983), .B(n17982), .ZN(
        P3_U2823) );
  NAND2_X1 U21144 ( .A1(n9772), .A2(n18753), .ZN(n17987) );
  NAND2_X1 U21145 ( .A1(n18049), .A2(n17987), .ZN(n18007) );
  OAI21_X1 U21146 ( .B1(n17986), .B2(n17985), .A(n17984), .ZN(n18293) );
  OAI22_X1 U21147 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17987), .B1(
        n18057), .B2(n18293), .ZN(n17988) );
  AOI21_X1 U21148 ( .B1(n18348), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17988), .ZN(
        n17993) );
  AOI21_X1 U21149 ( .B1(n18297), .B2(n17990), .A(n17989), .ZN(n18295) );
  AOI22_X1 U21150 ( .A1(n18047), .A2(n18295), .B1(n17991), .B2(n18048), .ZN(
        n17992) );
  OAI211_X1 U21151 ( .C1(n17994), .C2(n18007), .A(n17993), .B(n17992), .ZN(
        P3_U2824) );
  OAI21_X1 U21152 ( .B1(n17996), .B2(n18029), .A(n17995), .ZN(n17997) );
  INV_X1 U21153 ( .A(n17997), .ZN(n18008) );
  OAI21_X1 U21154 ( .B1(n18000), .B2(n17999), .A(n17998), .ZN(n18001) );
  INV_X1 U21155 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18305) );
  XOR2_X1 U21156 ( .A(n18001), .B(n18305), .Z(n18302) );
  NOR2_X1 U21157 ( .A1(n18358), .A2(n18922), .ZN(n18301) );
  OAI21_X1 U21158 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18003), .A(
        n18002), .ZN(n18299) );
  OAI22_X1 U21159 ( .A1(n18034), .A2(n18004), .B1(n18057), .B2(n18299), .ZN(
        n18005) );
  AOI211_X1 U21160 ( .C1(n18047), .C2(n18302), .A(n18301), .B(n18005), .ZN(
        n18006) );
  OAI21_X1 U21161 ( .B1(n18008), .B2(n18007), .A(n18006), .ZN(P3_U2825) );
  OAI21_X1 U21162 ( .B1(n18011), .B2(n18010), .A(n18009), .ZN(n18310) );
  AOI21_X1 U21163 ( .B1(n18014), .B2(n18013), .A(n18012), .ZN(n18307) );
  OAI22_X1 U21164 ( .A1(n18358), .A2(n18919), .B1(n18693), .B2(n18015), .ZN(
        n18016) );
  AOI21_X1 U21165 ( .B1(n18047), .B2(n18307), .A(n18016), .ZN(n18021) );
  OAI21_X1 U21166 ( .B1(n18018), .B2(n18017), .A(n18054), .ZN(n18030) );
  AOI22_X1 U21167 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18030), .B1(
        n18019), .B2(n18048), .ZN(n18020) );
  OAI211_X1 U21168 ( .C1(n18057), .C2(n18310), .A(n18021), .B(n18020), .ZN(
        P3_U2826) );
  AOI21_X1 U21169 ( .B1(n18024), .B2(n18023), .A(n18022), .ZN(n18323) );
  OAI21_X1 U21170 ( .B1(n18027), .B2(n18026), .A(n18025), .ZN(n18320) );
  OAI22_X1 U21171 ( .A1(n18057), .A2(n18320), .B1(n18358), .B2(n18917), .ZN(
        n18028) );
  AOI21_X1 U21172 ( .B1(n18047), .B2(n18323), .A(n18028), .ZN(n18032) );
  NOR2_X1 U21173 ( .A1(n18029), .A2(n18039), .ZN(n18038) );
  OAI21_X1 U21174 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18038), .A(
        n18030), .ZN(n18031) );
  OAI211_X1 U21175 ( .C1(n18034), .C2(n18033), .A(n18032), .B(n18031), .ZN(
        P3_U2827) );
  OAI21_X1 U21176 ( .B1(n18037), .B2(n18036), .A(n18035), .ZN(n18332) );
  AOI21_X1 U21177 ( .B1(n18039), .B2(n18693), .A(n18038), .ZN(n18041) );
  AOI211_X1 U21178 ( .C1(n18335), .C2(n18334), .A(n18333), .B(n18058), .ZN(
        n18040) );
  AOI211_X1 U21179 ( .C1(n18042), .C2(n18048), .A(n18041), .B(n18040), .ZN(
        n18043) );
  NAND2_X1 U21180 ( .A1(n18348), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18339) );
  OAI211_X1 U21181 ( .C1(n18057), .C2(n18332), .A(n18043), .B(n18339), .ZN(
        P3_U2828) );
  OAI21_X1 U21182 ( .B1(n18045), .B2(n18052), .A(n18044), .ZN(n18352) );
  NAND2_X1 U21183 ( .A1(n19011), .A2(n18053), .ZN(n18046) );
  XNOR2_X1 U21184 ( .A(n18046), .B(n18045), .ZN(n18347) );
  AOI22_X1 U21185 ( .A1(n18047), .A2(n18347), .B1(n18348), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18051) );
  AOI22_X1 U21186 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18049), .B1(
        n18048), .B2(n21104), .ZN(n18050) );
  OAI211_X1 U21187 ( .C1(n18057), .C2(n18352), .A(n18051), .B(n18050), .ZN(
        P3_U2829) );
  AOI21_X1 U21188 ( .B1(n18053), .B2(n19011), .A(n18052), .ZN(n18356) );
  INV_X1 U21189 ( .A(n18356), .ZN(n18354) );
  NAND3_X1 U21190 ( .A1(n18887), .A2(n18891), .A3(n18054), .ZN(n18055) );
  AOI22_X1 U21191 ( .A1(n18348), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18055), .ZN(n18056) );
  OAI221_X1 U21192 ( .B1(n18356), .B2(n18058), .C1(n18354), .C2(n18057), .A(
        n18056), .ZN(P3_U2830) );
  NOR2_X1 U21193 ( .A1(n18348), .A2(n18059), .ZN(n18068) );
  NAND2_X1 U21194 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18060), .ZN(
        n18119) );
  OAI21_X1 U21195 ( .B1(n18062), .B2(n18119), .A(n18061), .ZN(n18098) );
  OAI221_X1 U21196 ( .B1(n9863), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C1(
        n9863), .C2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n18098), .ZN(
        n18084) );
  NAND2_X1 U21197 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18076), .ZN(
        n18067) );
  AOI222_X1 U21198 ( .A1(n18068), .A2(n18067), .B1(n18068), .B2(n18359), .C1(
        n18067), .C2(n18066), .ZN(n18070) );
  NAND2_X1 U21199 ( .A1(n18348), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18069) );
  OAI211_X1 U21200 ( .C1(n18071), .C2(n18279), .A(n18070), .B(n18069), .ZN(
        P3_U2835) );
  INV_X1 U21201 ( .A(n18121), .ZN(n18073) );
  NOR3_X1 U21202 ( .A1(n18073), .A2(n18103), .A3(n18072), .ZN(n18078) );
  OAI22_X1 U21203 ( .A1(n18076), .A2(n21254), .B1(n18075), .B2(n18074), .ZN(
        n18077) );
  OAI21_X1 U21204 ( .B1(n18078), .B2(n18077), .A(n18338), .ZN(n18080) );
  OAI211_X1 U21205 ( .C1(n18343), .C2(n21254), .A(n18080), .B(n18079), .ZN(
        P3_U2836) );
  INV_X1 U21206 ( .A(n18081), .ZN(n18087) );
  NOR2_X1 U21207 ( .A1(n18103), .A2(n18082), .ZN(n18083) );
  AOI21_X1 U21208 ( .B1(n18116), .B2(n18083), .A(n18267), .ZN(n18085) );
  NOR2_X1 U21209 ( .A1(n18085), .A2(n18084), .ZN(n18086) );
  MUX2_X1 U21210 ( .A(n18087), .B(n18086), .S(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n18089) );
  OAI21_X1 U21211 ( .B1(n18359), .B2(n18089), .A(n18088), .ZN(n18093) );
  OAI22_X1 U21212 ( .A1(n18210), .A2(n18091), .B1(n18279), .B2(n18090), .ZN(
        n18092) );
  AOI211_X1 U21213 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18291), .A(
        n18093), .B(n18092), .ZN(n18094) );
  OAI21_X1 U21214 ( .B1(n18317), .B2(n18095), .A(n18094), .ZN(P3_U2837) );
  AOI22_X1 U21215 ( .A1(n18808), .A2(n18097), .B1(n18191), .B2(n18096), .ZN(
        n18099) );
  NAND3_X1 U21216 ( .A1(n18099), .A2(n18343), .A3(n18098), .ZN(n18102) );
  AOI211_X1 U21217 ( .C1(n18851), .C2(n18100), .A(n18113), .B(n18102), .ZN(
        n18101) );
  OR2_X1 U21218 ( .A1(n18348), .A2(n18101), .ZN(n18114) );
  OAI21_X1 U21219 ( .B1(n18270), .B2(n18102), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18108) );
  NOR3_X1 U21220 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18103), .A3(
        n18130), .ZN(n18104) );
  AOI21_X1 U21221 ( .B1(n18263), .B2(n18105), .A(n18104), .ZN(n18107) );
  OAI211_X1 U21222 ( .C1(n18114), .C2(n18108), .A(n18107), .B(n18106), .ZN(
        P3_U2838) );
  NAND3_X1 U21223 ( .A1(n18109), .A2(n18343), .A3(n18121), .ZN(n18112) );
  AOI22_X1 U21224 ( .A1(n18348), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18263), 
        .B2(n18110), .ZN(n18111) );
  OAI221_X1 U21225 ( .B1(n18114), .B2(n18113), .C1(n18114), .C2(n18112), .A(
        n18111), .ZN(P3_U2839) );
  AOI22_X1 U21226 ( .A1(n18808), .A2(n18115), .B1(n18191), .B2(n18190), .ZN(
        n18134) );
  AOI21_X1 U21227 ( .B1(n18137), .B2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n18237), .ZN(n18120) );
  INV_X1 U21228 ( .A(n18116), .ZN(n18156) );
  OAI21_X1 U21229 ( .B1(n18131), .B2(n18156), .A(n18851), .ZN(n18117) );
  OAI221_X1 U21230 ( .B1(n18832), .B2(n18155), .C1(n18832), .C2(n18145), .A(
        n18117), .ZN(n18135) );
  NOR2_X1 U21231 ( .A1(n18808), .A2(n18191), .ZN(n18246) );
  OAI22_X1 U21232 ( .A1(n18832), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18118), .B2(n18246), .ZN(n18139) );
  NOR4_X1 U21233 ( .A1(n18120), .A2(n18135), .A3(n18119), .A4(n18139), .ZN(
        n18124) );
  AOI21_X1 U21234 ( .B1(n18122), .B2(n18121), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18123) );
  AOI211_X1 U21235 ( .C1(n18134), .C2(n18124), .A(n18123), .B(n18359), .ZN(
        n18125) );
  AOI21_X1 U21236 ( .B1(n18126), .B2(n18263), .A(n18125), .ZN(n18128) );
  NAND2_X1 U21237 ( .A1(n18348), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18127) );
  OAI211_X1 U21238 ( .C1(n18343), .C2(n18129), .A(n18128), .B(n18127), .ZN(
        P3_U2840) );
  AOI22_X1 U21239 ( .A1(n18348), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18263), 
        .B2(n18132), .ZN(n18141) );
  NOR2_X1 U21240 ( .A1(n18851), .A2(n18828), .ZN(n18342) );
  NOR3_X1 U21241 ( .A1(n19011), .A2(n18163), .A3(n18201), .ZN(n18177) );
  AOI21_X1 U21242 ( .B1(n18133), .B2(n18177), .A(n18843), .ZN(n18136) );
  NAND2_X1 U21243 ( .A1(n18338), .A2(n18134), .ZN(n18181) );
  NOR3_X1 U21244 ( .A1(n18136), .A2(n18181), .A3(n18135), .ZN(n18144) );
  OAI21_X1 U21245 ( .B1(n18137), .B2(n18342), .A(n18144), .ZN(n18138) );
  OAI211_X1 U21246 ( .C1(n18139), .C2(n18138), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18358), .ZN(n18140) );
  OAI211_X1 U21247 ( .C1(n18142), .C2(n18154), .A(n18141), .B(n18140), .ZN(
        P3_U2841) );
  AOI22_X1 U21248 ( .A1(n18348), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18263), 
        .B2(n18143), .ZN(n18148) );
  AOI221_X1 U21249 ( .B1(n18145), .B2(n18144), .C1(n18246), .C2(n18144), .A(
        n18348), .ZN(n18151) );
  NOR3_X1 U21250 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18342), .A3(
        n18866), .ZN(n18146) );
  OAI21_X1 U21251 ( .B1(n18151), .B2(n18146), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18147) );
  OAI211_X1 U21252 ( .C1(n18154), .C2(n18149), .A(n18148), .B(n18147), .ZN(
        P3_U2842) );
  AOI22_X1 U21253 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18151), .B1(
        n18263), .B2(n18150), .ZN(n18153) );
  OAI211_X1 U21254 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18154), .A(
        n18153), .B(n18152), .ZN(P3_U2843) );
  AOI21_X1 U21255 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18155), .A(
        n9863), .ZN(n18160) );
  NAND2_X1 U21256 ( .A1(n18851), .A2(n18156), .ZN(n18157) );
  NAND2_X1 U21257 ( .A1(n18828), .A2(n19011), .ZN(n18325) );
  OAI211_X1 U21258 ( .C1(n18158), .C2(n18246), .A(n18157), .B(n18325), .ZN(
        n18159) );
  NOR3_X1 U21259 ( .A1(n18160), .A2(n18181), .A3(n18159), .ZN(n18170) );
  AOI221_X1 U21260 ( .B1(n9863), .B2(n18170), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18170), .A(n18348), .ZN(
        n18166) );
  AOI22_X1 U21261 ( .A1(n18851), .A2(n18161), .B1(n18308), .B2(n18329), .ZN(
        n18319) );
  NOR2_X1 U21262 ( .A1(n18319), .A2(n18162), .ZN(n18282) );
  NAND2_X1 U21263 ( .A1(n18217), .A2(n18282), .ZN(n18188) );
  AOI211_X1 U21264 ( .C1(n18164), .C2(n18188), .A(n18163), .B(n18359), .ZN(
        n18183) );
  AOI22_X1 U21265 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18166), .B1(
        n18165), .B2(n18183), .ZN(n18168) );
  NAND2_X1 U21266 ( .A1(n18348), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18167) );
  OAI211_X1 U21267 ( .C1(n18169), .C2(n18279), .A(n18168), .B(n18167), .ZN(
        P3_U2844) );
  NOR2_X1 U21268 ( .A1(n18348), .A2(n18170), .ZN(n18172) );
  OAI222_X1 U21269 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18183), .C1(n18172), .C2(
        n18171), .ZN(n18174) );
  OAI211_X1 U21270 ( .C1(n18175), .C2(n18279), .A(n18174), .B(n18173), .ZN(
        P3_U2845) );
  AOI22_X1 U21271 ( .A1(n18851), .A2(n18176), .B1(n18818), .B2(n18201), .ZN(
        n18241) );
  AOI21_X1 U21272 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18843), .A(
        n18177), .ZN(n18178) );
  INV_X1 U21273 ( .A(n18178), .ZN(n18179) );
  OAI211_X1 U21274 ( .C1(n18180), .C2(n18237), .A(n18241), .B(n18179), .ZN(
        n18189) );
  OAI221_X1 U21275 ( .B1(n18181), .B2(n18270), .C1(n18181), .C2(n18189), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18186) );
  AOI22_X1 U21276 ( .A1(n18263), .A2(n18184), .B1(n18183), .B2(n18182), .ZN(
        n18185) );
  OAI221_X1 U21277 ( .B1(n18348), .B2(n18186), .C1(n18358), .C2(n18940), .A(
        n18185), .ZN(P3_U2846) );
  INV_X1 U21278 ( .A(n18187), .ZN(n18200) );
  AOI22_X1 U21279 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18291), .B1(
        n18348), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18199) );
  NOR2_X1 U21280 ( .A1(n18204), .A2(n18188), .ZN(n18207) );
  OAI21_X1 U21281 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18207), .A(
        n18189), .ZN(n18194) );
  NAND2_X1 U21282 ( .A1(n18191), .A2(n18190), .ZN(n18192) );
  OAI22_X1 U21283 ( .A1(n18195), .A2(n18194), .B1(n18193), .B2(n18192), .ZN(
        n18197) );
  AOI22_X1 U21284 ( .A1(n18338), .A2(n18197), .B1(n18263), .B2(n18196), .ZN(
        n18198) );
  OAI211_X1 U21285 ( .C1(n18317), .C2(n18200), .A(n18199), .B(n18198), .ZN(
        P3_U2847) );
  NOR2_X1 U21286 ( .A1(n19011), .A2(n18201), .ZN(n18242) );
  OAI221_X1 U21287 ( .B1(n18843), .B2(n18202), .C1(n18843), .C2(n18242), .A(
        n18241), .ZN(n18221) );
  AOI211_X1 U21288 ( .C1(n18204), .C2(n18252), .A(n18203), .B(n18221), .ZN(
        n18205) );
  OAI21_X1 U21289 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18342), .A(
        n18205), .ZN(n18206) );
  OAI211_X1 U21290 ( .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18207), .A(
        n18338), .B(n18206), .ZN(n18208) );
  OAI21_X1 U21291 ( .B1(n18937), .B2(n18358), .A(n18208), .ZN(n18213) );
  OAI22_X1 U21292 ( .A1(n18317), .A2(n18211), .B1(n18210), .B2(n18209), .ZN(
        n18212) );
  AOI211_X1 U21293 ( .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18291), .A(
        n18213), .B(n18212), .ZN(n18214) );
  OAI21_X1 U21294 ( .B1(n18215), .B2(n18279), .A(n18214), .ZN(P3_U2848) );
  NAND2_X1 U21295 ( .A1(n18338), .A2(n18282), .ZN(n18298) );
  INV_X1 U21296 ( .A(n18298), .ZN(n18216) );
  AOI222_X1 U21297 ( .A1(n9878), .A2(n18355), .B1(n18240), .B2(n18275), .C1(
        n18217), .C2(n18216), .ZN(n18265) );
  AOI22_X1 U21298 ( .A1(n18348), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18263), 
        .B2(n18218), .ZN(n18225) );
  OAI22_X1 U21299 ( .A1(n18238), .A2(n18237), .B1(n18219), .B2(n18239), .ZN(
        n18220) );
  AOI211_X1 U21300 ( .C1(n18808), .C2(n18222), .A(n18221), .B(n18220), .ZN(
        n18229) );
  OAI211_X1 U21301 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18237), .A(
        n18338), .B(n18229), .ZN(n18223) );
  NAND3_X1 U21302 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18358), .A3(
        n18223), .ZN(n18224) );
  OAI211_X1 U21303 ( .C1(n18265), .C2(n18226), .A(n18225), .B(n18224), .ZN(
        P3_U2849) );
  OAI22_X1 U21304 ( .A1(n18265), .A2(n18228), .B1(n18227), .B2(n18359), .ZN(
        n18231) );
  NAND2_X1 U21305 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18229), .ZN(
        n18230) );
  AOI22_X1 U21306 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18291), .B1(
        n18231), .B2(n18230), .ZN(n18233) );
  OAI211_X1 U21307 ( .C1(n18234), .C2(n18279), .A(n18233), .B(n18232), .ZN(
        P3_U2850) );
  AOI21_X1 U21308 ( .B1(n18263), .B2(n18236), .A(n18235), .ZN(n18250) );
  NOR2_X1 U21309 ( .A1(n18238), .A2(n18237), .ZN(n18248) );
  NOR2_X1 U21310 ( .A1(n18240), .A2(n18239), .ZN(n18244) );
  OAI211_X1 U21311 ( .C1(n18843), .C2(n18242), .A(n18338), .B(n18241), .ZN(
        n18243) );
  AOI211_X1 U21312 ( .C1(n18245), .C2(n18808), .A(n18244), .B(n18243), .ZN(
        n18259) );
  OAI221_X1 U21313 ( .B1(n18247), .B2(n18843), .C1(n18247), .C2(n18246), .A(
        n18259), .ZN(n18253) );
  OAI211_X1 U21314 ( .C1(n18248), .C2(n18253), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18358), .ZN(n18249) );
  OAI211_X1 U21315 ( .C1(n18265), .C2(n18251), .A(n18250), .B(n18249), .ZN(
        P3_U2851) );
  OAI221_X1 U21316 ( .B1(n18253), .B2(n18258), .C1(n18253), .C2(n18252), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18257) );
  NOR3_X1 U21317 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18265), .A3(
        n18258), .ZN(n18254) );
  AOI21_X1 U21318 ( .B1(n18263), .B2(n18255), .A(n18254), .ZN(n18256) );
  OAI221_X1 U21319 ( .B1(n18348), .B2(n18257), .C1(n18358), .C2(n18929), .A(
        n18256), .ZN(P3_U2852) );
  NOR3_X1 U21320 ( .A1(n18348), .A2(n18259), .A3(n18258), .ZN(n18260) );
  AOI211_X1 U21321 ( .C1(n18263), .C2(n18262), .A(n18261), .B(n18260), .ZN(
        n18264) );
  OAI21_X1 U21322 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18265), .A(
        n18264), .ZN(P3_U2853) );
  NOR3_X1 U21323 ( .A1(n18285), .A2(n18297), .A3(n18298), .ZN(n18273) );
  AND2_X1 U21324 ( .A1(n18266), .A2(n18325), .ZN(n18269) );
  OAI22_X1 U21325 ( .A1(n9863), .A2(n18269), .B1(n18268), .B2(n18267), .ZN(
        n18292) );
  AOI211_X1 U21326 ( .C1(n18270), .C2(n18297), .A(n18285), .B(n18292), .ZN(
        n18283) );
  OAI21_X1 U21327 ( .B1(n18283), .B2(n18344), .A(n18343), .ZN(n18272) );
  NOR2_X1 U21328 ( .A1(n18358), .A2(n18927), .ZN(n18271) );
  AOI221_X1 U21329 ( .B1(n18273), .B2(n9918), .C1(n18272), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18271), .ZN(n18278) );
  AOI22_X1 U21330 ( .A1(n18355), .A2(n18276), .B1(n18275), .B2(n18274), .ZN(
        n18277) );
  OAI211_X1 U21331 ( .C1(n18280), .C2(n18279), .A(n18278), .B(n18277), .ZN(
        P3_U2854) );
  AOI21_X1 U21332 ( .B1(n18291), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18281), .ZN(n18289) );
  INV_X1 U21333 ( .A(n18282), .ZN(n18284) );
  AOI221_X1 U21334 ( .B1(n18297), .B2(n18285), .C1(n18284), .C2(n18285), .A(
        n18283), .ZN(n18287) );
  AOI22_X1 U21335 ( .A1(n18338), .A2(n18287), .B1(n18355), .B2(n18286), .ZN(
        n18288) );
  OAI211_X1 U21336 ( .C1(n18351), .C2(n18290), .A(n18289), .B(n18288), .ZN(
        P3_U2855) );
  AOI21_X1 U21337 ( .B1(n18338), .B2(n18292), .A(n18291), .ZN(n18304) );
  OAI22_X1 U21338 ( .A1(n18358), .A2(n18923), .B1(n18351), .B2(n18293), .ZN(
        n18294) );
  AOI21_X1 U21339 ( .B1(n18355), .B2(n18295), .A(n18294), .ZN(n18296) );
  OAI221_X1 U21340 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18298), .C1(
        n18297), .C2(n18304), .A(n18296), .ZN(P3_U2856) );
  NOR3_X1 U21341 ( .A1(n18319), .A2(n18359), .A3(n13167), .ZN(n18314) );
  NAND2_X1 U21342 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18314), .ZN(
        n18306) );
  NOR2_X1 U21343 ( .A1(n18351), .A2(n18299), .ZN(n18300) );
  AOI211_X1 U21344 ( .C1(n18355), .C2(n18302), .A(n18301), .B(n18300), .ZN(
        n18303) );
  OAI221_X1 U21345 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18306), .C1(
        n18305), .C2(n18304), .A(n18303), .ZN(P3_U2857) );
  INV_X1 U21346 ( .A(n18307), .ZN(n18316) );
  OAI211_X1 U21347 ( .C1(n9863), .C2(n18308), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18325), .ZN(n18309) );
  AOI21_X1 U21348 ( .B1(n18851), .B2(n18328), .A(n18309), .ZN(n18318) );
  OAI21_X1 U21349 ( .B1(n18318), .B2(n18344), .A(n18343), .ZN(n18312) );
  OAI22_X1 U21350 ( .A1(n18358), .A2(n18919), .B1(n18351), .B2(n18310), .ZN(
        n18311) );
  AOI221_X1 U21351 ( .B1(n18314), .B2(n18313), .C1(n18312), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18311), .ZN(n18315) );
  OAI21_X1 U21352 ( .B1(n18317), .B2(n18316), .A(n18315), .ZN(P3_U2858) );
  AOI211_X1 U21353 ( .C1(n18319), .C2(n13167), .A(n18318), .B(n18359), .ZN(
        n18322) );
  OAI22_X1 U21354 ( .A1(n18358), .A2(n18917), .B1(n18351), .B2(n18320), .ZN(
        n18321) );
  AOI211_X1 U21355 ( .C1(n18323), .C2(n18355), .A(n18322), .B(n18321), .ZN(
        n18324) );
  OAI21_X1 U21356 ( .B1(n13167), .B2(n18343), .A(n18324), .ZN(P3_U2859) );
  NAND3_X1 U21357 ( .A1(n18851), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18326) );
  OAI211_X1 U21358 ( .C1(n9863), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18326), .B(n18325), .ZN(n18327) );
  AOI22_X1 U21359 ( .A1(n18851), .A2(n18328), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18327), .ZN(n18331) );
  NAND3_X1 U21360 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18329), .A3(
        n18341), .ZN(n18330) );
  OAI211_X1 U21361 ( .C1(n18332), .C2(n18814), .A(n18331), .B(n18330), .ZN(
        n18337) );
  AOI21_X1 U21362 ( .B1(n18335), .B2(n18334), .A(n18333), .ZN(n18336) );
  AOI22_X1 U21363 ( .A1(n18338), .A2(n18337), .B1(n18355), .B2(n18336), .ZN(
        n18340) );
  OAI211_X1 U21364 ( .C1(n18343), .C2(n18341), .A(n18340), .B(n18339), .ZN(
        P3_U2860) );
  OR3_X1 U21365 ( .A1(n18359), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18342), .ZN(n18361) );
  AOI21_X1 U21366 ( .B1(n18343), .B2(n18361), .A(n18994), .ZN(n18346) );
  AOI211_X1 U21367 ( .C1(n18832), .C2(n19011), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18344), .ZN(n18345) );
  AOI211_X1 U21368 ( .C1(n18355), .C2(n18347), .A(n18346), .B(n18345), .ZN(
        n18350) );
  NAND2_X1 U21369 ( .A1(n18348), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18349) );
  OAI211_X1 U21370 ( .C1(n18352), .C2(n18351), .A(n18350), .B(n18349), .ZN(
        P3_U2861) );
  INV_X1 U21371 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19022) );
  NOR2_X1 U21372 ( .A1(n18358), .A2(n19022), .ZN(n18353) );
  AOI221_X1 U21373 ( .B1(n18357), .B2(n18356), .C1(n18355), .C2(n18354), .A(
        n18353), .ZN(n18362) );
  OAI211_X1 U21374 ( .C1(n18818), .C2(n18359), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18358), .ZN(n18360) );
  NAND3_X1 U21375 ( .A1(n18362), .A2(n18361), .A3(n18360), .ZN(P3_U2862) );
  AOI21_X1 U21376 ( .B1(n18365), .B2(n18364), .A(n18363), .ZN(n18877) );
  OAI21_X1 U21377 ( .B1(n18877), .B2(n18414), .A(n18370), .ZN(n18366) );
  OAI221_X1 U21378 ( .B1(n18834), .B2(n19028), .C1(n18834), .C2(n18370), .A(
        n18366), .ZN(P3_U2863) );
  INV_X1 U21379 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18858) );
  NAND2_X1 U21380 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18855), .ZN(
        n18618) );
  NAND2_X1 U21381 ( .A1(n18858), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18547) );
  AND2_X1 U21382 ( .A1(n18618), .A2(n18547), .ZN(n18368) );
  OAI22_X1 U21383 ( .A1(n18369), .A2(n18858), .B1(n18368), .B2(n18367), .ZN(
        P3_U2866) );
  NOR2_X1 U21384 ( .A1(n18859), .A2(n18370), .ZN(P3_U2867) );
  NAND2_X1 U21385 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18753), .ZN(n18697) );
  NAND2_X1 U21386 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18691) );
  NAND2_X1 U21387 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18833), .ZN(
        n18594) );
  NOR2_X2 U21388 ( .A1(n18691), .A2(n18594), .ZN(n18799) );
  INV_X1 U21389 ( .A(n18799), .ZN(n18769) );
  NOR2_X1 U21390 ( .A1(n18693), .A2(n18371), .ZN(n18689) );
  NOR2_X1 U21391 ( .A1(n18858), .A2(n18372), .ZN(n18751) );
  NAND2_X1 U21392 ( .A1(n18834), .A2(n18751), .ZN(n18737) );
  INV_X1 U21393 ( .A(n18737), .ZN(n18741) );
  NOR2_X2 U21394 ( .A1(n18620), .A2(n18373), .ZN(n18748) );
  NAND2_X1 U21395 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18751), .ZN(
        n18789) );
  NAND2_X1 U21396 ( .A1(n18833), .A2(n18834), .ZN(n18837) );
  NOR2_X1 U21397 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18459) );
  INV_X1 U21398 ( .A(n18459), .ZN(n18415) );
  NOR2_X2 U21399 ( .A1(n18837), .A2(n18415), .ZN(n18475) );
  INV_X1 U21400 ( .A(n18475), .ZN(n18474) );
  NAND2_X1 U21401 ( .A1(n18789), .A2(n18474), .ZN(n18374) );
  INV_X1 U21402 ( .A(n18374), .ZN(n18439) );
  NOR2_X1 U21403 ( .A1(n18747), .A2(n18439), .ZN(n18408) );
  AOI22_X1 U21404 ( .A1(n18689), .A2(n18741), .B1(n18748), .B2(n18408), .ZN(
        n18381) );
  NOR2_X1 U21405 ( .A1(n18799), .A2(n18741), .ZN(n18717) );
  INV_X1 U21406 ( .A(n18717), .ZN(n18376) );
  AOI21_X1 U21407 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18620), .ZN(n18375) );
  AOI22_X1 U21408 ( .A1(n18753), .A2(n18376), .B1(n18375), .B2(n18374), .ZN(
        n18411) );
  NAND2_X1 U21409 ( .A1(n18378), .A2(n18377), .ZN(n18409) );
  NOR2_X2 U21410 ( .A1(n18379), .A2(n18409), .ZN(n18754) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18411), .B1(
        n18754), .B2(n18475), .ZN(n18380) );
  OAI211_X1 U21412 ( .C1(n18697), .C2(n18769), .A(n18381), .B(n18380), .ZN(
        P3_U2868) );
  NOR2_X1 U21413 ( .A1(n18409), .A2(n19033), .ZN(n18598) );
  AND2_X1 U21414 ( .A1(n18753), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18759) );
  NOR2_X2 U21415 ( .A1(n18620), .A2(n18382), .ZN(n18758) );
  AOI22_X1 U21416 ( .A1(n18759), .A2(n18741), .B1(n18758), .B2(n18408), .ZN(
        n18384) );
  AND2_X1 U21417 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18753), .ZN(n18760) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18411), .B1(
        n18760), .B2(n18799), .ZN(n18383) );
  OAI211_X1 U21419 ( .C1(n18763), .C2(n18474), .A(n18384), .B(n18383), .ZN(
        P3_U2869) );
  NAND2_X1 U21420 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18753), .ZN(n18729) );
  NAND2_X1 U21421 ( .A1(n18753), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18770) );
  INV_X1 U21422 ( .A(n18770), .ZN(n18726) );
  NOR2_X2 U21423 ( .A1(n18620), .A2(n18385), .ZN(n18764) );
  AOI22_X1 U21424 ( .A1(n18726), .A2(n18741), .B1(n18764), .B2(n18408), .ZN(
        n18388) );
  NOR2_X2 U21425 ( .A1(n18386), .A2(n18409), .ZN(n18766) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18411), .B1(
        n18766), .B2(n18475), .ZN(n18387) );
  OAI211_X1 U21427 ( .C1(n18729), .C2(n18769), .A(n18388), .B(n18387), .ZN(
        P3_U2870) );
  INV_X1 U21428 ( .A(n18409), .ZN(n18399) );
  NAND2_X1 U21429 ( .A1(n18399), .A2(n18389), .ZN(n18776) );
  NOR2_X2 U21430 ( .A1(n18620), .A2(n18390), .ZN(n18772) );
  AND2_X1 U21431 ( .A1(n18753), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18771) );
  AOI22_X1 U21432 ( .A1(n18772), .A2(n18408), .B1(n18771), .B2(n18741), .ZN(
        n18392) );
  AND2_X1 U21433 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18753), .ZN(n18773) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18411), .B1(
        n18773), .B2(n18799), .ZN(n18391) );
  OAI211_X1 U21435 ( .C1(n18776), .C2(n18474), .A(n18392), .B(n18391), .ZN(
        P3_U2871) );
  NAND2_X1 U21436 ( .A1(n18399), .A2(n18393), .ZN(n18782) );
  AND2_X1 U21437 ( .A1(n18753), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18779) );
  NOR2_X2 U21438 ( .A1(n18620), .A2(n18394), .ZN(n18777) );
  AOI22_X1 U21439 ( .A1(n18779), .A2(n18741), .B1(n18777), .B2(n18408), .ZN(
        n18397) );
  NOR2_X2 U21440 ( .A1(n18395), .A2(n18693), .ZN(n18778) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18411), .B1(
        n18778), .B2(n18799), .ZN(n18396) );
  OAI211_X1 U21442 ( .C1(n18782), .C2(n18474), .A(n18397), .B(n18396), .ZN(
        P3_U2872) );
  NAND2_X1 U21443 ( .A1(n18399), .A2(n18398), .ZN(n18790) );
  AND2_X1 U21444 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18753), .ZN(n18784) );
  NOR2_X2 U21445 ( .A1(n18620), .A2(n18400), .ZN(n18783) );
  AOI22_X1 U21446 ( .A1(n18784), .A2(n18799), .B1(n18783), .B2(n18408), .ZN(
        n18402) );
  AND2_X1 U21447 ( .A1(n18753), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18786) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18411), .B1(
        n18786), .B2(n18741), .ZN(n18401) );
  OAI211_X1 U21449 ( .C1(n18790), .C2(n18474), .A(n18402), .B(n18401), .ZN(
        P3_U2873) );
  NOR2_X1 U21450 ( .A1(n18693), .A2(n14504), .ZN(n18792) );
  INV_X1 U21451 ( .A(n18792), .ZN(n18682) );
  NOR2_X2 U21452 ( .A1(n18620), .A2(n18403), .ZN(n18791) );
  NAND2_X1 U21453 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18753), .ZN(n18796) );
  INV_X1 U21454 ( .A(n18796), .ZN(n18679) );
  AOI22_X1 U21455 ( .A1(n18791), .A2(n18408), .B1(n18679), .B2(n18799), .ZN(
        n18406) );
  NOR2_X2 U21456 ( .A1(n18404), .A2(n18409), .ZN(n18793) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18411), .B1(
        n18793), .B2(n18475), .ZN(n18405) );
  OAI211_X1 U21458 ( .C1(n18682), .C2(n18737), .A(n18406), .B(n18405), .ZN(
        P3_U2874) );
  NAND2_X1 U21459 ( .A1(n18753), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18806) );
  NAND2_X1 U21460 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18753), .ZN(n18716) );
  INV_X1 U21461 ( .A(n18716), .ZN(n18800) );
  NOR2_X2 U21462 ( .A1(n18407), .A2(n18620), .ZN(n18798) );
  AOI22_X1 U21463 ( .A1(n18800), .A2(n18741), .B1(n18798), .B2(n18408), .ZN(
        n18413) );
  NOR2_X2 U21464 ( .A1(n18410), .A2(n18409), .ZN(n18802) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18411), .B1(
        n18802), .B2(n18475), .ZN(n18412) );
  OAI211_X1 U21466 ( .C1(n18806), .C2(n18769), .A(n18413), .B(n18412), .ZN(
        P3_U2875) );
  INV_X1 U21467 ( .A(n18751), .ZN(n18746) );
  NOR2_X1 U21468 ( .A1(n18414), .A2(n18620), .ZN(n18750) );
  NAND2_X1 U21469 ( .A1(n18750), .A2(n18833), .ZN(n18690) );
  OAI22_X1 U21470 ( .A1(n18693), .A2(n18746), .B1(n18415), .B2(n18690), .ZN(
        n18437) );
  OR2_X1 U21471 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18747), .ZN(
        n18688) );
  NOR2_X1 U21472 ( .A1(n18415), .A2(n18688), .ZN(n18434) );
  INV_X1 U21473 ( .A(n18697), .ZN(n18749) );
  AOI22_X1 U21474 ( .A1(n18748), .A2(n18434), .B1(n18749), .B2(n18741), .ZN(
        n18417) );
  INV_X1 U21475 ( .A(n18789), .ZN(n18801) );
  NOR2_X2 U21476 ( .A1(n18594), .A2(n18415), .ZN(n18494) );
  AOI22_X1 U21477 ( .A1(n18689), .A2(n18801), .B1(n18754), .B2(n18494), .ZN(
        n18416) );
  OAI211_X1 U21478 ( .C1(n18418), .C2(n18437), .A(n18417), .B(n18416), .ZN(
        P3_U2876) );
  AOI22_X1 U21479 ( .A1(n18759), .A2(n18801), .B1(n18758), .B2(n18434), .ZN(
        n18420) );
  AOI22_X1 U21480 ( .A1(n18760), .A2(n18741), .B1(n18598), .B2(n18494), .ZN(
        n18419) );
  OAI211_X1 U21481 ( .C1(n18421), .C2(n18437), .A(n18420), .B(n18419), .ZN(
        P3_U2877) );
  AOI22_X1 U21482 ( .A1(n18726), .A2(n18801), .B1(n18764), .B2(n18434), .ZN(
        n18423) );
  INV_X1 U21483 ( .A(n18729), .ZN(n18765) );
  AOI22_X1 U21484 ( .A1(n18766), .A2(n18494), .B1(n18765), .B2(n18741), .ZN(
        n18422) );
  OAI211_X1 U21485 ( .C1(n18424), .C2(n18437), .A(n18423), .B(n18422), .ZN(
        P3_U2878) );
  INV_X1 U21486 ( .A(n18494), .ZN(n18501) );
  AOI22_X1 U21487 ( .A1(n18773), .A2(n18741), .B1(n18772), .B2(n18434), .ZN(
        n18426) );
  INV_X1 U21488 ( .A(n18437), .ZN(n18431) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18431), .B1(
        n18771), .B2(n18801), .ZN(n18425) );
  OAI211_X1 U21490 ( .C1(n18776), .C2(n18501), .A(n18426), .B(n18425), .ZN(
        P3_U2879) );
  AOI22_X1 U21491 ( .A1(n18779), .A2(n18801), .B1(n18777), .B2(n18434), .ZN(
        n18428) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18431), .B1(
        n18778), .B2(n18741), .ZN(n18427) );
  OAI211_X1 U21493 ( .C1(n18782), .C2(n18501), .A(n18428), .B(n18427), .ZN(
        P3_U2880) );
  AOI22_X1 U21494 ( .A1(n18786), .A2(n18801), .B1(n18783), .B2(n18434), .ZN(
        n18430) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18431), .B1(
        n18784), .B2(n18741), .ZN(n18429) );
  OAI211_X1 U21496 ( .C1(n18790), .C2(n18501), .A(n18430), .B(n18429), .ZN(
        P3_U2881) );
  AOI22_X1 U21497 ( .A1(n18792), .A2(n18801), .B1(n18791), .B2(n18434), .ZN(
        n18433) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18431), .B1(
        n18793), .B2(n18494), .ZN(n18432) );
  OAI211_X1 U21499 ( .C1(n18796), .C2(n18737), .A(n18433), .B(n18432), .ZN(
        P3_U2882) );
  INV_X1 U21500 ( .A(n18806), .ZN(n18711) );
  AOI22_X1 U21501 ( .A1(n18798), .A2(n18434), .B1(n18711), .B2(n18741), .ZN(
        n18436) );
  AOI22_X1 U21502 ( .A1(n18800), .A2(n18801), .B1(n18802), .B2(n18494), .ZN(
        n18435) );
  OAI211_X1 U21503 ( .C1(n18438), .C2(n18437), .A(n18436), .B(n18435), .ZN(
        P3_U2883) );
  NAND2_X1 U21504 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18459), .ZN(
        n18502) );
  NOR2_X2 U21505 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18502), .ZN(
        n18519) );
  NOR2_X1 U21506 ( .A1(n18494), .A2(n18519), .ZN(n18480) );
  NOR2_X1 U21507 ( .A1(n18747), .A2(n18480), .ZN(n18455) );
  AOI22_X1 U21508 ( .A1(n18689), .A2(n18475), .B1(n18748), .B2(n18455), .ZN(
        n18442) );
  OAI22_X1 U21509 ( .A1(n18439), .A2(n18693), .B1(n18480), .B2(n18620), .ZN(
        n18440) );
  OAI21_X1 U21510 ( .B1(n18519), .B2(n18983), .A(n18440), .ZN(n18456) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18456), .B1(
        n18754), .B2(n18519), .ZN(n18441) );
  OAI211_X1 U21512 ( .C1(n18697), .C2(n18789), .A(n18442), .B(n18441), .ZN(
        P3_U2884) );
  INV_X1 U21513 ( .A(n18519), .ZN(n18518) );
  AOI22_X1 U21514 ( .A1(n18760), .A2(n18801), .B1(n18758), .B2(n18455), .ZN(
        n18444) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18456), .B1(
        n18759), .B2(n18475), .ZN(n18443) );
  OAI211_X1 U21516 ( .C1(n18763), .C2(n18518), .A(n18444), .B(n18443), .ZN(
        P3_U2885) );
  AOI22_X1 U21517 ( .A1(n18765), .A2(n18801), .B1(n18764), .B2(n18455), .ZN(
        n18446) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18456), .B1(
        n18766), .B2(n18519), .ZN(n18445) );
  OAI211_X1 U21519 ( .C1(n18770), .C2(n18474), .A(n18446), .B(n18445), .ZN(
        P3_U2886) );
  AOI22_X1 U21520 ( .A1(n18773), .A2(n18801), .B1(n18772), .B2(n18455), .ZN(
        n18448) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18456), .B1(
        n18771), .B2(n18475), .ZN(n18447) );
  OAI211_X1 U21522 ( .C1(n18776), .C2(n18518), .A(n18448), .B(n18447), .ZN(
        P3_U2887) );
  AOI22_X1 U21523 ( .A1(n18778), .A2(n18801), .B1(n18777), .B2(n18455), .ZN(
        n18450) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18456), .B1(
        n18779), .B2(n18475), .ZN(n18449) );
  OAI211_X1 U21525 ( .C1(n18782), .C2(n18518), .A(n18450), .B(n18449), .ZN(
        P3_U2888) );
  AOI22_X1 U21526 ( .A1(n18786), .A2(n18475), .B1(n18783), .B2(n18455), .ZN(
        n18452) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18456), .B1(
        n18784), .B2(n18801), .ZN(n18451) );
  OAI211_X1 U21528 ( .C1(n18790), .C2(n18518), .A(n18452), .B(n18451), .ZN(
        P3_U2889) );
  AOI22_X1 U21529 ( .A1(n18792), .A2(n18475), .B1(n18791), .B2(n18455), .ZN(
        n18454) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18456), .B1(
        n18793), .B2(n18519), .ZN(n18453) );
  OAI211_X1 U21531 ( .C1(n18796), .C2(n18789), .A(n18454), .B(n18453), .ZN(
        P3_U2890) );
  AOI22_X1 U21532 ( .A1(n18798), .A2(n18455), .B1(n18711), .B2(n18801), .ZN(
        n18458) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18456), .B1(
        n18802), .B2(n18519), .ZN(n18457) );
  OAI211_X1 U21534 ( .C1(n18716), .C2(n18474), .A(n18458), .B(n18457), .ZN(
        P3_U2891) );
  INV_X1 U21535 ( .A(n18689), .ZN(n18757) );
  NOR2_X1 U21536 ( .A1(n18747), .A2(n18502), .ZN(n18476) );
  AOI22_X1 U21537 ( .A1(n18748), .A2(n18476), .B1(n18749), .B2(n18475), .ZN(
        n18461) );
  NOR2_X2 U21538 ( .A1(n18834), .A2(n18502), .ZN(n18542) );
  AOI21_X1 U21539 ( .B1(n18833), .B2(n18718), .A(n18620), .ZN(n18548) );
  OAI211_X1 U21540 ( .C1(n18542), .C2(n18983), .A(n18459), .B(n18548), .ZN(
        n18477) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18477), .B1(
        n18754), .B2(n18542), .ZN(n18460) );
  OAI211_X1 U21542 ( .C1(n18757), .C2(n18501), .A(n18461), .B(n18460), .ZN(
        P3_U2892) );
  INV_X1 U21543 ( .A(n18542), .ZN(n18529) );
  AOI22_X1 U21544 ( .A1(n18760), .A2(n18475), .B1(n18758), .B2(n18476), .ZN(
        n18463) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18477), .B1(
        n18759), .B2(n18494), .ZN(n18462) );
  OAI211_X1 U21546 ( .C1(n18763), .C2(n18529), .A(n18463), .B(n18462), .ZN(
        P3_U2893) );
  AOI22_X1 U21547 ( .A1(n18765), .A2(n18475), .B1(n18764), .B2(n18476), .ZN(
        n18465) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18477), .B1(
        n18766), .B2(n18542), .ZN(n18464) );
  OAI211_X1 U21549 ( .C1(n18770), .C2(n18501), .A(n18465), .B(n18464), .ZN(
        P3_U2894) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18477), .B1(
        n18772), .B2(n18476), .ZN(n18467) );
  AOI22_X1 U21551 ( .A1(n18773), .A2(n18475), .B1(n18771), .B2(n18494), .ZN(
        n18466) );
  OAI211_X1 U21552 ( .C1(n18776), .C2(n18529), .A(n18467), .B(n18466), .ZN(
        P3_U2895) );
  AOI22_X1 U21553 ( .A1(n18778), .A2(n18475), .B1(n18777), .B2(n18476), .ZN(
        n18469) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18477), .B1(
        n18779), .B2(n18494), .ZN(n18468) );
  OAI211_X1 U21555 ( .C1(n18782), .C2(n18529), .A(n18469), .B(n18468), .ZN(
        P3_U2896) );
  AOI22_X1 U21556 ( .A1(n18784), .A2(n18475), .B1(n18783), .B2(n18476), .ZN(
        n18471) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18477), .B1(
        n18786), .B2(n18494), .ZN(n18470) );
  OAI211_X1 U21558 ( .C1(n18790), .C2(n18529), .A(n18471), .B(n18470), .ZN(
        P3_U2897) );
  AOI22_X1 U21559 ( .A1(n18792), .A2(n18494), .B1(n18791), .B2(n18476), .ZN(
        n18473) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18477), .B1(
        n18793), .B2(n18542), .ZN(n18472) );
  OAI211_X1 U21561 ( .C1(n18796), .C2(n18474), .A(n18473), .B(n18472), .ZN(
        P3_U2898) );
  AOI22_X1 U21562 ( .A1(n18798), .A2(n18476), .B1(n18711), .B2(n18475), .ZN(
        n18479) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18477), .B1(
        n18802), .B2(n18542), .ZN(n18478) );
  OAI211_X1 U21564 ( .C1(n18716), .C2(n18501), .A(n18479), .B(n18478), .ZN(
        P3_U2899) );
  NOR2_X2 U21565 ( .A1(n18837), .A2(n18547), .ZN(n18567) );
  NOR2_X1 U21566 ( .A1(n18542), .A2(n18567), .ZN(n18525) );
  NOR2_X1 U21567 ( .A1(n18747), .A2(n18525), .ZN(n18497) );
  AOI22_X1 U21568 ( .A1(n18748), .A2(n18497), .B1(n18749), .B2(n18494), .ZN(
        n18483) );
  OAI21_X1 U21569 ( .B1(n18480), .B2(n18718), .A(n18525), .ZN(n18481) );
  OAI211_X1 U21570 ( .C1(n18567), .C2(n18983), .A(n18721), .B(n18481), .ZN(
        n18498) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18498), .B1(
        n18754), .B2(n18567), .ZN(n18482) );
  OAI211_X1 U21572 ( .C1(n18757), .C2(n18518), .A(n18483), .B(n18482), .ZN(
        P3_U2900) );
  INV_X1 U21573 ( .A(n18567), .ZN(n18564) );
  AOI22_X1 U21574 ( .A1(n18759), .A2(n18519), .B1(n18758), .B2(n18497), .ZN(
        n18485) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18498), .B1(
        n18760), .B2(n18494), .ZN(n18484) );
  OAI211_X1 U21576 ( .C1(n18763), .C2(n18564), .A(n18485), .B(n18484), .ZN(
        P3_U2901) );
  AOI22_X1 U21577 ( .A1(n18726), .A2(n18519), .B1(n18764), .B2(n18497), .ZN(
        n18487) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18498), .B1(
        n18766), .B2(n18567), .ZN(n18486) );
  OAI211_X1 U21579 ( .C1(n18729), .C2(n18501), .A(n18487), .B(n18486), .ZN(
        P3_U2902) );
  AOI22_X1 U21580 ( .A1(n18773), .A2(n18494), .B1(n18772), .B2(n18497), .ZN(
        n18489) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18498), .B1(
        n18771), .B2(n18519), .ZN(n18488) );
  OAI211_X1 U21582 ( .C1(n18776), .C2(n18564), .A(n18489), .B(n18488), .ZN(
        P3_U2903) );
  AOI22_X1 U21583 ( .A1(n18778), .A2(n18494), .B1(n18777), .B2(n18497), .ZN(
        n18491) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18498), .B1(
        n18779), .B2(n18519), .ZN(n18490) );
  OAI211_X1 U21585 ( .C1(n18782), .C2(n18564), .A(n18491), .B(n18490), .ZN(
        P3_U2904) );
  AOI22_X1 U21586 ( .A1(n18786), .A2(n18519), .B1(n18783), .B2(n18497), .ZN(
        n18493) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18498), .B1(
        n18784), .B2(n18494), .ZN(n18492) );
  OAI211_X1 U21588 ( .C1(n18790), .C2(n18564), .A(n18493), .B(n18492), .ZN(
        P3_U2905) );
  AOI22_X1 U21589 ( .A1(n18791), .A2(n18497), .B1(n18679), .B2(n18494), .ZN(
        n18496) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18498), .B1(
        n18793), .B2(n18567), .ZN(n18495) );
  OAI211_X1 U21591 ( .C1(n18682), .C2(n18518), .A(n18496), .B(n18495), .ZN(
        P3_U2906) );
  AOI22_X1 U21592 ( .A1(n18800), .A2(n18519), .B1(n18798), .B2(n18497), .ZN(
        n18500) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18498), .B1(
        n18802), .B2(n18567), .ZN(n18499) );
  OAI211_X1 U21594 ( .C1(n18806), .C2(n18501), .A(n18500), .B(n18499), .ZN(
        P3_U2907) );
  NOR2_X1 U21595 ( .A1(n18547), .A2(n18688), .ZN(n18520) );
  AOI22_X1 U21596 ( .A1(n18689), .A2(n18542), .B1(n18748), .B2(n18520), .ZN(
        n18505) );
  OAI22_X1 U21597 ( .A1(n18693), .A2(n18502), .B1(n18547), .B2(n18690), .ZN(
        n18503) );
  INV_X1 U21598 ( .A(n18503), .ZN(n18521) );
  NOR2_X2 U21599 ( .A1(n18594), .A2(n18547), .ZN(n18584) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18521), .B1(
        n18754), .B2(n18584), .ZN(n18504) );
  OAI211_X1 U21601 ( .C1(n18697), .C2(n18518), .A(n18505), .B(n18504), .ZN(
        P3_U2908) );
  INV_X1 U21602 ( .A(n18584), .ZN(n18592) );
  AOI22_X1 U21603 ( .A1(n18760), .A2(n18519), .B1(n18758), .B2(n18520), .ZN(
        n18507) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18521), .B1(
        n18759), .B2(n18542), .ZN(n18506) );
  OAI211_X1 U21605 ( .C1(n18763), .C2(n18592), .A(n18507), .B(n18506), .ZN(
        P3_U2909) );
  AOI22_X1 U21606 ( .A1(n18726), .A2(n18542), .B1(n18764), .B2(n18520), .ZN(
        n18509) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18521), .B1(
        n18766), .B2(n18584), .ZN(n18508) );
  OAI211_X1 U21608 ( .C1(n18729), .C2(n18518), .A(n18509), .B(n18508), .ZN(
        P3_U2910) );
  AOI22_X1 U21609 ( .A1(n18772), .A2(n18520), .B1(n18771), .B2(n18542), .ZN(
        n18511) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18521), .B1(
        n18773), .B2(n18519), .ZN(n18510) );
  OAI211_X1 U21611 ( .C1(n18776), .C2(n18592), .A(n18511), .B(n18510), .ZN(
        P3_U2911) );
  AOI22_X1 U21612 ( .A1(n18778), .A2(n18519), .B1(n18777), .B2(n18520), .ZN(
        n18513) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18521), .B1(
        n18779), .B2(n18542), .ZN(n18512) );
  OAI211_X1 U21614 ( .C1(n18782), .C2(n18592), .A(n18513), .B(n18512), .ZN(
        P3_U2912) );
  AOI22_X1 U21615 ( .A1(n18784), .A2(n18519), .B1(n18783), .B2(n18520), .ZN(
        n18515) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18521), .B1(
        n18786), .B2(n18542), .ZN(n18514) );
  OAI211_X1 U21617 ( .C1(n18790), .C2(n18592), .A(n18515), .B(n18514), .ZN(
        P3_U2913) );
  AOI22_X1 U21618 ( .A1(n18792), .A2(n18542), .B1(n18791), .B2(n18520), .ZN(
        n18517) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18521), .B1(
        n18793), .B2(n18584), .ZN(n18516) );
  OAI211_X1 U21620 ( .C1(n18796), .C2(n18518), .A(n18517), .B(n18516), .ZN(
        P3_U2914) );
  AOI22_X1 U21621 ( .A1(n18798), .A2(n18520), .B1(n18711), .B2(n18519), .ZN(
        n18523) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18521), .B1(
        n18802), .B2(n18584), .ZN(n18522) );
  OAI211_X1 U21623 ( .C1(n18716), .C2(n18529), .A(n18523), .B(n18522), .ZN(
        P3_U2915) );
  NAND2_X1 U21624 ( .A1(n18524), .A2(n18858), .ZN(n18593) );
  NOR2_X1 U21625 ( .A1(n18584), .A2(n18608), .ZN(n18570) );
  NOR2_X1 U21626 ( .A1(n18747), .A2(n18570), .ZN(n18543) );
  AOI22_X1 U21627 ( .A1(n18689), .A2(n18567), .B1(n18748), .B2(n18543), .ZN(
        n18528) );
  OAI22_X1 U21628 ( .A1(n18525), .A2(n18693), .B1(n18570), .B2(n18620), .ZN(
        n18526) );
  OAI21_X1 U21629 ( .B1(n18608), .B2(n18983), .A(n18526), .ZN(n18544) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18544), .B1(
        n18754), .B2(n18608), .ZN(n18527) );
  OAI211_X1 U21631 ( .C1(n18697), .C2(n18529), .A(n18528), .B(n18527), .ZN(
        P3_U2916) );
  INV_X1 U21632 ( .A(n18608), .ZN(n18587) );
  AOI22_X1 U21633 ( .A1(n18760), .A2(n18542), .B1(n18758), .B2(n18543), .ZN(
        n18531) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18544), .B1(
        n18759), .B2(n18567), .ZN(n18530) );
  OAI211_X1 U21635 ( .C1(n18763), .C2(n18587), .A(n18531), .B(n18530), .ZN(
        P3_U2917) );
  AOI22_X1 U21636 ( .A1(n18765), .A2(n18542), .B1(n18764), .B2(n18543), .ZN(
        n18533) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18544), .B1(
        n18766), .B2(n18608), .ZN(n18532) );
  OAI211_X1 U21638 ( .C1(n18770), .C2(n18564), .A(n18533), .B(n18532), .ZN(
        P3_U2918) );
  AOI22_X1 U21639 ( .A1(n18772), .A2(n18543), .B1(n18771), .B2(n18567), .ZN(
        n18535) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18544), .B1(
        n18773), .B2(n18542), .ZN(n18534) );
  OAI211_X1 U21641 ( .C1(n18776), .C2(n18587), .A(n18535), .B(n18534), .ZN(
        P3_U2919) );
  AOI22_X1 U21642 ( .A1(n18778), .A2(n18542), .B1(n18777), .B2(n18543), .ZN(
        n18537) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18544), .B1(
        n18779), .B2(n18567), .ZN(n18536) );
  OAI211_X1 U21644 ( .C1(n18782), .C2(n18587), .A(n18537), .B(n18536), .ZN(
        P3_U2920) );
  AOI22_X1 U21645 ( .A1(n18786), .A2(n18567), .B1(n18783), .B2(n18543), .ZN(
        n18539) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18544), .B1(
        n18784), .B2(n18542), .ZN(n18538) );
  OAI211_X1 U21647 ( .C1(n18790), .C2(n18587), .A(n18539), .B(n18538), .ZN(
        P3_U2921) );
  AOI22_X1 U21648 ( .A1(n18791), .A2(n18543), .B1(n18679), .B2(n18542), .ZN(
        n18541) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18544), .B1(
        n18793), .B2(n18608), .ZN(n18540) );
  OAI211_X1 U21650 ( .C1(n18682), .C2(n18564), .A(n18541), .B(n18540), .ZN(
        P3_U2922) );
  AOI22_X1 U21651 ( .A1(n18798), .A2(n18543), .B1(n18711), .B2(n18542), .ZN(
        n18546) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18544), .B1(
        n18802), .B2(n18608), .ZN(n18545) );
  OAI211_X1 U21653 ( .C1(n18716), .C2(n18564), .A(n18546), .B(n18545), .ZN(
        P3_U2923) );
  NOR2_X1 U21654 ( .A1(n18747), .A2(n18593), .ZN(n18565) );
  AOI22_X1 U21655 ( .A1(n18689), .A2(n18584), .B1(n18748), .B2(n18565), .ZN(
        n18551) );
  NOR2_X2 U21656 ( .A1(n18834), .A2(n18593), .ZN(n18634) );
  INV_X1 U21657 ( .A(n18547), .ZN(n18549) );
  OAI211_X1 U21658 ( .C1(n18634), .C2(n18983), .A(n18549), .B(n18548), .ZN(
        n18566) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18566), .B1(
        n18754), .B2(n18634), .ZN(n18550) );
  OAI211_X1 U21660 ( .C1(n18697), .C2(n18564), .A(n18551), .B(n18550), .ZN(
        P3_U2924) );
  INV_X1 U21661 ( .A(n18634), .ZN(n18641) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18566), .B1(
        n18758), .B2(n18565), .ZN(n18553) );
  AOI22_X1 U21663 ( .A1(n18760), .A2(n18567), .B1(n18759), .B2(n18584), .ZN(
        n18552) );
  OAI211_X1 U21664 ( .C1(n18763), .C2(n18641), .A(n18553), .B(n18552), .ZN(
        P3_U2925) );
  AOI22_X1 U21665 ( .A1(n18726), .A2(n18584), .B1(n18764), .B2(n18565), .ZN(
        n18555) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18566), .B1(
        n18766), .B2(n18634), .ZN(n18554) );
  OAI211_X1 U21667 ( .C1(n18729), .C2(n18564), .A(n18555), .B(n18554), .ZN(
        P3_U2926) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18566), .B1(
        n18772), .B2(n18565), .ZN(n18557) );
  AOI22_X1 U21669 ( .A1(n18773), .A2(n18567), .B1(n18771), .B2(n18584), .ZN(
        n18556) );
  OAI211_X1 U21670 ( .C1(n18776), .C2(n18641), .A(n18557), .B(n18556), .ZN(
        P3_U2927) );
  AOI22_X1 U21671 ( .A1(n18779), .A2(n18584), .B1(n18777), .B2(n18565), .ZN(
        n18559) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18566), .B1(
        n18778), .B2(n18567), .ZN(n18558) );
  OAI211_X1 U21673 ( .C1(n18782), .C2(n18641), .A(n18559), .B(n18558), .ZN(
        P3_U2928) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18566), .B1(
        n18783), .B2(n18565), .ZN(n18561) );
  AOI22_X1 U21675 ( .A1(n18784), .A2(n18567), .B1(n18786), .B2(n18584), .ZN(
        n18560) );
  OAI211_X1 U21676 ( .C1(n18790), .C2(n18641), .A(n18561), .B(n18560), .ZN(
        P3_U2929) );
  AOI22_X1 U21677 ( .A1(n18792), .A2(n18584), .B1(n18791), .B2(n18565), .ZN(
        n18563) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18566), .B1(
        n18793), .B2(n18634), .ZN(n18562) );
  OAI211_X1 U21679 ( .C1(n18796), .C2(n18564), .A(n18563), .B(n18562), .ZN(
        P3_U2930) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18566), .B1(
        n18798), .B2(n18565), .ZN(n18569) );
  AOI22_X1 U21681 ( .A1(n18802), .A2(n18634), .B1(n18711), .B2(n18567), .ZN(
        n18568) );
  OAI211_X1 U21682 ( .C1(n18716), .C2(n18592), .A(n18569), .B(n18568), .ZN(
        P3_U2931) );
  NOR2_X2 U21683 ( .A1(n18837), .A2(n18618), .ZN(n18659) );
  NOR2_X1 U21684 ( .A1(n18634), .A2(n18659), .ZN(n18619) );
  NOR2_X1 U21685 ( .A1(n18747), .A2(n18619), .ZN(n18588) );
  AOI22_X1 U21686 ( .A1(n18689), .A2(n18608), .B1(n18748), .B2(n18588), .ZN(
        n18573) );
  OAI21_X1 U21687 ( .B1(n18570), .B2(n18718), .A(n18619), .ZN(n18571) );
  OAI211_X1 U21688 ( .C1(n18659), .C2(n18983), .A(n18721), .B(n18571), .ZN(
        n18589) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18589), .B1(
        n18754), .B2(n18659), .ZN(n18572) );
  OAI211_X1 U21690 ( .C1(n18697), .C2(n18592), .A(n18573), .B(n18572), .ZN(
        P3_U2932) );
  INV_X1 U21691 ( .A(n18659), .ZN(n18650) );
  AOI22_X1 U21692 ( .A1(n18760), .A2(n18584), .B1(n18758), .B2(n18588), .ZN(
        n18575) );
  AOI22_X1 U21693 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18589), .B1(
        n18759), .B2(n18608), .ZN(n18574) );
  OAI211_X1 U21694 ( .C1(n18763), .C2(n18650), .A(n18575), .B(n18574), .ZN(
        P3_U2933) );
  AOI22_X1 U21695 ( .A1(n18765), .A2(n18584), .B1(n18764), .B2(n18588), .ZN(
        n18577) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18589), .B1(
        n18766), .B2(n18659), .ZN(n18576) );
  OAI211_X1 U21697 ( .C1(n18770), .C2(n18587), .A(n18577), .B(n18576), .ZN(
        P3_U2934) );
  AOI22_X1 U21698 ( .A1(n18773), .A2(n18584), .B1(n18772), .B2(n18588), .ZN(
        n18579) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18589), .B1(
        n18771), .B2(n18608), .ZN(n18578) );
  OAI211_X1 U21700 ( .C1(n18776), .C2(n18650), .A(n18579), .B(n18578), .ZN(
        P3_U2935) );
  AOI22_X1 U21701 ( .A1(n18779), .A2(n18608), .B1(n18777), .B2(n18588), .ZN(
        n18581) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18589), .B1(
        n18778), .B2(n18584), .ZN(n18580) );
  OAI211_X1 U21703 ( .C1(n18782), .C2(n18650), .A(n18581), .B(n18580), .ZN(
        P3_U2936) );
  AOI22_X1 U21704 ( .A1(n18786), .A2(n18608), .B1(n18783), .B2(n18588), .ZN(
        n18583) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18589), .B1(
        n18784), .B2(n18584), .ZN(n18582) );
  OAI211_X1 U21706 ( .C1(n18790), .C2(n18650), .A(n18583), .B(n18582), .ZN(
        P3_U2937) );
  AOI22_X1 U21707 ( .A1(n18791), .A2(n18588), .B1(n18679), .B2(n18584), .ZN(
        n18586) );
  AOI22_X1 U21708 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18589), .B1(
        n18793), .B2(n18659), .ZN(n18585) );
  OAI211_X1 U21709 ( .C1(n18682), .C2(n18587), .A(n18586), .B(n18585), .ZN(
        P3_U2938) );
  AOI22_X1 U21710 ( .A1(n18800), .A2(n18608), .B1(n18798), .B2(n18588), .ZN(
        n18591) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18589), .B1(
        n18802), .B2(n18659), .ZN(n18590) );
  OAI211_X1 U21712 ( .C1(n18806), .C2(n18592), .A(n18591), .B(n18590), .ZN(
        P3_U2939) );
  OAI22_X1 U21713 ( .A1(n18693), .A2(n18593), .B1(n18618), .B2(n18690), .ZN(
        n18613) );
  NOR2_X1 U21714 ( .A1(n18618), .A2(n18688), .ZN(n18643) );
  AOI22_X1 U21715 ( .A1(n18748), .A2(n18643), .B1(n18749), .B2(n18608), .ZN(
        n18596) );
  NOR2_X2 U21716 ( .A1(n18618), .A2(n18594), .ZN(n18684) );
  AOI22_X1 U21717 ( .A1(n18689), .A2(n18634), .B1(n18684), .B2(n18754), .ZN(
        n18595) );
  OAI211_X1 U21718 ( .C1(n18597), .C2(n18613), .A(n18596), .B(n18595), .ZN(
        P3_U2940) );
  AOI22_X1 U21719 ( .A1(n18760), .A2(n18608), .B1(n18758), .B2(n18643), .ZN(
        n18600) );
  AOI22_X1 U21720 ( .A1(n18684), .A2(n18598), .B1(n18759), .B2(n18634), .ZN(
        n18599) );
  OAI211_X1 U21721 ( .C1(n18601), .C2(n18613), .A(n18600), .B(n18599), .ZN(
        P3_U2941) );
  AOI22_X1 U21722 ( .A1(n18765), .A2(n18608), .B1(n18764), .B2(n18643), .ZN(
        n18603) );
  INV_X1 U21723 ( .A(n18613), .ZN(n18615) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18615), .B1(
        n18684), .B2(n18766), .ZN(n18602) );
  OAI211_X1 U21725 ( .C1(n18770), .C2(n18641), .A(n18603), .B(n18602), .ZN(
        P3_U2942) );
  INV_X1 U21726 ( .A(n18684), .ZN(n18664) );
  AOI22_X1 U21727 ( .A1(n18773), .A2(n18608), .B1(n18772), .B2(n18643), .ZN(
        n18605) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18615), .B1(
        n18771), .B2(n18634), .ZN(n18604) );
  OAI211_X1 U21729 ( .C1(n18664), .C2(n18776), .A(n18605), .B(n18604), .ZN(
        P3_U2943) );
  AOI22_X1 U21730 ( .A1(n18778), .A2(n18608), .B1(n18777), .B2(n18643), .ZN(
        n18607) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18615), .B1(
        n18779), .B2(n18634), .ZN(n18606) );
  OAI211_X1 U21732 ( .C1(n18664), .C2(n18782), .A(n18607), .B(n18606), .ZN(
        P3_U2944) );
  AOI22_X1 U21733 ( .A1(n18786), .A2(n18634), .B1(n18783), .B2(n18643), .ZN(
        n18610) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18615), .B1(
        n18784), .B2(n18608), .ZN(n18609) );
  OAI211_X1 U21735 ( .C1(n18664), .C2(n18790), .A(n18610), .B(n18609), .ZN(
        P3_U2945) );
  AOI22_X1 U21736 ( .A1(n18792), .A2(n18634), .B1(n18791), .B2(n18643), .ZN(
        n18612) );
  AOI22_X1 U21737 ( .A1(n18684), .A2(n18793), .B1(n18679), .B2(n18608), .ZN(
        n18611) );
  OAI211_X1 U21738 ( .C1(n18614), .C2(n18613), .A(n18612), .B(n18611), .ZN(
        P3_U2946) );
  AOI22_X1 U21739 ( .A1(n18798), .A2(n18643), .B1(n18711), .B2(n18608), .ZN(
        n18617) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18615), .B1(
        n18684), .B2(n18802), .ZN(n18616) );
  OAI211_X1 U21741 ( .C1(n18716), .C2(n18641), .A(n18617), .B(n18616), .ZN(
        P3_U2947) );
  NOR2_X1 U21742 ( .A1(n18833), .A2(n18618), .ZN(n18642) );
  INV_X1 U21743 ( .A(n18642), .ZN(n18692) );
  NOR2_X2 U21744 ( .A1(n18692), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18712) );
  NOR2_X1 U21745 ( .A1(n18712), .A2(n18684), .ZN(n18665) );
  NOR2_X1 U21746 ( .A1(n18665), .A2(n18747), .ZN(n18637) );
  AOI22_X1 U21747 ( .A1(n18689), .A2(n18659), .B1(n18748), .B2(n18637), .ZN(
        n18623) );
  OAI22_X1 U21748 ( .A1(n18665), .A2(n18620), .B1(n18619), .B2(n18693), .ZN(
        n18621) );
  OAI21_X1 U21749 ( .B1(n18712), .B2(n18983), .A(n18621), .ZN(n18638) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18638), .B1(
        n18712), .B2(n18754), .ZN(n18622) );
  OAI211_X1 U21751 ( .C1(n18697), .C2(n18641), .A(n18623), .B(n18622), .ZN(
        P3_U2948) );
  INV_X1 U21752 ( .A(n18712), .ZN(n18710) );
  AOI22_X1 U21753 ( .A1(n18760), .A2(n18634), .B1(n18758), .B2(n18637), .ZN(
        n18625) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18638), .B1(
        n18759), .B2(n18659), .ZN(n18624) );
  OAI211_X1 U21755 ( .C1(n18710), .C2(n18763), .A(n18625), .B(n18624), .ZN(
        P3_U2949) );
  AOI22_X1 U21756 ( .A1(n18765), .A2(n18634), .B1(n18764), .B2(n18637), .ZN(
        n18627) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18638), .B1(
        n18712), .B2(n18766), .ZN(n18626) );
  OAI211_X1 U21758 ( .C1(n18770), .C2(n18650), .A(n18627), .B(n18626), .ZN(
        P3_U2950) );
  AOI22_X1 U21759 ( .A1(n18772), .A2(n18637), .B1(n18771), .B2(n18659), .ZN(
        n18629) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18638), .B1(
        n18773), .B2(n18634), .ZN(n18628) );
  OAI211_X1 U21761 ( .C1(n18710), .C2(n18776), .A(n18629), .B(n18628), .ZN(
        P3_U2951) );
  AOI22_X1 U21762 ( .A1(n18779), .A2(n18659), .B1(n18777), .B2(n18637), .ZN(
        n18631) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18638), .B1(
        n18778), .B2(n18634), .ZN(n18630) );
  OAI211_X1 U21764 ( .C1(n18710), .C2(n18782), .A(n18631), .B(n18630), .ZN(
        P3_U2952) );
  AOI22_X1 U21765 ( .A1(n18786), .A2(n18659), .B1(n18783), .B2(n18637), .ZN(
        n18633) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18638), .B1(
        n18784), .B2(n18634), .ZN(n18632) );
  OAI211_X1 U21767 ( .C1(n18710), .C2(n18790), .A(n18633), .B(n18632), .ZN(
        P3_U2953) );
  AOI22_X1 U21768 ( .A1(n18791), .A2(n18637), .B1(n18679), .B2(n18634), .ZN(
        n18636) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18638), .B1(
        n18712), .B2(n18793), .ZN(n18635) );
  OAI211_X1 U21770 ( .C1(n18682), .C2(n18650), .A(n18636), .B(n18635), .ZN(
        P3_U2954) );
  AOI22_X1 U21771 ( .A1(n18800), .A2(n18659), .B1(n18798), .B2(n18637), .ZN(
        n18640) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18638), .B1(
        n18712), .B2(n18802), .ZN(n18639) );
  OAI211_X1 U21773 ( .C1(n18806), .C2(n18641), .A(n18640), .B(n18639), .ZN(
        P3_U2955) );
  NOR2_X1 U21774 ( .A1(n18747), .A2(n18692), .ZN(n18660) );
  AOI22_X1 U21775 ( .A1(n18689), .A2(n18684), .B1(n18748), .B2(n18660), .ZN(
        n18645) );
  AOI22_X1 U21776 ( .A1(n18753), .A2(n18643), .B1(n18642), .B2(n18750), .ZN(
        n18661) );
  NOR2_X2 U21777 ( .A1(n18834), .A2(n18692), .ZN(n18734) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18661), .B1(
        n18734), .B2(n18754), .ZN(n18644) );
  OAI211_X1 U21779 ( .C1(n18697), .C2(n18650), .A(n18645), .B(n18644), .ZN(
        P3_U2956) );
  INV_X1 U21780 ( .A(n18734), .ZN(n18745) );
  AOI22_X1 U21781 ( .A1(n18684), .A2(n18759), .B1(n18758), .B2(n18660), .ZN(
        n18647) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18661), .B1(
        n18760), .B2(n18659), .ZN(n18646) );
  OAI211_X1 U21783 ( .C1(n18745), .C2(n18763), .A(n18647), .B(n18646), .ZN(
        P3_U2957) );
  AOI22_X1 U21784 ( .A1(n18684), .A2(n18726), .B1(n18764), .B2(n18660), .ZN(
        n18649) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18661), .B1(
        n18734), .B2(n18766), .ZN(n18648) );
  OAI211_X1 U21786 ( .C1(n18729), .C2(n18650), .A(n18649), .B(n18648), .ZN(
        P3_U2958) );
  AOI22_X1 U21787 ( .A1(n18773), .A2(n18659), .B1(n18772), .B2(n18660), .ZN(
        n18652) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18661), .B1(
        n18684), .B2(n18771), .ZN(n18651) );
  OAI211_X1 U21789 ( .C1(n18745), .C2(n18776), .A(n18652), .B(n18651), .ZN(
        P3_U2959) );
  AOI22_X1 U21790 ( .A1(n18684), .A2(n18779), .B1(n18777), .B2(n18660), .ZN(
        n18654) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18661), .B1(
        n18778), .B2(n18659), .ZN(n18653) );
  OAI211_X1 U21792 ( .C1(n18745), .C2(n18782), .A(n18654), .B(n18653), .ZN(
        P3_U2960) );
  AOI22_X1 U21793 ( .A1(n18784), .A2(n18659), .B1(n18783), .B2(n18660), .ZN(
        n18656) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18661), .B1(
        n18684), .B2(n18786), .ZN(n18655) );
  OAI211_X1 U21795 ( .C1(n18745), .C2(n18790), .A(n18656), .B(n18655), .ZN(
        P3_U2961) );
  AOI22_X1 U21796 ( .A1(n18791), .A2(n18660), .B1(n18679), .B2(n18659), .ZN(
        n18658) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18661), .B1(
        n18734), .B2(n18793), .ZN(n18657) );
  OAI211_X1 U21798 ( .C1(n18664), .C2(n18682), .A(n18658), .B(n18657), .ZN(
        P3_U2962) );
  AOI22_X1 U21799 ( .A1(n18798), .A2(n18660), .B1(n18711), .B2(n18659), .ZN(
        n18663) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18661), .B1(
        n18734), .B2(n18802), .ZN(n18662) );
  OAI211_X1 U21801 ( .C1(n18664), .C2(n18716), .A(n18663), .B(n18662), .ZN(
        P3_U2963) );
  NOR2_X2 U21802 ( .A1(n18837), .A2(n18691), .ZN(n18785) );
  INV_X1 U21803 ( .A(n18785), .ZN(n18807) );
  AOI21_X1 U21804 ( .B1(n18807), .B2(n18745), .A(n18747), .ZN(n18683) );
  AOI22_X1 U21805 ( .A1(n18684), .A2(n18749), .B1(n18748), .B2(n18683), .ZN(
        n18668) );
  AOI221_X1 U21806 ( .B1(n18665), .B2(n18745), .C1(n18718), .C2(n18745), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18666) );
  OAI21_X1 U21807 ( .B1(n18785), .B2(n18666), .A(n18721), .ZN(n18685) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18685), .B1(
        n18785), .B2(n18754), .ZN(n18667) );
  OAI211_X1 U21809 ( .C1(n18757), .C2(n18710), .A(n18668), .B(n18667), .ZN(
        P3_U2964) );
  AOI22_X1 U21810 ( .A1(n18712), .A2(n18759), .B1(n18683), .B2(n18758), .ZN(
        n18670) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18685), .B1(
        n18684), .B2(n18760), .ZN(n18669) );
  OAI211_X1 U21812 ( .C1(n18807), .C2(n18763), .A(n18670), .B(n18669), .ZN(
        P3_U2965) );
  AOI22_X1 U21813 ( .A1(n18684), .A2(n18765), .B1(n18683), .B2(n18764), .ZN(
        n18672) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18685), .B1(
        n18785), .B2(n18766), .ZN(n18671) );
  OAI211_X1 U21815 ( .C1(n18710), .C2(n18770), .A(n18672), .B(n18671), .ZN(
        P3_U2966) );
  AOI22_X1 U21816 ( .A1(n18712), .A2(n18771), .B1(n18683), .B2(n18772), .ZN(
        n18674) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18685), .B1(
        n18684), .B2(n18773), .ZN(n18673) );
  OAI211_X1 U21818 ( .C1(n18807), .C2(n18776), .A(n18674), .B(n18673), .ZN(
        P3_U2967) );
  AOI22_X1 U21819 ( .A1(n18712), .A2(n18779), .B1(n18683), .B2(n18777), .ZN(
        n18676) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18685), .B1(
        n18684), .B2(n18778), .ZN(n18675) );
  OAI211_X1 U21821 ( .C1(n18807), .C2(n18782), .A(n18676), .B(n18675), .ZN(
        P3_U2968) );
  AOI22_X1 U21822 ( .A1(n18712), .A2(n18786), .B1(n18683), .B2(n18783), .ZN(
        n18678) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18685), .B1(
        n18684), .B2(n18784), .ZN(n18677) );
  OAI211_X1 U21824 ( .C1(n18807), .C2(n18790), .A(n18678), .B(n18677), .ZN(
        P3_U2969) );
  AOI22_X1 U21825 ( .A1(n18684), .A2(n18679), .B1(n18683), .B2(n18791), .ZN(
        n18681) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18685), .B1(
        n18785), .B2(n18793), .ZN(n18680) );
  OAI211_X1 U21827 ( .C1(n18710), .C2(n18682), .A(n18681), .B(n18680), .ZN(
        P3_U2970) );
  AOI22_X1 U21828 ( .A1(n18684), .A2(n18711), .B1(n18683), .B2(n18798), .ZN(
        n18687) );
  AOI22_X1 U21829 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18685), .B1(
        n18785), .B2(n18802), .ZN(n18686) );
  OAI211_X1 U21830 ( .C1(n18710), .C2(n18716), .A(n18687), .B(n18686), .ZN(
        P3_U2971) );
  NOR2_X1 U21831 ( .A1(n18691), .A2(n18688), .ZN(n18752) );
  AOI22_X1 U21832 ( .A1(n18689), .A2(n18734), .B1(n18748), .B2(n18752), .ZN(
        n18696) );
  OAI22_X1 U21833 ( .A1(n18693), .A2(n18692), .B1(n18691), .B2(n18690), .ZN(
        n18694) );
  INV_X1 U21834 ( .A(n18694), .ZN(n18713) );
  AOI22_X1 U21835 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18713), .B1(
        n18754), .B2(n18799), .ZN(n18695) );
  OAI211_X1 U21836 ( .C1(n18710), .C2(n18697), .A(n18696), .B(n18695), .ZN(
        P3_U2972) );
  AOI22_X1 U21837 ( .A1(n18712), .A2(n18760), .B1(n18758), .B2(n18752), .ZN(
        n18699) );
  AOI22_X1 U21838 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18713), .B1(
        n18734), .B2(n18759), .ZN(n18698) );
  OAI211_X1 U21839 ( .C1(n18763), .C2(n18769), .A(n18699), .B(n18698), .ZN(
        P3_U2973) );
  AOI22_X1 U21840 ( .A1(n18734), .A2(n18726), .B1(n18764), .B2(n18752), .ZN(
        n18701) );
  AOI22_X1 U21841 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18713), .B1(
        n18766), .B2(n18799), .ZN(n18700) );
  OAI211_X1 U21842 ( .C1(n18710), .C2(n18729), .A(n18701), .B(n18700), .ZN(
        P3_U2974) );
  AOI22_X1 U21843 ( .A1(n18734), .A2(n18771), .B1(n18772), .B2(n18752), .ZN(
        n18703) );
  AOI22_X1 U21844 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18713), .B1(
        n18712), .B2(n18773), .ZN(n18702) );
  OAI211_X1 U21845 ( .C1(n18776), .C2(n18769), .A(n18703), .B(n18702), .ZN(
        P3_U2975) );
  AOI22_X1 U21846 ( .A1(n18734), .A2(n18779), .B1(n18777), .B2(n18752), .ZN(
        n18705) );
  AOI22_X1 U21847 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18713), .B1(
        n18712), .B2(n18778), .ZN(n18704) );
  OAI211_X1 U21848 ( .C1(n18782), .C2(n18769), .A(n18705), .B(n18704), .ZN(
        P3_U2976) );
  AOI22_X1 U21849 ( .A1(n18712), .A2(n18784), .B1(n18783), .B2(n18752), .ZN(
        n18707) );
  AOI22_X1 U21850 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18713), .B1(
        n18734), .B2(n18786), .ZN(n18706) );
  OAI211_X1 U21851 ( .C1(n18790), .C2(n18769), .A(n18707), .B(n18706), .ZN(
        P3_U2977) );
  AOI22_X1 U21852 ( .A1(n18734), .A2(n18792), .B1(n18791), .B2(n18752), .ZN(
        n18709) );
  AOI22_X1 U21853 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18713), .B1(
        n18793), .B2(n18799), .ZN(n18708) );
  OAI211_X1 U21854 ( .C1(n18710), .C2(n18796), .A(n18709), .B(n18708), .ZN(
        P3_U2978) );
  AOI22_X1 U21855 ( .A1(n18712), .A2(n18711), .B1(n18798), .B2(n18752), .ZN(
        n18715) );
  AOI22_X1 U21856 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18713), .B1(
        n18802), .B2(n18799), .ZN(n18714) );
  OAI211_X1 U21857 ( .C1(n18745), .C2(n18716), .A(n18715), .B(n18714), .ZN(
        P3_U2979) );
  NOR2_X1 U21858 ( .A1(n18747), .A2(n18717), .ZN(n18740) );
  AOI22_X1 U21859 ( .A1(n18734), .A2(n18749), .B1(n18748), .B2(n18740), .ZN(
        n18723) );
  NOR2_X1 U21860 ( .A1(n18785), .A2(n18734), .ZN(n18719) );
  OAI21_X1 U21861 ( .B1(n18719), .B2(n18718), .A(n18717), .ZN(n18720) );
  OAI211_X1 U21862 ( .C1(n18741), .C2(n18983), .A(n18721), .B(n18720), .ZN(
        n18742) );
  AOI22_X1 U21863 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18742), .B1(
        n18754), .B2(n18741), .ZN(n18722) );
  OAI211_X1 U21864 ( .C1(n18757), .C2(n18807), .A(n18723), .B(n18722), .ZN(
        P3_U2980) );
  AOI22_X1 U21865 ( .A1(n18785), .A2(n18759), .B1(n18758), .B2(n18740), .ZN(
        n18725) );
  AOI22_X1 U21866 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18742), .B1(
        n18734), .B2(n18760), .ZN(n18724) );
  OAI211_X1 U21867 ( .C1(n18763), .C2(n18737), .A(n18725), .B(n18724), .ZN(
        P3_U2981) );
  AOI22_X1 U21868 ( .A1(n18785), .A2(n18726), .B1(n18764), .B2(n18740), .ZN(
        n18728) );
  AOI22_X1 U21869 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18742), .B1(
        n18766), .B2(n18741), .ZN(n18727) );
  OAI211_X1 U21870 ( .C1(n18745), .C2(n18729), .A(n18728), .B(n18727), .ZN(
        P3_U2982) );
  AOI22_X1 U21871 ( .A1(n18734), .A2(n18773), .B1(n18772), .B2(n18740), .ZN(
        n18731) );
  AOI22_X1 U21872 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18742), .B1(
        n18785), .B2(n18771), .ZN(n18730) );
  OAI211_X1 U21873 ( .C1(n18776), .C2(n18737), .A(n18731), .B(n18730), .ZN(
        P3_U2983) );
  AOI22_X1 U21874 ( .A1(n18785), .A2(n18779), .B1(n18777), .B2(n18740), .ZN(
        n18733) );
  AOI22_X1 U21875 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18742), .B1(
        n18734), .B2(n18778), .ZN(n18732) );
  OAI211_X1 U21876 ( .C1(n18782), .C2(n18737), .A(n18733), .B(n18732), .ZN(
        P3_U2984) );
  AOI22_X1 U21877 ( .A1(n18785), .A2(n18786), .B1(n18783), .B2(n18740), .ZN(
        n18736) );
  AOI22_X1 U21878 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18742), .B1(
        n18734), .B2(n18784), .ZN(n18735) );
  OAI211_X1 U21879 ( .C1(n18790), .C2(n18737), .A(n18736), .B(n18735), .ZN(
        P3_U2985) );
  AOI22_X1 U21880 ( .A1(n18785), .A2(n18792), .B1(n18791), .B2(n18740), .ZN(
        n18739) );
  AOI22_X1 U21881 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18742), .B1(
        n18793), .B2(n18741), .ZN(n18738) );
  OAI211_X1 U21882 ( .C1(n18745), .C2(n18796), .A(n18739), .B(n18738), .ZN(
        P3_U2986) );
  AOI22_X1 U21883 ( .A1(n18785), .A2(n18800), .B1(n18798), .B2(n18740), .ZN(
        n18744) );
  AOI22_X1 U21884 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18742), .B1(
        n18802), .B2(n18741), .ZN(n18743) );
  OAI211_X1 U21885 ( .C1(n18745), .C2(n18806), .A(n18744), .B(n18743), .ZN(
        P3_U2987) );
  NOR2_X1 U21886 ( .A1(n18747), .A2(n18746), .ZN(n18797) );
  AOI22_X1 U21887 ( .A1(n18785), .A2(n18749), .B1(n18748), .B2(n18797), .ZN(
        n18756) );
  AOI22_X1 U21888 ( .A1(n18753), .A2(n18752), .B1(n18751), .B2(n18750), .ZN(
        n18803) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18803), .B1(
        n18754), .B2(n18801), .ZN(n18755) );
  OAI211_X1 U21890 ( .C1(n18757), .C2(n18769), .A(n18756), .B(n18755), .ZN(
        P3_U2988) );
  AOI22_X1 U21891 ( .A1(n18759), .A2(n18799), .B1(n18758), .B2(n18797), .ZN(
        n18762) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18803), .B1(
        n18785), .B2(n18760), .ZN(n18761) );
  OAI211_X1 U21893 ( .C1(n18763), .C2(n18789), .A(n18762), .B(n18761), .ZN(
        P3_U2989) );
  AOI22_X1 U21894 ( .A1(n18785), .A2(n18765), .B1(n18764), .B2(n18797), .ZN(
        n18768) );
  AOI22_X1 U21895 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18803), .B1(
        n18766), .B2(n18801), .ZN(n18767) );
  OAI211_X1 U21896 ( .C1(n18770), .C2(n18769), .A(n18768), .B(n18767), .ZN(
        P3_U2990) );
  AOI22_X1 U21897 ( .A1(n18772), .A2(n18797), .B1(n18771), .B2(n18799), .ZN(
        n18775) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18803), .B1(
        n18785), .B2(n18773), .ZN(n18774) );
  OAI211_X1 U21899 ( .C1(n18776), .C2(n18789), .A(n18775), .B(n18774), .ZN(
        P3_U2991) );
  AOI22_X1 U21900 ( .A1(n18785), .A2(n18778), .B1(n18777), .B2(n18797), .ZN(
        n18781) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18803), .B1(
        n18779), .B2(n18799), .ZN(n18780) );
  OAI211_X1 U21902 ( .C1(n18782), .C2(n18789), .A(n18781), .B(n18780), .ZN(
        P3_U2992) );
  AOI22_X1 U21903 ( .A1(n18785), .A2(n18784), .B1(n18783), .B2(n18797), .ZN(
        n18788) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18803), .B1(
        n18786), .B2(n18799), .ZN(n18787) );
  OAI211_X1 U21905 ( .C1(n18790), .C2(n18789), .A(n18788), .B(n18787), .ZN(
        P3_U2993) );
  AOI22_X1 U21906 ( .A1(n18792), .A2(n18799), .B1(n18791), .B2(n18797), .ZN(
        n18795) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18803), .B1(
        n18793), .B2(n18801), .ZN(n18794) );
  OAI211_X1 U21908 ( .C1(n18807), .C2(n18796), .A(n18795), .B(n18794), .ZN(
        P3_U2994) );
  AOI22_X1 U21909 ( .A1(n18800), .A2(n18799), .B1(n18798), .B2(n18797), .ZN(
        n18805) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18803), .B1(
        n18802), .B2(n18801), .ZN(n18804) );
  OAI211_X1 U21911 ( .C1(n18807), .C2(n18806), .A(n18805), .B(n18804), .ZN(
        P3_U2995) );
  NOR2_X1 U21912 ( .A1(n18851), .A2(n18808), .ZN(n18810) );
  OAI222_X1 U21913 ( .A1(n18814), .A2(n18813), .B1(n18812), .B2(n18811), .C1(
        n18810), .C2(n18809), .ZN(n19027) );
  OAI21_X1 U21914 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18815), .ZN(n18816) );
  OAI211_X1 U21915 ( .C1(n21141), .C2(n18852), .A(n18817), .B(n18816), .ZN(
        n18864) );
  NOR2_X1 U21916 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18818), .ZN(
        n18830) );
  INV_X1 U21917 ( .A(n18830), .ZN(n18819) );
  AOI22_X1 U21918 ( .A1(n18851), .A2(n18823), .B1(n18840), .B2(n18819), .ZN(
        n18989) );
  NOR2_X1 U21919 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18989), .ZN(
        n18827) );
  OAI21_X1 U21920 ( .B1(n18822), .B2(n18821), .A(n18820), .ZN(n18838) );
  OAI21_X1 U21921 ( .B1(n18832), .B2(n18840), .A(n18823), .ZN(n18824) );
  AOI21_X1 U21922 ( .B1(n18825), .B2(n18838), .A(n18824), .ZN(n18985) );
  NAND2_X1 U21923 ( .A1(n18852), .A2(n18985), .ZN(n18826) );
  AOI22_X1 U21924 ( .A1(n18852), .A2(n18827), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18826), .ZN(n18862) );
  NOR2_X1 U21925 ( .A1(n18829), .A2(n18828), .ZN(n18831) );
  OAI22_X1 U21926 ( .A1(n18831), .A2(n19001), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18830), .ZN(n19006) );
  AOI22_X1 U21927 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18832), .B1(
        n18831), .B2(n19014), .ZN(n19009) );
  OAI221_X1 U21928 ( .B1(n19006), .B2(n19009), .C1(n19006), .C2(n18833), .A(
        n18852), .ZN(n18836) );
  NOR3_X1 U21929 ( .A1(n19009), .A2(n18834), .A3(n18833), .ZN(n18835) );
  AOI21_X1 U21930 ( .B1(n18837), .B2(n18836), .A(n18835), .ZN(n18856) );
  INV_X1 U21931 ( .A(n18852), .ZN(n18853) );
  AOI21_X1 U21932 ( .B1(n9732), .B2(n18844), .A(n18838), .ZN(n18849) );
  NAND2_X1 U21933 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18839), .ZN(
        n18848) );
  AOI211_X1 U21934 ( .C1(n13063), .C2(n13208), .A(n18841), .B(n18840), .ZN(
        n18842) );
  INV_X1 U21935 ( .A(n18842), .ZN(n18847) );
  NOR2_X1 U21936 ( .A1(n18843), .A2(n19014), .ZN(n18845) );
  OAI211_X1 U21937 ( .C1(n18845), .C2(n18844), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n13063), .ZN(n18846) );
  OAI211_X1 U21938 ( .C1(n18849), .C2(n18848), .A(n18847), .B(n18846), .ZN(
        n18850) );
  AOI21_X1 U21939 ( .B1(n18851), .B2(n18995), .A(n18850), .ZN(n18997) );
  AOI22_X1 U21940 ( .A1(n18853), .A2(n13063), .B1(n18997), .B2(n18852), .ZN(
        n18857) );
  AND2_X1 U21941 ( .A1(n18856), .A2(n18857), .ZN(n18854) );
  OAI221_X1 U21942 ( .B1(n18856), .B2(n18857), .C1(n18855), .C2(n18854), .A(
        n18859), .ZN(n18861) );
  AOI21_X1 U21943 ( .B1(n18859), .B2(n18858), .A(n18857), .ZN(n18860) );
  AOI222_X1 U21944 ( .A1(n18862), .A2(n18861), .B1(n18862), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18861), .C2(n18860), .ZN(
        n18863) );
  NOR4_X1 U21945 ( .A1(n18865), .A2(n19027), .A3(n18864), .A4(n18863), .ZN(
        n18879) );
  NAND3_X1 U21946 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18894), .A3(n18866), 
        .ZN(n18888) );
  OAI211_X1 U21947 ( .C1(n18869), .C2(n18868), .A(n18867), .B(n18879), .ZN(
        n18870) );
  INV_X1 U21948 ( .A(n18870), .ZN(n18881) );
  NOR2_X1 U21949 ( .A1(n18881), .A2(n18871), .ZN(n18984) );
  NAND2_X1 U21950 ( .A1(n18984), .A2(n18872), .ZN(n18876) );
  INV_X1 U21951 ( .A(n18872), .ZN(n18873) );
  AOI22_X1 U21952 ( .A1(n18874), .A2(n18894), .B1(n18873), .B2(n21141), .ZN(
        n18875) );
  OAI22_X1 U21953 ( .A1(n18877), .A2(n18876), .B1(P3_STATE2_REG_0__SCAN_IN), 
        .B2(n18875), .ZN(n18878) );
  OAI211_X1 U21954 ( .C1(n18879), .C2(n18883), .A(n18888), .B(n18878), .ZN(
        P3_U2996) );
  NOR2_X1 U21955 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19034), .ZN(n18880) );
  AOI211_X1 U21956 ( .C1(n18883), .C2(n18882), .A(n18881), .B(n18880), .ZN(
        n18884) );
  AOI211_X1 U21957 ( .C1(n18894), .C2(n19030), .A(n18885), .B(n18884), .ZN(
        n18886) );
  OAI21_X1 U21958 ( .B1(n18887), .B2(n18888), .A(n18886), .ZN(P3_U2997) );
  NOR2_X1 U21959 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATEBS16_REG_SCAN_IN), .ZN(n18892) );
  INV_X1 U21960 ( .A(n18888), .ZN(n18889) );
  AOI221_X1 U21961 ( .B1(n18892), .B2(n18891), .C1(n18890), .C2(n18891), .A(
        n18889), .ZN(P3_U2998) );
  INV_X1 U21962 ( .A(n18981), .ZN(n18893) );
  AND2_X1 U21963 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18893), .ZN(
        P3_U2999) );
  AND2_X1 U21964 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18893), .ZN(
        P3_U3000) );
  AND2_X1 U21965 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18893), .ZN(
        P3_U3001) );
  AND2_X1 U21966 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18893), .ZN(
        P3_U3002) );
  AND2_X1 U21967 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18893), .ZN(
        P3_U3003) );
  AND2_X1 U21968 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18893), .ZN(
        P3_U3004) );
  AND2_X1 U21969 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18893), .ZN(
        P3_U3005) );
  AND2_X1 U21970 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18893), .ZN(
        P3_U3006) );
  AND2_X1 U21971 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18893), .ZN(
        P3_U3007) );
  AND2_X1 U21972 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18893), .ZN(
        P3_U3008) );
  AND2_X1 U21973 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18893), .ZN(
        P3_U3009) );
  AND2_X1 U21974 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18893), .ZN(
        P3_U3010) );
  AND2_X1 U21975 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18893), .ZN(
        P3_U3011) );
  AND2_X1 U21976 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18893), .ZN(
        P3_U3012) );
  AND2_X1 U21977 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18893), .ZN(
        P3_U3013) );
  AND2_X1 U21978 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18893), .ZN(
        P3_U3014) );
  AND2_X1 U21979 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18893), .ZN(
        P3_U3015) );
  AND2_X1 U21980 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18893), .ZN(
        P3_U3016) );
  AND2_X1 U21981 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18893), .ZN(
        P3_U3017) );
  AND2_X1 U21982 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18893), .ZN(
        P3_U3018) );
  AND2_X1 U21983 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18893), .ZN(
        P3_U3019) );
  AND2_X1 U21984 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18893), .ZN(
        P3_U3020) );
  AND2_X1 U21985 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18893), .ZN(P3_U3021) );
  AND2_X1 U21986 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18893), .ZN(P3_U3022) );
  AND2_X1 U21987 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18893), .ZN(P3_U3023) );
  AND2_X1 U21988 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18893), .ZN(P3_U3024) );
  AND2_X1 U21989 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18893), .ZN(P3_U3025) );
  AND2_X1 U21990 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18893), .ZN(P3_U3026) );
  AND2_X1 U21991 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18893), .ZN(P3_U3027) );
  AND2_X1 U21992 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18893), .ZN(P3_U3028) );
  NOR2_X1 U21993 ( .A1(n18903), .A2(n20937), .ZN(n18901) );
  NOR2_X1 U21994 ( .A1(n18913), .A2(n20937), .ZN(n18908) );
  INV_X1 U21995 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18898) );
  NOR3_X1 U21996 ( .A1(n18901), .A2(n18908), .A3(n18898), .ZN(n18897) );
  NAND2_X1 U21997 ( .A1(n18894), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18906) );
  AND2_X1 U21998 ( .A1(n18906), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18912) );
  INV_X1 U21999 ( .A(NA), .ZN(n20930) );
  OAI21_X1 U22000 ( .B1(n20930), .B2(n18895), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18911) );
  INV_X1 U22001 ( .A(n18911), .ZN(n18896) );
  OAI22_X1 U22002 ( .A1(n19041), .A2(n18897), .B1(n18912), .B2(n18896), .ZN(
        P3_U3029) );
  AOI21_X1 U22003 ( .B1(n18899), .B2(HOLD), .A(n18898), .ZN(n18900) );
  AOI21_X1 U22004 ( .B1(n18913), .B2(n18901), .A(n18900), .ZN(n18902) );
  OAI22_X1 U22005 ( .A1(n19034), .A2(n18903), .B1(n18910), .B2(n18902), .ZN(
        n18904) );
  INV_X1 U22006 ( .A(n18904), .ZN(n18905) );
  NAND2_X1 U22007 ( .A1(n18905), .A2(n19031), .ZN(P3_U3030) );
  OAI22_X1 U22008 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18906), .ZN(n18907) );
  OAI22_X1 U22009 ( .A1(n18908), .A2(n18907), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18909) );
  OAI22_X1 U22010 ( .A1(n18912), .A2(n18911), .B1(n18910), .B2(n18909), .ZN(
        P3_U3031) );
  OAI222_X1 U22011 ( .A1(n19016), .A2(n18967), .B1(n18914), .B2(n19041), .C1(
        n18915), .C2(n18964), .ZN(P3_U3032) );
  OAI222_X1 U22012 ( .A1(n18964), .A2(n18917), .B1(n18916), .B2(n19041), .C1(
        n18915), .C2(n18973), .ZN(P3_U3033) );
  OAI222_X1 U22013 ( .A1(n18964), .A2(n18919), .B1(n18918), .B2(n19041), .C1(
        n18917), .C2(n18967), .ZN(P3_U3034) );
  OAI222_X1 U22014 ( .A1(n18964), .A2(n18922), .B1(n18920), .B2(n19041), .C1(
        n18919), .C2(n18967), .ZN(P3_U3035) );
  OAI222_X1 U22015 ( .A1(n18922), .A2(n18967), .B1(n18921), .B2(n19041), .C1(
        n18923), .C2(n18964), .ZN(P3_U3036) );
  OAI222_X1 U22016 ( .A1(n18964), .A2(n18925), .B1(n18924), .B2(n19041), .C1(
        n18923), .C2(n18967), .ZN(P3_U3037) );
  OAI222_X1 U22017 ( .A1(n18964), .A2(n18927), .B1(n18926), .B2(n19041), .C1(
        n18925), .C2(n18967), .ZN(P3_U3038) );
  OAI222_X1 U22018 ( .A1(n18927), .A2(n18967), .B1(n21321), .B2(n19041), .C1(
        n21094), .C2(n18964), .ZN(P3_U3039) );
  OAI222_X1 U22019 ( .A1(n21094), .A2(n18967), .B1(n18928), .B2(n19041), .C1(
        n18929), .C2(n18964), .ZN(P3_U3040) );
  OAI222_X1 U22020 ( .A1(n18964), .A2(n21241), .B1(n18930), .B2(n19041), .C1(
        n18929), .C2(n18967), .ZN(P3_U3041) );
  OAI222_X1 U22021 ( .A1(n18964), .A2(n18932), .B1(n18931), .B2(n19041), .C1(
        n21241), .C2(n18967), .ZN(P3_U3042) );
  OAI222_X1 U22022 ( .A1(n18964), .A2(n18934), .B1(n18933), .B2(n19041), .C1(
        n18932), .C2(n18967), .ZN(P3_U3043) );
  OAI222_X1 U22023 ( .A1(n18964), .A2(n18937), .B1(n18935), .B2(n19041), .C1(
        n18934), .C2(n18967), .ZN(P3_U3044) );
  OAI222_X1 U22024 ( .A1(n18937), .A2(n18967), .B1(n18936), .B2(n19041), .C1(
        n18938), .C2(n18964), .ZN(P3_U3045) );
  OAI222_X1 U22025 ( .A1(n18964), .A2(n18940), .B1(n18939), .B2(n19041), .C1(
        n18938), .C2(n18967), .ZN(P3_U3046) );
  OAI222_X1 U22026 ( .A1(n18964), .A2(n18943), .B1(n18941), .B2(n19041), .C1(
        n18940), .C2(n18973), .ZN(P3_U3047) );
  OAI222_X1 U22027 ( .A1(n18943), .A2(n18967), .B1(n18942), .B2(n19041), .C1(
        n18944), .C2(n18964), .ZN(P3_U3048) );
  OAI222_X1 U22028 ( .A1(n18964), .A2(n18946), .B1(n18945), .B2(n19041), .C1(
        n18944), .C2(n18973), .ZN(P3_U3049) );
  OAI222_X1 U22029 ( .A1(n18964), .A2(n18948), .B1(n18947), .B2(n19041), .C1(
        n18946), .C2(n18973), .ZN(P3_U3050) );
  OAI222_X1 U22030 ( .A1(n18964), .A2(n18950), .B1(n18949), .B2(n19041), .C1(
        n18948), .C2(n18973), .ZN(P3_U3051) );
  INV_X1 U22031 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18952) );
  OAI222_X1 U22032 ( .A1(n18964), .A2(n18952), .B1(n18951), .B2(n19041), .C1(
        n18950), .C2(n18973), .ZN(P3_U3052) );
  OAI222_X1 U22033 ( .A1(n18964), .A2(n18955), .B1(n18953), .B2(n19041), .C1(
        n18952), .C2(n18973), .ZN(P3_U3053) );
  OAI222_X1 U22034 ( .A1(n18955), .A2(n18967), .B1(n18954), .B2(n19041), .C1(
        n18956), .C2(n18964), .ZN(P3_U3054) );
  OAI222_X1 U22035 ( .A1(n18964), .A2(n18958), .B1(n18957), .B2(n19041), .C1(
        n18956), .C2(n18973), .ZN(P3_U3055) );
  INV_X1 U22036 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18960) );
  OAI222_X1 U22037 ( .A1(n18964), .A2(n18960), .B1(n18959), .B2(n19041), .C1(
        n18958), .C2(n18973), .ZN(P3_U3056) );
  OAI222_X1 U22038 ( .A1(n18964), .A2(n18962), .B1(n18961), .B2(n19041), .C1(
        n18960), .C2(n18967), .ZN(P3_U3057) );
  INV_X1 U22039 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18966) );
  OAI222_X1 U22040 ( .A1(n18964), .A2(n18966), .B1(n18963), .B2(n19041), .C1(
        n18962), .C2(n18967), .ZN(P3_U3058) );
  OAI222_X1 U22041 ( .A1(n18966), .A2(n18967), .B1(n18965), .B2(n19041), .C1(
        n18968), .C2(n18964), .ZN(P3_U3059) );
  OAI222_X1 U22042 ( .A1(n18964), .A2(n18972), .B1(n18969), .B2(n19041), .C1(
        n18968), .C2(n18967), .ZN(P3_U3060) );
  OAI222_X1 U22043 ( .A1(n18973), .A2(n18972), .B1(n18971), .B2(n19041), .C1(
        n18970), .C2(n18964), .ZN(P3_U3061) );
  OAI22_X1 U22044 ( .A1(n19042), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19041), .ZN(n18974) );
  INV_X1 U22045 ( .A(n18974), .ZN(P3_U3274) );
  OAI22_X1 U22046 ( .A1(n19042), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19041), .ZN(n18975) );
  INV_X1 U22047 ( .A(n18975), .ZN(P3_U3275) );
  OAI22_X1 U22048 ( .A1(n19042), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19041), .ZN(n18976) );
  INV_X1 U22049 ( .A(n18976), .ZN(P3_U3276) );
  OAI22_X1 U22050 ( .A1(n19042), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19041), .ZN(n18977) );
  INV_X1 U22051 ( .A(n18977), .ZN(P3_U3277) );
  OAI21_X1 U22052 ( .B1(n18981), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18979), 
        .ZN(n18978) );
  INV_X1 U22053 ( .A(n18978), .ZN(P3_U3280) );
  OAI21_X1 U22054 ( .B1(n18981), .B2(n18980), .A(n18979), .ZN(P3_U3281) );
  OAI21_X1 U22055 ( .B1(n18984), .B2(n18983), .A(n18982), .ZN(P3_U3282) );
  OAI21_X1 U22056 ( .B1(n18985), .B2(n18996), .A(n19012), .ZN(n18991) );
  NAND2_X1 U22057 ( .A1(n19010), .A2(n18986), .ZN(n18988) );
  OAI22_X1 U22058 ( .A1(n18989), .A2(n18988), .B1(n19002), .B2(n18987), .ZN(
        n18990) );
  AOI22_X1 U22059 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18991), .B1(
        n19012), .B2(n18990), .ZN(n18992) );
  INV_X1 U22060 ( .A(n18992), .ZN(P3_U3285) );
  AOI22_X1 U22061 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18994), .B2(n18993), .ZN(
        n19004) );
  NAND2_X1 U22062 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19003) );
  INV_X1 U22063 ( .A(n19003), .ZN(n18999) );
  OAI22_X1 U22064 ( .A1(n18997), .A2(n18996), .B1(n19002), .B2(n18995), .ZN(
        n18998) );
  AOI21_X1 U22065 ( .B1(n19004), .B2(n18999), .A(n18998), .ZN(n19000) );
  AOI22_X1 U22066 ( .A1(n19015), .A2(n13063), .B1(n19000), .B2(n19012), .ZN(
        P3_U3288) );
  OAI22_X1 U22067 ( .A1(n19004), .A2(n19003), .B1(n19002), .B2(n19001), .ZN(
        n19005) );
  AOI21_X1 U22068 ( .B1(n19010), .B2(n19006), .A(n19005), .ZN(n19007) );
  AOI22_X1 U22069 ( .A1(n19015), .A2(n13208), .B1(n19007), .B2(n19012), .ZN(
        P3_U3289) );
  AOI222_X1 U22070 ( .A1(n19011), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19010), 
        .B2(n19009), .C1(n19014), .C2(n19008), .ZN(n19013) );
  AOI22_X1 U22071 ( .A1(n19015), .A2(n19014), .B1(n19013), .B2(n19012), .ZN(
        P3_U3290) );
  AOI21_X1 U22072 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19017) );
  AOI22_X1 U22073 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19017), .B2(n19016), .ZN(n19019) );
  INV_X1 U22074 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19018) );
  AOI22_X1 U22075 ( .A1(n19020), .A2(n19019), .B1(n19018), .B2(n19023), .ZN(
        P3_U3292) );
  INV_X1 U22076 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19024) );
  NOR2_X1 U22077 ( .A1(n19023), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19021) );
  AOI22_X1 U22078 ( .A1(n19024), .A2(n19023), .B1(n19022), .B2(n19021), .ZN(
        P3_U3293) );
  INV_X1 U22079 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19025) );
  AOI22_X1 U22080 ( .A1(n19041), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19025), 
        .B2(n19042), .ZN(P3_U3294) );
  MUX2_X1 U22081 ( .A(P3_MORE_REG_SCAN_IN), .B(n19027), .S(n19026), .Z(
        P3_U3295) );
  AOI21_X1 U22082 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n19028), .ZN(n19029) );
  AOI211_X1 U22083 ( .C1(n19030), .C2(n19034), .A(n19029), .B(n19044), .ZN(
        n19040) );
  AOI21_X1 U22084 ( .B1(n19033), .B2(n19032), .A(n19031), .ZN(n19035) );
  OAI211_X1 U22085 ( .C1(n19035), .C2(n19047), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19034), .ZN(n19037) );
  AOI21_X1 U22086 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19037), .A(n19036), 
        .ZN(n19039) );
  NAND2_X1 U22087 ( .A1(n19040), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19038) );
  OAI21_X1 U22088 ( .B1(n19040), .B2(n19039), .A(n19038), .ZN(P3_U3296) );
  OAI22_X1 U22089 ( .A1(n19042), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19041), .ZN(n19043) );
  INV_X1 U22090 ( .A(n19043), .ZN(P3_U3297) );
  OR2_X1 U22091 ( .A1(n19045), .A2(n19044), .ZN(n19050) );
  OAI22_X1 U22092 ( .A1(n19047), .A2(n19046), .B1(n19050), .B2(
        P3_READREQUEST_REG_SCAN_IN), .ZN(n19048) );
  INV_X1 U22093 ( .A(n19048), .ZN(P3_U3298) );
  OAI21_X1 U22094 ( .B1(n19050), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n19049), 
        .ZN(n19051) );
  INV_X1 U22095 ( .A(n19051), .ZN(P3_U3299) );
  INV_X1 U22096 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19058) );
  NAND2_X1 U22097 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19950), .ZN(n19939) );
  NAND2_X1 U22098 ( .A1(n19058), .A2(n19052), .ZN(n19936) );
  OAI21_X1 U22099 ( .B1(n19058), .B2(n19939), .A(n19936), .ZN(n20002) );
  AOI21_X1 U22100 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20002), .ZN(n19053) );
  INV_X1 U22101 ( .A(n19053), .ZN(P2_U2815) );
  INV_X1 U22102 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19056) );
  NAND2_X1 U22103 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20033), .ZN(n19054) );
  OAI22_X1 U22104 ( .A1(n19057), .A2(n19056), .B1(n19055), .B2(n19054), .ZN(
        P2_U2816) );
  NAND2_X1 U22105 ( .A1(n19058), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20053) );
  AOI21_X1 U22106 ( .B1(n19058), .B2(n19950), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19059) );
  AOI22_X1 U22107 ( .A1(n20052), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19059), 
        .B2(n20053), .ZN(P2_U2817) );
  OAI21_X1 U22108 ( .B1(n19943), .B2(BS16), .A(n20002), .ZN(n20000) );
  OAI21_X1 U22109 ( .B1(n20002), .B2(n19691), .A(n20000), .ZN(P2_U2818) );
  NOR4_X1 U22110 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19063) );
  NOR4_X1 U22111 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19062) );
  NOR4_X1 U22112 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19061) );
  NOR4_X1 U22113 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19060) );
  NAND4_X1 U22114 ( .A1(n19063), .A2(n19062), .A3(n19061), .A4(n19060), .ZN(
        n19069) );
  NOR4_X1 U22115 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19067) );
  AOI211_X1 U22116 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_11__SCAN_IN), .B(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19066) );
  NOR4_X1 U22117 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19065) );
  NOR4_X1 U22118 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19064) );
  NAND4_X1 U22119 ( .A1(n19067), .A2(n19066), .A3(n19065), .A4(n19064), .ZN(
        n19068) );
  NOR2_X1 U22120 ( .A1(n19069), .A2(n19068), .ZN(n19080) );
  INV_X1 U22121 ( .A(n19080), .ZN(n19078) );
  NOR2_X1 U22122 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19078), .ZN(n19072) );
  INV_X1 U22123 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19070) );
  AOI22_X1 U22124 ( .A1(n19072), .A2(n19073), .B1(n19078), .B2(n19070), .ZN(
        P2_U2820) );
  OR3_X1 U22125 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19077) );
  INV_X1 U22126 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19071) );
  AOI22_X1 U22127 ( .A1(n19072), .A2(n19077), .B1(n19078), .B2(n19071), .ZN(
        P2_U2821) );
  INV_X1 U22128 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20001) );
  NAND2_X1 U22129 ( .A1(n19072), .A2(n20001), .ZN(n19076) );
  OAI21_X1 U22130 ( .B1(n19951), .B2(n19073), .A(n19080), .ZN(n19074) );
  OAI21_X1 U22131 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19080), .A(n19074), 
        .ZN(n19075) );
  OAI221_X1 U22132 ( .B1(n19076), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19076), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19075), .ZN(P2_U2822) );
  INV_X1 U22133 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19079) );
  OAI221_X1 U22134 ( .B1(n19080), .B2(n19079), .C1(n19078), .C2(n19077), .A(
        n19076), .ZN(P2_U2823) );
  NOR2_X1 U22135 ( .A1(n19242), .A2(n19081), .ZN(n19082) );
  XOR2_X1 U22136 ( .A(n19083), .B(n19082), .Z(n19093) );
  INV_X1 U22137 ( .A(n19084), .ZN(n19086) );
  AOI22_X1 U22138 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19279), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n19265), .ZN(n19085) );
  OAI21_X1 U22139 ( .B1(n19086), .B2(n19270), .A(n19085), .ZN(n19087) );
  AOI211_X1 U22140 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19264), .A(n19399), .B(
        n19087), .ZN(n19092) );
  INV_X1 U22141 ( .A(n19088), .ZN(n19090) );
  AOI22_X1 U22142 ( .A1(n19090), .A2(n19273), .B1(n19089), .B2(n19266), .ZN(
        n19091) );
  OAI211_X1 U22143 ( .C1(n19928), .C2(n19093), .A(n19092), .B(n19091), .ZN(
        P2_U2836) );
  NAND2_X1 U22144 ( .A1(n19226), .A2(n19094), .ZN(n19095) );
  XOR2_X1 U22145 ( .A(n19096), .B(n19095), .Z(n19106) );
  AOI22_X1 U22146 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19279), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19265), .ZN(n19097) );
  OAI21_X1 U22147 ( .B1(n19098), .B2(n19270), .A(n19097), .ZN(n19099) );
  AOI211_X1 U22148 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n19264), .A(n19399), .B(
        n19099), .ZN(n19105) );
  INV_X1 U22149 ( .A(n19100), .ZN(n19101) );
  OAI22_X1 U22150 ( .A1(n19102), .A2(n19230), .B1(n19258), .B2(n19101), .ZN(
        n19103) );
  INV_X1 U22151 ( .A(n19103), .ZN(n19104) );
  OAI211_X1 U22152 ( .C1(n19928), .C2(n19106), .A(n19105), .B(n19104), .ZN(
        P2_U2837) );
  NOR2_X1 U22153 ( .A1(n19242), .A2(n19107), .ZN(n19108) );
  XOR2_X1 U22154 ( .A(n19109), .B(n19108), .Z(n19117) );
  AOI22_X1 U22155 ( .A1(n19110), .A2(n19255), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19279), .ZN(n19111) );
  OAI21_X1 U22156 ( .B1(n15436), .B2(n19222), .A(n19111), .ZN(n19112) );
  AOI211_X1 U22157 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19264), .A(n19399), .B(
        n19112), .ZN(n19116) );
  AOI22_X1 U22158 ( .A1(n19114), .A2(n19273), .B1(n19266), .B2(n19113), .ZN(
        n19115) );
  OAI211_X1 U22159 ( .C1(n19928), .C2(n19117), .A(n19116), .B(n19115), .ZN(
        P2_U2838) );
  NAND2_X1 U22160 ( .A1(n19226), .A2(n19118), .ZN(n19119) );
  XOR2_X1 U22161 ( .A(n19120), .B(n19119), .Z(n19128) );
  AOI22_X1 U22162 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19279), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19265), .ZN(n19121) );
  OAI21_X1 U22163 ( .B1(n19122), .B2(n19270), .A(n19121), .ZN(n19123) );
  AOI211_X1 U22164 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19264), .A(n19399), .B(
        n19123), .ZN(n19127) );
  INV_X1 U22165 ( .A(n19124), .ZN(n19292) );
  AOI22_X1 U22166 ( .A1(n19125), .A2(n19273), .B1(n19266), .B2(n19292), .ZN(
        n19126) );
  OAI211_X1 U22167 ( .C1(n19928), .C2(n19128), .A(n19127), .B(n19126), .ZN(
        P2_U2839) );
  NOR2_X1 U22168 ( .A1(n19242), .A2(n19129), .ZN(n19130) );
  XOR2_X1 U22169 ( .A(n19131), .B(n19130), .Z(n19139) );
  OAI21_X1 U22170 ( .B1(n10707), .B2(n19252), .A(n19214), .ZN(n19134) );
  OAI22_X1 U22171 ( .A1(n19132), .A2(n19270), .B1(n19250), .B2(n21179), .ZN(
        n19133) );
  AOI211_X1 U22172 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19265), .A(n19134), 
        .B(n19133), .ZN(n19138) );
  INV_X1 U22173 ( .A(n19299), .ZN(n19135) );
  AOI22_X1 U22174 ( .A1(n19136), .A2(n19273), .B1(n19266), .B2(n19135), .ZN(
        n19137) );
  OAI211_X1 U22175 ( .C1(n19928), .C2(n19139), .A(n19138), .B(n19137), .ZN(
        P2_U2840) );
  NAND2_X1 U22176 ( .A1(n19226), .A2(n19140), .ZN(n19141) );
  XOR2_X1 U22177 ( .A(n19142), .B(n19141), .Z(n19150) );
  INV_X1 U22178 ( .A(n19143), .ZN(n19145) );
  AOI22_X1 U22179 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19279), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19265), .ZN(n19144) );
  OAI21_X1 U22180 ( .B1(n19145), .B2(n19270), .A(n19144), .ZN(n19146) );
  AOI211_X1 U22181 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n19264), .A(n19399), .B(
        n19146), .ZN(n19149) );
  AOI22_X1 U22182 ( .A1(n19147), .A2(n19273), .B1(n19266), .B2(n19300), .ZN(
        n19148) );
  OAI211_X1 U22183 ( .C1(n19928), .C2(n19150), .A(n19149), .B(n19148), .ZN(
        P2_U2841) );
  OAI22_X1 U22184 ( .A1(n19151), .A2(n19270), .B1(n21161), .B2(n19222), .ZN(
        n19152) );
  AOI211_X1 U22185 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n19264), .A(n19399), .B(
        n19152), .ZN(n19160) );
  NOR2_X1 U22186 ( .A1(n19242), .A2(n19153), .ZN(n19154) );
  XOR2_X1 U22187 ( .A(n19155), .B(n19154), .Z(n19158) );
  OAI22_X1 U22188 ( .A1(n19156), .A2(n19230), .B1(n19258), .B2(n19303), .ZN(
        n19157) );
  AOI21_X1 U22189 ( .B1(n19158), .B2(n19246), .A(n19157), .ZN(n19159) );
  OAI211_X1 U22190 ( .C1(n19161), .C2(n19250), .A(n19160), .B(n19159), .ZN(
        P2_U2842) );
  NAND2_X1 U22191 ( .A1(n19226), .A2(n19162), .ZN(n19164) );
  XNOR2_X1 U22192 ( .A(n19164), .B(n19163), .ZN(n19173) );
  INV_X1 U22193 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n19168) );
  OAI22_X1 U22194 ( .A1(n19165), .A2(n19270), .B1(n19967), .B2(n19222), .ZN(
        n19166) );
  INV_X1 U22195 ( .A(n19166), .ZN(n19167) );
  OAI211_X1 U22196 ( .C1(n19168), .C2(n19252), .A(n19167), .B(n19214), .ZN(
        n19171) );
  OAI22_X1 U22197 ( .A1(n19169), .A2(n19230), .B1(n19306), .B2(n19258), .ZN(
        n19170) );
  AOI211_X1 U22198 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n19279), .A(
        n19171), .B(n19170), .ZN(n19172) );
  OAI21_X1 U22199 ( .B1(n19173), .B2(n19928), .A(n19172), .ZN(P2_U2843) );
  OAI22_X1 U22200 ( .A1(n19174), .A2(n19270), .B1(n19965), .B2(n19222), .ZN(
        n19175) );
  AOI211_X1 U22201 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n19264), .A(n19399), .B(
        n19175), .ZN(n19183) );
  NOR2_X1 U22202 ( .A1(n19242), .A2(n19176), .ZN(n19177) );
  XOR2_X1 U22203 ( .A(n19178), .B(n19177), .Z(n19181) );
  OAI22_X1 U22204 ( .A1(n19179), .A2(n19230), .B1(n19258), .B2(n19308), .ZN(
        n19180) );
  AOI21_X1 U22205 ( .B1(n19181), .B2(n19246), .A(n19180), .ZN(n19182) );
  OAI211_X1 U22206 ( .C1(n19184), .C2(n19250), .A(n19183), .B(n19182), .ZN(
        P2_U2844) );
  NAND2_X1 U22207 ( .A1(n19226), .A2(n19185), .ZN(n19187) );
  XNOR2_X1 U22208 ( .A(n19187), .B(n19186), .ZN(n19197) );
  OAI22_X1 U22209 ( .A1(n19189), .A2(n19270), .B1(n19188), .B2(n19222), .ZN(
        n19190) );
  INV_X1 U22210 ( .A(n19190), .ZN(n19191) );
  OAI211_X1 U22211 ( .C1(n19192), .C2(n19252), .A(n19191), .B(n19214), .ZN(
        n19195) );
  OAI22_X1 U22212 ( .A1(n19193), .A2(n19230), .B1(n19258), .B2(n19311), .ZN(
        n19194) );
  AOI211_X1 U22213 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19279), .A(
        n19195), .B(n19194), .ZN(n19196) );
  OAI21_X1 U22214 ( .B1(n19197), .B2(n19928), .A(n19196), .ZN(P2_U2845) );
  INV_X1 U22215 ( .A(n19198), .ZN(n19199) );
  OAI22_X1 U22216 ( .A1(n19199), .A2(n19270), .B1(n19962), .B2(n19222), .ZN(
        n19200) );
  AOI211_X1 U22217 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19264), .A(n19399), .B(
        n19200), .ZN(n19208) );
  NOR2_X1 U22218 ( .A1(n19242), .A2(n19201), .ZN(n19202) );
  XOR2_X1 U22219 ( .A(n19203), .B(n19202), .Z(n19206) );
  OAI22_X1 U22220 ( .A1(n19204), .A2(n19230), .B1(n19258), .B2(n19313), .ZN(
        n19205) );
  AOI21_X1 U22221 ( .B1(n19206), .B2(n19246), .A(n19205), .ZN(n19207) );
  OAI211_X1 U22222 ( .C1(n19209), .C2(n19250), .A(n19208), .B(n19207), .ZN(
        P2_U2846) );
  NOR2_X1 U22223 ( .A1(n19242), .A2(n19210), .ZN(n19211) );
  XOR2_X1 U22224 ( .A(n19212), .B(n19211), .Z(n19221) );
  AOI22_X1 U22225 ( .A1(n19213), .A2(n19255), .B1(P2_REIP_REG_7__SCAN_IN), 
        .B2(n19265), .ZN(n19215) );
  OAI211_X1 U22226 ( .C1(n19216), .C2(n19252), .A(n19215), .B(n19214), .ZN(
        n19219) );
  OAI22_X1 U22227 ( .A1(n19319), .A2(n19258), .B1(n19230), .B2(n19217), .ZN(
        n19218) );
  AOI211_X1 U22228 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19279), .A(
        n19219), .B(n19218), .ZN(n19220) );
  OAI21_X1 U22229 ( .B1(n19928), .B2(n19221), .A(n19220), .ZN(P2_U2848) );
  OAI22_X1 U22230 ( .A1(n19223), .A2(n19270), .B1(n19958), .B2(n19222), .ZN(
        n19224) );
  AOI211_X1 U22231 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19264), .A(n19399), .B(
        n19224), .ZN(n19234) );
  NAND2_X1 U22232 ( .A1(n19226), .A2(n19225), .ZN(n19227) );
  XNOR2_X1 U22233 ( .A(n19228), .B(n19227), .ZN(n19232) );
  OAI22_X1 U22234 ( .A1(n19321), .A2(n19258), .B1(n19230), .B2(n19229), .ZN(
        n19231) );
  AOI21_X1 U22235 ( .B1(n19246), .B2(n19232), .A(n19231), .ZN(n19233) );
  OAI211_X1 U22236 ( .C1(n19235), .C2(n19250), .A(n19234), .B(n19233), .ZN(
        P2_U2849) );
  INV_X1 U22237 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19236) );
  OAI21_X1 U22238 ( .B1(n19236), .B2(n19252), .A(n19214), .ZN(n19240) );
  OAI22_X1 U22239 ( .A1(n19238), .A2(n19270), .B1(n19250), .B2(n19237), .ZN(
        n19239) );
  AOI211_X1 U22240 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19265), .A(n19240), .B(
        n19239), .ZN(n19249) );
  NOR2_X1 U22241 ( .A1(n19242), .A2(n19241), .ZN(n19244) );
  XNOR2_X1 U22242 ( .A(n19244), .B(n19243), .ZN(n19247) );
  AOI22_X1 U22243 ( .A1(n19247), .A2(n19246), .B1(n19273), .B2(n19245), .ZN(
        n19248) );
  OAI211_X1 U22244 ( .C1(n19258), .C2(n19329), .A(n19249), .B(n19248), .ZN(
        P2_U2850) );
  INV_X1 U22245 ( .A(n20030), .ZN(n19259) );
  OAI22_X1 U22246 ( .A1(n19252), .A2(n19251), .B1(n19250), .B2(n12933), .ZN(
        n19253) );
  AOI21_X1 U22247 ( .B1(n19255), .B2(n19254), .A(n19253), .ZN(n19257) );
  NAND2_X1 U22248 ( .A1(n19265), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19256) );
  OAI211_X1 U22249 ( .C1(n19259), .C2(n19258), .A(n19257), .B(n19256), .ZN(
        n19260) );
  AOI21_X1 U22250 ( .B1(n11288), .B2(n19273), .A(n19260), .ZN(n19262) );
  AOI22_X1 U22251 ( .A1(n20026), .A2(n19276), .B1(n19278), .B2(n12933), .ZN(
        n19261) );
  OAI211_X1 U22252 ( .C1(n19928), .C2(n19263), .A(n19262), .B(n19261), .ZN(
        P2_U2854) );
  AOI22_X1 U22253 ( .A1(n19265), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19264), 
        .B2(P2_EBX_REG_0__SCAN_IN), .ZN(n19269) );
  NAND2_X1 U22254 ( .A1(n19267), .A2(n19266), .ZN(n19268) );
  OAI211_X1 U22255 ( .C1(n19271), .C2(n19270), .A(n19269), .B(n19268), .ZN(
        n19272) );
  AOI21_X1 U22256 ( .B1(n11289), .B2(n19273), .A(n19272), .ZN(n19282) );
  AOI22_X1 U22257 ( .A1(n19277), .A2(n19276), .B1(n19275), .B2(n19274), .ZN(
        n19281) );
  OAI21_X1 U22258 ( .B1(n19279), .B2(n19278), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19280) );
  NAND3_X1 U22259 ( .A1(n19282), .A2(n19281), .A3(n19280), .ZN(P2_U2855) );
  INV_X1 U22260 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19283) );
  OAI22_X1 U22261 ( .A1(n14528), .A2(n19297), .B1(n19284), .B2(n19283), .ZN(
        n19285) );
  INV_X1 U22262 ( .A(n19285), .ZN(n19287) );
  AOI22_X1 U22263 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19338), .B1(n19291), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19286) );
  NAND2_X1 U22264 ( .A1(n19287), .A2(n19286), .ZN(P2_U2888) );
  AOI22_X1 U22265 ( .A1(n19289), .A2(n19288), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19338), .ZN(n19296) );
  AOI22_X1 U22266 ( .A1(n19291), .A2(BUF1_REG_16__SCAN_IN), .B1(n19290), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19295) );
  AOI22_X1 U22267 ( .A1(n19293), .A2(n19343), .B1(n19339), .B2(n19292), .ZN(
        n19294) );
  NAND3_X1 U22268 ( .A1(n19296), .A2(n19295), .A3(n19294), .ZN(P2_U2903) );
  OAI222_X1 U22269 ( .A1(n19299), .A2(n19330), .B1(n13539), .B2(n19322), .C1(
        n19298), .C2(n19347), .ZN(P2_U2904) );
  INV_X1 U22270 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n21151) );
  INV_X1 U22271 ( .A(n19330), .ZN(n19315) );
  AOI22_X1 U22272 ( .A1(n19300), .A2(n19315), .B1(n19388), .B2(n19314), .ZN(
        n19301) );
  OAI21_X1 U22273 ( .B1(n19322), .B2(n21151), .A(n19301), .ZN(P2_U2905) );
  OAI222_X1 U22274 ( .A1(n19303), .A2(n19330), .B1(n13491), .B2(n19322), .C1(
        n19347), .C2(n19302), .ZN(P2_U2906) );
  AOI22_X1 U22275 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19338), .B1(n19304), 
        .B2(n19314), .ZN(n19305) );
  OAI21_X1 U22276 ( .B1(n19330), .B2(n19306), .A(n19305), .ZN(P2_U2907) );
  OAI222_X1 U22277 ( .A1(n19308), .A2(n19330), .B1(n13496), .B2(n19322), .C1(
        n19347), .C2(n19307), .ZN(P2_U2908) );
  AOI22_X1 U22278 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19338), .B1(n19309), 
        .B2(n19314), .ZN(n19310) );
  OAI21_X1 U22279 ( .B1(n19330), .B2(n19311), .A(n19310), .ZN(P2_U2909) );
  OAI222_X1 U22280 ( .A1(n19313), .A2(n19330), .B1(n13484), .B2(n19322), .C1(
        n19347), .C2(n19312), .ZN(P2_U2910) );
  INV_X1 U22281 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19369) );
  AOI22_X1 U22282 ( .A1(n19316), .A2(n19315), .B1(n19386), .B2(n19314), .ZN(
        n19317) );
  OAI21_X1 U22283 ( .B1(n19322), .B2(n19369), .A(n19317), .ZN(P2_U2911) );
  INV_X1 U22284 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n21250) );
  OAI222_X1 U22285 ( .A1(n19319), .A2(n19330), .B1(n21250), .B2(n19322), .C1(
        n19347), .C2(n19318), .ZN(P2_U2912) );
  INV_X1 U22286 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19372) );
  OAI222_X1 U22287 ( .A1(n19321), .A2(n19330), .B1(n19372), .B2(n19322), .C1(
        n19347), .C2(n19320), .ZN(P2_U2913) );
  INV_X1 U22288 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n21296) );
  OAI22_X1 U22289 ( .A1(n21296), .A2(n19322), .B1(n19436), .B2(n19347), .ZN(
        n19323) );
  INV_X1 U22290 ( .A(n19323), .ZN(n19328) );
  OR3_X1 U22291 ( .A1(n19326), .A2(n19325), .A3(n19324), .ZN(n19327) );
  OAI211_X1 U22292 ( .C1(n19330), .C2(n19329), .A(n19328), .B(n19327), .ZN(
        P2_U2914) );
  INV_X1 U22293 ( .A(n19331), .ZN(n20009) );
  AOI22_X1 U22294 ( .A1(n20009), .A2(n19339), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19338), .ZN(n19337) );
  OAI21_X1 U22295 ( .B1(n19334), .B2(n19333), .A(n19332), .ZN(n19335) );
  NAND2_X1 U22296 ( .A1(n19335), .A2(n19343), .ZN(n19336) );
  OAI211_X1 U22297 ( .C1(n19426), .C2(n19347), .A(n19337), .B(n19336), .ZN(
        P2_U2916) );
  AOI22_X1 U22298 ( .A1(n19339), .A2(n20030), .B1(n19338), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19346) );
  OAI21_X1 U22299 ( .B1(n19342), .B2(n19341), .A(n19340), .ZN(n19344) );
  NAND2_X1 U22300 ( .A1(n19344), .A2(n19343), .ZN(n19345) );
  OAI211_X1 U22301 ( .C1(n19348), .C2(n19347), .A(n19346), .B(n19345), .ZN(
        P2_U2918) );
  NOR2_X1 U22302 ( .A1(n19357), .A2(n19349), .ZN(P2_U2920) );
  INV_X1 U22303 ( .A(n19350), .ZN(n19355) );
  AOI22_X1 U22304 ( .A1(n19355), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19383), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19351) );
  OAI21_X1 U22305 ( .B1(n19357), .B2(n19352), .A(n19351), .ZN(P2_U2921) );
  INV_X1 U22306 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n19354) );
  AOI22_X1 U22307 ( .A1(n19355), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n19383), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n19353) );
  OAI21_X1 U22308 ( .B1(n19354), .B2(n19357), .A(n19353), .ZN(P2_U2927) );
  AOI22_X1 U22309 ( .A1(n19355), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19383), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n19356) );
  OAI21_X1 U22310 ( .B1(n19358), .B2(n19357), .A(n19356), .ZN(P2_U2935) );
  AOI22_X1 U22311 ( .A1(n19383), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19359) );
  OAI21_X1 U22312 ( .B1(n19385), .B2(n13539), .A(n19359), .ZN(P2_U2936) );
  AOI22_X1 U22313 ( .A1(n19383), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19360) );
  OAI21_X1 U22314 ( .B1(n19385), .B2(n21151), .A(n19360), .ZN(P2_U2937) );
  AOI22_X1 U22315 ( .A1(n19383), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19361) );
  OAI21_X1 U22316 ( .B1(n19385), .B2(n13491), .A(n19361), .ZN(P2_U2938) );
  AOI22_X1 U22317 ( .A1(n19383), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19362) );
  OAI21_X1 U22318 ( .B1(n19385), .B2(n19363), .A(n19362), .ZN(P2_U2939) );
  AOI22_X1 U22319 ( .A1(n19383), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19364) );
  OAI21_X1 U22320 ( .B1(n19385), .B2(n13496), .A(n19364), .ZN(P2_U2940) );
  AOI22_X1 U22321 ( .A1(n19383), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19365) );
  OAI21_X1 U22322 ( .B1(n19385), .B2(n19366), .A(n19365), .ZN(P2_U2941) );
  AOI22_X1 U22323 ( .A1(n19383), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19367) );
  OAI21_X1 U22324 ( .B1(n19385), .B2(n13484), .A(n19367), .ZN(P2_U2942) );
  AOI22_X1 U22325 ( .A1(n19383), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19368) );
  OAI21_X1 U22326 ( .B1(n19385), .B2(n19369), .A(n19368), .ZN(P2_U2943) );
  AOI22_X1 U22327 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n19382), .B1(n19383), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n19370) );
  OAI21_X1 U22328 ( .B1(n19385), .B2(n21250), .A(n19370), .ZN(P2_U2944) );
  AOI22_X1 U22329 ( .A1(n19383), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19371) );
  OAI21_X1 U22330 ( .B1(n19385), .B2(n19372), .A(n19371), .ZN(P2_U2945) );
  AOI22_X1 U22331 ( .A1(n19383), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19373) );
  OAI21_X1 U22332 ( .B1(n19385), .B2(n21296), .A(n19373), .ZN(P2_U2946) );
  INV_X1 U22333 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19375) );
  AOI22_X1 U22334 ( .A1(n19383), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19374) );
  OAI21_X1 U22335 ( .B1(n19385), .B2(n19375), .A(n19374), .ZN(P2_U2947) );
  INV_X1 U22336 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19377) );
  AOI22_X1 U22337 ( .A1(n19383), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19376) );
  OAI21_X1 U22338 ( .B1(n19385), .B2(n19377), .A(n19376), .ZN(P2_U2948) );
  INV_X1 U22339 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19379) );
  AOI22_X1 U22340 ( .A1(n19383), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19378) );
  OAI21_X1 U22341 ( .B1(n19385), .B2(n19379), .A(n19378), .ZN(P2_U2949) );
  INV_X1 U22342 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19381) );
  AOI22_X1 U22343 ( .A1(n19383), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19380) );
  OAI21_X1 U22344 ( .B1(n19385), .B2(n19381), .A(n19380), .ZN(P2_U2950) );
  AOI22_X1 U22345 ( .A1(n19383), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19382), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19384) );
  OAI21_X1 U22346 ( .B1(n19385), .B2(n13499), .A(n19384), .ZN(P2_U2951) );
  AOI22_X1 U22347 ( .A1(n19394), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19393), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n19387) );
  NAND2_X1 U22348 ( .A1(n19389), .A2(n19386), .ZN(n19391) );
  NAND2_X1 U22349 ( .A1(n19387), .A2(n19391), .ZN(P2_U2960) );
  AOI22_X1 U22350 ( .A1(n19394), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19393), 
        .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n19390) );
  NAND2_X1 U22351 ( .A1(n19389), .A2(n19388), .ZN(n19395) );
  NAND2_X1 U22352 ( .A1(n19390), .A2(n19395), .ZN(P2_U2966) );
  AOI22_X1 U22353 ( .A1(n19394), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19393), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n19392) );
  NAND2_X1 U22354 ( .A1(n19392), .A2(n19391), .ZN(P2_U2975) );
  AOI22_X1 U22355 ( .A1(n19394), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19393), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n19396) );
  NAND2_X1 U22356 ( .A1(n19396), .A2(n19395), .ZN(P2_U2981) );
  AOI22_X1 U22357 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19399), .B1(n19398), 
        .B2(n19397), .ZN(n19407) );
  AOI222_X1 U22358 ( .A1(n19405), .A2(n19404), .B1(n19403), .B2(n19402), .C1(
        n19401), .C2(n19400), .ZN(n19406) );
  OAI211_X1 U22359 ( .C1(n19409), .C2(n19408), .A(n19407), .B(n19406), .ZN(
        P2_U3010) );
  NOR2_X1 U22360 ( .A1(n19410), .A2(n19504), .ZN(n19441) );
  AOI22_X1 U22361 ( .A1(n19854), .A2(n19442), .B1(n19842), .B2(n19441), .ZN(
        n19419) );
  AOI21_X1 U22362 ( .B1(n19919), .B2(n19475), .A(n19691), .ZN(n19411) );
  NOR2_X1 U22363 ( .A1(n19411), .A2(n20013), .ZN(n19414) );
  INV_X1 U22364 ( .A(n19853), .ZN(n19910) );
  AOI21_X1 U22365 ( .B1(n19415), .B2(n20033), .A(n20004), .ZN(n19412) );
  AOI21_X1 U22366 ( .B1(n19414), .B2(n19910), .A(n19412), .ZN(n19413) );
  OAI21_X1 U22367 ( .B1(n19413), .B2(n19441), .A(n19851), .ZN(n19444) );
  OAI21_X1 U22368 ( .B1(n19853), .B2(n19441), .A(n19414), .ZN(n19417) );
  OAI21_X1 U22369 ( .B1(n19415), .B2(n19441), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19416) );
  NAND2_X1 U22370 ( .A1(n19417), .A2(n19416), .ZN(n19443) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19444), .B1(
        n19791), .B2(n19443), .ZN(n19418) );
  OAI211_X1 U22372 ( .C1(n19857), .C2(n19475), .A(n19419), .B(n19418), .ZN(
        P2_U3048) );
  AOI22_X1 U22373 ( .A1(n19863), .A2(n19442), .B1(n19859), .B2(n19441), .ZN(
        n19421) );
  AOI22_X1 U22374 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19444), .B1(
        n19858), .B2(n19443), .ZN(n19420) );
  OAI211_X1 U22375 ( .C1(n19866), .C2(n19475), .A(n19421), .B(n19420), .ZN(
        P2_U3049) );
  AOI22_X1 U22376 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19433), .ZN(n21353) );
  AOI22_X1 U22377 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19433), .ZN(n19739) );
  AND2_X1 U22378 ( .A1(n10240), .A2(n19434), .ZN(n21344) );
  AOI22_X1 U22379 ( .A1(n21346), .A2(n19442), .B1(n21344), .B2(n19441), .ZN(
        n19424) );
  NOR2_X2 U22380 ( .A1(n19422), .A2(n19765), .ZN(n21348) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19444), .B1(
        n21348), .B2(n19443), .ZN(n19423) );
  OAI211_X1 U22382 ( .C1(n21353), .C2(n19475), .A(n19424), .B(n19423), .ZN(
        P2_U3050) );
  AOI22_X1 U22383 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19433), .ZN(n19880) );
  AOI22_X1 U22384 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19433), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19432), .ZN(n19802) );
  AND2_X1 U22385 ( .A1(n19425), .A2(n19434), .ZN(n19873) );
  AOI22_X1 U22386 ( .A1(n19877), .A2(n19442), .B1(n19873), .B2(n19441), .ZN(
        n19428) );
  NOR2_X2 U22387 ( .A1(n19426), .A2(n19765), .ZN(n19872) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19444), .B1(
        n19872), .B2(n19443), .ZN(n19427) );
  OAI211_X1 U22389 ( .C1(n19880), .C2(n19475), .A(n19428), .B(n19427), .ZN(
        P2_U3051) );
  AOI22_X1 U22390 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19433), .ZN(n19889) );
  AOI22_X1 U22391 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19433), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19432), .ZN(n19744) );
  AOI22_X1 U22392 ( .A1(n19886), .A2(n19442), .B1(n19882), .B2(n19441), .ZN(
        n19431) );
  NOR2_X2 U22393 ( .A1(n19429), .A2(n19765), .ZN(n19881) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19444), .B1(
        n19881), .B2(n19443), .ZN(n19430) );
  OAI211_X1 U22395 ( .C1(n19889), .C2(n19475), .A(n19431), .B(n19430), .ZN(
        P2_U3052) );
  AOI22_X1 U22396 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19432), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19433), .ZN(n19898) );
  AOI22_X1 U22397 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19433), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19432), .ZN(n19747) );
  AOI22_X1 U22398 ( .A1(n19895), .A2(n19442), .B1(n19891), .B2(n19441), .ZN(
        n19438) );
  NOR2_X2 U22399 ( .A1(n19436), .A2(n19765), .ZN(n19890) );
  AOI22_X1 U22400 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19444), .B1(
        n19890), .B2(n19443), .ZN(n19437) );
  OAI211_X1 U22401 ( .C1(n19898), .C2(n19475), .A(n19438), .B(n19437), .ZN(
        P2_U3053) );
  AOI22_X1 U22402 ( .A1(n19903), .A2(n19442), .B1(n9707), .B2(n19441), .ZN(
        n19440) );
  AOI22_X1 U22403 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19444), .B1(
        n19782), .B2(n19443), .ZN(n19439) );
  OAI211_X1 U22404 ( .C1(n19906), .C2(n19475), .A(n19440), .B(n19439), .ZN(
        P2_U3054) );
  AOI22_X1 U22405 ( .A1(n19914), .A2(n19442), .B1(n19908), .B2(n19441), .ZN(
        n19446) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19444), .B1(
        n19907), .B2(n19443), .ZN(n19445) );
  OAI211_X1 U22407 ( .C1(n19920), .C2(n19475), .A(n19446), .B(n19445), .ZN(
        P2_U3055) );
  NOR2_X1 U22408 ( .A1(n19504), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19453) );
  INV_X1 U22409 ( .A(n19453), .ZN(n19448) );
  NOR3_X2 U22410 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20040), .A3(
        n19504), .ZN(n19470) );
  OAI21_X1 U22411 ( .B1(n10485), .B2(n19470), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19447) );
  OAI21_X1 U22412 ( .B1(n19448), .B2(n20013), .A(n19447), .ZN(n19471) );
  AOI22_X1 U22413 ( .A1(n19471), .A2(n19791), .B1(n19842), .B2(n19470), .ZN(
        n19457) );
  NOR2_X1 U22414 ( .A1(n20011), .A2(n19449), .ZN(n19454) );
  INV_X1 U22415 ( .A(n19470), .ZN(n19450) );
  OAI211_X1 U22416 ( .C1(n19451), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19450), 
        .B(n20013), .ZN(n19452) );
  OAI211_X1 U22417 ( .C1(n19454), .C2(n19453), .A(n19851), .B(n19452), .ZN(
        n19472) );
  NOR2_X2 U22418 ( .A1(n19455), .A2(n19609), .ZN(n19499) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19472), .B1(
        n19499), .B2(n19792), .ZN(n19456) );
  OAI211_X1 U22420 ( .C1(n19733), .C2(n19475), .A(n19457), .B(n19456), .ZN(
        P2_U3056) );
  AOI22_X1 U22421 ( .A1(n19471), .A2(n19858), .B1(n19859), .B2(n19470), .ZN(
        n19459) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19472), .B1(
        n19499), .B2(n19811), .ZN(n19458) );
  OAI211_X1 U22423 ( .C1(n19736), .C2(n19475), .A(n19459), .B(n19458), .ZN(
        P2_U3057) );
  AOI22_X1 U22424 ( .A1(n19471), .A2(n21348), .B1(n21344), .B2(n19470), .ZN(
        n19461) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19472), .B1(
        n19499), .B2(n19815), .ZN(n19460) );
  OAI211_X1 U22426 ( .C1(n19739), .C2(n19475), .A(n19461), .B(n19460), .ZN(
        P2_U3058) );
  AOI22_X1 U22427 ( .A1(n19471), .A2(n19872), .B1(n19873), .B2(n19470), .ZN(
        n19463) );
  INV_X1 U22428 ( .A(n19880), .ZN(n19819) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19472), .B1(
        n19499), .B2(n19819), .ZN(n19462) );
  OAI211_X1 U22430 ( .C1(n19802), .C2(n19475), .A(n19463), .B(n19462), .ZN(
        P2_U3059) );
  AOI22_X1 U22431 ( .A1(n19471), .A2(n19881), .B1(n19882), .B2(n19470), .ZN(
        n19465) );
  INV_X1 U22432 ( .A(n19889), .ZN(n19822) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19472), .B1(
        n19499), .B2(n19822), .ZN(n19464) );
  OAI211_X1 U22434 ( .C1(n19744), .C2(n19475), .A(n19465), .B(n19464), .ZN(
        P2_U3060) );
  AOI22_X1 U22435 ( .A1(n19471), .A2(n19890), .B1(n19891), .B2(n19470), .ZN(
        n19467) );
  INV_X1 U22436 ( .A(n19898), .ZN(n19826) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19472), .B1(
        n19499), .B2(n19826), .ZN(n19466) );
  OAI211_X1 U22438 ( .C1(n19747), .C2(n19475), .A(n19467), .B(n19466), .ZN(
        P2_U3061) );
  AOI22_X1 U22439 ( .A1(n19471), .A2(n19782), .B1(n9707), .B2(n19470), .ZN(
        n19469) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19472), .B1(
        n19499), .B2(n19748), .ZN(n19468) );
  OAI211_X1 U22441 ( .C1(n19751), .C2(n19475), .A(n19469), .B(n19468), .ZN(
        P2_U3062) );
  AOI22_X1 U22442 ( .A1(n19471), .A2(n19907), .B1(n19908), .B2(n19470), .ZN(
        n19474) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19472), .B1(
        n19499), .B2(n19831), .ZN(n19473) );
  OAI211_X1 U22444 ( .C1(n19758), .C2(n19475), .A(n19474), .B(n19473), .ZN(
        P2_U3063) );
  INV_X1 U22445 ( .A(n19504), .ZN(n19476) );
  NAND2_X1 U22446 ( .A1(n19694), .A2(n19476), .ZN(n19480) );
  NOR3_X2 U22447 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20032), .A3(
        n19504), .ZN(n19497) );
  OAI21_X1 U22448 ( .B1(n10475), .B2(n19497), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19477) );
  OAI21_X1 U22449 ( .B1(n19480), .B2(n20013), .A(n19477), .ZN(n19498) );
  AOI22_X1 U22450 ( .A1(n19498), .A2(n19791), .B1(n19842), .B2(n19497), .ZN(
        n19484) );
  AOI21_X1 U22451 ( .B1(n19478), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19482) );
  OAI21_X1 U22452 ( .B1(n19499), .B2(n19524), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19479) );
  NAND2_X1 U22453 ( .A1(n19480), .A2(n19479), .ZN(n19481) );
  OAI211_X1 U22454 ( .C1(n19497), .C2(n19482), .A(n19481), .B(n19851), .ZN(
        n19500) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19854), .ZN(n19483) );
  OAI211_X1 U22456 ( .C1(n19857), .C2(n19533), .A(n19484), .B(n19483), .ZN(
        P2_U3064) );
  AOI22_X1 U22457 ( .A1(n19498), .A2(n19858), .B1(n19859), .B2(n19497), .ZN(
        n19486) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19863), .ZN(n19485) );
  OAI211_X1 U22459 ( .C1(n19866), .C2(n19533), .A(n19486), .B(n19485), .ZN(
        P2_U3065) );
  AOI22_X1 U22460 ( .A1(n19498), .A2(n21348), .B1(n21344), .B2(n19497), .ZN(
        n19488) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n21346), .ZN(n19487) );
  OAI211_X1 U22462 ( .C1(n21353), .C2(n19533), .A(n19488), .B(n19487), .ZN(
        P2_U3066) );
  AOI22_X1 U22463 ( .A1(n19498), .A2(n19872), .B1(n19873), .B2(n19497), .ZN(
        n19490) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19877), .ZN(n19489) );
  OAI211_X1 U22465 ( .C1(n19880), .C2(n19533), .A(n19490), .B(n19489), .ZN(
        P2_U3067) );
  AOI22_X1 U22466 ( .A1(n19498), .A2(n19881), .B1(n19882), .B2(n19497), .ZN(
        n19492) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19886), .ZN(n19491) );
  OAI211_X1 U22468 ( .C1(n19889), .C2(n19533), .A(n19492), .B(n19491), .ZN(
        P2_U3068) );
  AOI22_X1 U22469 ( .A1(n19498), .A2(n19890), .B1(n19891), .B2(n19497), .ZN(
        n19494) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19895), .ZN(n19493) );
  OAI211_X1 U22471 ( .C1(n19898), .C2(n19533), .A(n19494), .B(n19493), .ZN(
        P2_U3069) );
  AOI22_X1 U22472 ( .A1(n19498), .A2(n19782), .B1(n9707), .B2(n19497), .ZN(
        n19496) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19903), .ZN(n19495) );
  OAI211_X1 U22474 ( .C1(n19906), .C2(n19533), .A(n19496), .B(n19495), .ZN(
        P2_U3070) );
  AOI22_X1 U22475 ( .A1(n19498), .A2(n19907), .B1(n19908), .B2(n19497), .ZN(
        n19502) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19914), .ZN(n19501) );
  OAI211_X1 U22477 ( .C1(n19920), .C2(n19533), .A(n19502), .B(n19501), .ZN(
        P2_U3071) );
  NOR2_X1 U22478 ( .A1(n19611), .A2(n19504), .ZN(n19528) );
  AOI22_X1 U22479 ( .A1(n19854), .A2(n19524), .B1(n19842), .B2(n19528), .ZN(
        n19513) );
  NAND2_X1 U22480 ( .A1(n19503), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19614) );
  OAI21_X1 U22481 ( .B1(n19614), .B2(n20003), .A(n20004), .ZN(n19511) );
  NOR2_X1 U22482 ( .A1(n20032), .A2(n19504), .ZN(n19508) );
  OAI21_X1 U22483 ( .B1(n10515), .B2(n19763), .A(n20033), .ZN(n19506) );
  INV_X1 U22484 ( .A(n19528), .ZN(n19505) );
  AOI21_X1 U22485 ( .B1(n19506), .B2(n19505), .A(n19765), .ZN(n19507) );
  OAI21_X1 U22486 ( .B1(n19511), .B2(n19508), .A(n19507), .ZN(n19530) );
  INV_X1 U22487 ( .A(n19508), .ZN(n19510) );
  OAI21_X1 U22488 ( .B1(n10515), .B2(n19528), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19509) );
  OAI21_X1 U22489 ( .B1(n19511), .B2(n19510), .A(n19509), .ZN(n19529) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19530), .B1(
        n19791), .B2(n19529), .ZN(n19512) );
  OAI211_X1 U22491 ( .C1(n19857), .C2(n19527), .A(n19513), .B(n19512), .ZN(
        P2_U3072) );
  AOI22_X1 U22492 ( .A1(n19863), .A2(n19524), .B1(n19859), .B2(n19528), .ZN(
        n19515) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19530), .B1(
        n19858), .B2(n19529), .ZN(n19514) );
  OAI211_X1 U22494 ( .C1(n19866), .C2(n19527), .A(n19515), .B(n19514), .ZN(
        P2_U3073) );
  AOI22_X1 U22495 ( .A1(n19815), .A2(n19545), .B1(n19528), .B2(n21344), .ZN(
        n19517) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19530), .B1(
        n21348), .B2(n19529), .ZN(n19516) );
  OAI211_X1 U22497 ( .C1(n19739), .C2(n19533), .A(n19517), .B(n19516), .ZN(
        P2_U3074) );
  AOI22_X1 U22498 ( .A1(n19877), .A2(n19524), .B1(n19528), .B2(n19873), .ZN(
        n19519) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19530), .B1(
        n19872), .B2(n19529), .ZN(n19518) );
  OAI211_X1 U22500 ( .C1(n19880), .C2(n19527), .A(n19519), .B(n19518), .ZN(
        P2_U3075) );
  AOI22_X1 U22501 ( .A1(n19886), .A2(n19524), .B1(n19528), .B2(n19882), .ZN(
        n19521) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19530), .B1(
        n19881), .B2(n19529), .ZN(n19520) );
  OAI211_X1 U22503 ( .C1(n19889), .C2(n19527), .A(n19521), .B(n19520), .ZN(
        P2_U3076) );
  AOI22_X1 U22504 ( .A1(n19826), .A2(n19545), .B1(n19528), .B2(n19891), .ZN(
        n19523) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19530), .B1(
        n19890), .B2(n19529), .ZN(n19522) );
  OAI211_X1 U22506 ( .C1(n19747), .C2(n19533), .A(n19523), .B(n19522), .ZN(
        P2_U3077) );
  AOI22_X1 U22507 ( .A1(n19903), .A2(n19524), .B1(n9707), .B2(n19528), .ZN(
        n19526) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19530), .B1(
        n19782), .B2(n19529), .ZN(n19525) );
  OAI211_X1 U22509 ( .C1(n19906), .C2(n19527), .A(n19526), .B(n19525), .ZN(
        P2_U3078) );
  AOI22_X1 U22510 ( .A1(n19831), .A2(n19545), .B1(n19908), .B2(n19528), .ZN(
        n19532) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19530), .B1(
        n19907), .B2(n19529), .ZN(n19531) );
  OAI211_X1 U22512 ( .C1(n19758), .C2(n19533), .A(n19532), .B(n19531), .ZN(
        P2_U3079) );
  INV_X1 U22513 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19536) );
  AOI22_X1 U22514 ( .A1(n19815), .A2(n21345), .B1(n19544), .B2(n21344), .ZN(
        n19535) );
  AOI22_X1 U22515 ( .A1(n21348), .A2(n19546), .B1(n19545), .B2(n21346), .ZN(
        n19534) );
  OAI211_X1 U22516 ( .C1(n19549), .C2(n19536), .A(n19535), .B(n19534), .ZN(
        P2_U3082) );
  AOI22_X1 U22517 ( .A1(n19819), .A2(n21345), .B1(n19544), .B2(n19873), .ZN(
        n19538) );
  AOI22_X1 U22518 ( .A1(n19872), .A2(n19546), .B1(n19545), .B2(n19877), .ZN(
        n19537) );
  OAI211_X1 U22519 ( .C1(n19549), .C2(n10415), .A(n19538), .B(n19537), .ZN(
        P2_U3083) );
  INV_X1 U22520 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n19541) );
  AOI22_X1 U22521 ( .A1(n19822), .A2(n21345), .B1(n19544), .B2(n19882), .ZN(
        n19540) );
  AOI22_X1 U22522 ( .A1(n19881), .A2(n19546), .B1(n19545), .B2(n19886), .ZN(
        n19539) );
  OAI211_X1 U22523 ( .C1(n19549), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P2_U3084) );
  AOI22_X1 U22524 ( .A1(n19895), .A2(n19545), .B1(n19544), .B2(n19891), .ZN(
        n19543) );
  AOI22_X1 U22525 ( .A1(n19890), .A2(n19546), .B1(n21345), .B2(n19826), .ZN(
        n19542) );
  OAI211_X1 U22526 ( .C1(n19549), .C2(n10490), .A(n19543), .B(n19542), .ZN(
        P2_U3085) );
  AOI22_X1 U22527 ( .A1(n19748), .A2(n21345), .B1(n9707), .B2(n19544), .ZN(
        n19548) );
  AOI22_X1 U22528 ( .A1(n19782), .A2(n19546), .B1(n19545), .B2(n19903), .ZN(
        n19547) );
  OAI211_X1 U22529 ( .C1(n19549), .C2(n10523), .A(n19548), .B(n19547), .ZN(
        P2_U3086) );
  NOR2_X1 U22530 ( .A1(n19610), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19554) );
  INV_X1 U22531 ( .A(n19554), .ZN(n19557) );
  NOR2_X1 U22532 ( .A1(n20040), .A2(n19557), .ZN(n21343) );
  AOI22_X1 U22533 ( .A1(n19792), .A2(n19599), .B1(n19842), .B2(n21343), .ZN(
        n19560) );
  OAI21_X1 U22534 ( .B1(n19614), .B2(n19550), .A(n20004), .ZN(n19558) );
  OAI21_X1 U22535 ( .B1(n19555), .B2(n19763), .A(n20033), .ZN(n19552) );
  INV_X1 U22536 ( .A(n21343), .ZN(n19551) );
  AOI21_X1 U22537 ( .B1(n19552), .B2(n19551), .A(n19765), .ZN(n19553) );
  OAI21_X1 U22538 ( .B1(n19558), .B2(n19554), .A(n19553), .ZN(n21349) );
  OAI21_X1 U22539 ( .B1(n19555), .B2(n21343), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19556) );
  OAI21_X1 U22540 ( .B1(n19558), .B2(n19557), .A(n19556), .ZN(n21347) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21349), .B1(
        n19791), .B2(n21347), .ZN(n19559) );
  OAI211_X1 U22542 ( .C1(n19733), .C2(n19563), .A(n19560), .B(n19559), .ZN(
        P2_U3088) );
  AOI22_X1 U22543 ( .A1(n19811), .A2(n19599), .B1(n19859), .B2(n21343), .ZN(
        n19562) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21349), .B1(
        n19858), .B2(n21347), .ZN(n19561) );
  OAI211_X1 U22545 ( .C1(n19736), .C2(n19563), .A(n19562), .B(n19561), .ZN(
        P2_U3089) );
  AOI22_X1 U22546 ( .A1(n19877), .A2(n21345), .B1(n19873), .B2(n21343), .ZN(
        n19565) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21349), .B1(
        n19872), .B2(n21347), .ZN(n19564) );
  OAI211_X1 U22548 ( .C1(n19880), .C2(n21352), .A(n19565), .B(n19564), .ZN(
        P2_U3091) );
  AOI22_X1 U22549 ( .A1(n19886), .A2(n21345), .B1(n19882), .B2(n21343), .ZN(
        n19567) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21349), .B1(
        n19881), .B2(n21347), .ZN(n19566) );
  OAI211_X1 U22551 ( .C1(n19889), .C2(n21352), .A(n19567), .B(n19566), .ZN(
        P2_U3092) );
  AOI22_X1 U22552 ( .A1(n19895), .A2(n21345), .B1(n19891), .B2(n21343), .ZN(
        n19569) );
  AOI22_X1 U22553 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21349), .B1(
        n19890), .B2(n21347), .ZN(n19568) );
  OAI211_X1 U22554 ( .C1(n19898), .C2(n21352), .A(n19569), .B(n19568), .ZN(
        P2_U3093) );
  AOI22_X1 U22555 ( .A1(n19903), .A2(n21345), .B1(n9707), .B2(n21343), .ZN(
        n19571) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21349), .B1(
        n19782), .B2(n21347), .ZN(n19570) );
  OAI211_X1 U22557 ( .C1(n19906), .C2(n21352), .A(n19571), .B(n19570), .ZN(
        P2_U3094) );
  AOI22_X1 U22558 ( .A1(n19914), .A2(n21345), .B1(n19908), .B2(n21343), .ZN(
        n19573) );
  AOI22_X1 U22559 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21349), .B1(
        n19907), .B2(n21347), .ZN(n19572) );
  OAI211_X1 U22560 ( .C1(n19920), .C2(n21352), .A(n19573), .B(n19572), .ZN(
        P2_U3095) );
  OAI21_X1 U22561 ( .B1(n19599), .B2(n19631), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19577) );
  INV_X1 U22562 ( .A(n19610), .ZN(n19575) );
  NAND2_X1 U22563 ( .A1(n19694), .A2(n19575), .ZN(n19576) );
  NAND2_X1 U22564 ( .A1(n19577), .A2(n19576), .ZN(n19583) );
  NAND2_X1 U22565 ( .A1(n19584), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19578) );
  NAND2_X1 U22566 ( .A1(n19578), .A2(n20033), .ZN(n19581) );
  NAND2_X1 U22567 ( .A1(n19579), .A2(n20017), .ZN(n19615) );
  NOR2_X1 U22568 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19615), .ZN(
        n19604) );
  INV_X1 U22569 ( .A(n19604), .ZN(n19580) );
  AOI21_X1 U22570 ( .B1(n19581), .B2(n19580), .A(n19765), .ZN(n19582) );
  INV_X1 U22571 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n21277) );
  INV_X1 U22572 ( .A(n19584), .ZN(n19585) );
  OAI21_X1 U22573 ( .B1(n19585), .B2(n19604), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19586) );
  OAI21_X1 U22574 ( .B1(n19610), .B2(n19587), .A(n19586), .ZN(n19605) );
  AOI22_X1 U22575 ( .A1(n19605), .A2(n19791), .B1(n19842), .B2(n19604), .ZN(
        n19589) );
  AOI22_X1 U22576 ( .A1(n19599), .A2(n19854), .B1(n19631), .B2(n19792), .ZN(
        n19588) );
  OAI211_X1 U22577 ( .C1(n19592), .C2(n21277), .A(n19589), .B(n19588), .ZN(
        P2_U3096) );
  AOI22_X1 U22578 ( .A1(n19605), .A2(n19858), .B1(n19859), .B2(n19604), .ZN(
        n19591) );
  AOI22_X1 U22579 ( .A1(n19599), .A2(n19863), .B1(n19631), .B2(n19811), .ZN(
        n19590) );
  OAI211_X1 U22580 ( .C1(n19592), .C2(n11082), .A(n19591), .B(n19590), .ZN(
        P2_U3097) );
  AOI22_X1 U22581 ( .A1(n19605), .A2(n21348), .B1(n21344), .B2(n19604), .ZN(
        n19594) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19606), .B1(
        n19631), .B2(n19815), .ZN(n19593) );
  OAI211_X1 U22583 ( .C1(n19739), .C2(n21352), .A(n19594), .B(n19593), .ZN(
        P2_U3098) );
  AOI22_X1 U22584 ( .A1(n19605), .A2(n19872), .B1(n19873), .B2(n19604), .ZN(
        n19596) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19606), .B1(
        n19599), .B2(n19877), .ZN(n19595) );
  OAI211_X1 U22586 ( .C1(n19880), .C2(n19638), .A(n19596), .B(n19595), .ZN(
        P2_U3099) );
  AOI22_X1 U22587 ( .A1(n19605), .A2(n19881), .B1(n19882), .B2(n19604), .ZN(
        n19598) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19606), .B1(
        n19599), .B2(n19886), .ZN(n19597) );
  OAI211_X1 U22589 ( .C1(n19889), .C2(n19638), .A(n19598), .B(n19597), .ZN(
        P2_U3100) );
  AOI22_X1 U22590 ( .A1(n19605), .A2(n19890), .B1(n19891), .B2(n19604), .ZN(
        n19601) );
  AOI22_X1 U22591 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19606), .B1(
        n19599), .B2(n19895), .ZN(n19600) );
  OAI211_X1 U22592 ( .C1(n19898), .C2(n19638), .A(n19601), .B(n19600), .ZN(
        P2_U3101) );
  AOI22_X1 U22593 ( .A1(n19605), .A2(n19782), .B1(n9707), .B2(n19604), .ZN(
        n19603) );
  AOI22_X1 U22594 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19606), .B1(
        n19631), .B2(n19748), .ZN(n19602) );
  OAI211_X1 U22595 ( .C1(n19751), .C2(n21352), .A(n19603), .B(n19602), .ZN(
        P2_U3102) );
  AOI22_X1 U22596 ( .A1(n19605), .A2(n19907), .B1(n19908), .B2(n19604), .ZN(
        n19608) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19606), .B1(
        n19631), .B2(n19831), .ZN(n19607) );
  OAI211_X1 U22598 ( .C1(n19758), .C2(n21352), .A(n19608), .B(n19607), .ZN(
        P2_U3103) );
  NOR2_X1 U22599 ( .A1(n19611), .A2(n19610), .ZN(n19646) );
  OAI21_X1 U22600 ( .B1(n19612), .B2(n19646), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19613) );
  OAI21_X1 U22601 ( .B1(n19615), .B2(n20013), .A(n19613), .ZN(n19634) );
  AOI22_X1 U22602 ( .A1(n19634), .A2(n19791), .B1(n19842), .B2(n19646), .ZN(
        n19620) );
  OR2_X1 U22603 ( .A1(n19614), .A2(n19846), .ZN(n20014) );
  INV_X1 U22604 ( .A(n20014), .ZN(n19618) );
  INV_X1 U22605 ( .A(n19615), .ZN(n19617) );
  INV_X1 U22606 ( .A(n19646), .ZN(n19643) );
  OAI211_X1 U22607 ( .C1(n10480), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19643), 
        .B(n20013), .ZN(n19616) );
  OAI211_X1 U22608 ( .C1(n19618), .C2(n19617), .A(n19851), .B(n19616), .ZN(
        n19635) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19635), .B1(
        n19631), .B2(n19854), .ZN(n19619) );
  OAI211_X1 U22610 ( .C1(n19857), .C2(n19663), .A(n19620), .B(n19619), .ZN(
        P2_U3104) );
  AOI22_X1 U22611 ( .A1(n19634), .A2(n19858), .B1(n19859), .B2(n19646), .ZN(
        n19622) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19635), .B1(
        n19665), .B2(n19811), .ZN(n19621) );
  OAI211_X1 U22613 ( .C1(n19736), .C2(n19638), .A(n19622), .B(n19621), .ZN(
        P2_U3105) );
  AOI22_X1 U22614 ( .A1(n19634), .A2(n21348), .B1(n19646), .B2(n21344), .ZN(
        n19624) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19635), .B1(
        n19665), .B2(n19815), .ZN(n19623) );
  OAI211_X1 U22616 ( .C1(n19739), .C2(n19638), .A(n19624), .B(n19623), .ZN(
        P2_U3106) );
  AOI22_X1 U22617 ( .A1(n19634), .A2(n19872), .B1(n19646), .B2(n19873), .ZN(
        n19626) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19635), .B1(
        n19631), .B2(n19877), .ZN(n19625) );
  OAI211_X1 U22619 ( .C1(n19880), .C2(n19663), .A(n19626), .B(n19625), .ZN(
        P2_U3107) );
  AOI22_X1 U22620 ( .A1(n19634), .A2(n19881), .B1(n19646), .B2(n19882), .ZN(
        n19628) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19635), .B1(
        n19665), .B2(n19822), .ZN(n19627) );
  OAI211_X1 U22622 ( .C1(n19744), .C2(n19638), .A(n19628), .B(n19627), .ZN(
        P2_U3108) );
  AOI22_X1 U22623 ( .A1(n19634), .A2(n19890), .B1(n19646), .B2(n19891), .ZN(
        n19630) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19635), .B1(
        n19631), .B2(n19895), .ZN(n19629) );
  OAI211_X1 U22625 ( .C1(n19898), .C2(n19663), .A(n19630), .B(n19629), .ZN(
        P2_U3109) );
  AOI22_X1 U22626 ( .A1(n19634), .A2(n19782), .B1(n9707), .B2(n19646), .ZN(
        n19633) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19635), .B1(
        n19631), .B2(n19903), .ZN(n19632) );
  OAI211_X1 U22628 ( .C1(n19906), .C2(n19663), .A(n19633), .B(n19632), .ZN(
        P2_U3110) );
  AOI22_X1 U22629 ( .A1(n19634), .A2(n19907), .B1(n19908), .B2(n19646), .ZN(
        n19637) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19635), .B1(
        n19665), .B2(n19831), .ZN(n19636) );
  OAI211_X1 U22631 ( .C1(n19758), .C2(n19638), .A(n19637), .B(n19636), .ZN(
        P2_U3111) );
  NOR2_X1 U22632 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19639), .ZN(
        n19664) );
  AOI22_X1 U22633 ( .A1(n19854), .A2(n19665), .B1(n19842), .B2(n19664), .ZN(
        n19650) );
  AOI21_X1 U22634 ( .B1(n19683), .B2(n19663), .A(n19691), .ZN(n19640) );
  NOR2_X1 U22635 ( .A1(n19640), .A2(n20013), .ZN(n19645) );
  OAI21_X1 U22636 ( .B1(n10522), .B2(n19763), .A(n20033), .ZN(n19642) );
  AOI21_X1 U22637 ( .B1(n19645), .B2(n19643), .A(n19642), .ZN(n19644) );
  OAI21_X1 U22638 ( .B1(n19664), .B2(n19644), .A(n19851), .ZN(n19667) );
  OAI21_X1 U22639 ( .B1(n19646), .B2(n19664), .A(n19645), .ZN(n19648) );
  OAI21_X1 U22640 ( .B1(n10522), .B2(n19664), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19647) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19667), .B1(
        n19791), .B2(n19666), .ZN(n19649) );
  OAI211_X1 U22642 ( .C1(n19857), .C2(n19683), .A(n19650), .B(n19649), .ZN(
        P2_U3112) );
  AOI22_X1 U22643 ( .A1(n19863), .A2(n19665), .B1(n19859), .B2(n19664), .ZN(
        n19652) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19667), .B1(
        n19858), .B2(n19666), .ZN(n19651) );
  OAI211_X1 U22645 ( .C1(n19866), .C2(n19683), .A(n19652), .B(n19651), .ZN(
        P2_U3113) );
  AOI22_X1 U22646 ( .A1(n21346), .A2(n19665), .B1(n21344), .B2(n19664), .ZN(
        n19654) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19667), .B1(
        n21348), .B2(n19666), .ZN(n19653) );
  OAI211_X1 U22648 ( .C1(n21353), .C2(n19683), .A(n19654), .B(n19653), .ZN(
        P2_U3114) );
  AOI22_X1 U22649 ( .A1(n19877), .A2(n19665), .B1(n19873), .B2(n19664), .ZN(
        n19656) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19667), .B1(
        n19872), .B2(n19666), .ZN(n19655) );
  OAI211_X1 U22651 ( .C1(n19880), .C2(n19683), .A(n19656), .B(n19655), .ZN(
        P2_U3115) );
  AOI22_X1 U22652 ( .A1(n19886), .A2(n19665), .B1(n19882), .B2(n19664), .ZN(
        n19658) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19667), .B1(
        n19881), .B2(n19666), .ZN(n19657) );
  OAI211_X1 U22654 ( .C1(n19889), .C2(n19683), .A(n19658), .B(n19657), .ZN(
        P2_U3116) );
  AOI22_X1 U22655 ( .A1(n19826), .A2(n19685), .B1(n19891), .B2(n19664), .ZN(
        n19660) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19667), .B1(
        n19890), .B2(n19666), .ZN(n19659) );
  OAI211_X1 U22657 ( .C1(n19747), .C2(n19663), .A(n19660), .B(n19659), .ZN(
        P2_U3117) );
  AOI22_X1 U22658 ( .A1(n19748), .A2(n19685), .B1(n9707), .B2(n19664), .ZN(
        n19662) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19667), .B1(
        n19782), .B2(n19666), .ZN(n19661) );
  OAI211_X1 U22660 ( .C1(n19751), .C2(n19663), .A(n19662), .B(n19661), .ZN(
        P2_U3118) );
  AOI22_X1 U22661 ( .A1(n19914), .A2(n19665), .B1(n19908), .B2(n19664), .ZN(
        n19669) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19667), .B1(
        n19907), .B2(n19666), .ZN(n19668) );
  OAI211_X1 U22663 ( .C1(n19920), .C2(n19683), .A(n19669), .B(n19668), .ZN(
        P2_U3119) );
  AOI22_X1 U22664 ( .A1(n19815), .A2(n19714), .B1(n19684), .B2(n21344), .ZN(
        n19671) );
  AOI22_X1 U22665 ( .A1(n19685), .A2(n21346), .B1(n21348), .B2(n19686), .ZN(
        n19670) );
  OAI211_X1 U22666 ( .C1(n19678), .C2(n11100), .A(n19671), .B(n19670), .ZN(
        P2_U3122) );
  INV_X1 U22667 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n19674) );
  AOI22_X1 U22668 ( .A1(n19819), .A2(n19714), .B1(n19684), .B2(n19873), .ZN(
        n19673) );
  AOI22_X1 U22669 ( .A1(n19685), .A2(n19877), .B1(n19872), .B2(n19686), .ZN(
        n19672) );
  OAI211_X1 U22670 ( .C1(n19678), .C2(n19674), .A(n19673), .B(n19672), .ZN(
        P2_U3123) );
  AOI22_X1 U22671 ( .A1(n19822), .A2(n19714), .B1(n19684), .B2(n19882), .ZN(
        n19676) );
  AOI22_X1 U22672 ( .A1(n19685), .A2(n19886), .B1(n19881), .B2(n19686), .ZN(
        n19675) );
  OAI211_X1 U22673 ( .C1(n19678), .C2(n19677), .A(n19676), .B(n19675), .ZN(
        P2_U3124) );
  AOI22_X1 U22674 ( .A1(n19826), .A2(n19714), .B1(n19684), .B2(n19891), .ZN(
        n19680) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19687), .B1(
        n19890), .B2(n19686), .ZN(n19679) );
  OAI211_X1 U22676 ( .C1(n19747), .C2(n19683), .A(n19680), .B(n19679), .ZN(
        P2_U3125) );
  AOI22_X1 U22677 ( .A1(n19748), .A2(n19714), .B1(n9707), .B2(n19684), .ZN(
        n19682) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19687), .B1(
        n19782), .B2(n19686), .ZN(n19681) );
  OAI211_X1 U22679 ( .C1(n19751), .C2(n19683), .A(n19682), .B(n19681), .ZN(
        P2_U3126) );
  AOI22_X1 U22680 ( .A1(n19914), .A2(n19685), .B1(n19908), .B2(n19684), .ZN(
        n19689) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19687), .B1(
        n19907), .B2(n19686), .ZN(n19688) );
  OAI211_X1 U22682 ( .C1(n19920), .C2(n19723), .A(n19689), .B(n19688), .ZN(
        P2_U3127) );
  NAND3_X1 U22683 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20024), .ZN(n19727) );
  NOR2_X1 U22684 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19727), .ZN(
        n19717) );
  AOI22_X1 U22685 ( .A1(n19854), .A2(n19714), .B1(n19842), .B2(n19717), .ZN(
        n19703) );
  AOI21_X1 U22686 ( .B1(n19723), .B2(n19757), .A(n19691), .ZN(n19692) );
  NOR2_X1 U22687 ( .A1(n19692), .A2(n20013), .ZN(n19697) );
  AND2_X1 U22688 ( .A1(n20024), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19693) );
  NAND2_X1 U22689 ( .A1(n19694), .A2(n19693), .ZN(n19700) );
  NAND2_X1 U22690 ( .A1(n19697), .A2(n19700), .ZN(n19695) );
  OAI211_X1 U22691 ( .C1(n19717), .C2(n19696), .A(n19695), .B(n19851), .ZN(
        n19720) );
  INV_X1 U22692 ( .A(n19697), .ZN(n19701) );
  OAI21_X1 U22693 ( .B1(n19698), .B2(n19717), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19699) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19720), .B1(
        n19791), .B2(n19719), .ZN(n19702) );
  OAI211_X1 U22695 ( .C1(n19857), .C2(n19757), .A(n19703), .B(n19702), .ZN(
        P2_U3128) );
  INV_X1 U22696 ( .A(n19757), .ZN(n19718) );
  AOI22_X1 U22697 ( .A1(n19811), .A2(n19718), .B1(n19859), .B2(n19717), .ZN(
        n19705) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19720), .B1(
        n19858), .B2(n19719), .ZN(n19704) );
  OAI211_X1 U22699 ( .C1(n19736), .C2(n19723), .A(n19705), .B(n19704), .ZN(
        P2_U3129) );
  AOI22_X1 U22700 ( .A1(n19815), .A2(n19718), .B1(n21344), .B2(n19717), .ZN(
        n19707) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19720), .B1(
        n21348), .B2(n19719), .ZN(n19706) );
  OAI211_X1 U22702 ( .C1(n19739), .C2(n19723), .A(n19707), .B(n19706), .ZN(
        P2_U3130) );
  AOI22_X1 U22703 ( .A1(n19877), .A2(n19714), .B1(n19873), .B2(n19717), .ZN(
        n19709) );
  AOI22_X1 U22704 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19720), .B1(
        n19872), .B2(n19719), .ZN(n19708) );
  OAI211_X1 U22705 ( .C1(n19880), .C2(n19757), .A(n19709), .B(n19708), .ZN(
        P2_U3131) );
  AOI22_X1 U22706 ( .A1(n19886), .A2(n19714), .B1(n19882), .B2(n19717), .ZN(
        n19711) );
  AOI22_X1 U22707 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19720), .B1(
        n19881), .B2(n19719), .ZN(n19710) );
  OAI211_X1 U22708 ( .C1(n19889), .C2(n19757), .A(n19711), .B(n19710), .ZN(
        P2_U3132) );
  AOI22_X1 U22709 ( .A1(n19895), .A2(n19714), .B1(n19891), .B2(n19717), .ZN(
        n19713) );
  AOI22_X1 U22710 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19720), .B1(
        n19890), .B2(n19719), .ZN(n19712) );
  OAI211_X1 U22711 ( .C1(n19898), .C2(n19757), .A(n19713), .B(n19712), .ZN(
        P2_U3133) );
  AOI22_X1 U22712 ( .A1(n19903), .A2(n19714), .B1(n9707), .B2(n19717), .ZN(
        n19716) );
  AOI22_X1 U22713 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19720), .B1(
        n19782), .B2(n19719), .ZN(n19715) );
  OAI211_X1 U22714 ( .C1(n19906), .C2(n19757), .A(n19716), .B(n19715), .ZN(
        P2_U3134) );
  AOI22_X1 U22715 ( .A1(n19831), .A2(n19718), .B1(n19908), .B2(n19717), .ZN(
        n19722) );
  AOI22_X1 U22716 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19720), .B1(
        n19907), .B2(n19719), .ZN(n19721) );
  OAI211_X1 U22717 ( .C1(n19758), .C2(n19723), .A(n19722), .B(n19721), .ZN(
        P2_U3135) );
  NOR2_X1 U22718 ( .A1(n20040), .A2(n19727), .ZN(n19752) );
  OAI21_X1 U22719 ( .B1(n19725), .B2(n19752), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19724) );
  OAI21_X1 U22720 ( .B1(n19727), .B2(n20013), .A(n19724), .ZN(n19753) );
  AOI22_X1 U22721 ( .A1(n19753), .A2(n19791), .B1(n19842), .B2(n19752), .ZN(
        n19732) );
  INV_X1 U22722 ( .A(n19725), .ZN(n19726) );
  AOI21_X1 U22723 ( .B1(n19726), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19729) );
  OAI21_X1 U22724 ( .B1(n19847), .B2(n20003), .A(n19727), .ZN(n19728) );
  OAI211_X1 U22725 ( .C1(n19752), .C2(n19729), .A(n19728), .B(n19851), .ZN(
        n19754) );
  NOR2_X2 U22726 ( .A1(n19730), .A2(n20003), .ZN(n19787) );
  AOI22_X1 U22727 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19754), .B1(
        n19787), .B2(n19792), .ZN(n19731) );
  OAI211_X1 U22728 ( .C1(n19733), .C2(n19757), .A(n19732), .B(n19731), .ZN(
        P2_U3136) );
  AOI22_X1 U22729 ( .A1(n19753), .A2(n19858), .B1(n19859), .B2(n19752), .ZN(
        n19735) );
  AOI22_X1 U22730 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19754), .B1(
        n19787), .B2(n19811), .ZN(n19734) );
  OAI211_X1 U22731 ( .C1(n19736), .C2(n19757), .A(n19735), .B(n19734), .ZN(
        P2_U3137) );
  AOI22_X1 U22732 ( .A1(n19753), .A2(n21348), .B1(n21344), .B2(n19752), .ZN(
        n19738) );
  AOI22_X1 U22733 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19754), .B1(
        n19787), .B2(n19815), .ZN(n19737) );
  OAI211_X1 U22734 ( .C1(n19739), .C2(n19757), .A(n19738), .B(n19737), .ZN(
        P2_U3138) );
  AOI22_X1 U22735 ( .A1(n19753), .A2(n19872), .B1(n19873), .B2(n19752), .ZN(
        n19741) );
  AOI22_X1 U22736 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19754), .B1(
        n19787), .B2(n19819), .ZN(n19740) );
  OAI211_X1 U22737 ( .C1(n19802), .C2(n19757), .A(n19741), .B(n19740), .ZN(
        P2_U3139) );
  AOI22_X1 U22738 ( .A1(n19753), .A2(n19881), .B1(n19882), .B2(n19752), .ZN(
        n19743) );
  AOI22_X1 U22739 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19754), .B1(
        n19787), .B2(n19822), .ZN(n19742) );
  OAI211_X1 U22740 ( .C1(n19744), .C2(n19757), .A(n19743), .B(n19742), .ZN(
        P2_U3140) );
  AOI22_X1 U22741 ( .A1(n19753), .A2(n19890), .B1(n19891), .B2(n19752), .ZN(
        n19746) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19754), .B1(
        n19787), .B2(n19826), .ZN(n19745) );
  OAI211_X1 U22743 ( .C1(n19747), .C2(n19757), .A(n19746), .B(n19745), .ZN(
        P2_U3141) );
  AOI22_X1 U22744 ( .A1(n19753), .A2(n19782), .B1(n9707), .B2(n19752), .ZN(
        n19750) );
  AOI22_X1 U22745 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19754), .B1(
        n19787), .B2(n19748), .ZN(n19749) );
  OAI211_X1 U22746 ( .C1(n19751), .C2(n19757), .A(n19750), .B(n19749), .ZN(
        P2_U3142) );
  AOI22_X1 U22747 ( .A1(n19753), .A2(n19907), .B1(n19908), .B2(n19752), .ZN(
        n19756) );
  AOI22_X1 U22748 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19754), .B1(
        n19787), .B2(n19831), .ZN(n19755) );
  OAI211_X1 U22749 ( .C1(n19758), .C2(n19757), .A(n19756), .B(n19755), .ZN(
        P2_U3143) );
  NAND3_X1 U22750 ( .A1(n19764), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n20033), .ZN(n19762) );
  INV_X1 U22751 ( .A(n19759), .ZN(n19761) );
  NOR2_X1 U22752 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19760), .ZN(
        n19785) );
  NOR3_X1 U22753 ( .A1(n19761), .A2(n19785), .A3(n19763), .ZN(n19766) );
  AOI21_X1 U22754 ( .B1(n19763), .B2(n19762), .A(n19766), .ZN(n19786) );
  AOI22_X1 U22755 ( .A1(n19786), .A2(n19791), .B1(n19842), .B2(n19785), .ZN(
        n19771) );
  OAI21_X1 U22756 ( .B1(n19787), .B2(n19807), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19768) );
  NAND2_X1 U22757 ( .A1(n19764), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19767) );
  AOI211_X1 U22758 ( .C1(n19768), .C2(n19767), .A(n19766), .B(n19765), .ZN(
        n19769) );
  AOI22_X1 U22759 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19788), .B1(
        n19787), .B2(n19854), .ZN(n19770) );
  OAI211_X1 U22760 ( .C1(n19857), .C2(n19801), .A(n19771), .B(n19770), .ZN(
        P2_U3144) );
  AOI22_X1 U22761 ( .A1(n19786), .A2(n19858), .B1(n19859), .B2(n19785), .ZN(
        n19773) );
  AOI22_X1 U22762 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19788), .B1(
        n19787), .B2(n19863), .ZN(n19772) );
  OAI211_X1 U22763 ( .C1(n19866), .C2(n19801), .A(n19773), .B(n19772), .ZN(
        P2_U3145) );
  AOI22_X1 U22764 ( .A1(n19786), .A2(n21348), .B1(n21344), .B2(n19785), .ZN(
        n19775) );
  AOI22_X1 U22765 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19788), .B1(
        n19787), .B2(n21346), .ZN(n19774) );
  OAI211_X1 U22766 ( .C1(n21353), .C2(n19801), .A(n19775), .B(n19774), .ZN(
        P2_U3146) );
  AOI22_X1 U22767 ( .A1(n19786), .A2(n19872), .B1(n19873), .B2(n19785), .ZN(
        n19777) );
  AOI22_X1 U22768 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19788), .B1(
        n19787), .B2(n19877), .ZN(n19776) );
  OAI211_X1 U22769 ( .C1(n19880), .C2(n19801), .A(n19777), .B(n19776), .ZN(
        P2_U3147) );
  AOI22_X1 U22770 ( .A1(n19786), .A2(n19881), .B1(n19882), .B2(n19785), .ZN(
        n19779) );
  AOI22_X1 U22771 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19788), .B1(
        n19787), .B2(n19886), .ZN(n19778) );
  OAI211_X1 U22772 ( .C1(n19889), .C2(n19801), .A(n19779), .B(n19778), .ZN(
        P2_U3148) );
  AOI22_X1 U22773 ( .A1(n19786), .A2(n19890), .B1(n19891), .B2(n19785), .ZN(
        n19781) );
  AOI22_X1 U22774 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19788), .B1(
        n19787), .B2(n19895), .ZN(n19780) );
  OAI211_X1 U22775 ( .C1(n19898), .C2(n19801), .A(n19781), .B(n19780), .ZN(
        P2_U3149) );
  AOI22_X1 U22776 ( .A1(n19786), .A2(n19782), .B1(n9707), .B2(n19785), .ZN(
        n19784) );
  AOI22_X1 U22777 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19788), .B1(
        n19787), .B2(n19903), .ZN(n19783) );
  OAI211_X1 U22778 ( .C1(n19906), .C2(n19801), .A(n19784), .B(n19783), .ZN(
        P2_U3150) );
  AOI22_X1 U22779 ( .A1(n19786), .A2(n19907), .B1(n19908), .B2(n19785), .ZN(
        n19790) );
  AOI22_X1 U22780 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19788), .B1(
        n19787), .B2(n19914), .ZN(n19789) );
  OAI211_X1 U22781 ( .C1(n19920), .C2(n19801), .A(n19790), .B(n19789), .ZN(
        P2_U3151) );
  INV_X1 U22782 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n19795) );
  AOI22_X1 U22783 ( .A1(n19806), .A2(n19791), .B1(n19805), .B2(n19842), .ZN(
        n19794) );
  AOI22_X1 U22784 ( .A1(n19807), .A2(n19854), .B1(n19832), .B2(n19792), .ZN(
        n19793) );
  OAI211_X1 U22785 ( .C1(n19810), .C2(n19795), .A(n19794), .B(n19793), .ZN(
        P2_U3152) );
  AOI22_X1 U22786 ( .A1(n19806), .A2(n21348), .B1(n19805), .B2(n21344), .ZN(
        n19797) );
  AOI22_X1 U22787 ( .A1(n19807), .A2(n21346), .B1(n19832), .B2(n19815), .ZN(
        n19796) );
  OAI211_X1 U22788 ( .C1(n19810), .C2(n11099), .A(n19797), .B(n19796), .ZN(
        P2_U3154) );
  AOI22_X1 U22789 ( .A1(n19806), .A2(n19872), .B1(n19805), .B2(n19873), .ZN(
        n19800) );
  AOI22_X1 U22790 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19798), .B1(
        n19832), .B2(n19819), .ZN(n19799) );
  OAI211_X1 U22791 ( .C1(n19802), .C2(n19801), .A(n19800), .B(n19799), .ZN(
        P2_U3155) );
  INV_X1 U22792 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n21275) );
  AOI22_X1 U22793 ( .A1(n19806), .A2(n19881), .B1(n19805), .B2(n19882), .ZN(
        n19804) );
  AOI22_X1 U22794 ( .A1(n19807), .A2(n19886), .B1(n19832), .B2(n19822), .ZN(
        n19803) );
  OAI211_X1 U22795 ( .C1(n19810), .C2(n21275), .A(n19804), .B(n19803), .ZN(
        P2_U3156) );
  AOI22_X1 U22796 ( .A1(n19806), .A2(n19890), .B1(n19805), .B2(n19891), .ZN(
        n19809) );
  AOI22_X1 U22797 ( .A1(n19832), .A2(n19826), .B1(n19807), .B2(n19895), .ZN(
        n19808) );
  OAI211_X1 U22798 ( .C1(n19810), .C2(n11156), .A(n19809), .B(n19808), .ZN(
        P2_U3157) );
  INV_X1 U22799 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n19814) );
  AOI22_X1 U22800 ( .A1(n19863), .A2(n19832), .B1(n19859), .B2(n19830), .ZN(
        n19813) );
  AOI22_X1 U22801 ( .A1(n19858), .A2(n19833), .B1(n19915), .B2(n19811), .ZN(
        n19812) );
  OAI211_X1 U22802 ( .C1(n19837), .C2(n19814), .A(n19813), .B(n19812), .ZN(
        P2_U3161) );
  INV_X1 U22803 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19818) );
  AOI22_X1 U22804 ( .A1(n21346), .A2(n19832), .B1(n19830), .B2(n21344), .ZN(
        n19817) );
  AOI22_X1 U22805 ( .A1(n21348), .A2(n19833), .B1(n19915), .B2(n19815), .ZN(
        n19816) );
  OAI211_X1 U22806 ( .C1(n19837), .C2(n19818), .A(n19817), .B(n19816), .ZN(
        P2_U3162) );
  AOI22_X1 U22807 ( .A1(n19819), .A2(n19915), .B1(n19830), .B2(n19873), .ZN(
        n19821) );
  AOI22_X1 U22808 ( .A1(n19872), .A2(n19833), .B1(n19832), .B2(n19877), .ZN(
        n19820) );
  OAI211_X1 U22809 ( .C1(n19837), .C2(n10417), .A(n19821), .B(n19820), .ZN(
        P2_U3163) );
  INV_X1 U22810 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U22811 ( .A1(n19886), .A2(n19832), .B1(n19830), .B2(n19882), .ZN(
        n19824) );
  AOI22_X1 U22812 ( .A1(n19881), .A2(n19833), .B1(n19915), .B2(n19822), .ZN(
        n19823) );
  OAI211_X1 U22813 ( .C1(n19837), .C2(n19825), .A(n19824), .B(n19823), .ZN(
        P2_U3164) );
  INV_X1 U22814 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n19829) );
  AOI22_X1 U22815 ( .A1(n19826), .A2(n19915), .B1(n19830), .B2(n19891), .ZN(
        n19828) );
  AOI22_X1 U22816 ( .A1(n19890), .A2(n19833), .B1(n19832), .B2(n19895), .ZN(
        n19827) );
  OAI211_X1 U22817 ( .C1(n19837), .C2(n19829), .A(n19828), .B(n19827), .ZN(
        P2_U3165) );
  INV_X1 U22818 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19836) );
  AOI22_X1 U22819 ( .A1(n19831), .A2(n19915), .B1(n19908), .B2(n19830), .ZN(
        n19835) );
  AOI22_X1 U22820 ( .A1(n19907), .A2(n19833), .B1(n19832), .B2(n19914), .ZN(
        n19834) );
  OAI211_X1 U22821 ( .C1(n19837), .C2(n19836), .A(n19835), .B(n19834), .ZN(
        P2_U3167) );
  NAND2_X1 U22822 ( .A1(n19910), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19838) );
  NOR2_X1 U22823 ( .A1(n19839), .A2(n19838), .ZN(n19848) );
  INV_X1 U22824 ( .A(n19849), .ZN(n19840) );
  AOI21_X1 U22825 ( .B1(n20033), .B2(n19840), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19841) );
  INV_X1 U22826 ( .A(n19842), .ZN(n19843) );
  OAI22_X1 U22827 ( .A1(n19912), .A2(n19844), .B1(n19910), .B2(n19843), .ZN(
        n19845) );
  INV_X1 U22828 ( .A(n19845), .ZN(n19856) );
  OR2_X1 U22829 ( .A1(n19847), .A2(n19846), .ZN(n19850) );
  AOI21_X1 U22830 ( .B1(n19850), .B2(n19849), .A(n19848), .ZN(n19852) );
  OAI211_X1 U22831 ( .C1(n19853), .C2(n20033), .A(n19852), .B(n19851), .ZN(
        n19916) );
  AOI22_X1 U22832 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n19854), .ZN(n19855) );
  OAI211_X1 U22833 ( .C1(n19857), .C2(n19919), .A(n19856), .B(n19855), .ZN(
        P2_U3168) );
  INV_X1 U22834 ( .A(n19858), .ZN(n19861) );
  INV_X1 U22835 ( .A(n19859), .ZN(n19860) );
  OAI22_X1 U22836 ( .A1(n19912), .A2(n19861), .B1(n19910), .B2(n19860), .ZN(
        n19862) );
  INV_X1 U22837 ( .A(n19862), .ZN(n19865) );
  AOI22_X1 U22838 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n19863), .ZN(n19864) );
  OAI211_X1 U22839 ( .C1(n19866), .C2(n19919), .A(n19865), .B(n19864), .ZN(
        P2_U3169) );
  INV_X1 U22840 ( .A(n21348), .ZN(n19868) );
  INV_X1 U22841 ( .A(n21344), .ZN(n19867) );
  OAI22_X1 U22842 ( .A1(n19912), .A2(n19868), .B1(n19910), .B2(n19867), .ZN(
        n19869) );
  INV_X1 U22843 ( .A(n19869), .ZN(n19871) );
  AOI22_X1 U22844 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n21346), .ZN(n19870) );
  OAI211_X1 U22845 ( .C1(n21353), .C2(n19919), .A(n19871), .B(n19870), .ZN(
        P2_U3170) );
  INV_X1 U22846 ( .A(n19872), .ZN(n19875) );
  INV_X1 U22847 ( .A(n19873), .ZN(n19874) );
  OAI22_X1 U22848 ( .A1(n19912), .A2(n19875), .B1(n19910), .B2(n19874), .ZN(
        n19876) );
  INV_X1 U22849 ( .A(n19876), .ZN(n19879) );
  AOI22_X1 U22850 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n19877), .ZN(n19878) );
  OAI211_X1 U22851 ( .C1(n19880), .C2(n19919), .A(n19879), .B(n19878), .ZN(
        P2_U3171) );
  INV_X1 U22852 ( .A(n19881), .ZN(n19884) );
  INV_X1 U22853 ( .A(n19882), .ZN(n19883) );
  OAI22_X1 U22854 ( .A1(n19912), .A2(n19884), .B1(n19910), .B2(n19883), .ZN(
        n19885) );
  INV_X1 U22855 ( .A(n19885), .ZN(n19888) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n19886), .ZN(n19887) );
  OAI211_X1 U22857 ( .C1(n19889), .C2(n19919), .A(n19888), .B(n19887), .ZN(
        P2_U3172) );
  INV_X1 U22858 ( .A(n19890), .ZN(n19893) );
  INV_X1 U22859 ( .A(n19891), .ZN(n19892) );
  OAI22_X1 U22860 ( .A1(n19912), .A2(n19893), .B1(n19910), .B2(n19892), .ZN(
        n19894) );
  INV_X1 U22861 ( .A(n19894), .ZN(n19897) );
  AOI22_X1 U22862 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n19895), .ZN(n19896) );
  OAI211_X1 U22863 ( .C1(n19898), .C2(n19919), .A(n19897), .B(n19896), .ZN(
        P2_U3173) );
  OAI22_X1 U22865 ( .A1(n19912), .A2(n19901), .B1(n19910), .B2(n21356), .ZN(
        n19902) );
  INV_X1 U22866 ( .A(n19902), .ZN(n19905) );
  AOI22_X1 U22867 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n19903), .ZN(n19904) );
  OAI211_X1 U22868 ( .C1(n19906), .C2(n19919), .A(n19905), .B(n19904), .ZN(
        P2_U3174) );
  INV_X1 U22869 ( .A(n19907), .ZN(n19911) );
  INV_X1 U22870 ( .A(n19908), .ZN(n19909) );
  OAI22_X1 U22871 ( .A1(n19912), .A2(n19911), .B1(n19910), .B2(n19909), .ZN(
        n19913) );
  INV_X1 U22872 ( .A(n19913), .ZN(n19918) );
  AOI22_X1 U22873 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19916), .B1(
        n19915), .B2(n19914), .ZN(n19917) );
  OAI211_X1 U22874 ( .C1(n19920), .C2(n19919), .A(n19918), .B(n19917), .ZN(
        P2_U3175) );
  NOR3_X1 U22875 ( .A1(n19942), .A2(n20006), .A3(n12955), .ZN(n19925) );
  AOI211_X1 U22876 ( .C1(n19923), .C2(n19926), .A(n19922), .B(n19921), .ZN(
        n19924) );
  AOI221_X1 U22877 ( .B1(n19927), .B2(n19926), .C1(n19925), .C2(n19926), .A(
        n19924), .ZN(n19929) );
  NAND2_X1 U22878 ( .A1(n19929), .A2(n19928), .ZN(P2_U3177) );
  AND2_X1 U22879 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19930), .ZN(
        P2_U3179) );
  AND2_X1 U22880 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19930), .ZN(
        P2_U3180) );
  AND2_X1 U22881 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19930), .ZN(
        P2_U3181) );
  AND2_X1 U22882 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19930), .ZN(
        P2_U3182) );
  AND2_X1 U22883 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19930), .ZN(
        P2_U3183) );
  AND2_X1 U22884 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19930), .ZN(
        P2_U3184) );
  AND2_X1 U22885 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19930), .ZN(
        P2_U3185) );
  AND2_X1 U22886 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19930), .ZN(
        P2_U3186) );
  AND2_X1 U22887 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19930), .ZN(
        P2_U3187) );
  AND2_X1 U22888 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19930), .ZN(
        P2_U3188) );
  AND2_X1 U22889 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19930), .ZN(
        P2_U3189) );
  AND2_X1 U22890 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19930), .ZN(
        P2_U3190) );
  AND2_X1 U22891 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19930), .ZN(
        P2_U3191) );
  AND2_X1 U22892 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19930), .ZN(
        P2_U3192) );
  AND2_X1 U22893 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19930), .ZN(
        P2_U3193) );
  AND2_X1 U22894 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19930), .ZN(
        P2_U3194) );
  AND2_X1 U22895 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19930), .ZN(
        P2_U3195) );
  AND2_X1 U22896 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19930), .ZN(
        P2_U3196) );
  AND2_X1 U22897 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19930), .ZN(
        P2_U3197) );
  AND2_X1 U22898 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19930), .ZN(
        P2_U3198) );
  AND2_X1 U22899 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19930), .ZN(
        P2_U3199) );
  AND2_X1 U22900 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19930), .ZN(
        P2_U3200) );
  AND2_X1 U22901 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19930), .ZN(P2_U3201) );
  AND2_X1 U22902 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19930), .ZN(P2_U3202) );
  AND2_X1 U22903 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19930), .ZN(P2_U3203) );
  AND2_X1 U22904 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19930), .ZN(P2_U3204) );
  AND2_X1 U22905 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19930), .ZN(P2_U3205) );
  AND2_X1 U22906 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19930), .ZN(P2_U3206) );
  AND2_X1 U22907 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19930), .ZN(P2_U3207) );
  AND2_X1 U22908 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19930), .ZN(P2_U3208) );
  NAND2_X1 U22909 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19942), .ZN(n19944) );
  NAND3_X1 U22910 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19944), .ZN(n19932) );
  AOI211_X1 U22911 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20937), .A(
        n19943), .B(n20052), .ZN(n19931) );
  NOR2_X1 U22912 ( .A1(n20930), .A2(n19936), .ZN(n19949) );
  AOI211_X1 U22913 ( .C1(n19950), .C2(n19932), .A(n19931), .B(n19949), .ZN(
        n19933) );
  INV_X1 U22914 ( .A(n19933), .ZN(P2_U3209) );
  INV_X1 U22915 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19934) );
  AOI21_X1 U22916 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20937), .A(n19950), 
        .ZN(n19940) );
  NOR2_X1 U22917 ( .A1(n19934), .A2(n19940), .ZN(n19937) );
  AOI21_X1 U22918 ( .B1(n19937), .B2(n19936), .A(n19935), .ZN(n19938) );
  OAI211_X1 U22919 ( .C1(n20937), .C2(n19939), .A(n19938), .B(n19944), .ZN(
        P2_U3210) );
  AOI21_X1 U22920 ( .B1(n19942), .B2(n19941), .A(n19940), .ZN(n19948) );
  INV_X1 U22921 ( .A(n19943), .ZN(n19945) );
  OAI22_X1 U22922 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19945), .B1(NA), 
        .B2(n19944), .ZN(n19946) );
  OAI211_X1 U22923 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19946), .ZN(n19947) );
  OAI21_X1 U22924 ( .B1(n19949), .B2(n19948), .A(n19947), .ZN(P2_U3211) );
  OAI222_X1 U22925 ( .A1(n19995), .A2(n19953), .B1(n19952), .B2(n20052), .C1(
        n19951), .C2(n19993), .ZN(P2_U3212) );
  OAI222_X1 U22926 ( .A1(n19995), .A2(n14174), .B1(n21183), .B2(n20052), .C1(
        n19953), .C2(n19993), .ZN(P2_U3213) );
  OAI222_X1 U22927 ( .A1(n19995), .A2(n19955), .B1(n19954), .B2(n20052), .C1(
        n14174), .C2(n19993), .ZN(P2_U3214) );
  OAI222_X1 U22928 ( .A1(n19995), .A2(n14307), .B1(n19956), .B2(n20052), .C1(
        n19955), .C2(n19993), .ZN(P2_U3215) );
  OAI222_X1 U22929 ( .A1(n19995), .A2(n19958), .B1(n19957), .B2(n20052), .C1(
        n14307), .C2(n19993), .ZN(P2_U3216) );
  OAI222_X1 U22930 ( .A1(n19995), .A2(n15508), .B1(n19959), .B2(n20052), .C1(
        n19958), .C2(n19993), .ZN(P2_U3217) );
  OAI222_X1 U22931 ( .A1(n19995), .A2(n14269), .B1(n19960), .B2(n20052), .C1(
        n15508), .C2(n19993), .ZN(P2_U3218) );
  OAI222_X1 U22932 ( .A1(n19995), .A2(n19962), .B1(n19961), .B2(n20052), .C1(
        n14269), .C2(n19993), .ZN(P2_U3219) );
  OAI222_X1 U22933 ( .A1(n19995), .A2(n19188), .B1(n19963), .B2(n20052), .C1(
        n19962), .C2(n19993), .ZN(P2_U3220) );
  OAI222_X1 U22934 ( .A1(n19995), .A2(n19965), .B1(n19964), .B2(n20052), .C1(
        n19188), .C2(n19993), .ZN(P2_U3221) );
  OAI222_X1 U22935 ( .A1(n19995), .A2(n19967), .B1(n19966), .B2(n20052), .C1(
        n19965), .C2(n19993), .ZN(P2_U3222) );
  OAI222_X1 U22936 ( .A1(n19995), .A2(n21161), .B1(n19968), .B2(n20052), .C1(
        n19967), .C2(n19993), .ZN(P2_U3223) );
  INV_X1 U22937 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19969) );
  OAI222_X1 U22938 ( .A1(n19995), .A2(n19969), .B1(n21157), .B2(n20052), .C1(
        n21161), .C2(n19993), .ZN(P2_U3224) );
  INV_X1 U22939 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19971) );
  OAI222_X1 U22940 ( .A1(n19995), .A2(n19971), .B1(n19970), .B2(n20052), .C1(
        n19969), .C2(n19993), .ZN(P2_U3225) );
  OAI222_X1 U22941 ( .A1(n19995), .A2(n10855), .B1(n19972), .B2(n20052), .C1(
        n19971), .C2(n19993), .ZN(P2_U3226) );
  OAI222_X1 U22942 ( .A1(n19995), .A2(n15436), .B1(n19973), .B2(n20052), .C1(
        n10855), .C2(n19993), .ZN(P2_U3227) );
  OAI222_X1 U22943 ( .A1(n19995), .A2(n19974), .B1(n21304), .B2(n20052), .C1(
        n15436), .C2(n19993), .ZN(P2_U3228) );
  OAI222_X1 U22944 ( .A1(n19995), .A2(n19976), .B1(n19975), .B2(n20052), .C1(
        n19974), .C2(n19993), .ZN(P2_U3229) );
  OAI222_X1 U22945 ( .A1(n19995), .A2(n19978), .B1(n19977), .B2(n20052), .C1(
        n19976), .C2(n19993), .ZN(P2_U3230) );
  OAI222_X1 U22946 ( .A1(n19995), .A2(n19979), .B1(n21121), .B2(n20052), .C1(
        n19978), .C2(n19993), .ZN(P2_U3231) );
  OAI222_X1 U22947 ( .A1(n19995), .A2(n19980), .B1(n21186), .B2(n20052), .C1(
        n19979), .C2(n19993), .ZN(P2_U3232) );
  OAI222_X1 U22948 ( .A1(n19995), .A2(n19982), .B1(n19981), .B2(n20052), .C1(
        n19980), .C2(n19993), .ZN(P2_U3233) );
  OAI222_X1 U22949 ( .A1(n19995), .A2(n19984), .B1(n19983), .B2(n20052), .C1(
        n19982), .C2(n19993), .ZN(P2_U3234) );
  OAI222_X1 U22950 ( .A1(n19995), .A2(n19986), .B1(n19985), .B2(n20052), .C1(
        n19984), .C2(n19993), .ZN(P2_U3235) );
  OAI222_X1 U22951 ( .A1(n19995), .A2(n15333), .B1(n19987), .B2(n20052), .C1(
        n19986), .C2(n19993), .ZN(P2_U3236) );
  OAI222_X1 U22952 ( .A1(n19995), .A2(n19989), .B1(n19988), .B2(n20052), .C1(
        n15333), .C2(n19993), .ZN(P2_U3237) );
  OAI222_X1 U22953 ( .A1(n19993), .A2(n19989), .B1(n21152), .B2(n20052), .C1(
        n21168), .C2(n19995), .ZN(P2_U3238) );
  OAI222_X1 U22954 ( .A1(n19995), .A2(n19991), .B1(n19990), .B2(n20052), .C1(
        n21168), .C2(n19993), .ZN(P2_U3239) );
  INV_X1 U22955 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n21173) );
  OAI222_X1 U22956 ( .A1(n19995), .A2(n21173), .B1(n19992), .B2(n20052), .C1(
        n19991), .C2(n19993), .ZN(P2_U3240) );
  OAI222_X1 U22957 ( .A1(n19995), .A2(n11266), .B1(n19994), .B2(n20052), .C1(
        n21173), .C2(n19993), .ZN(P2_U3241) );
  OAI22_X1 U22958 ( .A1(n20053), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20052), .ZN(n19996) );
  INV_X1 U22959 ( .A(n19996), .ZN(P2_U3585) );
  MUX2_X1 U22960 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20053), .Z(P2_U3586) );
  OAI22_X1 U22961 ( .A1(n20053), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20052), .ZN(n19997) );
  INV_X1 U22962 ( .A(n19997), .ZN(P2_U3587) );
  OAI22_X1 U22963 ( .A1(n20053), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20052), .ZN(n19998) );
  INV_X1 U22964 ( .A(n19998), .ZN(P2_U3588) );
  OAI21_X1 U22965 ( .B1(n20002), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20000), 
        .ZN(n19999) );
  INV_X1 U22966 ( .A(n19999), .ZN(P2_U3591) );
  OAI21_X1 U22967 ( .B1(n20002), .B2(n20001), .A(n20000), .ZN(P2_U3592) );
  INV_X1 U22968 ( .A(n20003), .ZN(n20005) );
  AND2_X1 U22969 ( .A1(n20004), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20028) );
  NAND2_X1 U22970 ( .A1(n20005), .A2(n20028), .ZN(n20018) );
  NAND3_X1 U22971 ( .A1(n20026), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20006), 
        .ZN(n20008) );
  NAND2_X1 U22972 ( .A1(n20008), .A2(n20007), .ZN(n20019) );
  NAND2_X1 U22973 ( .A1(n20018), .A2(n20019), .ZN(n20010) );
  AOI22_X1 U22974 ( .A1(n20011), .A2(n20010), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20009), .ZN(n20012) );
  OAI21_X1 U22975 ( .B1(n20014), .B2(n20013), .A(n20012), .ZN(n20015) );
  INV_X1 U22976 ( .A(n20015), .ZN(n20016) );
  AOI22_X1 U22977 ( .A1(n20041), .A2(n20017), .B1(n20016), .B2(n20038), .ZN(
        P2_U3602) );
  OAI21_X1 U22978 ( .B1(n20020), .B2(n20019), .A(n20018), .ZN(n20021) );
  AOI21_X1 U22979 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20022), .A(n20021), 
        .ZN(n20023) );
  AOI22_X1 U22980 ( .A1(n20041), .A2(n20024), .B1(n20023), .B2(n20038), .ZN(
        P2_U3603) );
  NOR2_X1 U22981 ( .A1(n20034), .A2(n20025), .ZN(n20027) );
  MUX2_X1 U22982 ( .A(n20028), .B(n20027), .S(n20026), .Z(n20029) );
  AOI21_X1 U22983 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20030), .A(n20029), 
        .ZN(n20031) );
  AOI22_X1 U22984 ( .A1(n20041), .A2(n20032), .B1(n20031), .B2(n20038), .ZN(
        P2_U3604) );
  OAI22_X1 U22985 ( .A1(n20035), .A2(n20034), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20033), .ZN(n20036) );
  AOI21_X1 U22986 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20037), .A(n20036), 
        .ZN(n20039) );
  AOI22_X1 U22987 ( .A1(n20041), .A2(n20040), .B1(n20039), .B2(n20038), .ZN(
        P2_U3605) );
  INV_X1 U22988 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20042) );
  AOI22_X1 U22989 ( .A1(n20052), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20042), 
        .B2(n20053), .ZN(P2_U3608) );
  INV_X1 U22990 ( .A(n20043), .ZN(n20047) );
  NAND2_X1 U22991 ( .A1(n20045), .A2(n20044), .ZN(n20046) );
  OAI211_X1 U22992 ( .C1(n20049), .C2(n20048), .A(n20047), .B(n20046), .ZN(
        n20051) );
  MUX2_X1 U22993 ( .A(P2_MORE_REG_SCAN_IN), .B(n20051), .S(n20050), .Z(
        P2_U3609) );
  OAI22_X1 U22994 ( .A1(n20053), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20052), .ZN(n20054) );
  INV_X1 U22995 ( .A(n20054), .ZN(P2_U3611) );
  AOI21_X1 U22996 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20940), .A(n20932), 
        .ZN(n20935) );
  INV_X1 U22997 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20055) );
  AOI21_X1 U22998 ( .B1(n20935), .B2(n20055), .A(n21009), .ZN(P1_U2802) );
  INV_X1 U22999 ( .A(n20056), .ZN(n20058) );
  OAI21_X1 U23000 ( .B1(n20058), .B2(n20057), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20059) );
  OAI21_X1 U23001 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20060), .A(n20059), 
        .ZN(P1_U2803) );
  INV_X2 U23002 ( .A(n21009), .ZN(n21022) );
  NOR2_X1 U23003 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20062) );
  OAI21_X1 U23004 ( .B1(n20062), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21022), .ZN(
        n20061) );
  OAI21_X1 U23005 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21022), .A(n20061), 
        .ZN(P1_U2804) );
  NOR2_X1 U23006 ( .A1(n21009), .A2(n20935), .ZN(n20990) );
  OAI21_X1 U23007 ( .B1(BS16), .B2(n20062), .A(n20990), .ZN(n20988) );
  OAI21_X1 U23008 ( .B1(n20990), .B2(n21012), .A(n20988), .ZN(P1_U2805) );
  OAI21_X1 U23009 ( .B1(n20064), .B2(n20063), .A(n20220), .ZN(P1_U2806) );
  NOR4_X1 U23010 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20068) );
  NOR4_X1 U23011 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20067) );
  NOR4_X1 U23012 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20066) );
  NOR4_X1 U23013 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20065) );
  NAND4_X1 U23014 ( .A1(n20068), .A2(n20067), .A3(n20066), .A4(n20065), .ZN(
        n20074) );
  NOR4_X1 U23015 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20072) );
  AOI211_X1 U23016 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20071) );
  NOR4_X1 U23017 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20070) );
  NOR4_X1 U23018 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20069) );
  NAND4_X1 U23019 ( .A1(n20072), .A2(n20071), .A3(n20070), .A4(n20069), .ZN(
        n20073) );
  NOR2_X1 U23020 ( .A1(n20074), .A2(n20073), .ZN(n21007) );
  INV_X1 U23021 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20076) );
  NOR3_X1 U23022 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20077) );
  OAI21_X1 U23023 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20077), .A(n21007), .ZN(
        n20075) );
  OAI21_X1 U23024 ( .B1(n21007), .B2(n20076), .A(n20075), .ZN(P1_U2807) );
  INV_X1 U23025 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20989) );
  AOI21_X1 U23026 ( .B1(n21000), .B2(n20989), .A(n20077), .ZN(n20079) );
  INV_X1 U23027 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20078) );
  INV_X1 U23028 ( .A(n21007), .ZN(n21002) );
  AOI22_X1 U23029 ( .A1(n21007), .A2(n20079), .B1(n20078), .B2(n21002), .ZN(
        P1_U2808) );
  NAND2_X1 U23030 ( .A1(n20080), .A2(n20106), .ZN(n20088) );
  AOI22_X1 U23031 ( .A1(n20081), .A2(n20131), .B1(n20127), .B2(n20144), .ZN(
        n20082) );
  OAI211_X1 U23032 ( .C1(n20094), .C2(n20083), .A(n20082), .B(n20100), .ZN(
        n20084) );
  AOI21_X1 U23033 ( .B1(n20133), .B2(P1_EBX_REG_9__SCAN_IN), .A(n20084), .ZN(
        n20087) );
  AOI22_X1 U23034 ( .A1(n20145), .A2(n20099), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n20085), .ZN(n20086) );
  OAI211_X1 U23035 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n20088), .A(n20087), .B(
        n20086), .ZN(P1_U2831) );
  INV_X1 U23036 ( .A(n20089), .ZN(n20090) );
  AOI22_X1 U23037 ( .A1(n20090), .A2(n20131), .B1(n20127), .B2(n9822), .ZN(
        n20103) );
  INV_X1 U23038 ( .A(n20091), .ZN(n20092) );
  NOR2_X1 U23039 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20092), .ZN(n20097) );
  OAI22_X1 U23040 ( .A1(n20095), .A2(n20152), .B1(n20094), .B2(n20093), .ZN(
        n20096) );
  AOI21_X1 U23041 ( .B1(n20097), .B2(n20106), .A(n20096), .ZN(n20102) );
  AOI22_X1 U23042 ( .A1(n20150), .A2(n20099), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n20098), .ZN(n20101) );
  NAND4_X1 U23043 ( .A1(n20103), .A2(n20102), .A3(n20101), .A4(n20100), .ZN(
        P1_U2833) );
  AOI22_X1 U23044 ( .A1(n20105), .A2(n20131), .B1(n20127), .B2(n20104), .ZN(
        n20112) );
  AOI22_X1 U23045 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20128), .B1(
        n20106), .B2(n20946), .ZN(n20111) );
  AOI21_X1 U23046 ( .B1(n20133), .B2(P1_EBX_REG_5__SCAN_IN), .A(n20232), .ZN(
        n20110) );
  AOI22_X1 U23047 ( .A1(n20108), .A2(n20136), .B1(n20107), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20109) );
  NAND4_X1 U23048 ( .A1(n20112), .A2(n20111), .A3(n20110), .A4(n20109), .ZN(
        P1_U2835) );
  AOI222_X1 U23049 ( .A1(n20563), .A2(n20129), .B1(n20127), .B2(n20113), .C1(
        n20128), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20124) );
  INV_X1 U23050 ( .A(n20114), .ZN(n20115) );
  AOI22_X1 U23051 ( .A1(n20133), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20115), .B2(
        n20131), .ZN(n20123) );
  OR2_X1 U23052 ( .A1(n20118), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20117) );
  AND2_X1 U23053 ( .A1(n20117), .A2(n20116), .ZN(n20134) );
  OAI21_X1 U23054 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n20118), .A(n20134), .ZN(
        n20119) );
  AOI22_X1 U23055 ( .A1(n20120), .A2(n20136), .B1(P1_REIP_REG_3__SCAN_IN), 
        .B2(n20119), .ZN(n20122) );
  NAND4_X1 U23056 ( .A1(n20139), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .A4(n13943), .ZN(n20121) );
  NAND4_X1 U23057 ( .A1(n20124), .A2(n20123), .A3(n20122), .A4(n20121), .ZN(
        P1_U2837) );
  INV_X1 U23058 ( .A(n13861), .ZN(n20247) );
  INV_X1 U23059 ( .A(n20125), .ZN(n20126) );
  AOI222_X1 U23060 ( .A1(n20247), .A2(n20129), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20128), .C1(n20127), .C2(
        n20126), .ZN(n20143) );
  INV_X1 U23061 ( .A(n20130), .ZN(n20132) );
  AOI22_X1 U23062 ( .A1(n20133), .A2(P1_EBX_REG_2__SCAN_IN), .B1(n20132), .B2(
        n20131), .ZN(n20142) );
  NOR2_X1 U23063 ( .A1(n20134), .A2(n20138), .ZN(n20135) );
  AOI21_X1 U23064 ( .B1(n20137), .B2(n20136), .A(n20135), .ZN(n20141) );
  NAND3_X1 U23065 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n20139), .A3(n20138), 
        .ZN(n20140) );
  NAND4_X1 U23066 ( .A1(n20143), .A2(n20142), .A3(n20141), .A4(n20140), .ZN(
        P1_U2838) );
  AOI22_X1 U23067 ( .A1(n20145), .A2(n20149), .B1(n20148), .B2(n20144), .ZN(
        n20146) );
  OAI21_X1 U23068 ( .B1(n20153), .B2(n20147), .A(n20146), .ZN(P1_U2863) );
  AOI22_X1 U23069 ( .A1(n20150), .A2(n20149), .B1(n20148), .B2(n9822), .ZN(
        n20151) );
  OAI21_X1 U23070 ( .B1(n20153), .B2(n20152), .A(n20151), .ZN(P1_U2865) );
  AOI22_X1 U23071 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20155) );
  OAI21_X1 U23072 ( .B1(n13597), .B2(n20179), .A(n20155), .ZN(P1_U2921) );
  AOI22_X1 U23073 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20156) );
  OAI21_X1 U23074 ( .B1(n14373), .B2(n20179), .A(n20156), .ZN(P1_U2922) );
  AOI22_X1 U23075 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20157) );
  OAI21_X1 U23076 ( .B1(n14429), .B2(n20179), .A(n20157), .ZN(P1_U2923) );
  AOI22_X1 U23077 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20158) );
  OAI21_X1 U23078 ( .B1(n14366), .B2(n20179), .A(n20158), .ZN(P1_U2924) );
  AOI22_X1 U23079 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20159) );
  OAI21_X1 U23080 ( .B1(n14426), .B2(n20179), .A(n20159), .ZN(P1_U2925) );
  INV_X1 U23081 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20161) );
  AOI22_X1 U23082 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20160) );
  OAI21_X1 U23083 ( .B1(n20161), .B2(n20179), .A(n20160), .ZN(P1_U2926) );
  AOI22_X1 U23084 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21019), .B1(n20163), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20162) );
  OAI21_X1 U23085 ( .B1(n14234), .B2(n20179), .A(n20162), .ZN(P1_U2927) );
  AOI22_X1 U23086 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21019), .B1(n20163), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20164) );
  OAI21_X1 U23087 ( .B1(n14215), .B2(n20179), .A(n20164), .ZN(P1_U2928) );
  AOI22_X1 U23088 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20165) );
  OAI21_X1 U23089 ( .B1(n14123), .B2(n20179), .A(n20165), .ZN(P1_U2929) );
  AOI22_X1 U23090 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20166) );
  OAI21_X1 U23091 ( .B1(n12454), .B2(n20179), .A(n20166), .ZN(P1_U2930) );
  AOI22_X1 U23092 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20167) );
  OAI21_X1 U23093 ( .B1(n20168), .B2(n20179), .A(n20167), .ZN(P1_U2931) );
  AOI22_X1 U23094 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20169) );
  OAI21_X1 U23095 ( .B1(n20170), .B2(n20179), .A(n20169), .ZN(P1_U2932) );
  AOI22_X1 U23096 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20171) );
  OAI21_X1 U23097 ( .B1(n20172), .B2(n20179), .A(n20171), .ZN(P1_U2933) );
  AOI22_X1 U23098 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20173) );
  OAI21_X1 U23099 ( .B1(n20174), .B2(n20179), .A(n20173), .ZN(P1_U2934) );
  AOI22_X1 U23100 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20175) );
  OAI21_X1 U23101 ( .B1(n20176), .B2(n20179), .A(n20175), .ZN(P1_U2935) );
  AOI22_X1 U23102 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21019), .B1(n20177), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20178) );
  OAI21_X1 U23103 ( .B1(n20180), .B2(n20179), .A(n20178), .ZN(P1_U2936) );
  AOI22_X1 U23104 ( .A1(n20216), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20215), .ZN(n20183) );
  INV_X1 U23105 ( .A(n20181), .ZN(n20182) );
  NAND2_X1 U23106 ( .A1(n20201), .A2(n20182), .ZN(n20203) );
  NAND2_X1 U23107 ( .A1(n20183), .A2(n20203), .ZN(P1_U2945) );
  AOI22_X1 U23108 ( .A1(n20216), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20186) );
  INV_X1 U23109 ( .A(n20184), .ZN(n20185) );
  NAND2_X1 U23110 ( .A1(n20201), .A2(n20185), .ZN(n20205) );
  NAND2_X1 U23111 ( .A1(n20186), .A2(n20205), .ZN(P1_U2946) );
  AOI22_X1 U23112 ( .A1(n20187), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20189) );
  NAND2_X1 U23113 ( .A1(n20201), .A2(n20188), .ZN(n20207) );
  NAND2_X1 U23114 ( .A1(n20189), .A2(n20207), .ZN(P1_U2947) );
  AOI22_X1 U23115 ( .A1(n20216), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20192) );
  INV_X1 U23116 ( .A(n20190), .ZN(n20191) );
  NAND2_X1 U23117 ( .A1(n20201), .A2(n20191), .ZN(n20209) );
  NAND2_X1 U23118 ( .A1(n20192), .A2(n20209), .ZN(P1_U2948) );
  AOI22_X1 U23119 ( .A1(n20216), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20195) );
  INV_X1 U23120 ( .A(n20193), .ZN(n20194) );
  NAND2_X1 U23121 ( .A1(n20201), .A2(n20194), .ZN(n20211) );
  NAND2_X1 U23122 ( .A1(n20195), .A2(n20211), .ZN(P1_U2949) );
  AOI22_X1 U23123 ( .A1(n20216), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20198) );
  INV_X1 U23124 ( .A(n20196), .ZN(n20197) );
  NAND2_X1 U23125 ( .A1(n20201), .A2(n20197), .ZN(n20213) );
  NAND2_X1 U23126 ( .A1(n20198), .A2(n20213), .ZN(P1_U2950) );
  AOI22_X1 U23127 ( .A1(n20216), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20215), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20202) );
  INV_X1 U23128 ( .A(n20199), .ZN(n20200) );
  NAND2_X1 U23129 ( .A1(n20201), .A2(n20200), .ZN(n20217) );
  NAND2_X1 U23130 ( .A1(n20202), .A2(n20217), .ZN(P1_U2951) );
  AOI22_X1 U23131 ( .A1(n20216), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20215), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20204) );
  NAND2_X1 U23132 ( .A1(n20204), .A2(n20203), .ZN(P1_U2960) );
  AOI22_X1 U23133 ( .A1(n20216), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20215), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20206) );
  NAND2_X1 U23134 ( .A1(n20206), .A2(n20205), .ZN(P1_U2961) );
  AOI22_X1 U23135 ( .A1(n20216), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20215), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20208) );
  NAND2_X1 U23136 ( .A1(n20208), .A2(n20207), .ZN(P1_U2962) );
  AOI22_X1 U23137 ( .A1(n20216), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20215), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20210) );
  NAND2_X1 U23138 ( .A1(n20210), .A2(n20209), .ZN(P1_U2963) );
  AOI22_X1 U23139 ( .A1(n20216), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20215), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20212) );
  NAND2_X1 U23140 ( .A1(n20212), .A2(n20211), .ZN(P1_U2964) );
  AOI22_X1 U23141 ( .A1(n20216), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20215), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20214) );
  NAND2_X1 U23142 ( .A1(n20214), .A2(n20213), .ZN(P1_U2965) );
  AOI22_X1 U23143 ( .A1(n20216), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20215), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20218) );
  NAND2_X1 U23144 ( .A1(n20218), .A2(n20217), .ZN(P1_U2966) );
  OAI22_X1 U23145 ( .A1(n20221), .A2(n20220), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20219), .ZN(n20222) );
  AOI211_X1 U23146 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20228), .A(
        n20223), .B(n20222), .ZN(n20224) );
  OAI21_X1 U23147 ( .B1(n20238), .B2(n20225), .A(n20224), .ZN(P1_U2998) );
  INV_X1 U23148 ( .A(n20226), .ZN(n20231) );
  OR2_X1 U23149 ( .A1(n20228), .A2(n20227), .ZN(n20229) );
  AOI22_X1 U23150 ( .A1(n20231), .A2(n20230), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20229), .ZN(n20234) );
  NAND2_X1 U23151 ( .A1(n20232), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20233) );
  OAI211_X1 U23152 ( .C1(n20235), .C2(n20238), .A(n20234), .B(n20233), .ZN(
        P1_U2999) );
  NOR2_X1 U23153 ( .A1(n20236), .A2(n20996), .ZN(P1_U3032) );
  NOR2_X2 U23154 ( .A1(n20238), .A2(n20237), .ZN(n20288) );
  AOI22_X1 U23155 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20288), .B1(DATAI_16_), 
        .B2(n20240), .ZN(n20814) );
  NAND2_X1 U23156 ( .A1(n20287), .A2(n20243), .ZN(n20855) );
  NAND2_X1 U23157 ( .A1(n21136), .A2(n20562), .ZN(n20367) );
  OR2_X1 U23158 ( .A1(n20720), .A2(n20367), .ZN(n20289) );
  AOI22_X1 U23159 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20288), .B1(DATAI_24_), 
        .B2(n20240), .ZN(n20864) );
  OAI22_X1 U23160 ( .A1(n20855), .A2(n20289), .B1(n20864), .B2(n20906), .ZN(
        n20244) );
  INV_X1 U23161 ( .A(n20244), .ZN(n20256) );
  INV_X1 U23162 ( .A(n20332), .ZN(n20245) );
  OAI21_X1 U23163 ( .B1(n20245), .B2(n20914), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20246) );
  NAND2_X1 U23164 ( .A1(n20246), .A2(n20689), .ZN(n20254) );
  OR2_X1 U23165 ( .A1(n20563), .A2(n20247), .ZN(n20373) );
  NOR2_X1 U23166 ( .A1(n20373), .A2(n20804), .ZN(n20251) );
  INV_X1 U23167 ( .A(n20565), .ZN(n20248) );
  NAND2_X1 U23168 ( .A1(n20248), .A2(n20642), .ZN(n20407) );
  AOI22_X1 U23169 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20407), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20289), .ZN(n20249) );
  AND2_X1 U23170 ( .A1(n20252), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20796) );
  OAI211_X1 U23171 ( .C1(n20254), .C2(n20251), .A(n20249), .B(n20643), .ZN(
        n20293) );
  INV_X1 U23172 ( .A(n20251), .ZN(n20253) );
  OR2_X1 U23173 ( .A1(n20252), .A2(n21011), .ZN(n20647) );
  OAI22_X1 U23174 ( .A1(n20254), .A2(n20253), .B1(n20647), .B2(n20407), .ZN(
        n20292) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20293), .B1(
        n20800), .B2(n20292), .ZN(n20255) );
  OAI211_X1 U23176 ( .C1(n20814), .C2(n20332), .A(n20256), .B(n20255), .ZN(
        P1_U3033) );
  AOI22_X1 U23177 ( .A1(DATAI_17_), .A2(n20240), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20288), .ZN(n20818) );
  NOR2_X2 U23178 ( .A1(n20281), .A2(n20257), .ZN(n20866) );
  INV_X1 U23179 ( .A(n20289), .ZN(n20282) );
  AOI22_X1 U23180 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20288), .B1(DATAI_25_), 
        .B2(n20240), .ZN(n20870) );
  INV_X1 U23181 ( .A(n20870), .ZN(n20815) );
  AOI22_X1 U23182 ( .A1(n20866), .A2(n20282), .B1(n20914), .B2(n20815), .ZN(
        n20260) );
  NOR2_X2 U23183 ( .A1(n20258), .A2(n20412), .ZN(n20865) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20293), .B1(
        n20865), .B2(n20292), .ZN(n20259) );
  OAI211_X1 U23185 ( .C1(n20818), .C2(n20332), .A(n20260), .B(n20259), .ZN(
        P1_U3034) );
  AOI22_X1 U23186 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20288), .B1(DATAI_18_), 
        .B2(n20240), .ZN(n20877) );
  NAND2_X1 U23187 ( .A1(n20287), .A2(n20261), .ZN(n20872) );
  OAI22_X1 U23188 ( .A1(n20872), .A2(n20289), .B1(n20739), .B2(n20906), .ZN(
        n20262) );
  INV_X1 U23189 ( .A(n20262), .ZN(n20265) );
  AOI22_X1 U23190 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20293), .B1(
        n20819), .B2(n20292), .ZN(n20264) );
  OAI211_X1 U23191 ( .C1(n20877), .C2(n20332), .A(n20265), .B(n20264), .ZN(
        P1_U3035) );
  AOI22_X1 U23192 ( .A1(DATAI_19_), .A2(n20240), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20288), .ZN(n20826) );
  NOR2_X2 U23193 ( .A1(n20281), .A2(n20266), .ZN(n20879) );
  INV_X1 U23194 ( .A(n20883), .ZN(n20823) );
  AOI22_X1 U23195 ( .A1(n20879), .A2(n20282), .B1(n20914), .B2(n20823), .ZN(
        n20269) );
  NOR2_X2 U23196 ( .A1(n20267), .A2(n20412), .ZN(n20878) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20293), .B1(
        n20878), .B2(n20292), .ZN(n20268) );
  OAI211_X1 U23198 ( .C1(n20826), .C2(n20332), .A(n20269), .B(n20268), .ZN(
        P1_U3036) );
  AOI22_X1 U23199 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20288), .B1(DATAI_20_), 
        .B2(n20240), .ZN(n20832) );
  NAND2_X1 U23200 ( .A1(n20287), .A2(n20270), .ZN(n20885) );
  OAI22_X1 U23201 ( .A1(n20885), .A2(n20289), .B1(n20890), .B2(n20906), .ZN(
        n20271) );
  INV_X1 U23202 ( .A(n20271), .ZN(n20274) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20293), .B1(
        n20827), .B2(n20292), .ZN(n20273) );
  OAI211_X1 U23204 ( .C1(n20832), .C2(n20332), .A(n20274), .B(n20273), .ZN(
        P1_U3037) );
  NAND2_X1 U23205 ( .A1(n20287), .A2(n20275), .ZN(n20892) );
  AOI22_X1 U23206 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20288), .B1(DATAI_29_), 
        .B2(n20240), .ZN(n20747) );
  OAI22_X1 U23207 ( .A1(n20892), .A2(n20289), .B1(n20747), .B2(n20906), .ZN(
        n20276) );
  INV_X1 U23208 ( .A(n20276), .ZN(n20279) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20293), .B1(
        n20833), .B2(n20292), .ZN(n20278) );
  OAI211_X1 U23210 ( .C1(n20897), .C2(n20332), .A(n20279), .B(n20278), .ZN(
        P1_U3038) );
  AOI22_X1 U23211 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20288), .B1(DATAI_22_), 
        .B2(n20240), .ZN(n20907) );
  NOR2_X2 U23212 ( .A1(n20281), .A2(n20280), .ZN(n20901) );
  AOI22_X1 U23213 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20288), .B1(DATAI_30_), 
        .B2(n20240), .ZN(n20751) );
  INV_X1 U23214 ( .A(n20751), .ZN(n20902) );
  AOI22_X1 U23215 ( .A1(n20901), .A2(n20282), .B1(n20914), .B2(n20902), .ZN(
        n20285) );
  NOR2_X2 U23216 ( .A1(n20283), .A2(n20412), .ZN(n20899) );
  AOI22_X1 U23217 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20293), .B1(
        n20899), .B2(n20292), .ZN(n20284) );
  OAI211_X1 U23218 ( .C1(n20907), .C2(n20332), .A(n20285), .B(n20284), .ZN(
        P1_U3039) );
  AOI22_X1 U23219 ( .A1(DATAI_23_), .A2(n20240), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20288), .ZN(n20848) );
  NAND2_X1 U23220 ( .A1(n20287), .A2(n20286), .ZN(n20911) );
  OAI22_X1 U23221 ( .A1(n20911), .A2(n20289), .B1(n20919), .B2(n20906), .ZN(
        n20290) );
  INV_X1 U23222 ( .A(n20290), .ZN(n20295) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20293), .B1(
        n20840), .B2(n20292), .ZN(n20294) );
  OAI211_X1 U23224 ( .C1(n20848), .C2(n20332), .A(n20295), .B(n20294), .ZN(
        P1_U3040) );
  NOR2_X1 U23225 ( .A1(n20367), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20305) );
  INV_X1 U23226 ( .A(n20305), .ZN(n20296) );
  NOR2_X1 U23227 ( .A1(n20759), .A2(n20296), .ZN(n20323) );
  INV_X1 U23228 ( .A(n20323), .ZN(n20327) );
  OR2_X1 U23229 ( .A1(n20373), .A2(n20297), .ZN(n20298) );
  NAND2_X1 U23230 ( .A1(n20298), .A2(n20327), .ZN(n20302) );
  NAND2_X1 U23231 ( .A1(n20302), .A2(n20689), .ZN(n20300) );
  NAND2_X1 U23232 ( .A1(n20305), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20299) );
  OAI22_X1 U23233 ( .A1(n20855), .A2(n20327), .B1(n20326), .B2(n20854), .ZN(
        n20301) );
  INV_X1 U23234 ( .A(n20301), .ZN(n20308) );
  INV_X1 U23235 ( .A(n20302), .ZN(n20303) );
  OAI211_X1 U23236 ( .C1(n20370), .C2(n21012), .A(n20689), .B(n20303), .ZN(
        n20304) );
  OAI211_X1 U23237 ( .C1(n20689), .C2(n20305), .A(n20859), .B(n20304), .ZN(
        n20329) );
  INV_X1 U23238 ( .A(n20814), .ZN(n20861) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20329), .B1(
        n20335), .B2(n20861), .ZN(n20307) );
  OAI211_X1 U23240 ( .C1(n20864), .C2(n20332), .A(n20308), .B(n20307), .ZN(
        P1_U3041) );
  INV_X1 U23241 ( .A(n20326), .ZN(n20322) );
  AOI22_X1 U23242 ( .A1(n20866), .A2(n20323), .B1(n20865), .B2(n20322), .ZN(
        n20310) );
  INV_X1 U23243 ( .A(n20818), .ZN(n20867) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20329), .B1(
        n20335), .B2(n20867), .ZN(n20309) );
  OAI211_X1 U23245 ( .C1(n20870), .C2(n20332), .A(n20310), .B(n20309), .ZN(
        P1_U3042) );
  OAI22_X1 U23246 ( .A1(n20872), .A2(n20327), .B1(n20326), .B2(n20871), .ZN(
        n20311) );
  INV_X1 U23247 ( .A(n20311), .ZN(n20313) );
  INV_X1 U23248 ( .A(n20877), .ZN(n20736) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20329), .B1(
        n20335), .B2(n20736), .ZN(n20312) );
  OAI211_X1 U23250 ( .C1(n20739), .C2(n20332), .A(n20313), .B(n20312), .ZN(
        P1_U3043) );
  AOI22_X1 U23251 ( .A1(n20879), .A2(n20323), .B1(n20878), .B2(n20322), .ZN(
        n20315) );
  INV_X1 U23252 ( .A(n20826), .ZN(n20880) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20329), .B1(
        n20335), .B2(n20880), .ZN(n20314) );
  OAI211_X1 U23254 ( .C1(n20883), .C2(n20332), .A(n20315), .B(n20314), .ZN(
        P1_U3044) );
  OAI22_X1 U23255 ( .A1(n20885), .A2(n20327), .B1(n20326), .B2(n20884), .ZN(
        n20316) );
  INV_X1 U23256 ( .A(n20316), .ZN(n20318) );
  INV_X1 U23257 ( .A(n20832), .ZN(n20887) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20329), .B1(
        n20335), .B2(n20887), .ZN(n20317) );
  OAI211_X1 U23259 ( .C1(n20890), .C2(n20332), .A(n20318), .B(n20317), .ZN(
        P1_U3045) );
  OAI22_X1 U23260 ( .A1(n20892), .A2(n20327), .B1(n20326), .B2(n20891), .ZN(
        n20319) );
  INV_X1 U23261 ( .A(n20319), .ZN(n20321) );
  INV_X1 U23262 ( .A(n20897), .ZN(n20744) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20329), .B1(
        n20335), .B2(n20744), .ZN(n20320) );
  OAI211_X1 U23264 ( .C1(n20747), .C2(n20332), .A(n20321), .B(n20320), .ZN(
        P1_U3046) );
  AOI22_X1 U23265 ( .A1(n20901), .A2(n20323), .B1(n20899), .B2(n20322), .ZN(
        n20325) );
  INV_X1 U23266 ( .A(n20907), .ZN(n20748) );
  AOI22_X1 U23267 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20329), .B1(
        n20335), .B2(n20748), .ZN(n20324) );
  OAI211_X1 U23268 ( .C1(n20751), .C2(n20332), .A(n20325), .B(n20324), .ZN(
        P1_U3047) );
  OAI22_X1 U23269 ( .A1(n20911), .A2(n20327), .B1(n20326), .B2(n20908), .ZN(
        n20328) );
  INV_X1 U23270 ( .A(n20328), .ZN(n20331) );
  INV_X1 U23271 ( .A(n20848), .ZN(n20913) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20329), .B1(
        n20335), .B2(n20913), .ZN(n20330) );
  OAI211_X1 U23273 ( .C1(n20919), .C2(n20332), .A(n20331), .B(n20330), .ZN(
        P1_U3048) );
  NAND2_X1 U23274 ( .A1(n13889), .A2(n12423), .ZN(n20638) );
  INV_X1 U23275 ( .A(n20367), .ZN(n20333) );
  NAND2_X1 U23276 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20333), .ZN(
        n20377) );
  NOR2_X1 U23277 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20377), .ZN(
        n20357) );
  INV_X1 U23278 ( .A(n20357), .ZN(n20360) );
  OAI22_X1 U23279 ( .A1(n20366), .A2(n20864), .B1(n20855), .B2(n20360), .ZN(
        n20334) );
  INV_X1 U23280 ( .A(n20334), .ZN(n20343) );
  OAI21_X1 U23281 ( .B1(n20335), .B2(n20387), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20336) );
  NAND2_X1 U23282 ( .A1(n20336), .A2(n20689), .ZN(n20341) );
  NOR2_X1 U23283 ( .A1(n20373), .A2(n14101), .ZN(n20339) );
  OR2_X1 U23284 ( .A1(n20642), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20488) );
  NAND2_X1 U23285 ( .A1(n20488), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20484) );
  OAI211_X1 U23286 ( .C1(n20726), .C2(n20357), .A(n20484), .B(n20643), .ZN(
        n20337) );
  INV_X1 U23287 ( .A(n20337), .ZN(n20338) );
  INV_X1 U23288 ( .A(n20339), .ZN(n20340) );
  OAI22_X1 U23289 ( .A1(n20341), .A2(n20340), .B1(n20647), .B2(n20488), .ZN(
        n20362) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20363), .B1(
        n20800), .B2(n20362), .ZN(n20342) );
  OAI211_X1 U23291 ( .C1(n20814), .C2(n20399), .A(n20343), .B(n20342), .ZN(
        P1_U3049) );
  AOI22_X1 U23292 ( .A1(n20387), .A2(n20867), .B1(n20866), .B2(n20357), .ZN(
        n20345) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20363), .B1(
        n20865), .B2(n20362), .ZN(n20344) );
  OAI211_X1 U23294 ( .C1(n20870), .C2(n20366), .A(n20345), .B(n20344), .ZN(
        P1_U3050) );
  OAI22_X1 U23295 ( .A1(n20366), .A2(n20739), .B1(n20360), .B2(n20872), .ZN(
        n20346) );
  INV_X1 U23296 ( .A(n20346), .ZN(n20348) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20363), .B1(
        n20819), .B2(n20362), .ZN(n20347) );
  OAI211_X1 U23298 ( .C1(n20877), .C2(n20399), .A(n20348), .B(n20347), .ZN(
        P1_U3051) );
  AOI22_X1 U23299 ( .A1(n20387), .A2(n20880), .B1(n20879), .B2(n20357), .ZN(
        n20350) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20363), .B1(
        n20878), .B2(n20362), .ZN(n20349) );
  OAI211_X1 U23301 ( .C1(n20883), .C2(n20366), .A(n20350), .B(n20349), .ZN(
        P1_U3052) );
  OAI22_X1 U23302 ( .A1(n20885), .A2(n20360), .B1(n20399), .B2(n20832), .ZN(
        n20351) );
  INV_X1 U23303 ( .A(n20351), .ZN(n20353) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20363), .B1(
        n20827), .B2(n20362), .ZN(n20352) );
  OAI211_X1 U23305 ( .C1(n20890), .C2(n20366), .A(n20353), .B(n20352), .ZN(
        P1_U3053) );
  OAI22_X1 U23306 ( .A1(n20892), .A2(n20360), .B1(n20399), .B2(n20897), .ZN(
        n20354) );
  INV_X1 U23307 ( .A(n20354), .ZN(n20356) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20363), .B1(
        n20833), .B2(n20362), .ZN(n20355) );
  OAI211_X1 U23309 ( .C1(n20747), .C2(n20366), .A(n20356), .B(n20355), .ZN(
        P1_U3054) );
  AOI22_X1 U23310 ( .A1(n20387), .A2(n20748), .B1(n20901), .B2(n20357), .ZN(
        n20359) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20363), .B1(
        n20899), .B2(n20362), .ZN(n20358) );
  OAI211_X1 U23312 ( .C1(n20751), .C2(n20366), .A(n20359), .B(n20358), .ZN(
        P1_U3055) );
  OAI22_X1 U23313 ( .A1(n20911), .A2(n20360), .B1(n20399), .B2(n20848), .ZN(
        n20361) );
  INV_X1 U23314 ( .A(n20361), .ZN(n20365) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20363), .B1(
        n20840), .B2(n20362), .ZN(n20364) );
  OAI211_X1 U23316 ( .C1(n20919), .C2(n20366), .A(n20365), .B(n20364), .ZN(
        P1_U3056) );
  INV_X1 U23317 ( .A(n20690), .ZN(n20531) );
  NOR2_X1 U23318 ( .A1(n20368), .A2(n20367), .ZN(n20396) );
  INV_X1 U23319 ( .A(n20396), .ZN(n20400) );
  OAI22_X1 U23320 ( .A1(n20855), .A2(n20400), .B1(n20399), .B2(n20864), .ZN(
        n20369) );
  INV_X1 U23321 ( .A(n20369), .ZN(n20381) );
  AOI21_X1 U23322 ( .B1(n20370), .B2(n20689), .A(n20685), .ZN(n20379) );
  NAND2_X1 U23323 ( .A1(n20372), .A2(n20371), .ZN(n20849) );
  OR2_X1 U23324 ( .A1(n20373), .A2(n20849), .ZN(n20374) );
  AND2_X1 U23325 ( .A1(n20374), .A2(n20400), .ZN(n20378) );
  INV_X1 U23326 ( .A(n20378), .ZN(n20376) );
  INV_X1 U23327 ( .A(n20859), .ZN(n20764) );
  AOI21_X1 U23328 ( .B1(n20760), .B2(n20377), .A(n20764), .ZN(n20375) );
  OAI21_X1 U23329 ( .B1(n20379), .B2(n20376), .A(n20375), .ZN(n20403) );
  OAI22_X1 U23330 ( .A1(n20379), .A2(n20378), .B1(n21011), .B2(n20377), .ZN(
        n20402) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20403), .B1(
        n20800), .B2(n20402), .ZN(n20380) );
  OAI211_X1 U23332 ( .C1(n20814), .C2(n20440), .A(n20381), .B(n20380), .ZN(
        P1_U3057) );
  AOI22_X1 U23333 ( .A1(n20387), .A2(n20815), .B1(n20866), .B2(n20396), .ZN(
        n20383) );
  AOI22_X1 U23334 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20403), .B1(
        n20865), .B2(n20402), .ZN(n20382) );
  OAI211_X1 U23335 ( .C1(n20818), .C2(n20440), .A(n20383), .B(n20382), .ZN(
        P1_U3058) );
  OAI22_X1 U23336 ( .A1(n20872), .A2(n20400), .B1(n20440), .B2(n20877), .ZN(
        n20384) );
  INV_X1 U23337 ( .A(n20384), .ZN(n20386) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20403), .B1(
        n20819), .B2(n20402), .ZN(n20385) );
  OAI211_X1 U23339 ( .C1(n20739), .C2(n20399), .A(n20386), .B(n20385), .ZN(
        P1_U3059) );
  AOI22_X1 U23340 ( .A1(n20387), .A2(n20823), .B1(n20879), .B2(n20396), .ZN(
        n20389) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20403), .B1(
        n20878), .B2(n20402), .ZN(n20388) );
  OAI211_X1 U23342 ( .C1(n20826), .C2(n20440), .A(n20389), .B(n20388), .ZN(
        P1_U3060) );
  OAI22_X1 U23343 ( .A1(n20885), .A2(n20400), .B1(n20440), .B2(n20832), .ZN(
        n20390) );
  INV_X1 U23344 ( .A(n20390), .ZN(n20392) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20403), .B1(
        n20827), .B2(n20402), .ZN(n20391) );
  OAI211_X1 U23346 ( .C1(n20890), .C2(n20399), .A(n20392), .B(n20391), .ZN(
        P1_U3061) );
  OAI22_X1 U23347 ( .A1(n20892), .A2(n20400), .B1(n20399), .B2(n20747), .ZN(
        n20393) );
  INV_X1 U23348 ( .A(n20393), .ZN(n20395) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20403), .B1(
        n20833), .B2(n20402), .ZN(n20394) );
  OAI211_X1 U23350 ( .C1(n20897), .C2(n20440), .A(n20395), .B(n20394), .ZN(
        P1_U3062) );
  AOI22_X1 U23351 ( .A1(n20419), .A2(n20748), .B1(n20901), .B2(n20396), .ZN(
        n20398) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20403), .B1(
        n20899), .B2(n20402), .ZN(n20397) );
  OAI211_X1 U23353 ( .C1(n20751), .C2(n20399), .A(n20398), .B(n20397), .ZN(
        P1_U3063) );
  OAI22_X1 U23354 ( .A1(n20911), .A2(n20400), .B1(n20399), .B2(n20919), .ZN(
        n20401) );
  INV_X1 U23355 ( .A(n20401), .ZN(n20405) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20403), .B1(
        n20840), .B2(n20402), .ZN(n20404) );
  OAI211_X1 U23357 ( .C1(n20848), .C2(n20440), .A(n20405), .B(n20404), .ZN(
        P1_U3064) );
  NAND2_X1 U23358 ( .A1(n20441), .A2(n12423), .ZN(n20463) );
  OR2_X1 U23359 ( .A1(n20720), .A2(n20478), .ZN(n20435) );
  OR2_X1 U23360 ( .A1(n13861), .A2(n20406), .ZN(n20522) );
  OR3_X1 U23361 ( .A1(n20522), .A2(n20804), .A3(n20760), .ZN(n20409) );
  INV_X1 U23362 ( .A(n20796), .ZN(n20729) );
  OR2_X1 U23363 ( .A1(n20407), .A2(n20729), .ZN(n20408) );
  OAI22_X1 U23364 ( .A1(n20855), .A2(n20435), .B1(n20434), .B2(n20854), .ZN(
        n20410) );
  INV_X1 U23365 ( .A(n20410), .ZN(n20415) );
  INV_X1 U23366 ( .A(n20435), .ZN(n20431) );
  OAI21_X1 U23367 ( .B1(n20474), .B2(n20419), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20411) );
  OAI21_X1 U23368 ( .B1(n20804), .B2(n20522), .A(n20411), .ZN(n20413) );
  INV_X1 U23369 ( .A(n20647), .ZN(n20566) );
  OAI221_X1 U23370 ( .B1(n20431), .B2(n20726), .C1(n20431), .C2(n20413), .A(
        n20808), .ZN(n20437) );
  INV_X1 U23371 ( .A(n20864), .ZN(n20811) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20437), .B1(
        n20419), .B2(n20811), .ZN(n20414) );
  OAI211_X1 U23373 ( .C1(n20814), .C2(n20463), .A(n20415), .B(n20414), .ZN(
        P1_U3065) );
  INV_X1 U23374 ( .A(n20434), .ZN(n20430) );
  AOI22_X1 U23375 ( .A1(n20866), .A2(n20431), .B1(n20865), .B2(n20430), .ZN(
        n20417) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20437), .B1(
        n20474), .B2(n20867), .ZN(n20416) );
  OAI211_X1 U23377 ( .C1(n20870), .C2(n20440), .A(n20417), .B(n20416), .ZN(
        P1_U3066) );
  OAI22_X1 U23378 ( .A1(n20872), .A2(n20435), .B1(n20434), .B2(n20871), .ZN(
        n20418) );
  INV_X1 U23379 ( .A(n20418), .ZN(n20421) );
  INV_X1 U23380 ( .A(n20739), .ZN(n20874) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20437), .B1(
        n20419), .B2(n20874), .ZN(n20420) );
  OAI211_X1 U23382 ( .C1(n20877), .C2(n20463), .A(n20421), .B(n20420), .ZN(
        P1_U3067) );
  AOI22_X1 U23383 ( .A1(n20879), .A2(n20431), .B1(n20878), .B2(n20430), .ZN(
        n20423) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20437), .B1(
        n20474), .B2(n20880), .ZN(n20422) );
  OAI211_X1 U23385 ( .C1(n20883), .C2(n20440), .A(n20423), .B(n20422), .ZN(
        P1_U3068) );
  OAI22_X1 U23386 ( .A1(n20885), .A2(n20435), .B1(n20434), .B2(n20884), .ZN(
        n20424) );
  INV_X1 U23387 ( .A(n20424), .ZN(n20426) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20437), .B1(
        n20474), .B2(n20887), .ZN(n20425) );
  OAI211_X1 U23389 ( .C1(n20890), .C2(n20440), .A(n20426), .B(n20425), .ZN(
        P1_U3069) );
  OAI22_X1 U23390 ( .A1(n20892), .A2(n20435), .B1(n20434), .B2(n20891), .ZN(
        n20427) );
  INV_X1 U23391 ( .A(n20427), .ZN(n20429) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20437), .B1(
        n20474), .B2(n20744), .ZN(n20428) );
  OAI211_X1 U23393 ( .C1(n20747), .C2(n20440), .A(n20429), .B(n20428), .ZN(
        P1_U3070) );
  AOI22_X1 U23394 ( .A1(n20901), .A2(n20431), .B1(n20899), .B2(n20430), .ZN(
        n20433) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20437), .B1(
        n20474), .B2(n20748), .ZN(n20432) );
  OAI211_X1 U23396 ( .C1(n20751), .C2(n20440), .A(n20433), .B(n20432), .ZN(
        P1_U3071) );
  OAI22_X1 U23397 ( .A1(n20911), .A2(n20435), .B1(n20434), .B2(n20908), .ZN(
        n20436) );
  INV_X1 U23398 ( .A(n20436), .ZN(n20439) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20437), .B1(
        n20474), .B2(n20913), .ZN(n20438) );
  OAI211_X1 U23400 ( .C1(n20919), .C2(n20440), .A(n20439), .B(n20438), .ZN(
        P1_U3072) );
  NOR2_X1 U23401 ( .A1(n20478), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20450) );
  INV_X1 U23402 ( .A(n20450), .ZN(n20442) );
  NOR2_X1 U23403 ( .A1(n20759), .A2(n20442), .ZN(n20468) );
  INV_X1 U23404 ( .A(n20468), .ZN(n20472) );
  OR2_X1 U23405 ( .A1(n20522), .A2(n20297), .ZN(n20443) );
  NAND2_X1 U23406 ( .A1(n20443), .A2(n20472), .ZN(n20447) );
  NAND2_X1 U23407 ( .A1(n20447), .A2(n20689), .ZN(n20445) );
  NAND2_X1 U23408 ( .A1(n20450), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20444) );
  AND2_X1 U23409 ( .A1(n20445), .A2(n20444), .ZN(n20471) );
  OAI22_X1 U23410 ( .A1(n20855), .A2(n20472), .B1(n20471), .B2(n20854), .ZN(
        n20446) );
  INV_X1 U23411 ( .A(n20446), .ZN(n20452) );
  INV_X1 U23412 ( .A(n20447), .ZN(n20448) );
  OAI211_X1 U23413 ( .C1(n20532), .C2(n21012), .A(n20689), .B(n20448), .ZN(
        n20449) );
  OAI211_X1 U23414 ( .C1(n20689), .C2(n20450), .A(n20859), .B(n20449), .ZN(
        n20475) );
  AOI22_X1 U23415 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20475), .B1(
        n20474), .B2(n20811), .ZN(n20451) );
  OAI211_X1 U23416 ( .C1(n20814), .C2(n20513), .A(n20452), .B(n20451), .ZN(
        P1_U3073) );
  INV_X1 U23417 ( .A(n20471), .ZN(n20467) );
  AOI22_X1 U23418 ( .A1(n20866), .A2(n20468), .B1(n20865), .B2(n20467), .ZN(
        n20454) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20475), .B1(
        n20474), .B2(n20815), .ZN(n20453) );
  OAI211_X1 U23420 ( .C1(n20818), .C2(n20513), .A(n20454), .B(n20453), .ZN(
        P1_U3074) );
  OAI22_X1 U23421 ( .A1(n20872), .A2(n20472), .B1(n20471), .B2(n20871), .ZN(
        n20455) );
  INV_X1 U23422 ( .A(n20455), .ZN(n20457) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20475), .B1(
        n20510), .B2(n20736), .ZN(n20456) );
  OAI211_X1 U23424 ( .C1(n20739), .C2(n20463), .A(n20457), .B(n20456), .ZN(
        P1_U3075) );
  AOI22_X1 U23425 ( .A1(n20879), .A2(n20468), .B1(n20878), .B2(n20467), .ZN(
        n20459) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20475), .B1(
        n20510), .B2(n20880), .ZN(n20458) );
  OAI211_X1 U23427 ( .C1(n20883), .C2(n20463), .A(n20459), .B(n20458), .ZN(
        P1_U3076) );
  OAI22_X1 U23428 ( .A1(n20885), .A2(n20472), .B1(n20471), .B2(n20884), .ZN(
        n20460) );
  INV_X1 U23429 ( .A(n20460), .ZN(n20462) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20475), .B1(
        n20510), .B2(n20887), .ZN(n20461) );
  OAI211_X1 U23431 ( .C1(n20890), .C2(n20463), .A(n20462), .B(n20461), .ZN(
        P1_U3077) );
  OAI22_X1 U23432 ( .A1(n20892), .A2(n20472), .B1(n20471), .B2(n20891), .ZN(
        n20464) );
  INV_X1 U23433 ( .A(n20464), .ZN(n20466) );
  INV_X1 U23434 ( .A(n20747), .ZN(n20894) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20475), .B1(
        n20474), .B2(n20894), .ZN(n20465) );
  OAI211_X1 U23436 ( .C1(n20897), .C2(n20513), .A(n20466), .B(n20465), .ZN(
        P1_U3078) );
  AOI22_X1 U23437 ( .A1(n20901), .A2(n20468), .B1(n20899), .B2(n20467), .ZN(
        n20470) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20475), .B1(
        n20474), .B2(n20902), .ZN(n20469) );
  OAI211_X1 U23439 ( .C1(n20907), .C2(n20513), .A(n20470), .B(n20469), .ZN(
        P1_U3079) );
  OAI22_X1 U23440 ( .A1(n20911), .A2(n20472), .B1(n20471), .B2(n20908), .ZN(
        n20473) );
  INV_X1 U23441 ( .A(n20473), .ZN(n20477) );
  INV_X1 U23442 ( .A(n20919), .ZN(n20843) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20475), .B1(
        n20474), .B2(n20843), .ZN(n20476) );
  OAI211_X1 U23444 ( .C1(n20848), .C2(n20513), .A(n20477), .B(n20476), .ZN(
        P1_U3080) );
  NOR2_X1 U23445 ( .A1(n20998), .A2(n20478), .ZN(n20527) );
  INV_X1 U23446 ( .A(n20527), .ZN(n20479) );
  NOR2_X1 U23447 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20479), .ZN(
        n20509) );
  INV_X1 U23448 ( .A(n20509), .ZN(n20515) );
  OR2_X1 U23449 ( .A1(n20561), .A2(n20814), .ZN(n20481) );
  OAI21_X1 U23450 ( .B1(n20855), .B2(n20515), .A(n20481), .ZN(n20482) );
  INV_X1 U23451 ( .A(n20482), .ZN(n20492) );
  OAI21_X1 U23452 ( .B1(n20551), .B2(n20510), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20483) );
  NAND2_X1 U23453 ( .A1(n20483), .A2(n20689), .ZN(n20490) );
  INV_X1 U23454 ( .A(n20490), .ZN(n20486) );
  OR2_X1 U23455 ( .A1(n20522), .A2(n14101), .ZN(n20489) );
  INV_X1 U23456 ( .A(n20484), .ZN(n20485) );
  AOI21_X1 U23457 ( .B1(n20486), .B2(n20489), .A(n20485), .ZN(n20487) );
  OAI211_X1 U23458 ( .C1(n20509), .C2(n20726), .A(n20808), .B(n20487), .ZN(
        n20518) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20518), .B1(
        n20800), .B2(n20517), .ZN(n20491) );
  OAI211_X1 U23460 ( .C1(n20864), .C2(n20513), .A(n20492), .B(n20491), .ZN(
        P1_U3081) );
  AOI22_X1 U23461 ( .A1(n20510), .A2(n20815), .B1(n20866), .B2(n20509), .ZN(
        n20494) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20518), .B1(
        n20865), .B2(n20517), .ZN(n20493) );
  OAI211_X1 U23463 ( .C1(n20818), .C2(n20561), .A(n20494), .B(n20493), .ZN(
        P1_U3082) );
  OR2_X1 U23464 ( .A1(n20513), .A2(n20739), .ZN(n20495) );
  OAI21_X1 U23465 ( .B1(n20872), .B2(n20515), .A(n20495), .ZN(n20496) );
  INV_X1 U23466 ( .A(n20496), .ZN(n20498) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20518), .B1(
        n20819), .B2(n20517), .ZN(n20497) );
  OAI211_X1 U23468 ( .C1(n20877), .C2(n20561), .A(n20498), .B(n20497), .ZN(
        P1_U3083) );
  AOI22_X1 U23469 ( .A1(n20551), .A2(n20880), .B1(n20879), .B2(n20509), .ZN(
        n20500) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20518), .B1(
        n20878), .B2(n20517), .ZN(n20499) );
  OAI211_X1 U23471 ( .C1(n20883), .C2(n20513), .A(n20500), .B(n20499), .ZN(
        P1_U3084) );
  OR2_X1 U23472 ( .A1(n20513), .A2(n20890), .ZN(n20501) );
  OAI21_X1 U23473 ( .B1(n20885), .B2(n20515), .A(n20501), .ZN(n20502) );
  INV_X1 U23474 ( .A(n20502), .ZN(n20504) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20518), .B1(
        n20827), .B2(n20517), .ZN(n20503) );
  OAI211_X1 U23476 ( .C1(n20832), .C2(n20561), .A(n20504), .B(n20503), .ZN(
        P1_U3085) );
  OR2_X1 U23477 ( .A1(n20561), .A2(n20897), .ZN(n20505) );
  OAI21_X1 U23478 ( .B1(n20892), .B2(n20515), .A(n20505), .ZN(n20506) );
  INV_X1 U23479 ( .A(n20506), .ZN(n20508) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20518), .B1(
        n20833), .B2(n20517), .ZN(n20507) );
  OAI211_X1 U23481 ( .C1(n20747), .C2(n20513), .A(n20508), .B(n20507), .ZN(
        P1_U3086) );
  AOI22_X1 U23482 ( .A1(n20510), .A2(n20902), .B1(n20901), .B2(n20509), .ZN(
        n20512) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20518), .B1(
        n20899), .B2(n20517), .ZN(n20511) );
  OAI211_X1 U23484 ( .C1(n20907), .C2(n20561), .A(n20512), .B(n20511), .ZN(
        P1_U3087) );
  OR2_X1 U23485 ( .A1(n20513), .A2(n20919), .ZN(n20514) );
  OAI21_X1 U23486 ( .B1(n20911), .B2(n20515), .A(n20514), .ZN(n20516) );
  INV_X1 U23487 ( .A(n20516), .ZN(n20520) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20518), .B1(
        n20840), .B2(n20517), .ZN(n20519) );
  OAI211_X1 U23489 ( .C1(n20848), .C2(n20561), .A(n20520), .B(n20519), .ZN(
        P1_U3088) );
  INV_X1 U23490 ( .A(n20532), .ZN(n20521) );
  NOR2_X1 U23491 ( .A1(n20521), .A2(n20760), .ZN(n20524) );
  OR2_X1 U23492 ( .A1(n20522), .A2(n20849), .ZN(n20523) );
  AND2_X1 U23493 ( .A1(n20523), .A2(n20556), .ZN(n20526) );
  OAI21_X1 U23494 ( .B1(n20685), .B2(n20524), .A(n20526), .ZN(n20525) );
  OAI211_X1 U23495 ( .C1(n20689), .C2(n20527), .A(n20525), .B(n20859), .ZN(
        n20558) );
  INV_X1 U23496 ( .A(n20558), .ZN(n20535) );
  INV_X1 U23497 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n21253) );
  OR2_X1 U23498 ( .A1(n20526), .A2(n20760), .ZN(n20529) );
  NAND2_X1 U23499 ( .A1(n20527), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20528) );
  NAND2_X1 U23500 ( .A1(n20529), .A2(n20528), .ZN(n20549) );
  INV_X1 U23501 ( .A(n20549), .ZN(n20555) );
  OAI22_X1 U23502 ( .A1(n20855), .A2(n20556), .B1(n20555), .B2(n20854), .ZN(
        n20530) );
  INV_X1 U23503 ( .A(n20530), .ZN(n20534) );
  AOI22_X1 U23504 ( .A1(n20551), .A2(n20811), .B1(n20597), .B2(n20861), .ZN(
        n20533) );
  OAI211_X1 U23505 ( .C1(n20535), .C2(n21253), .A(n20534), .B(n20533), .ZN(
        P1_U3089) );
  INV_X1 U23506 ( .A(n20556), .ZN(n20550) );
  AOI22_X1 U23507 ( .A1(n20866), .A2(n20550), .B1(n20865), .B2(n20549), .ZN(
        n20537) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20558), .B1(
        n20551), .B2(n20815), .ZN(n20536) );
  OAI211_X1 U23509 ( .C1(n20818), .C2(n20554), .A(n20537), .B(n20536), .ZN(
        P1_U3090) );
  OAI22_X1 U23510 ( .A1(n20872), .A2(n20556), .B1(n20555), .B2(n20871), .ZN(
        n20538) );
  INV_X1 U23511 ( .A(n20538), .ZN(n20540) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20558), .B1(
        n20597), .B2(n20736), .ZN(n20539) );
  OAI211_X1 U23513 ( .C1(n20739), .C2(n20561), .A(n20540), .B(n20539), .ZN(
        P1_U3091) );
  AOI22_X1 U23514 ( .A1(n20879), .A2(n20550), .B1(n20878), .B2(n20549), .ZN(
        n20542) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20558), .B1(
        n20597), .B2(n20880), .ZN(n20541) );
  OAI211_X1 U23516 ( .C1(n20883), .C2(n20561), .A(n20542), .B(n20541), .ZN(
        P1_U3092) );
  OAI22_X1 U23517 ( .A1(n20885), .A2(n20556), .B1(n20555), .B2(n20884), .ZN(
        n20543) );
  INV_X1 U23518 ( .A(n20543), .ZN(n20545) );
  INV_X1 U23519 ( .A(n20890), .ZN(n20829) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20558), .B1(
        n20551), .B2(n20829), .ZN(n20544) );
  OAI211_X1 U23521 ( .C1(n20832), .C2(n20554), .A(n20545), .B(n20544), .ZN(
        P1_U3093) );
  OAI22_X1 U23522 ( .A1(n20892), .A2(n20556), .B1(n20555), .B2(n20891), .ZN(
        n20546) );
  INV_X1 U23523 ( .A(n20546), .ZN(n20548) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20558), .B1(
        n20597), .B2(n20744), .ZN(n20547) );
  OAI211_X1 U23525 ( .C1(n20747), .C2(n20561), .A(n20548), .B(n20547), .ZN(
        P1_U3094) );
  AOI22_X1 U23526 ( .A1(n20901), .A2(n20550), .B1(n20899), .B2(n20549), .ZN(
        n20553) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20558), .B1(
        n20551), .B2(n20902), .ZN(n20552) );
  OAI211_X1 U23528 ( .C1(n20907), .C2(n20554), .A(n20553), .B(n20552), .ZN(
        P1_U3095) );
  OAI22_X1 U23529 ( .A1(n20911), .A2(n20556), .B1(n20555), .B2(n20908), .ZN(
        n20557) );
  INV_X1 U23530 ( .A(n20557), .ZN(n20560) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20558), .B1(
        n20597), .B2(n20913), .ZN(n20559) );
  OAI211_X1 U23532 ( .C1(n20919), .C2(n20561), .A(n20560), .B(n20559), .ZN(
        P1_U3096) );
  NAND2_X1 U23533 ( .A1(n20562), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20676) );
  OR2_X1 U23534 ( .A1(n20720), .A2(n20676), .ZN(n20595) );
  NAND2_X1 U23535 ( .A1(n20563), .A2(n13861), .ZN(n20679) );
  OR2_X1 U23536 ( .A1(n20679), .A2(n20804), .ZN(n20564) );
  OR2_X1 U23537 ( .A1(n20572), .A2(n20760), .ZN(n20569) );
  NAND2_X1 U23538 ( .A1(n20565), .A2(n20642), .ZN(n20728) );
  INV_X1 U23539 ( .A(n20728), .ZN(n20567) );
  NAND2_X1 U23540 ( .A1(n20567), .A2(n20566), .ZN(n20568) );
  AND2_X1 U23541 ( .A1(n20569), .A2(n20568), .ZN(n20594) );
  OAI22_X1 U23542 ( .A1(n20855), .A2(n20595), .B1(n20594), .B2(n20854), .ZN(
        n20570) );
  INV_X1 U23543 ( .A(n20570), .ZN(n20576) );
  INV_X1 U23544 ( .A(n20595), .ZN(n20591) );
  INV_X1 U23545 ( .A(n20636), .ZN(n20571) );
  OAI21_X1 U23546 ( .B1(n20571), .B2(n20597), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20573) );
  NAND2_X1 U23547 ( .A1(n20573), .A2(n20572), .ZN(n20574) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20811), .ZN(n20575) );
  OAI211_X1 U23549 ( .C1(n20814), .C2(n20636), .A(n20576), .B(n20575), .ZN(
        P1_U3097) );
  INV_X1 U23550 ( .A(n20594), .ZN(n20590) );
  AOI22_X1 U23551 ( .A1(n20866), .A2(n20591), .B1(n20865), .B2(n20590), .ZN(
        n20578) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20815), .ZN(n20577) );
  OAI211_X1 U23553 ( .C1(n20818), .C2(n20636), .A(n20578), .B(n20577), .ZN(
        P1_U3098) );
  OAI22_X1 U23554 ( .A1(n20872), .A2(n20595), .B1(n20594), .B2(n20871), .ZN(
        n20579) );
  INV_X1 U23555 ( .A(n20579), .ZN(n20581) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20874), .ZN(n20580) );
  OAI211_X1 U23557 ( .C1(n20877), .C2(n20636), .A(n20581), .B(n20580), .ZN(
        P1_U3099) );
  AOI22_X1 U23558 ( .A1(n20879), .A2(n20591), .B1(n20878), .B2(n20590), .ZN(
        n20583) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20823), .ZN(n20582) );
  OAI211_X1 U23560 ( .C1(n20826), .C2(n20636), .A(n20583), .B(n20582), .ZN(
        P1_U3100) );
  OAI22_X1 U23561 ( .A1(n20885), .A2(n20595), .B1(n20594), .B2(n20884), .ZN(
        n20584) );
  INV_X1 U23562 ( .A(n20584), .ZN(n20586) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20829), .ZN(n20585) );
  OAI211_X1 U23564 ( .C1(n20832), .C2(n20636), .A(n20586), .B(n20585), .ZN(
        P1_U3101) );
  OAI22_X1 U23565 ( .A1(n20892), .A2(n20595), .B1(n20594), .B2(n20891), .ZN(
        n20587) );
  INV_X1 U23566 ( .A(n20587), .ZN(n20589) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20894), .ZN(n20588) );
  OAI211_X1 U23568 ( .C1(n20897), .C2(n20636), .A(n20589), .B(n20588), .ZN(
        P1_U3102) );
  AOI22_X1 U23569 ( .A1(n20901), .A2(n20591), .B1(n20899), .B2(n20590), .ZN(
        n20593) );
  AOI22_X1 U23570 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20902), .ZN(n20592) );
  OAI211_X1 U23571 ( .C1(n20907), .C2(n20636), .A(n20593), .B(n20592), .ZN(
        P1_U3103) );
  OAI22_X1 U23572 ( .A1(n20911), .A2(n20595), .B1(n20594), .B2(n20908), .ZN(
        n20596) );
  INV_X1 U23573 ( .A(n20596), .ZN(n20600) );
  AOI22_X1 U23574 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20843), .ZN(n20599) );
  OAI211_X1 U23575 ( .C1(n20848), .C2(n20636), .A(n20600), .B(n20599), .ZN(
        P1_U3104) );
  NOR2_X1 U23576 ( .A1(n20676), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20608) );
  INV_X1 U23577 ( .A(n20608), .ZN(n20602) );
  NOR2_X1 U23578 ( .A1(n20759), .A2(n20602), .ZN(n20626) );
  INV_X1 U23579 ( .A(n20626), .ZN(n20630) );
  OR2_X1 U23580 ( .A1(n20679), .A2(n20297), .ZN(n20601) );
  NAND2_X1 U23581 ( .A1(n20601), .A2(n20630), .ZN(n20605) );
  NOR2_X1 U23582 ( .A1(n20602), .A2(n21011), .ZN(n20603) );
  AOI21_X1 U23583 ( .B1(n20605), .B2(n20689), .A(n20603), .ZN(n20629) );
  OAI22_X1 U23584 ( .A1(n20855), .A2(n20630), .B1(n20629), .B2(n20854), .ZN(
        n20604) );
  INV_X1 U23585 ( .A(n20604), .ZN(n20611) );
  INV_X1 U23586 ( .A(n20605), .ZN(n20606) );
  OAI211_X1 U23587 ( .C1(n20637), .C2(n21012), .A(n20689), .B(n20606), .ZN(
        n20607) );
  OAI211_X1 U23588 ( .C1(n20689), .C2(n20608), .A(n20859), .B(n20607), .ZN(
        n20633) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20633), .B1(
        n20632), .B2(n20861), .ZN(n20610) );
  OAI211_X1 U23590 ( .C1(n20864), .C2(n20636), .A(n20611), .B(n20610), .ZN(
        P1_U3105) );
  INV_X1 U23591 ( .A(n20629), .ZN(n20625) );
  AOI22_X1 U23592 ( .A1(n20866), .A2(n20626), .B1(n20865), .B2(n20625), .ZN(
        n20613) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20633), .B1(
        n20632), .B2(n20867), .ZN(n20612) );
  OAI211_X1 U23594 ( .C1(n20870), .C2(n20636), .A(n20613), .B(n20612), .ZN(
        P1_U3106) );
  OAI22_X1 U23595 ( .A1(n20872), .A2(n20630), .B1(n20629), .B2(n20871), .ZN(
        n20614) );
  INV_X1 U23596 ( .A(n20614), .ZN(n20616) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20633), .B1(
        n20632), .B2(n20736), .ZN(n20615) );
  OAI211_X1 U23598 ( .C1(n20739), .C2(n20636), .A(n20616), .B(n20615), .ZN(
        P1_U3107) );
  AOI22_X1 U23599 ( .A1(n20879), .A2(n20626), .B1(n20878), .B2(n20625), .ZN(
        n20618) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20633), .B1(
        n20632), .B2(n20880), .ZN(n20617) );
  OAI211_X1 U23601 ( .C1(n20883), .C2(n20636), .A(n20618), .B(n20617), .ZN(
        P1_U3108) );
  OAI22_X1 U23602 ( .A1(n20885), .A2(n20630), .B1(n20629), .B2(n20884), .ZN(
        n20619) );
  INV_X1 U23603 ( .A(n20619), .ZN(n20621) );
  AOI22_X1 U23604 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20633), .B1(
        n20632), .B2(n20887), .ZN(n20620) );
  OAI211_X1 U23605 ( .C1(n20890), .C2(n20636), .A(n20621), .B(n20620), .ZN(
        P1_U3109) );
  OAI22_X1 U23606 ( .A1(n20892), .A2(n20630), .B1(n20629), .B2(n20891), .ZN(
        n20622) );
  INV_X1 U23607 ( .A(n20622), .ZN(n20624) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20633), .B1(
        n20632), .B2(n20744), .ZN(n20623) );
  OAI211_X1 U23609 ( .C1(n20747), .C2(n20636), .A(n20624), .B(n20623), .ZN(
        P1_U3110) );
  AOI22_X1 U23610 ( .A1(n20901), .A2(n20626), .B1(n20899), .B2(n20625), .ZN(
        n20628) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20633), .B1(
        n20632), .B2(n20748), .ZN(n20627) );
  OAI211_X1 U23612 ( .C1(n20751), .C2(n20636), .A(n20628), .B(n20627), .ZN(
        P1_U3111) );
  OAI22_X1 U23613 ( .A1(n20911), .A2(n20630), .B1(n20629), .B2(n20908), .ZN(
        n20631) );
  INV_X1 U23614 ( .A(n20631), .ZN(n20635) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20633), .B1(
        n20632), .B2(n20913), .ZN(n20634) );
  OAI211_X1 U23616 ( .C1(n20919), .C2(n20636), .A(n20635), .B(n20634), .ZN(
        P1_U3112) );
  INV_X1 U23617 ( .A(n20638), .ZN(n20794) );
  NOR2_X1 U23618 ( .A1(n20998), .A2(n20676), .ZN(n20688) );
  INV_X1 U23619 ( .A(n20688), .ZN(n20639) );
  NOR2_X1 U23620 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20639), .ZN(
        n20666) );
  INV_X1 U23621 ( .A(n20666), .ZN(n20669) );
  OAI22_X1 U23622 ( .A1(n20670), .A2(n20864), .B1(n20855), .B2(n20669), .ZN(
        n20640) );
  INV_X1 U23623 ( .A(n20640), .ZN(n20651) );
  AOI21_X1 U23624 ( .B1(n20670), .B2(n20702), .A(n21012), .ZN(n20641) );
  NOR2_X1 U23625 ( .A1(n20641), .A2(n20760), .ZN(n20646) );
  OR2_X1 U23626 ( .A1(n20679), .A2(n14101), .ZN(n20648) );
  OR2_X1 U23627 ( .A1(n20642), .A2(n21136), .ZN(n20795) );
  NAND2_X1 U23628 ( .A1(n20795), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20807) );
  OAI211_X1 U23629 ( .C1(n20726), .C2(n20666), .A(n20807), .B(n20643), .ZN(
        n20644) );
  AOI21_X1 U23630 ( .B1(n20646), .B2(n20648), .A(n20644), .ZN(n20645) );
  INV_X1 U23631 ( .A(n20646), .ZN(n20649) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20673), .B1(
        n20800), .B2(n20672), .ZN(n20650) );
  OAI211_X1 U23633 ( .C1(n20814), .C2(n20702), .A(n20651), .B(n20650), .ZN(
        P1_U3113) );
  AOI22_X1 U23634 ( .A1(n20716), .A2(n20867), .B1(n20666), .B2(n20866), .ZN(
        n20653) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20673), .B1(
        n20865), .B2(n20672), .ZN(n20652) );
  OAI211_X1 U23636 ( .C1(n20870), .C2(n20670), .A(n20653), .B(n20652), .ZN(
        P1_U3114) );
  OR2_X1 U23637 ( .A1(n20872), .A2(n20669), .ZN(n20654) );
  OAI21_X1 U23638 ( .B1(n20702), .B2(n20877), .A(n20654), .ZN(n20655) );
  INV_X1 U23639 ( .A(n20655), .ZN(n20657) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20673), .B1(
        n20819), .B2(n20672), .ZN(n20656) );
  OAI211_X1 U23641 ( .C1(n20739), .C2(n20670), .A(n20657), .B(n20656), .ZN(
        P1_U3115) );
  AOI22_X1 U23642 ( .A1(n20716), .A2(n20880), .B1(n20666), .B2(n20879), .ZN(
        n20659) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20673), .B1(
        n20878), .B2(n20672), .ZN(n20658) );
  OAI211_X1 U23644 ( .C1(n20883), .C2(n20670), .A(n20659), .B(n20658), .ZN(
        P1_U3116) );
  OAI22_X1 U23645 ( .A1(n20670), .A2(n20890), .B1(n20669), .B2(n20885), .ZN(
        n20660) );
  INV_X1 U23646 ( .A(n20660), .ZN(n20662) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20673), .B1(
        n20827), .B2(n20672), .ZN(n20661) );
  OAI211_X1 U23648 ( .C1(n20832), .C2(n20702), .A(n20662), .B(n20661), .ZN(
        P1_U3117) );
  OAI22_X1 U23649 ( .A1(n20670), .A2(n20747), .B1(n20669), .B2(n20892), .ZN(
        n20663) );
  INV_X1 U23650 ( .A(n20663), .ZN(n20665) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20673), .B1(
        n20833), .B2(n20672), .ZN(n20664) );
  OAI211_X1 U23652 ( .C1(n20897), .C2(n20702), .A(n20665), .B(n20664), .ZN(
        P1_U3118) );
  AOI22_X1 U23653 ( .A1(n20716), .A2(n20748), .B1(n20666), .B2(n20901), .ZN(
        n20668) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20673), .B1(
        n20899), .B2(n20672), .ZN(n20667) );
  OAI211_X1 U23655 ( .C1(n20751), .C2(n20670), .A(n20668), .B(n20667), .ZN(
        P1_U3119) );
  OAI22_X1 U23656 ( .A1(n20670), .A2(n20919), .B1(n20669), .B2(n20911), .ZN(
        n20671) );
  INV_X1 U23657 ( .A(n20671), .ZN(n20675) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20673), .B1(
        n20840), .B2(n20672), .ZN(n20674) );
  OAI211_X1 U23659 ( .C1(n20848), .C2(n20702), .A(n20675), .B(n20674), .ZN(
        P1_U3120) );
  INV_X1 U23660 ( .A(n20676), .ZN(n20677) );
  NAND2_X1 U23661 ( .A1(n20678), .A2(n20677), .ZN(n20714) );
  OR2_X1 U23662 ( .A1(n20679), .A2(n20849), .ZN(n20680) );
  OR2_X1 U23663 ( .A1(n20684), .A2(n20760), .ZN(n20682) );
  NAND2_X1 U23664 ( .A1(n20688), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20681) );
  AND2_X1 U23665 ( .A1(n20682), .A2(n20681), .ZN(n20713) );
  OAI22_X1 U23666 ( .A1(n20855), .A2(n20714), .B1(n20713), .B2(n20854), .ZN(
        n20683) );
  INV_X1 U23667 ( .A(n20683), .ZN(n20693) );
  NOR2_X1 U23668 ( .A1(n20691), .A2(n20760), .ZN(n20686) );
  OAI21_X1 U23669 ( .B1(n20686), .B2(n20685), .A(n20684), .ZN(n20687) );
  OAI211_X1 U23670 ( .C1(n20689), .C2(n20688), .A(n20859), .B(n20687), .ZN(
        n20717) );
  INV_X1 U23671 ( .A(n20756), .ZN(n20699) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20717), .B1(
        n20699), .B2(n20861), .ZN(n20692) );
  OAI211_X1 U23673 ( .C1(n20864), .C2(n20702), .A(n20693), .B(n20692), .ZN(
        P1_U3121) );
  INV_X1 U23674 ( .A(n20714), .ZN(n20710) );
  INV_X1 U23675 ( .A(n20713), .ZN(n20709) );
  AOI22_X1 U23676 ( .A1(n20866), .A2(n20710), .B1(n20865), .B2(n20709), .ZN(
        n20695) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20717), .B1(
        n20699), .B2(n20867), .ZN(n20694) );
  OAI211_X1 U23678 ( .C1(n20870), .C2(n20702), .A(n20695), .B(n20694), .ZN(
        P1_U3122) );
  OAI22_X1 U23679 ( .A1(n20872), .A2(n20714), .B1(n20713), .B2(n20871), .ZN(
        n20696) );
  INV_X1 U23680 ( .A(n20696), .ZN(n20698) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20717), .B1(
        n20699), .B2(n20736), .ZN(n20697) );
  OAI211_X1 U23682 ( .C1(n20739), .C2(n20702), .A(n20698), .B(n20697), .ZN(
        P1_U3123) );
  AOI22_X1 U23683 ( .A1(n20879), .A2(n20710), .B1(n20878), .B2(n20709), .ZN(
        n20701) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20717), .B1(
        n20699), .B2(n20880), .ZN(n20700) );
  OAI211_X1 U23685 ( .C1(n20883), .C2(n20702), .A(n20701), .B(n20700), .ZN(
        P1_U3124) );
  OAI22_X1 U23686 ( .A1(n20885), .A2(n20714), .B1(n20713), .B2(n20884), .ZN(
        n20703) );
  INV_X1 U23687 ( .A(n20703), .ZN(n20705) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n20829), .ZN(n20704) );
  OAI211_X1 U23689 ( .C1(n20832), .C2(n20756), .A(n20705), .B(n20704), .ZN(
        P1_U3125) );
  OAI22_X1 U23690 ( .A1(n20892), .A2(n20714), .B1(n20713), .B2(n20891), .ZN(
        n20706) );
  INV_X1 U23691 ( .A(n20706), .ZN(n20708) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n20894), .ZN(n20707) );
  OAI211_X1 U23693 ( .C1(n20897), .C2(n20756), .A(n20708), .B(n20707), .ZN(
        P1_U3126) );
  AOI22_X1 U23694 ( .A1(n20901), .A2(n20710), .B1(n20899), .B2(n20709), .ZN(
        n20712) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n20902), .ZN(n20711) );
  OAI211_X1 U23696 ( .C1(n20907), .C2(n20756), .A(n20712), .B(n20711), .ZN(
        P1_U3127) );
  OAI22_X1 U23697 ( .A1(n20911), .A2(n20714), .B1(n20713), .B2(n20908), .ZN(
        n20715) );
  INV_X1 U23698 ( .A(n20715), .ZN(n20719) );
  AOI22_X1 U23699 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n20843), .ZN(n20718) );
  OAI211_X1 U23700 ( .C1(n20848), .C2(n20756), .A(n20719), .B(n20718), .ZN(
        P1_U3128) );
  INV_X1 U23701 ( .A(n20855), .ZN(n20801) );
  AOI22_X1 U23702 ( .A1(n20801), .A2(n10110), .B1(n20790), .B2(n20861), .ZN(
        n20733) );
  INV_X1 U23703 ( .A(n20790), .ZN(n20722) );
  AOI21_X1 U23704 ( .B1(n20722), .B2(n20756), .A(n21012), .ZN(n20723) );
  NOR2_X1 U23705 ( .A1(n20723), .A2(n20760), .ZN(n20727) );
  OR2_X1 U23706 ( .A1(n13861), .A2(n20724), .ZN(n20802) );
  OR2_X1 U23707 ( .A1(n20802), .A2(n20804), .ZN(n20730) );
  AOI22_X1 U23708 ( .A1(n20727), .A2(n20730), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20728), .ZN(n20725) );
  OAI211_X1 U23709 ( .C1(n10110), .C2(n20726), .A(n20808), .B(n20725), .ZN(
        n20753) );
  INV_X1 U23710 ( .A(n20727), .ZN(n20731) );
  AOI22_X1 U23711 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20753), .B1(
        n20800), .B2(n20752), .ZN(n20732) );
  OAI211_X1 U23712 ( .C1(n20864), .C2(n20756), .A(n20733), .B(n20732), .ZN(
        P1_U3129) );
  AOI22_X1 U23713 ( .A1(n20790), .A2(n20867), .B1(n20866), .B2(n10110), .ZN(
        n20735) );
  AOI22_X1 U23714 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20753), .B1(
        n20865), .B2(n20752), .ZN(n20734) );
  OAI211_X1 U23715 ( .C1(n20870), .C2(n20756), .A(n20735), .B(n20734), .ZN(
        P1_U3130) );
  INV_X1 U23716 ( .A(n20872), .ZN(n20820) );
  AOI22_X1 U23717 ( .A1(n20820), .A2(n10110), .B1(n20790), .B2(n20736), .ZN(
        n20738) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20753), .B1(
        n20819), .B2(n20752), .ZN(n20737) );
  OAI211_X1 U23719 ( .C1(n20739), .C2(n20756), .A(n20738), .B(n20737), .ZN(
        P1_U3131) );
  AOI22_X1 U23720 ( .A1(n20790), .A2(n20880), .B1(n20879), .B2(n10110), .ZN(
        n20741) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20753), .B1(
        n20878), .B2(n20752), .ZN(n20740) );
  OAI211_X1 U23722 ( .C1(n20883), .C2(n20756), .A(n20741), .B(n20740), .ZN(
        P1_U3132) );
  INV_X1 U23723 ( .A(n20885), .ZN(n20828) );
  AOI22_X1 U23724 ( .A1(n20828), .A2(n10110), .B1(n20790), .B2(n20887), .ZN(
        n20743) );
  AOI22_X1 U23725 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20753), .B1(
        n20827), .B2(n20752), .ZN(n20742) );
  OAI211_X1 U23726 ( .C1(n20890), .C2(n20756), .A(n20743), .B(n20742), .ZN(
        P1_U3133) );
  INV_X1 U23727 ( .A(n20892), .ZN(n20834) );
  AOI22_X1 U23728 ( .A1(n20834), .A2(n10110), .B1(n20790), .B2(n20744), .ZN(
        n20746) );
  AOI22_X1 U23729 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20753), .B1(
        n20833), .B2(n20752), .ZN(n20745) );
  OAI211_X1 U23730 ( .C1(n20747), .C2(n20756), .A(n20746), .B(n20745), .ZN(
        P1_U3134) );
  AOI22_X1 U23731 ( .A1(n20790), .A2(n20748), .B1(n20901), .B2(n10110), .ZN(
        n20750) );
  AOI22_X1 U23732 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20753), .B1(
        n20899), .B2(n20752), .ZN(n20749) );
  OAI211_X1 U23733 ( .C1(n20751), .C2(n20756), .A(n20750), .B(n20749), .ZN(
        P1_U3135) );
  INV_X1 U23734 ( .A(n20911), .ZN(n20842) );
  AOI22_X1 U23735 ( .A1(n20842), .A2(n10110), .B1(n20790), .B2(n20913), .ZN(
        n20755) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20753), .B1(
        n20840), .B2(n20752), .ZN(n20754) );
  OAI211_X1 U23737 ( .C1(n20919), .C2(n20756), .A(n20755), .B(n20754), .ZN(
        P1_U3136) );
  NOR3_X1 U23738 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20759), .A3(
        n20851), .ZN(n20784) );
  OR2_X1 U23739 ( .A1(n20802), .A2(n20760), .ZN(n20850) );
  OR2_X1 U23740 ( .A1(n20850), .A2(n20297), .ZN(n20763) );
  OR2_X1 U23741 ( .A1(n20851), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20765) );
  INV_X1 U23742 ( .A(n20765), .ZN(n20761) );
  AOI22_X1 U23743 ( .A1(n20689), .A2(n20784), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20761), .ZN(n20762) );
  NAND2_X1 U23744 ( .A1(n20763), .A2(n20762), .ZN(n20783) );
  AOI22_X1 U23745 ( .A1(n20801), .A2(n20784), .B1(n20800), .B2(n20783), .ZN(
        n20769) );
  AOI21_X1 U23746 ( .B1(n20766), .B2(n20765), .A(n20764), .ZN(n20767) );
  AOI22_X1 U23747 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20811), .ZN(n20768) );
  OAI211_X1 U23748 ( .C1(n20814), .C2(n20810), .A(n20769), .B(n20768), .ZN(
        P1_U3137) );
  AOI22_X1 U23749 ( .A1(n20866), .A2(n20784), .B1(n20865), .B2(n20783), .ZN(
        n20771) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20815), .ZN(n20770) );
  OAI211_X1 U23751 ( .C1(n20818), .C2(n20810), .A(n20771), .B(n20770), .ZN(
        P1_U3138) );
  INV_X1 U23752 ( .A(n20784), .ZN(n20788) );
  INV_X1 U23753 ( .A(n20783), .ZN(n20787) );
  OAI22_X1 U23754 ( .A1(n20872), .A2(n20788), .B1(n20787), .B2(n20871), .ZN(
        n20772) );
  INV_X1 U23755 ( .A(n20772), .ZN(n20774) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20874), .ZN(n20773) );
  OAI211_X1 U23757 ( .C1(n20877), .C2(n20810), .A(n20774), .B(n20773), .ZN(
        P1_U3139) );
  AOI22_X1 U23758 ( .A1(n20879), .A2(n20784), .B1(n20878), .B2(n20783), .ZN(
        n20776) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20823), .ZN(n20775) );
  OAI211_X1 U23760 ( .C1(n20826), .C2(n20810), .A(n20776), .B(n20775), .ZN(
        P1_U3140) );
  OAI22_X1 U23761 ( .A1(n20885), .A2(n20788), .B1(n20787), .B2(n20884), .ZN(
        n20777) );
  INV_X1 U23762 ( .A(n20777), .ZN(n20779) );
  AOI22_X1 U23763 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20829), .ZN(n20778) );
  OAI211_X1 U23764 ( .C1(n20832), .C2(n20810), .A(n20779), .B(n20778), .ZN(
        P1_U3141) );
  OAI22_X1 U23765 ( .A1(n20892), .A2(n20788), .B1(n20787), .B2(n20891), .ZN(
        n20780) );
  INV_X1 U23766 ( .A(n20780), .ZN(n20782) );
  AOI22_X1 U23767 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20894), .ZN(n20781) );
  OAI211_X1 U23768 ( .C1(n20897), .C2(n20810), .A(n20782), .B(n20781), .ZN(
        P1_U3142) );
  AOI22_X1 U23769 ( .A1(n20901), .A2(n20784), .B1(n20899), .B2(n20783), .ZN(
        n20786) );
  AOI22_X1 U23770 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20902), .ZN(n20785) );
  OAI211_X1 U23771 ( .C1(n20907), .C2(n20810), .A(n20786), .B(n20785), .ZN(
        P1_U3143) );
  OAI22_X1 U23772 ( .A1(n20911), .A2(n20788), .B1(n20787), .B2(n20908), .ZN(
        n20789) );
  INV_X1 U23773 ( .A(n20789), .ZN(n20793) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20791), .B1(
        n20790), .B2(n20843), .ZN(n20792) );
  OAI211_X1 U23775 ( .C1(n20848), .C2(n20810), .A(n20793), .B(n20792), .ZN(
        P1_U3144) );
  NOR3_X2 U23776 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20998), .A3(
        n20851), .ZN(n20841) );
  OR2_X1 U23777 ( .A1(n20850), .A2(n14101), .ZN(n20799) );
  INV_X1 U23778 ( .A(n20795), .ZN(n20797) );
  NAND2_X1 U23779 ( .A1(n20797), .A2(n20796), .ZN(n20798) );
  NAND2_X1 U23780 ( .A1(n20799), .A2(n20798), .ZN(n20839) );
  AOI22_X1 U23781 ( .A1(n20801), .A2(n20841), .B1(n20800), .B2(n20839), .ZN(
        n20813) );
  INV_X1 U23782 ( .A(n20802), .ZN(n20805) );
  AOI21_X1 U23783 ( .B1(n20810), .B2(n20918), .A(n21012), .ZN(n20803) );
  AOI21_X1 U23784 ( .B1(n20805), .B2(n20804), .A(n20803), .ZN(n20806) );
  NOR2_X1 U23785 ( .A1(n20806), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20809) );
  AOI22_X1 U23786 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20845), .B1(
        n20844), .B2(n20811), .ZN(n20812) );
  OAI211_X1 U23787 ( .C1(n20814), .C2(n20918), .A(n20813), .B(n20812), .ZN(
        P1_U3145) );
  AOI22_X1 U23788 ( .A1(n20866), .A2(n20841), .B1(n20865), .B2(n20839), .ZN(
        n20817) );
  AOI22_X1 U23789 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20845), .B1(
        n20844), .B2(n20815), .ZN(n20816) );
  OAI211_X1 U23790 ( .C1(n20818), .C2(n20918), .A(n20817), .B(n20816), .ZN(
        P1_U3146) );
  AOI22_X1 U23791 ( .A1(n20820), .A2(n20841), .B1(n20819), .B2(n20839), .ZN(
        n20822) );
  AOI22_X1 U23792 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20845), .B1(
        n20844), .B2(n20874), .ZN(n20821) );
  OAI211_X1 U23793 ( .C1(n20877), .C2(n20918), .A(n20822), .B(n20821), .ZN(
        P1_U3147) );
  AOI22_X1 U23794 ( .A1(n20879), .A2(n20841), .B1(n20878), .B2(n20839), .ZN(
        n20825) );
  AOI22_X1 U23795 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20845), .B1(
        n20844), .B2(n20823), .ZN(n20824) );
  OAI211_X1 U23796 ( .C1(n20826), .C2(n20918), .A(n20825), .B(n20824), .ZN(
        P1_U3148) );
  AOI22_X1 U23797 ( .A1(n20828), .A2(n20841), .B1(n20827), .B2(n20839), .ZN(
        n20831) );
  AOI22_X1 U23798 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20845), .B1(
        n20844), .B2(n20829), .ZN(n20830) );
  OAI211_X1 U23799 ( .C1(n20832), .C2(n20918), .A(n20831), .B(n20830), .ZN(
        P1_U3149) );
  AOI22_X1 U23800 ( .A1(n20834), .A2(n20841), .B1(n20833), .B2(n20839), .ZN(
        n20836) );
  AOI22_X1 U23801 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20845), .B1(
        n20844), .B2(n20894), .ZN(n20835) );
  OAI211_X1 U23802 ( .C1(n20897), .C2(n20918), .A(n20836), .B(n20835), .ZN(
        P1_U3150) );
  AOI22_X1 U23803 ( .A1(n20901), .A2(n20841), .B1(n20899), .B2(n20839), .ZN(
        n20838) );
  AOI22_X1 U23804 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20845), .B1(
        n20844), .B2(n20902), .ZN(n20837) );
  OAI211_X1 U23805 ( .C1(n20907), .C2(n20918), .A(n20838), .B(n20837), .ZN(
        P1_U3151) );
  AOI22_X1 U23806 ( .A1(n20842), .A2(n20841), .B1(n20840), .B2(n20839), .ZN(
        n20847) );
  AOI22_X1 U23807 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20845), .B1(
        n20844), .B2(n20843), .ZN(n20846) );
  OAI211_X1 U23808 ( .C1(n20848), .C2(n20918), .A(n20847), .B(n20846), .ZN(
        P1_U3152) );
  OR2_X1 U23809 ( .A1(n20850), .A2(n20849), .ZN(n20853) );
  INV_X1 U23810 ( .A(n20910), .ZN(n20900) );
  AOI22_X1 U23811 ( .A1(n20900), .A2(n20689), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n10091), .ZN(n20852) );
  NAND2_X1 U23812 ( .A1(n20853), .A2(n20852), .ZN(n20898) );
  INV_X1 U23813 ( .A(n20898), .ZN(n20909) );
  OAI22_X1 U23814 ( .A1(n20855), .A2(n20910), .B1(n20909), .B2(n20854), .ZN(
        n20856) );
  INV_X1 U23815 ( .A(n20856), .ZN(n20863) );
  INV_X1 U23816 ( .A(n20857), .ZN(n20858) );
  NOR3_X1 U23817 ( .A1(n20858), .A2(n21012), .A3(n20991), .ZN(n20860) );
  OAI21_X1 U23818 ( .B1(n20860), .B2(n10091), .A(n20859), .ZN(n20915) );
  AOI22_X1 U23819 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20861), .ZN(n20862) );
  OAI211_X1 U23820 ( .C1(n20864), .C2(n20918), .A(n20863), .B(n20862), .ZN(
        P1_U3153) );
  AOI22_X1 U23821 ( .A1(n20866), .A2(n20900), .B1(n20865), .B2(n20898), .ZN(
        n20869) );
  AOI22_X1 U23822 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20867), .ZN(n20868) );
  OAI211_X1 U23823 ( .C1(n20870), .C2(n20918), .A(n20869), .B(n20868), .ZN(
        P1_U3154) );
  OAI22_X1 U23824 ( .A1(n20872), .A2(n20910), .B1(n20909), .B2(n20871), .ZN(
        n20873) );
  INV_X1 U23825 ( .A(n20873), .ZN(n20876) );
  INV_X1 U23826 ( .A(n20918), .ZN(n20903) );
  AOI22_X1 U23827 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20915), .B1(
        n20903), .B2(n20874), .ZN(n20875) );
  OAI211_X1 U23828 ( .C1(n20877), .C2(n20906), .A(n20876), .B(n20875), .ZN(
        P1_U3155) );
  AOI22_X1 U23829 ( .A1(n20879), .A2(n20900), .B1(n20878), .B2(n20898), .ZN(
        n20882) );
  AOI22_X1 U23830 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20880), .ZN(n20881) );
  OAI211_X1 U23831 ( .C1(n20883), .C2(n20918), .A(n20882), .B(n20881), .ZN(
        P1_U3156) );
  OAI22_X1 U23832 ( .A1(n20885), .A2(n20910), .B1(n20909), .B2(n20884), .ZN(
        n20886) );
  INV_X1 U23833 ( .A(n20886), .ZN(n20889) );
  AOI22_X1 U23834 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20887), .ZN(n20888) );
  OAI211_X1 U23835 ( .C1(n20890), .C2(n20918), .A(n20889), .B(n20888), .ZN(
        P1_U3157) );
  OAI22_X1 U23836 ( .A1(n20892), .A2(n20910), .B1(n20909), .B2(n20891), .ZN(
        n20893) );
  INV_X1 U23837 ( .A(n20893), .ZN(n20896) );
  AOI22_X1 U23838 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20915), .B1(
        n20903), .B2(n20894), .ZN(n20895) );
  OAI211_X1 U23839 ( .C1(n20897), .C2(n20906), .A(n20896), .B(n20895), .ZN(
        P1_U3158) );
  AOI22_X1 U23840 ( .A1(n20901), .A2(n20900), .B1(n20899), .B2(n20898), .ZN(
        n20905) );
  AOI22_X1 U23841 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20915), .B1(
        n20903), .B2(n20902), .ZN(n20904) );
  OAI211_X1 U23842 ( .C1(n20907), .C2(n20906), .A(n20905), .B(n20904), .ZN(
        P1_U3159) );
  OAI22_X1 U23843 ( .A1(n20911), .A2(n20910), .B1(n20909), .B2(n20908), .ZN(
        n20912) );
  INV_X1 U23844 ( .A(n20912), .ZN(n20917) );
  AOI22_X1 U23845 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20913), .ZN(n20916) );
  OAI211_X1 U23846 ( .C1(n20919), .C2(n20918), .A(n20917), .B(n20916), .ZN(
        P1_U3160) );
  NOR2_X1 U23847 ( .A1(n11887), .A2(n14021), .ZN(n20922) );
  INV_X1 U23848 ( .A(n20920), .ZN(n20921) );
  OAI21_X1 U23849 ( .B1(n20922), .B2(n21011), .A(n20921), .ZN(P1_U3163) );
  AND2_X1 U23850 ( .A1(n20923), .A2(P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(
        P1_U3164) );
  AND2_X1 U23851 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20923), .ZN(
        P1_U3165) );
  AND2_X1 U23852 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20923), .ZN(
        P1_U3166) );
  AND2_X1 U23853 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20923), .ZN(
        P1_U3167) );
  AND2_X1 U23854 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20923), .ZN(
        P1_U3168) );
  AND2_X1 U23855 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20923), .ZN(
        P1_U3169) );
  AND2_X1 U23856 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20923), .ZN(
        P1_U3170) );
  AND2_X1 U23857 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20923), .ZN(
        P1_U3171) );
  AND2_X1 U23858 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20923), .ZN(
        P1_U3172) );
  AND2_X1 U23859 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20923), .ZN(
        P1_U3173) );
  AND2_X1 U23860 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20923), .ZN(
        P1_U3174) );
  AND2_X1 U23861 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20923), .ZN(
        P1_U3175) );
  AND2_X1 U23862 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20923), .ZN(
        P1_U3176) );
  AND2_X1 U23863 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20923), .ZN(
        P1_U3177) );
  AND2_X1 U23864 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20923), .ZN(
        P1_U3178) );
  AND2_X1 U23865 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20923), .ZN(
        P1_U3179) );
  AND2_X1 U23866 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20923), .ZN(
        P1_U3180) );
  AND2_X1 U23867 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20923), .ZN(
        P1_U3181) );
  AND2_X1 U23868 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20923), .ZN(
        P1_U3182) );
  AND2_X1 U23869 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20923), .ZN(
        P1_U3183) );
  AND2_X1 U23870 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20923), .ZN(
        P1_U3184) );
  AND2_X1 U23871 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20923), .ZN(
        P1_U3185) );
  AND2_X1 U23872 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20923), .ZN(P1_U3186) );
  AND2_X1 U23873 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20923), .ZN(P1_U3187) );
  INV_X1 U23874 ( .A(P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n21291) );
  NOR2_X1 U23875 ( .A1(n20990), .A2(n21291), .ZN(P1_U3188) );
  AND2_X1 U23876 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20923), .ZN(P1_U3189) );
  AND2_X1 U23877 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20923), .ZN(P1_U3190) );
  AND2_X1 U23878 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20923), .ZN(P1_U3191) );
  AND2_X1 U23879 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20923), .ZN(P1_U3192) );
  AND2_X1 U23880 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20923), .ZN(P1_U3193) );
  AOI21_X1 U23881 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20924), .A(n20932), 
        .ZN(n20939) );
  NOR2_X1 U23882 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20925) );
  OAI21_X1 U23883 ( .B1(n20925), .B2(n20937), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20926) );
  AOI21_X1 U23884 ( .B1(NA), .B2(n20932), .A(n20926), .ZN(n20927) );
  OAI22_X1 U23885 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20939), .B1(n21009), 
        .B2(n20927), .ZN(P1_U3194) );
  INV_X1 U23886 ( .A(n20928), .ZN(n20931) );
  INV_X1 U23887 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20933) );
  NOR2_X1 U23888 ( .A1(n20932), .A2(n20933), .ZN(n20929) );
  OAI22_X1 U23889 ( .A1(n20931), .A2(n20930), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20929), .ZN(n20938) );
  NOR3_X1 U23890 ( .A1(NA), .A2(n20932), .A3(n21018), .ZN(n20934) );
  OAI22_X1 U23891 ( .A1(n20935), .A2(n20934), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20933), .ZN(n20936) );
  OAI22_X1 U23892 ( .A1(n20939), .A2(n20938), .B1(n20937), .B2(n20936), .ZN(
        P1_U3196) );
  NOR2_X2 U23893 ( .A1(n20940), .A2(n21022), .ZN(n20981) );
  AOI222_X1 U23894 ( .A1(n20980), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20981), .ZN(n20941) );
  INV_X1 U23895 ( .A(n20941), .ZN(P1_U3197) );
  AOI222_X1 U23896 ( .A1(n20981), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20980), .ZN(n20942) );
  INV_X1 U23897 ( .A(n20942), .ZN(P1_U3198) );
  INV_X1 U23898 ( .A(n20981), .ZN(n20974) );
  INV_X1 U23899 ( .A(n20980), .ZN(n20972) );
  OAI222_X1 U23900 ( .A1(n20974), .A2(n13943), .B1(n20943), .B2(n21009), .C1(
        n20944), .C2(n20972), .ZN(P1_U3199) );
  INV_X1 U23901 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21111) );
  OAI222_X1 U23902 ( .A1(n20972), .A2(n20946), .B1(n21111), .B2(n21009), .C1(
        n20944), .C2(n20974), .ZN(P1_U3200) );
  AOI22_X1 U23903 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n21022), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20980), .ZN(n20945) );
  OAI21_X1 U23904 ( .B1(n20946), .B2(n20974), .A(n20945), .ZN(P1_U3201) );
  AOI22_X1 U23905 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n21022), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20980), .ZN(n20947) );
  OAI21_X1 U23906 ( .B1(n20948), .B2(n20974), .A(n20947), .ZN(P1_U3202) );
  AOI222_X1 U23907 ( .A1(n20981), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20980), .ZN(n20949) );
  INV_X1 U23908 ( .A(n20949), .ZN(P1_U3203) );
  AOI22_X1 U23909 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n21022), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20980), .ZN(n20950) );
  OAI21_X1 U23910 ( .B1(n20951), .B2(n20974), .A(n20950), .ZN(P1_U3204) );
  AOI22_X1 U23911 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n21022), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20981), .ZN(n20952) );
  OAI21_X1 U23912 ( .B1(n14909), .B2(n20972), .A(n20952), .ZN(P1_U3205) );
  AOI222_X1 U23913 ( .A1(n20980), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20981), .ZN(n20953) );
  INV_X1 U23914 ( .A(n20953), .ZN(P1_U3206) );
  AOI22_X1 U23915 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21022), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20980), .ZN(n20954) );
  OAI21_X1 U23916 ( .B1(n20955), .B2(n20974), .A(n20954), .ZN(P1_U3207) );
  AOI22_X1 U23917 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21022), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20981), .ZN(n20956) );
  OAI21_X1 U23918 ( .B1(n20957), .B2(n20972), .A(n20956), .ZN(P1_U3208) );
  AOI222_X1 U23919 ( .A1(n20981), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20980), .ZN(n20958) );
  INV_X1 U23920 ( .A(n20958), .ZN(P1_U3209) );
  AOI222_X1 U23921 ( .A1(n20980), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20981), .ZN(n20959) );
  INV_X1 U23922 ( .A(n20959), .ZN(P1_U3210) );
  AOI222_X1 U23923 ( .A1(n20980), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20981), .ZN(n20960) );
  INV_X1 U23924 ( .A(n20960), .ZN(P1_U3211) );
  AOI22_X1 U23925 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21022), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20980), .ZN(n20961) );
  OAI21_X1 U23926 ( .B1(n21097), .B2(n20974), .A(n20961), .ZN(P1_U3212) );
  AOI22_X1 U23927 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21022), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20981), .ZN(n20962) );
  OAI21_X1 U23928 ( .B1(n20963), .B2(n20972), .A(n20962), .ZN(P1_U3213) );
  AOI222_X1 U23929 ( .A1(n20981), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20980), .ZN(n20964) );
  INV_X1 U23930 ( .A(n20964), .ZN(P1_U3214) );
  INV_X1 U23931 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n21303) );
  OAI222_X1 U23932 ( .A1(n20974), .A2(n20966), .B1(n21303), .B2(n21009), .C1(
        n20965), .C2(n20972), .ZN(P1_U3215) );
  AOI222_X1 U23933 ( .A1(n20980), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20981), .ZN(n20967) );
  INV_X1 U23934 ( .A(n20967), .ZN(P1_U3216) );
  AOI222_X1 U23935 ( .A1(n20981), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20980), .ZN(n20968) );
  INV_X1 U23936 ( .A(n20968), .ZN(P1_U3217) );
  AOI22_X1 U23937 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21022), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20980), .ZN(n20969) );
  OAI21_X1 U23938 ( .B1(n20970), .B2(n20974), .A(n20969), .ZN(P1_U3218) );
  AOI22_X1 U23939 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21022), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20981), .ZN(n20971) );
  OAI21_X1 U23940 ( .B1(n14644), .B2(n20972), .A(n20971), .ZN(P1_U3219) );
  INV_X1 U23941 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21260) );
  OAI222_X1 U23942 ( .A1(n20974), .A2(n14644), .B1(n21260), .B2(n21009), .C1(
        n20973), .C2(n20972), .ZN(P1_U3220) );
  AOI222_X1 U23943 ( .A1(n20981), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20980), .ZN(n20975) );
  INV_X1 U23944 ( .A(n20975), .ZN(P1_U3221) );
  AOI222_X1 U23945 ( .A1(n20981), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20980), .ZN(n20976) );
  INV_X1 U23946 ( .A(n20976), .ZN(P1_U3222) );
  AOI222_X1 U23947 ( .A1(n20981), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20980), .ZN(n20977) );
  INV_X1 U23948 ( .A(n20977), .ZN(P1_U3223) );
  AOI222_X1 U23949 ( .A1(n20981), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20980), .ZN(n20978) );
  INV_X1 U23950 ( .A(n20978), .ZN(P1_U3224) );
  AOI222_X1 U23951 ( .A1(n20981), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20980), .ZN(n20979) );
  INV_X1 U23952 ( .A(n20979), .ZN(P1_U3225) );
  AOI222_X1 U23953 ( .A1(n20981), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21022), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20980), .ZN(n20982) );
  INV_X1 U23954 ( .A(n20982), .ZN(P1_U3226) );
  OAI22_X1 U23955 ( .A1(n21022), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21009), .ZN(n20983) );
  INV_X1 U23956 ( .A(n20983), .ZN(P1_U3458) );
  OAI22_X1 U23957 ( .A1(n21022), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21009), .ZN(n20984) );
  INV_X1 U23958 ( .A(n20984), .ZN(P1_U3459) );
  OAI22_X1 U23959 ( .A1(n21022), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21009), .ZN(n20985) );
  INV_X1 U23960 ( .A(n20985), .ZN(P1_U3460) );
  OAI22_X1 U23961 ( .A1(n21022), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21009), .ZN(n20986) );
  INV_X1 U23962 ( .A(n20986), .ZN(P1_U3461) );
  OAI21_X1 U23963 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20990), .A(n20988), 
        .ZN(n20987) );
  INV_X1 U23964 ( .A(n20987), .ZN(P1_U3464) );
  OAI21_X1 U23965 ( .B1(n20990), .B2(n20989), .A(n20988), .ZN(P1_U3465) );
  INV_X1 U23966 ( .A(n20996), .ZN(n20999) );
  OR2_X1 U23967 ( .A1(n20991), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20993) );
  OAI211_X1 U23968 ( .C1(n20994), .C2(n14101), .A(n20993), .B(n20992), .ZN(
        n20995) );
  INV_X1 U23969 ( .A(n20995), .ZN(n20997) );
  AOI22_X1 U23970 ( .A1(n20999), .A2(n20998), .B1(n20997), .B2(n20996), .ZN(
        P1_U3477) );
  AOI21_X1 U23971 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21001) );
  AOI22_X1 U23972 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21001), .B2(n21000), .ZN(n21004) );
  INV_X1 U23973 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21003) );
  AOI22_X1 U23974 ( .A1(n21007), .A2(n21004), .B1(n21003), .B2(n21002), .ZN(
        P1_U3481) );
  INV_X1 U23975 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21006) );
  OAI21_X1 U23976 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21007), .ZN(n21005) );
  OAI21_X1 U23977 ( .B1(n21007), .B2(n21006), .A(n21005), .ZN(P1_U3482) );
  AOI22_X1 U23978 ( .A1(n21009), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21008), 
        .B2(n21022), .ZN(P1_U3483) );
  AOI211_X1 U23979 ( .C1(n21013), .C2(n21012), .A(n21011), .B(n21010), .ZN(
        n21015) );
  OAI21_X1 U23980 ( .B1(n21015), .B2(n11887), .A(n21014), .ZN(n21021) );
  AOI211_X1 U23981 ( .C1(n21019), .C2(n21018), .A(n21017), .B(n21016), .ZN(
        n21020) );
  MUX2_X1 U23982 ( .A(n21021), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21020), 
        .Z(P1_U3485) );
  MUX2_X1 U23983 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21022), .Z(P1_U3486) );
  INV_X1 U23984 ( .A(keyinput13), .ZN(n21023) );
  NOR4_X1 U23985 ( .A1(keyinput57), .A2(keyinput53), .A3(keyinput40), .A4(
        n21023), .ZN(n21084) );
  NAND2_X1 U23986 ( .A1(keyinput19), .A2(keyinput25), .ZN(n21024) );
  NOR3_X1 U23987 ( .A1(keyinput113), .A2(keyinput91), .A3(n21024), .ZN(n21083)
         );
  NAND2_X1 U23988 ( .A1(keyinput20), .A2(keyinput31), .ZN(n21025) );
  NOR3_X1 U23989 ( .A1(keyinput70), .A2(keyinput90), .A3(n21025), .ZN(n21026)
         );
  NAND3_X1 U23990 ( .A1(keyinput7), .A2(keyinput101), .A3(n21026), .ZN(n21034)
         );
  NOR3_X1 U23991 ( .A1(keyinput117), .A2(keyinput86), .A3(keyinput51), .ZN(
        n21027) );
  NAND2_X1 U23992 ( .A1(keyinput52), .A2(n21027), .ZN(n21028) );
  NOR4_X1 U23993 ( .A1(keyinput69), .A2(keyinput112), .A3(keyinput24), .A4(
        n21028), .ZN(n21032) );
  NOR2_X1 U23994 ( .A1(keyinput114), .A2(keyinput54), .ZN(n21029) );
  NAND3_X1 U23995 ( .A1(keyinput124), .A2(keyinput32), .A3(n21029), .ZN(n21030) );
  NOR3_X1 U23996 ( .A1(keyinput38), .A2(keyinput115), .A3(n21030), .ZN(n21031)
         );
  NAND4_X1 U23997 ( .A1(n21032), .A2(keyinput119), .A3(keyinput71), .A4(n21031), .ZN(n21033) );
  NOR4_X1 U23998 ( .A1(keyinput81), .A2(keyinput49), .A3(n21034), .A4(n21033), 
        .ZN(n21082) );
  NAND4_X1 U23999 ( .A1(keyinput110), .A2(keyinput95), .A3(keyinput48), .A4(
        keyinput122), .ZN(n21035) );
  NOR3_X1 U24000 ( .A1(keyinput120), .A2(keyinput47), .A3(n21035), .ZN(n21049)
         );
  NAND2_X1 U24001 ( .A1(keyinput39), .A2(keyinput22), .ZN(n21036) );
  NOR3_X1 U24002 ( .A1(keyinput27), .A2(keyinput10), .A3(n21036), .ZN(n21037)
         );
  NAND3_X1 U24003 ( .A1(keyinput17), .A2(keyinput6), .A3(n21037), .ZN(n21046)
         );
  INV_X1 U24004 ( .A(keyinput96), .ZN(n21038) );
  NOR4_X1 U24005 ( .A1(keyinput42), .A2(keyinput89), .A3(keyinput36), .A4(
        n21038), .ZN(n21044) );
  NOR4_X1 U24006 ( .A1(keyinput85), .A2(keyinput106), .A3(keyinput56), .A4(
        keyinput63), .ZN(n21043) );
  NAND3_X1 U24007 ( .A1(keyinput8), .A2(keyinput44), .A3(keyinput121), .ZN(
        n21039) );
  NOR2_X1 U24008 ( .A1(keyinput66), .A2(n21039), .ZN(n21042) );
  INV_X1 U24009 ( .A(keyinput64), .ZN(n21040) );
  NOR4_X1 U24010 ( .A1(keyinput50), .A2(keyinput98), .A3(keyinput0), .A4(
        n21040), .ZN(n21041) );
  NAND4_X1 U24011 ( .A1(n21044), .A2(n21043), .A3(n21042), .A4(n21041), .ZN(
        n21045) );
  NOR4_X1 U24012 ( .A1(keyinput107), .A2(keyinput33), .A3(n21046), .A4(n21045), 
        .ZN(n21048) );
  INV_X1 U24013 ( .A(keyinput83), .ZN(n21047) );
  NAND4_X1 U24014 ( .A1(keyinput26), .A2(n21049), .A3(n21048), .A4(n21047), 
        .ZN(n21080) );
  NOR2_X1 U24015 ( .A1(keyinput104), .A2(keyinput14), .ZN(n21050) );
  NAND3_X1 U24016 ( .A1(keyinput88), .A2(keyinput125), .A3(n21050), .ZN(n21051) );
  NOR3_X1 U24017 ( .A1(keyinput23), .A2(keyinput55), .A3(n21051), .ZN(n21063)
         );
  NAND2_X1 U24018 ( .A1(keyinput15), .A2(keyinput93), .ZN(n21052) );
  NOR3_X1 U24019 ( .A1(keyinput9), .A2(keyinput84), .A3(n21052), .ZN(n21053)
         );
  NAND3_X1 U24020 ( .A1(keyinput41), .A2(keyinput79), .A3(n21053), .ZN(n21061)
         );
  INV_X1 U24021 ( .A(keyinput58), .ZN(n21096) );
  NOR4_X1 U24022 ( .A1(keyinput67), .A2(keyinput43), .A3(keyinput108), .A4(
        n21096), .ZN(n21059) );
  NOR4_X1 U24023 ( .A1(keyinput118), .A2(keyinput35), .A3(keyinput28), .A4(
        keyinput78), .ZN(n21058) );
  INV_X1 U24024 ( .A(keyinput109), .ZN(n21054) );
  NOR4_X1 U24025 ( .A1(keyinput127), .A2(keyinput21), .A3(keyinput116), .A4(
        n21054), .ZN(n21057) );
  NAND3_X1 U24026 ( .A1(keyinput45), .A2(keyinput77), .A3(keyinput11), .ZN(
        n21055) );
  NOR2_X1 U24027 ( .A1(keyinput60), .A2(n21055), .ZN(n21056) );
  NAND4_X1 U24028 ( .A1(n21059), .A2(n21058), .A3(n21057), .A4(n21056), .ZN(
        n21060) );
  NOR4_X1 U24029 ( .A1(keyinput18), .A2(keyinput4), .A3(n21061), .A4(n21060), 
        .ZN(n21062) );
  NAND4_X1 U24030 ( .A1(keyinput12), .A2(keyinput1), .A3(n21063), .A4(n21062), 
        .ZN(n21079) );
  NOR4_X1 U24031 ( .A1(keyinput74), .A2(keyinput3), .A3(keyinput76), .A4(
        keyinput30), .ZN(n21069) );
  NAND2_X1 U24032 ( .A1(keyinput82), .A2(keyinput59), .ZN(n21064) );
  NOR3_X1 U24033 ( .A1(keyinput87), .A2(keyinput29), .A3(n21064), .ZN(n21068)
         );
  NAND2_X1 U24034 ( .A1(keyinput2), .A2(keyinput126), .ZN(n21065) );
  NOR3_X1 U24035 ( .A1(keyinput94), .A2(keyinput105), .A3(n21065), .ZN(n21067)
         );
  INV_X1 U24036 ( .A(keyinput65), .ZN(n21197) );
  NOR4_X1 U24037 ( .A1(keyinput75), .A2(keyinput37), .A3(keyinput111), .A4(
        n21197), .ZN(n21066) );
  NAND4_X1 U24038 ( .A1(n21069), .A2(n21068), .A3(n21067), .A4(n21066), .ZN(
        n21078) );
  NOR4_X1 U24039 ( .A1(keyinput61), .A2(keyinput16), .A3(keyinput92), .A4(
        keyinput68), .ZN(n21076) );
  NAND3_X1 U24040 ( .A1(keyinput62), .A2(keyinput99), .A3(keyinput5), .ZN(
        n21070) );
  NOR2_X1 U24041 ( .A1(keyinput73), .A2(n21070), .ZN(n21075) );
  NAND2_X1 U24042 ( .A1(keyinput102), .A2(keyinput80), .ZN(n21071) );
  NOR3_X1 U24043 ( .A1(keyinput72), .A2(keyinput103), .A3(n21071), .ZN(n21074)
         );
  NAND2_X1 U24044 ( .A1(keyinput97), .A2(keyinput34), .ZN(n21072) );
  NOR3_X1 U24045 ( .A1(keyinput100), .A2(keyinput123), .A3(n21072), .ZN(n21073) );
  NAND4_X1 U24046 ( .A1(n21076), .A2(n21075), .A3(n21074), .A4(n21073), .ZN(
        n21077) );
  NOR4_X1 U24047 ( .A1(n21080), .A2(n21079), .A3(n21078), .A4(n21077), .ZN(
        n21081) );
  NAND4_X1 U24048 ( .A1(n21084), .A2(n21083), .A3(n21082), .A4(n21081), .ZN(
        n21085) );
  AOI21_X1 U24049 ( .B1(keyinput46), .B2(n21085), .A(n21241), .ZN(n21342) );
  INV_X1 U24050 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n21088) );
  INV_X1 U24051 ( .A(keyinput78), .ZN(n21090) );
  AOI22_X1 U24052 ( .A1(n21091), .A2(keyinput67), .B1(
        P2_DATAWIDTH_REG_11__SCAN_IN), .B2(n21090), .ZN(n21089) );
  OAI221_X1 U24053 ( .B1(n21091), .B2(keyinput67), .C1(n21090), .C2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A(n21089), .ZN(n21100) );
  AOI22_X1 U24054 ( .A1(n21094), .A2(keyinput43), .B1(n21093), .B2(keyinput108), .ZN(n21092) );
  OAI221_X1 U24055 ( .B1(n21094), .B2(keyinput43), .C1(n21093), .C2(
        keyinput108), .A(n21092), .ZN(n21099) );
  AOI22_X1 U24056 ( .A1(n21097), .A2(keyinput104), .B1(
        P1_DATAWIDTH_REG_31__SCAN_IN), .B2(n21096), .ZN(n21095) );
  OAI221_X1 U24057 ( .B1(n21097), .B2(keyinput104), .C1(n21096), .C2(
        P1_DATAWIDTH_REG_31__SCAN_IN), .A(n21095), .ZN(n21098) );
  NOR4_X1 U24058 ( .A1(n21101), .A2(n21100), .A3(n21099), .A4(n21098), .ZN(
        n21149) );
  INV_X1 U24059 ( .A(keyinput125), .ZN(n21103) );
  AOI22_X1 U24060 ( .A1(n21104), .A2(keyinput88), .B1(P3_DATAO_REG_16__SCAN_IN), .B2(n21103), .ZN(n21102) );
  OAI221_X1 U24061 ( .B1(n21104), .B2(keyinput88), .C1(n21103), .C2(
        P3_DATAO_REG_16__SCAN_IN), .A(n21102), .ZN(n21116) );
  INV_X1 U24062 ( .A(keyinput12), .ZN(n21106) );
  AOI22_X1 U24063 ( .A1(n12972), .A2(keyinput14), .B1(P1_LWORD_REG_3__SCAN_IN), 
        .B2(n21106), .ZN(n21105) );
  OAI221_X1 U24064 ( .B1(n12972), .B2(keyinput14), .C1(n21106), .C2(
        P1_LWORD_REG_3__SCAN_IN), .A(n21105), .ZN(n21115) );
  INV_X1 U24065 ( .A(keyinput23), .ZN(n21108) );
  AOI22_X1 U24066 ( .A1(n21109), .A2(keyinput1), .B1(P3_BE_N_REG_2__SCAN_IN), 
        .B2(n21108), .ZN(n21107) );
  OAI221_X1 U24067 ( .B1(n21109), .B2(keyinput1), .C1(n21108), .C2(
        P3_BE_N_REG_2__SCAN_IN), .A(n21107), .ZN(n21114) );
  AOI22_X1 U24068 ( .A1(n21112), .A2(keyinput55), .B1(keyinput41), .B2(n21111), 
        .ZN(n21110) );
  OAI221_X1 U24069 ( .B1(n21112), .B2(keyinput55), .C1(n21111), .C2(keyinput41), .A(n21110), .ZN(n21113) );
  NOR4_X1 U24070 ( .A1(n21116), .A2(n21115), .A3(n21114), .A4(n21113), .ZN(
        n21148) );
  INV_X1 U24071 ( .A(keyinput79), .ZN(n21119) );
  INV_X1 U24072 ( .A(keyinput93), .ZN(n21118) );
  AOI22_X1 U24073 ( .A1(n21119), .A2(P3_EAX_REG_18__SCAN_IN), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n21118), .ZN(n21117) );
  OAI221_X1 U24074 ( .B1(n21119), .B2(P3_EAX_REG_18__SCAN_IN), .C1(n21118), 
        .C2(P1_DATAO_REG_20__SCAN_IN), .A(n21117), .ZN(n21131) );
  AOI22_X1 U24075 ( .A1(n21122), .A2(keyinput84), .B1(n21121), .B2(keyinput9), 
        .ZN(n21120) );
  OAI221_X1 U24076 ( .B1(n21122), .B2(keyinput84), .C1(n21121), .C2(keyinput9), 
        .A(n21120), .ZN(n21130) );
  INV_X1 U24077 ( .A(keyinput18), .ZN(n21124) );
  AOI22_X1 U24078 ( .A1(n9747), .A2(keyinput15), .B1(
        P2_BYTEENABLE_REG_3__SCAN_IN), .B2(n21124), .ZN(n21123) );
  OAI221_X1 U24079 ( .B1(n9747), .B2(keyinput15), .C1(n21124), .C2(
        P2_BYTEENABLE_REG_3__SCAN_IN), .A(n21123), .ZN(n21129) );
  AOI22_X1 U24080 ( .A1(n21127), .A2(keyinput4), .B1(n21126), .B2(keyinput77), 
        .ZN(n21125) );
  OAI221_X1 U24081 ( .B1(n21127), .B2(keyinput4), .C1(n21126), .C2(keyinput77), 
        .A(n21125), .ZN(n21128) );
  NOR4_X1 U24082 ( .A1(n21131), .A2(n21130), .A3(n21129), .A4(n21128), .ZN(
        n21147) );
  INV_X1 U24083 ( .A(DATAI_29_), .ZN(n21133) );
  AOI22_X1 U24084 ( .A1(n21133), .A2(keyinput11), .B1(n11100), .B2(keyinput127), .ZN(n21132) );
  OAI221_X1 U24085 ( .B1(n21133), .B2(keyinput11), .C1(n11100), .C2(
        keyinput127), .A(n21132), .ZN(n21145) );
  INV_X1 U24086 ( .A(keyinput21), .ZN(n21135) );
  AOI22_X1 U24087 ( .A1(n21136), .A2(keyinput45), .B1(P1_DATAO_REG_24__SCAN_IN), .B2(n21135), .ZN(n21134) );
  OAI221_X1 U24088 ( .B1(n21136), .B2(keyinput45), .C1(n21135), .C2(
        P1_DATAO_REG_24__SCAN_IN), .A(n21134), .ZN(n21144) );
  AOI22_X1 U24089 ( .A1(n21138), .A2(keyinput60), .B1(n14505), .B2(keyinput116), .ZN(n21137) );
  OAI221_X1 U24090 ( .B1(n21138), .B2(keyinput60), .C1(n14505), .C2(
        keyinput116), .A(n21137), .ZN(n21143) );
  INV_X1 U24091 ( .A(keyinput5), .ZN(n21140) );
  AOI22_X1 U24092 ( .A1(n21141), .A2(keyinput109), .B1(
        P3_DATAO_REG_26__SCAN_IN), .B2(n21140), .ZN(n21139) );
  OAI221_X1 U24093 ( .B1(n21141), .B2(keyinput109), .C1(n21140), .C2(
        P3_DATAO_REG_26__SCAN_IN), .A(n21139), .ZN(n21142) );
  NOR4_X1 U24094 ( .A1(n21145), .A2(n21144), .A3(n21143), .A4(n21142), .ZN(
        n21146) );
  NAND4_X1 U24095 ( .A1(n21149), .A2(n21148), .A3(n21147), .A4(n21146), .ZN(
        n21341) );
  AOI22_X1 U24096 ( .A1(n21152), .A2(keyinput73), .B1(n21151), .B2(keyinput99), 
        .ZN(n21150) );
  OAI221_X1 U24097 ( .B1(n21152), .B2(keyinput73), .C1(n21151), .C2(keyinput99), .A(n21150), .ZN(n21165) );
  INV_X1 U24098 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n21154) );
  AOI22_X1 U24099 ( .A1(n21155), .A2(keyinput62), .B1(n21154), .B2(keyinput61), 
        .ZN(n21153) );
  OAI221_X1 U24100 ( .B1(n21155), .B2(keyinput62), .C1(n21154), .C2(keyinput61), .A(n21153), .ZN(n21164) );
  AOI22_X1 U24101 ( .A1(n21158), .A2(keyinput16), .B1(keyinput92), .B2(n21157), 
        .ZN(n21156) );
  OAI221_X1 U24102 ( .B1(n21158), .B2(keyinput16), .C1(n21157), .C2(keyinput92), .A(n21156), .ZN(n21163) );
  INV_X1 U24103 ( .A(keyinput100), .ZN(n21160) );
  AOI22_X1 U24104 ( .A1(n21161), .A2(keyinput68), .B1(P3_EAX_REG_30__SCAN_IN), 
        .B2(n21160), .ZN(n21159) );
  OAI221_X1 U24105 ( .B1(n21161), .B2(keyinput68), .C1(n21160), .C2(
        P3_EAX_REG_30__SCAN_IN), .A(n21159), .ZN(n21162) );
  NOR4_X1 U24106 ( .A1(n21165), .A2(n21164), .A3(n21163), .A4(n21162), .ZN(
        n21210) );
  INV_X1 U24107 ( .A(keyinput34), .ZN(n21167) );
  AOI22_X1 U24108 ( .A1(n21168), .A2(keyinput97), .B1(
        P2_READREQUEST_REG_SCAN_IN), .B2(n21167), .ZN(n21166) );
  OAI221_X1 U24109 ( .B1(n21168), .B2(keyinput97), .C1(n21167), .C2(
        P2_READREQUEST_REG_SCAN_IN), .A(n21166), .ZN(n21177) );
  INV_X1 U24110 ( .A(keyinput72), .ZN(n21170) );
  AOI22_X1 U24111 ( .A1(n16390), .A2(keyinput123), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n21170), .ZN(n21169) );
  OAI221_X1 U24112 ( .B1(n16390), .B2(keyinput123), .C1(n21170), .C2(
        P2_DATAO_REG_16__SCAN_IN), .A(n21169), .ZN(n21176) );
  AOI22_X1 U24113 ( .A1(n11099), .A2(keyinput80), .B1(keyinput102), .B2(n16391), .ZN(n21171) );
  OAI221_X1 U24114 ( .B1(n11099), .B2(keyinput80), .C1(n16391), .C2(
        keyinput102), .A(n21171), .ZN(n21175) );
  AOI22_X1 U24115 ( .A1(n19251), .A2(keyinput103), .B1(keyinput87), .B2(n21173), .ZN(n21172) );
  OAI221_X1 U24116 ( .B1(n19251), .B2(keyinput103), .C1(n21173), .C2(
        keyinput87), .A(n21172), .ZN(n21174) );
  NOR4_X1 U24117 ( .A1(n21177), .A2(n21176), .A3(n21175), .A4(n21174), .ZN(
        n21209) );
  INV_X1 U24118 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n21180) );
  AOI22_X1 U24119 ( .A1(n21180), .A2(keyinput59), .B1(keyinput74), .B2(n21179), 
        .ZN(n21178) );
  OAI221_X1 U24120 ( .B1(n21180), .B2(keyinput59), .C1(n21179), .C2(keyinput74), .A(n21178), .ZN(n21193) );
  INV_X1 U24121 ( .A(keyinput82), .ZN(n21182) );
  AOI22_X1 U24122 ( .A1(n21183), .A2(keyinput3), .B1(P2_DATAO_REG_7__SCAN_IN), 
        .B2(n21182), .ZN(n21181) );
  OAI221_X1 U24123 ( .B1(n21183), .B2(keyinput3), .C1(n21182), .C2(
        P2_DATAO_REG_7__SCAN_IN), .A(n21181), .ZN(n21192) );
  INV_X1 U24124 ( .A(keyinput29), .ZN(n21185) );
  AOI22_X1 U24125 ( .A1(n21186), .A2(keyinput76), .B1(P2_UWORD_REG_10__SCAN_IN), .B2(n21185), .ZN(n21184) );
  OAI221_X1 U24126 ( .B1(n21186), .B2(keyinput76), .C1(n21185), .C2(
        P2_UWORD_REG_10__SCAN_IN), .A(n21184), .ZN(n21191) );
  INV_X1 U24127 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n21189) );
  INV_X1 U24128 ( .A(keyinput75), .ZN(n21188) );
  AOI22_X1 U24129 ( .A1(n21189), .A2(keyinput30), .B1(
        P3_ADDRESS_REG_25__SCAN_IN), .B2(n21188), .ZN(n21187) );
  OAI221_X1 U24130 ( .B1(n21189), .B2(keyinput30), .C1(n21188), .C2(
        P3_ADDRESS_REG_25__SCAN_IN), .A(n21187), .ZN(n21190) );
  NOR4_X1 U24131 ( .A1(n21193), .A2(n21192), .A3(n21191), .A4(n21190), .ZN(
        n21208) );
  AOI22_X1 U24132 ( .A1(n21195), .A2(keyinput37), .B1(keyinput111), .B2(n14034), .ZN(n21194) );
  OAI221_X1 U24133 ( .B1(n21195), .B2(keyinput37), .C1(n14034), .C2(
        keyinput111), .A(n21194), .ZN(n21206) );
  AOI22_X1 U24134 ( .A1(n21198), .A2(keyinput94), .B1(
        P2_DATAWIDTH_REG_4__SCAN_IN), .B2(n21197), .ZN(n21196) );
  OAI221_X1 U24135 ( .B1(n21198), .B2(keyinput94), .C1(n21197), .C2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A(n21196), .ZN(n21205) );
  AOI22_X1 U24136 ( .A1(n10017), .A2(keyinput126), .B1(n21200), .B2(keyinput2), 
        .ZN(n21199) );
  OAI221_X1 U24137 ( .B1(n10017), .B2(keyinput126), .C1(n21200), .C2(keyinput2), .A(n21199), .ZN(n21204) );
  INV_X1 U24138 ( .A(keyinput69), .ZN(n21202) );
  AOI22_X1 U24139 ( .A1(n9905), .A2(keyinput105), .B1(P3_LWORD_REG_9__SCAN_IN), 
        .B2(n21202), .ZN(n21201) );
  OAI221_X1 U24140 ( .B1(n9905), .B2(keyinput105), .C1(n21202), .C2(
        P3_LWORD_REG_9__SCAN_IN), .A(n21201), .ZN(n21203) );
  NOR4_X1 U24141 ( .A1(n21206), .A2(n21205), .A3(n21204), .A4(n21203), .ZN(
        n21207) );
  NAND4_X1 U24142 ( .A1(n21210), .A2(n21209), .A3(n21208), .A4(n21207), .ZN(
        n21340) );
  INV_X1 U24143 ( .A(keyinput24), .ZN(n21215) );
  INV_X1 U24144 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n21212) );
  OAI22_X1 U24145 ( .A1(n10621), .A2(keyinput112), .B1(n21212), .B2(keyinput52), .ZN(n21211) );
  AOI221_X1 U24146 ( .B1(n10621), .B2(keyinput112), .C1(keyinput52), .C2(
        n21212), .A(n21211), .ZN(n21213) );
  OAI221_X1 U24147 ( .B1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n21215), .C1(
        n21214), .C2(keyinput24), .A(n21213), .ZN(n21240) );
  INV_X1 U24148 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21217) );
  OAI22_X1 U24149 ( .A1(n21218), .A2(keyinput90), .B1(n21217), .B2(keyinput70), 
        .ZN(n21216) );
  AOI221_X1 U24150 ( .B1(n21218), .B2(keyinput90), .C1(keyinput70), .C2(n21217), .A(n21216), .ZN(n21238) );
  OAI22_X1 U24151 ( .A1(n21221), .A2(keyinput49), .B1(n21220), .B2(keyinput31), 
        .ZN(n21219) );
  AOI221_X1 U24152 ( .B1(n21221), .B2(keyinput49), .C1(keyinput31), .C2(n21220), .A(n21219), .ZN(n21237) );
  INV_X1 U24153 ( .A(keyinput7), .ZN(n21223) );
  AOI22_X1 U24154 ( .A1(n21224), .A2(keyinput20), .B1(P3_LWORD_REG_12__SCAN_IN), .B2(n21223), .ZN(n21222) );
  OAI221_X1 U24155 ( .B1(n21224), .B2(keyinput20), .C1(n21223), .C2(
        P3_LWORD_REG_12__SCAN_IN), .A(n21222), .ZN(n21235) );
  INV_X1 U24156 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n21227) );
  AOI22_X1 U24157 ( .A1(n21227), .A2(keyinput51), .B1(keyinput117), .B2(n21226), .ZN(n21225) );
  OAI221_X1 U24158 ( .B1(n21227), .B2(keyinput51), .C1(n21226), .C2(
        keyinput117), .A(n21225), .ZN(n21234) );
  INV_X1 U24159 ( .A(keyinput113), .ZN(n21229) );
  AOI22_X1 U24160 ( .A1(n11254), .A2(keyinput101), .B1(P3_DATAO_REG_4__SCAN_IN), .B2(n21229), .ZN(n21228) );
  OAI221_X1 U24161 ( .B1(n11254), .B2(keyinput101), .C1(n21229), .C2(
        P3_DATAO_REG_4__SCAN_IN), .A(n21228), .ZN(n21233) );
  XNOR2_X1 U24162 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(keyinput81), 
        .ZN(n21231) );
  XNOR2_X1 U24163 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B(keyinput86), .ZN(
        n21230) );
  NAND2_X1 U24164 ( .A1(n21231), .A2(n21230), .ZN(n21232) );
  NOR4_X1 U24165 ( .A1(n21235), .A2(n21234), .A3(n21233), .A4(n21232), .ZN(
        n21236) );
  NAND3_X1 U24166 ( .A1(n21238), .A2(n21237), .A3(n21236), .ZN(n21239) );
  AOI211_X1 U24167 ( .C1(keyinput46), .C2(n21241), .A(n21240), .B(n21239), 
        .ZN(n21338) );
  XOR2_X1 U24168 ( .A(keyinput98), .B(n21242), .Z(n21248) );
  INV_X1 U24169 ( .A(keyinput66), .ZN(n21243) );
  XOR2_X1 U24170 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n21243), .Z(n21247)
         );
  XNOR2_X1 U24171 ( .A(n21244), .B(keyinput0), .ZN(n21246) );
  XNOR2_X1 U24172 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B(keyinput64), .ZN(
        n21245) );
  NAND4_X1 U24173 ( .A1(n21248), .A2(n21247), .A3(n21246), .A4(n21245), .ZN(
        n21257) );
  AOI22_X1 U24174 ( .A1(n21251), .A2(keyinput121), .B1(keyinput44), .B2(n21250), .ZN(n21249) );
  OAI221_X1 U24175 ( .B1(n21251), .B2(keyinput121), .C1(n21250), .C2(
        keyinput44), .A(n21249), .ZN(n21256) );
  AOI22_X1 U24176 ( .A1(n21254), .A2(keyinput8), .B1(n21253), .B2(keyinput118), 
        .ZN(n21252) );
  OAI221_X1 U24177 ( .B1(n21254), .B2(keyinput8), .C1(n21253), .C2(keyinput118), .A(n21252), .ZN(n21255) );
  NOR3_X1 U24178 ( .A1(n21257), .A2(n21256), .A3(n21255), .ZN(n21337) );
  INV_X1 U24179 ( .A(keyinput39), .ZN(n21259) );
  AOI22_X1 U24180 ( .A1(n21260), .A2(keyinput17), .B1(P3_EAX_REG_4__SCAN_IN), 
        .B2(n21259), .ZN(n21258) );
  OAI221_X1 U24181 ( .B1(n21260), .B2(keyinput17), .C1(n21259), .C2(
        P3_EAX_REG_4__SCAN_IN), .A(n21258), .ZN(n21264) );
  XNOR2_X1 U24182 ( .A(n21261), .B(keyinput33), .ZN(n21263) );
  XOR2_X1 U24183 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B(keyinput50), .Z(
        n21262) );
  OR3_X1 U24184 ( .A1(n21264), .A2(n21263), .A3(n21262), .ZN(n21272) );
  AOI22_X1 U24185 ( .A1(n21267), .A2(keyinput22), .B1(keyinput10), .B2(n21266), 
        .ZN(n21265) );
  OAI221_X1 U24186 ( .B1(n21267), .B2(keyinput22), .C1(n21266), .C2(keyinput10), .A(n21265), .ZN(n21271) );
  INV_X1 U24187 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21269) );
  AOI22_X1 U24188 ( .A1(n11613), .A2(keyinput6), .B1(keyinput107), .B2(n21269), 
        .ZN(n21268) );
  OAI221_X1 U24189 ( .B1(n11613), .B2(keyinput6), .C1(n21269), .C2(keyinput107), .A(n21268), .ZN(n21270) );
  NOR3_X1 U24190 ( .A1(n21272), .A2(n21271), .A3(n21270), .ZN(n21336) );
  INV_X1 U24191 ( .A(keyinput119), .ZN(n21274) );
  OAI22_X1 U24192 ( .A1(n21275), .A2(keyinput114), .B1(n21274), .B2(
        P2_DATAO_REG_24__SCAN_IN), .ZN(n21273) );
  AOI221_X1 U24193 ( .B1(n21275), .B2(keyinput114), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(n21274), .A(n21273), .ZN(n21286) );
  OAI22_X1 U24194 ( .A1(n21277), .A2(keyinput115), .B1(n11156), .B2(
        keyinput124), .ZN(n21276) );
  AOI221_X1 U24195 ( .B1(n21277), .B2(keyinput115), .C1(keyinput124), .C2(
        n11156), .A(n21276), .ZN(n21285) );
  OAI22_X1 U24196 ( .A1(n21279), .A2(keyinput54), .B1(n10831), .B2(keyinput83), 
        .ZN(n21278) );
  AOI221_X1 U24197 ( .B1(n21279), .B2(keyinput54), .C1(keyinput83), .C2(n10831), .A(n21278), .ZN(n21284) );
  INV_X1 U24198 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n21282) );
  INV_X1 U24199 ( .A(keyinput32), .ZN(n21281) );
  OAI22_X1 U24200 ( .A1(n21282), .A2(keyinput71), .B1(n21281), .B2(
        P3_DATAO_REG_31__SCAN_IN), .ZN(n21280) );
  AOI221_X1 U24201 ( .B1(n21282), .B2(keyinput71), .C1(
        P3_DATAO_REG_31__SCAN_IN), .C2(n21281), .A(n21280), .ZN(n21283) );
  NAND4_X1 U24202 ( .A1(n21286), .A2(n21285), .A3(n21284), .A4(n21283), .ZN(
        n21334) );
  OAI22_X1 U24203 ( .A1(n11440), .A2(keyinput91), .B1(n21288), .B2(keyinput19), 
        .ZN(n21287) );
  AOI221_X1 U24204 ( .B1(n11440), .B2(keyinput91), .C1(keyinput19), .C2(n21288), .A(n21287), .ZN(n21301) );
  INV_X1 U24205 ( .A(keyinput57), .ZN(n21290) );
  OAI22_X1 U24206 ( .A1(keyinput25), .A2(n21291), .B1(n21290), .B2(
        P1_DATAO_REG_25__SCAN_IN), .ZN(n21289) );
  AOI221_X1 U24207 ( .B1(n21291), .B2(keyinput25), .C1(n21290), .C2(
        P1_DATAO_REG_25__SCAN_IN), .A(n21289), .ZN(n21300) );
  OAI22_X1 U24208 ( .A1(n21294), .A2(keyinput13), .B1(n21293), .B2(keyinput40), 
        .ZN(n21292) );
  AOI221_X1 U24209 ( .B1(n21294), .B2(keyinput13), .C1(keyinput40), .C2(n21293), .A(n21292), .ZN(n21299) );
  OAI22_X1 U24210 ( .A1(n21297), .A2(keyinput53), .B1(n21296), .B2(keyinput38), 
        .ZN(n21295) );
  AOI221_X1 U24211 ( .B1(n21297), .B2(keyinput53), .C1(keyinput38), .C2(n21296), .A(n21295), .ZN(n21298) );
  NAND4_X1 U24212 ( .A1(n21301), .A2(n21300), .A3(n21299), .A4(n21298), .ZN(
        n21333) );
  OAI22_X1 U24213 ( .A1(n21304), .A2(keyinput63), .B1(n21303), .B2(keyinput96), 
        .ZN(n21302) );
  AOI221_X1 U24214 ( .B1(n21304), .B2(keyinput63), .C1(keyinput96), .C2(n21303), .A(n21302), .ZN(n21316) );
  INV_X1 U24215 ( .A(keyinput56), .ZN(n21306) );
  OAI22_X1 U24216 ( .A1(n14906), .A2(keyinput106), .B1(n21306), .B2(
        P3_READREQUEST_REG_SCAN_IN), .ZN(n21305) );
  AOI221_X1 U24217 ( .B1(n14906), .B2(keyinput106), .C1(
        P3_READREQUEST_REG_SCAN_IN), .C2(n21306), .A(n21305), .ZN(n21315) );
  INV_X1 U24218 ( .A(keyinput36), .ZN(n21308) );
  OAI22_X1 U24219 ( .A1(n21309), .A2(keyinput27), .B1(n21308), .B2(
        P3_DATAO_REG_0__SCAN_IN), .ZN(n21307) );
  AOI221_X1 U24220 ( .B1(n21309), .B2(keyinput27), .C1(P3_DATAO_REG_0__SCAN_IN), .C2(n21308), .A(n21307), .ZN(n21314) );
  INV_X1 U24221 ( .A(keyinput89), .ZN(n21311) );
  OAI22_X1 U24222 ( .A1(n21312), .A2(keyinput42), .B1(n21311), .B2(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n21310) );
  AOI221_X1 U24223 ( .B1(n21312), .B2(keyinput42), .C1(
        P2_DATAWIDTH_REG_26__SCAN_IN), .C2(n21311), .A(n21310), .ZN(n21313) );
  NAND4_X1 U24224 ( .A1(n21316), .A2(n21315), .A3(n21314), .A4(n21313), .ZN(
        n21332) );
  INV_X1 U24225 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n21318) );
  OAI22_X1 U24226 ( .A1(n21318), .A2(keyinput95), .B1(n10020), .B2(keyinput120), .ZN(n21317) );
  AOI221_X1 U24227 ( .B1(n21318), .B2(keyinput95), .C1(keyinput120), .C2(
        n10020), .A(n21317), .ZN(n21330) );
  INV_X1 U24228 ( .A(keyinput110), .ZN(n21320) );
  OAI22_X1 U24229 ( .A1(keyinput26), .A2(n21321), .B1(n21320), .B2(
        P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21319) );
  AOI221_X1 U24230 ( .B1(n21321), .B2(keyinput26), .C1(n21320), .C2(
        P3_BYTEENABLE_REG_0__SCAN_IN), .A(n21319), .ZN(n21329) );
  OAI22_X1 U24231 ( .A1(n11948), .A2(keyinput122), .B1(n21323), .B2(keyinput85), .ZN(n21322) );
  AOI221_X1 U24232 ( .B1(n11948), .B2(keyinput122), .C1(keyinput85), .C2(
        n21323), .A(n21322), .ZN(n21328) );
  INV_X1 U24233 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21326) );
  INV_X1 U24234 ( .A(keyinput48), .ZN(n21325) );
  OAI22_X1 U24235 ( .A1(n21326), .A2(keyinput47), .B1(n21325), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n21324) );
  AOI221_X1 U24236 ( .B1(n21326), .B2(keyinput47), .C1(
        P1_DATAO_REG_31__SCAN_IN), .C2(n21325), .A(n21324), .ZN(n21327) );
  NAND4_X1 U24237 ( .A1(n21330), .A2(n21329), .A3(n21328), .A4(n21327), .ZN(
        n21331) );
  NOR4_X1 U24238 ( .A1(n21334), .A2(n21333), .A3(n21332), .A4(n21331), .ZN(
        n21335) );
  NAND4_X1 U24239 ( .A1(n21338), .A2(n21337), .A3(n21336), .A4(n21335), .ZN(
        n21339) );
  NOR4_X1 U24240 ( .A1(n21342), .A2(n21341), .A3(n21340), .A4(n21339), .ZN(
        n21355) );
  AOI22_X1 U24241 ( .A1(n21346), .A2(n21345), .B1(n21344), .B2(n21343), .ZN(
        n21351) );
  AOI22_X1 U24242 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21349), .B1(
        n21348), .B2(n21347), .ZN(n21350) );
  OAI211_X1 U24243 ( .C1(n21353), .C2(n21352), .A(n21351), .B(n21350), .ZN(
        n21354) );
  XOR2_X1 U24244 ( .A(n21355), .B(n21354), .Z(P2_U3090) );
  INV_X1 U11156 ( .A(n18398), .ZN(n17435) );
  CLKBUF_X1 U11153 ( .A(n10305), .Z(n9771) );
  CLKBUF_X1 U11159 ( .A(n11754), .Z(n12818) );
  CLKBUF_X1 U11173 ( .A(n11740), .Z(n12791) );
  CLKBUF_X1 U11176 ( .A(n11859), .Z(n12771) );
  CLKBUF_X1 U11177 ( .A(n11913), .Z(n11914) );
  CLKBUF_X2 U11191 ( .A(n10203), .Z(n11605) );
  CLKBUF_X1 U11202 ( .A(n10288), .Z(n9737) );
  AOI22_X1 U11204 ( .A1(n21088), .A2(keyinput35), .B1(keyinput28), .B2(n21087), 
        .ZN(n21086) );
  CLKBUF_X2 U11234 ( .A(n11814), .Z(n20261) );
  CLKBUF_X1 U11256 ( .A(n10484), .Z(n19555) );
  NOR2_X2 U11323 ( .A1(n9864), .A2(n15835), .ZN(n19698) );
  CLKBUF_X1 U11387 ( .A(n11842), .Z(n13591) );
  CLKBUF_X2 U11477 ( .A(n12358), .Z(n14841) );
  CLKBUF_X1 U11519 ( .A(n12398), .Z(n20280) );
  CLKBUF_X1 U11560 ( .A(n10111), .Z(n17210) );
  CLKBUF_X1 U11595 ( .A(n12425), .Z(n20372) );
  CLKBUF_X1 U11655 ( .A(n17628), .Z(n17634) );
  CLKBUF_X1 U11664 ( .A(n17659), .Z(n17690) );
  NOR2_X2 U12127 ( .A1(n17350), .A2(n17386), .ZN(n17366) );
  CLKBUF_X2 U12291 ( .A(n17559), .Z(n9718) );
  CLKBUF_X1 U12435 ( .A(n18973), .Z(n18967) );
  CLKBUF_X1 U12439 ( .A(n16653), .Z(n16664) );
  OR2_X1 U12469 ( .A1(n10187), .A2(n14010), .ZN(n21356) );
  CLKBUF_X1 U12471 ( .A(n19030), .Z(n18874) );
endmodule

