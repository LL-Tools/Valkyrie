

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, 
        P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, 
        P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, 
        P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, 
        P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, 
        P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, 
        P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, 
        P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, 
        P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, 
        P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, 
        P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN,
         P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN,
         P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN,
         P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN,
         P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN,
         P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN,
         P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN,
         P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN,
         P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN,
         P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN,
         P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
         P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
         P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
         P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
         P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
         P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
         P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN,
         P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN,
         P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
         P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN,
         P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
         P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
         P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
         P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
         P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
         P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
         P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
         P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
         P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
         P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
         P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
         P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
         P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
         P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
         P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
         P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
         P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
         P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
         P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
         P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
         P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
         P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
         P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
         P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN,
         P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN,
         P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
         P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN,
         P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN,
         P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN,
         P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN,
         P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN,
         P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN,
         P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN,
         P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN,
         P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN,
         P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN,
         P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN,
         P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN,
         P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN,
         P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
         P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN,
         P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN,
         P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
         P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
         P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
         P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
         P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
         P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
         P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
         P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
         P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
         P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
         P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
         P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
         P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
         P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN,
         P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN,
         P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
         P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN,
         P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN,
         P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN,
         P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN,
         P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN,
         P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN,
         P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN,
         P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN,
         P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN,
         P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN,
         P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN,
         P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN,
         P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN,
         P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN,
         P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN,
         P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN,
         P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN,
         P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032;

  INV_X2 U7265 ( .A(n15895), .ZN(n15898) );
  INV_X4 U7266 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X2 U7267 ( .A(n10054), .ZN(n10053) );
  INV_X2 U7268 ( .A(n14072), .ZN(n14038) );
  CLKBUF_X2 U7269 ( .A(n8383), .Z(n8765) );
  INV_X1 U7270 ( .A(n10680), .ZN(n7171) );
  INV_X1 U7271 ( .A(n9723), .ZN(n9893) );
  INV_X1 U7272 ( .A(n9088), .ZN(n10529) );
  CLKBUF_X3 U7273 ( .A(n10345), .Z(n10550) );
  INV_X1 U7274 ( .A(n8977), .ZN(n10755) );
  INV_X4 U7275 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14563) );
  AND2_X1 U7276 ( .A1(n13261), .A2(n13260), .ZN(n13272) );
  OAI211_X1 U7278 ( .C1(n7822), .C2(n7820), .A(n10597), .B(n7819), .ZN(n11670)
         );
  CLKBUF_X2 U7279 ( .A(n9890), .Z(n7210) );
  NOR2_X1 U7280 ( .A1(n12273), .A2(n12013), .ZN(n12349) );
  INV_X1 U7281 ( .A(n7210), .ZN(n9832) );
  CLKBUF_X2 U7282 ( .A(n8403), .Z(n10126) );
  CLKBUF_X2 U7283 ( .A(n13789), .Z(n7206) );
  NAND2_X1 U7284 ( .A1(n8495), .A2(n11279), .ZN(n8511) );
  AND2_X1 U7286 ( .A1(n14570), .A2(n8935), .ZN(n7237) );
  INV_X1 U7287 ( .A(n9722), .ZN(n9860) );
  OR2_X1 U7288 ( .A1(n11509), .A2(n14849), .ZN(n15063) );
  NAND2_X1 U7289 ( .A1(n15210), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9542) );
  OAI21_X1 U7290 ( .B1(n8107), .B2(n7814), .A(n7812), .ZN(n15053) );
  XOR2_X1 U7291 ( .A(n15436), .B(n15435), .Z(n15608) );
  AOI211_X1 U7292 ( .C1(n11423), .C2(n14102), .A(n11416), .B(n11415), .ZN(
        n11417) );
  INV_X1 U7293 ( .A(n11429), .ZN(n14190) );
  AND2_X1 U7294 ( .A1(n8238), .A2(n10344), .ZN(n7164) );
  BUF_X1 U7295 ( .A(n13789), .Z(n7165) );
  OAI211_X2 U7297 ( .C1(n8224), .C2(n7544), .A(n7543), .B(n7542), .ZN(n14706)
         );
  INV_X2 U7298 ( .A(n8918), .ZN(n8915) );
  NAND2_X2 U7299 ( .A1(n10186), .A2(n10185), .ZN(n12123) );
  NAND2_X2 U7300 ( .A1(n14162), .A2(n7417), .ZN(n14042) );
  NAND2_X2 U7301 ( .A1(n14145), .A2(n14035), .ZN(n14162) );
  NAND2_X1 U7302 ( .A1(n11299), .A2(n7245), .ZN(n7167) );
  NAND2_X2 U7303 ( .A1(n7747), .A2(n8661), .ZN(n7404) );
  INV_X2 U7304 ( .A(n8398), .ZN(n13221) );
  NOR2_X2 U7305 ( .A1(n15634), .A2(n15635), .ZN(n15633) );
  NOR2_X2 U7306 ( .A1(n11193), .A2(n15768), .ZN(n13231) );
  AOI21_X2 U7307 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(n10152) );
  AOI21_X1 U7308 ( .B1(n8175), .B2(n7215), .A(n7330), .ZN(n7524) );
  OR2_X2 U7309 ( .A1(n9543), .A2(n9537), .ZN(n9545) );
  XNOR2_X2 U7310 ( .A(n7970), .B(n9904), .ZN(n12729) );
  OR2_X2 U7311 ( .A1(n11635), .A2(n9433), .ZN(n7822) );
  XNOR2_X2 U7312 ( .A(n9542), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9552) );
  OAI22_X2 U7313 ( .A1(n14307), .A2(n9355), .B1(n7634), .B2(n14168), .ZN(
        n14290) );
  XNOR2_X2 U7314 ( .A(n14024), .B(n14025), .ZN(n14057) );
  OAI21_X2 U7315 ( .B1(n15547), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n15546), .ZN(
        n15554) );
  AOI21_X2 U7316 ( .B1(n11182), .B2(n11181), .A(n7492), .ZN(n11762) );
  INV_X2 U7317 ( .A(n8368), .ZN(n11371) );
  AND4_X2 U7318 ( .A1(n8354), .A2(n8355), .A3(n8353), .A4(n8352), .ZN(n8368)
         );
  XNOR2_X1 U7319 ( .A(n11036), .B(n7493), .ZN(n11115) );
  XNOR2_X2 U7320 ( .A(n7176), .B(n9536), .ZN(n15223) );
  NAND2_X2 U7321 ( .A1(n7177), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7176) );
  NAND2_X1 U7322 ( .A1(n13558), .A2(n13552), .ZN(n7743) );
  OR2_X2 U7324 ( .A1(n8496), .A2(n11278), .ZN(n8512) );
  BUF_X4 U7325 ( .A(n7359), .Z(n7170) );
  INV_X1 U7326 ( .A(n9757), .ZN(n7359) );
  XNOR2_X2 U7327 ( .A(n14023), .B(n7235), .ZN(n14127) );
  NAND2_X2 U7328 ( .A1(n14080), .A2(n14021), .ZN(n14023) );
  OAI22_X2 U7329 ( .A1(n11163), .A2(n11164), .B1(n11039), .B2(n11173), .ZN(
        n11182) );
  AOI22_X2 U7330 ( .A1(n11132), .A2(n11133), .B1(n7409), .B2(n11038), .ZN(
        n11163) );
  XNOR2_X2 U7331 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n15435) );
  NAND2_X1 U7332 ( .A1(n8164), .A2(n10581), .ZN(n10591) );
  NAND2_X1 U7333 ( .A1(n10106), .A2(n10266), .ZN(n10634) );
  AOI21_X1 U7334 ( .B1(n7908), .B2(n7172), .A(n7274), .ZN(n7173) );
  NAND2_X1 U7335 ( .A1(n7743), .A2(n7273), .ZN(n13529) );
  NAND2_X1 U7336 ( .A1(n7430), .A2(n8582), .ZN(n13605) );
  NAND2_X1 U7337 ( .A1(n9084), .A2(n9083), .ZN(n15831) );
  INV_X1 U7338 ( .A(n11383), .ZN(n15708) );
  NAND2_X1 U7339 ( .A1(n8345), .A2(n8344), .ZN(n8463) );
  NAND2_X1 U7340 ( .A1(n10160), .A2(n10165), .ZN(n11818) );
  INV_X2 U7341 ( .A(n12247), .ZN(n13216) );
  NAND2_X1 U7342 ( .A1(n11371), .A2(n11941), .ZN(n10157) );
  INV_X2 U7343 ( .A(n10550), .ZN(n10545) );
  INV_X1 U7344 ( .A(n10396), .ZN(n10372) );
  CLKBUF_X2 U7345 ( .A(n9195), .Z(n10534) );
  INV_X1 U7346 ( .A(n11292), .ZN(n7629) );
  AND2_X2 U7348 ( .A1(n8260), .A2(n8261), .ZN(n8383) );
  INV_X1 U7349 ( .A(n14743), .ZN(n7516) );
  CLKBUF_X2 U7350 ( .A(n10140), .Z(n7486) );
  NAND4_X1 U7351 ( .A1(n9700), .A2(n9699), .A3(n9698), .A4(n9697), .ZN(n14742)
         );
  NAND2_X2 U7352 ( .A1(n10770), .A2(n14580), .ZN(n8977) );
  NAND2_X1 U7354 ( .A1(n11042), .A2(n10801), .ZN(n10140) );
  INV_X2 U7355 ( .A(n9898), .ZN(n9721) );
  NAND2_X2 U7356 ( .A1(n12903), .A2(n13789), .ZN(n11042) );
  CLKBUF_X2 U7357 ( .A(n9723), .Z(n9882) );
  XNOR2_X1 U7358 ( .A(n8934), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8935) );
  INV_X2 U7359 ( .A(n10719), .ZN(n12485) );
  NAND2_X1 U7360 ( .A1(n8254), .A2(n8253), .ZN(n8272) );
  NAND2_X1 U7361 ( .A1(n8252), .A2(n8141), .ZN(n8801) );
  AND3_X1 U7362 ( .A1(n7624), .A2(n7623), .A3(n7622), .ZN(n9134) );
  NOR2_X1 U7363 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n8904) );
  AOI21_X1 U7364 ( .B1(n7395), .B2(n11967), .A(n10616), .ZN(n10618) );
  OAI21_X1 U7365 ( .B1(n9517), .B2(n15968), .A(n7854), .ZN(n9515) );
  MUX2_X1 U7366 ( .A(n10295), .B(n10294), .S(n11040), .Z(n10297) );
  XNOR2_X1 U7367 ( .A(n10634), .B(n10285), .ZN(n13435) );
  AND2_X1 U7368 ( .A1(n10072), .A2(n7448), .ZN(n10057) );
  NAND2_X1 U7369 ( .A1(n13457), .A2(n7752), .ZN(n10627) );
  OAI21_X1 U7370 ( .B1(n9922), .B2(n10058), .A(n9921), .ZN(n10066) );
  NAND2_X1 U7371 ( .A1(n9458), .A2(n9457), .ZN(n14302) );
  INV_X1 U7372 ( .A(n9903), .ZN(n15091) );
  AOI21_X1 U7373 ( .B1(n14883), .B2(n8234), .A(n7474), .ZN(n14863) );
  NAND2_X1 U7374 ( .A1(n8075), .A2(n7244), .ZN(n14913) );
  NAND2_X1 U7375 ( .A1(n13496), .A2(n10272), .ZN(n13480) );
  NAND2_X1 U7376 ( .A1(n14355), .A2(n9452), .ZN(n14343) );
  AOI21_X1 U7377 ( .B1(n7213), .B2(n14289), .A(n7285), .ZN(n8024) );
  OAI21_X1 U7378 ( .B1(n7412), .B2(n7174), .A(n7173), .ZN(n14883) );
  XNOR2_X1 U7379 ( .A(n13062), .B(n13060), .ZN(n13162) );
  CLKBUF_X1 U7380 ( .A(n13497), .Z(n13659) );
  INV_X1 U7381 ( .A(n7908), .ZN(n7174) );
  INV_X1 U7382 ( .A(n7403), .ZN(n7744) );
  NAND2_X1 U7383 ( .A1(n12886), .A2(n9562), .ZN(n14871) );
  NOR2_X1 U7384 ( .A1(n14928), .A2(n14929), .ZN(n7412) );
  AND2_X1 U7385 ( .A1(n7775), .A2(n7773), .ZN(n13421) );
  OR2_X1 U7386 ( .A1(n15105), .A2(n14887), .ZN(n12886) );
  NOR2_X1 U7387 ( .A1(n7774), .A2(n13418), .ZN(n7773) );
  NAND2_X1 U7388 ( .A1(n14678), .A2(n8220), .ZN(n14636) );
  NAND2_X1 U7389 ( .A1(n15016), .A2(n12868), .ZN(n15010) );
  AOI211_X1 U7390 ( .C1(n15618), .C2(n13407), .A(n13393), .B(n13392), .ZN(
        n13402) );
  NAND2_X1 U7391 ( .A1(n7402), .A2(n12883), .ZN(n15016) );
  NOR2_X1 U7392 ( .A1(n14724), .A2(n14729), .ZN(n7274) );
  OAI22_X1 U7393 ( .A1(n14968), .A2(n9599), .B1(n14699), .B2(n15154), .ZN(
        n14954) );
  NAND2_X2 U7394 ( .A1(n9564), .A2(n9563), .ZN(n15114) );
  XNOR2_X1 U7395 ( .A(n9395), .B(n9394), .ZN(n14574) );
  INV_X1 U7396 ( .A(n8231), .ZN(n7172) );
  AOI21_X1 U7397 ( .B1(n14410), .B2(n9446), .A(n7282), .ZN(n14386) );
  OAI22_X1 U7398 ( .A1(n9395), .A2(n9394), .B1(SI_28_), .B2(n9393), .ZN(n9519)
         );
  NAND2_X1 U7399 ( .A1(n13596), .A2(n8153), .ZN(n8152) );
  NAND2_X1 U7400 ( .A1(n15975), .A2(n7257), .ZN(n7543) );
  XNOR2_X1 U7401 ( .A(n12938), .B(n12937), .ZN(n15975) );
  NAND2_X1 U7402 ( .A1(n8677), .A2(n15234), .ZN(n8689) );
  AOI21_X1 U7403 ( .B1(n7189), .B2(n12882), .A(n12881), .ZN(n15027) );
  NOR2_X1 U7404 ( .A1(n14063), .A2(n7880), .ZN(n7879) );
  NAND2_X1 U7405 ( .A1(n14601), .A2(n12933), .ZN(n12938) );
  OAI21_X1 U7406 ( .B1(n8664), .B2(n8051), .A(n8050), .ZN(n8055) );
  AND2_X1 U7407 ( .A1(n15054), .A2(n12879), .ZN(n7189) );
  NAND2_X1 U7408 ( .A1(n7782), .A2(n8103), .ZN(n12420) );
  AND2_X1 U7409 ( .A1(n7566), .A2(n15555), .ZN(n15561) );
  NAND2_X1 U7410 ( .A1(n14645), .A2(n12919), .ZN(n14686) );
  NAND2_X1 U7411 ( .A1(n12630), .A2(n12629), .ZN(n12877) );
  OAI21_X1 U7412 ( .B1(n12630), .B2(n7188), .A(n7185), .ZN(n15054) );
  NAND2_X1 U7413 ( .A1(n8925), .A2(n8924), .ZN(n14500) );
  AND2_X1 U7414 ( .A1(n7911), .A2(n7186), .ZN(n7185) );
  NAND2_X1 U7415 ( .A1(n9228), .A2(n9227), .ZN(n14405) );
  INV_X1 U7416 ( .A(n7238), .ZN(n7188) );
  NAND2_X1 U7417 ( .A1(n7238), .A2(n7187), .ZN(n7186) );
  NAND2_X1 U7418 ( .A1(n12422), .A2(n12419), .ZN(n12412) );
  NOR2_X2 U7419 ( .A1(n15960), .A2(n12444), .ZN(n12597) );
  NAND2_X1 U7420 ( .A1(n12367), .A2(n12366), .ZN(n12557) );
  NAND2_X1 U7421 ( .A1(n12347), .A2(n12346), .ZN(n12409) );
  OAI21_X1 U7422 ( .B1(n12347), .B2(n7184), .A(n7181), .ZN(n12422) );
  NAND2_X1 U7423 ( .A1(n15536), .A2(n15537), .ZN(n15545) );
  NAND2_X1 U7424 ( .A1(n8619), .A2(n8618), .ZN(n8620) );
  NAND2_X1 U7425 ( .A1(n9223), .A2(n9222), .ZN(n9241) );
  INV_X1 U7426 ( .A(n12629), .ZN(n7187) );
  NAND2_X1 U7427 ( .A1(n8604), .A2(n8603), .ZN(n8619) );
  XNOR2_X1 U7428 ( .A(n7571), .B(n15534), .ZN(n15533) );
  AND2_X1 U7429 ( .A1(n7182), .A2(n12410), .ZN(n7181) );
  NAND2_X1 U7430 ( .A1(n7191), .A2(n7897), .ZN(n12007) );
  NAND2_X1 U7431 ( .A1(n7191), .A2(n7190), .ZN(n12095) );
  AND2_X1 U7432 ( .A1(n12707), .A2(n12706), .ZN(n13257) );
  NAND2_X1 U7433 ( .A1(n9786), .A2(n9785), .ZN(n15950) );
  NAND2_X1 U7434 ( .A1(n9168), .A2(n9167), .ZN(n12655) );
  AOI21_X1 U7435 ( .B1(n8104), .B2(n8105), .A(n7283), .ZN(n8103) );
  NAND2_X1 U7436 ( .A1(n12408), .A2(n7183), .ZN(n7182) );
  INV_X1 U7437 ( .A(n12346), .ZN(n7183) );
  NAND2_X1 U7438 ( .A1(n11861), .A2(n7898), .ZN(n7191) );
  INV_X1 U7439 ( .A(n12408), .ZN(n7184) );
  NAND2_X1 U7440 ( .A1(n11707), .A2(n11706), .ZN(n11861) );
  NAND2_X1 U7441 ( .A1(n12327), .A2(n12326), .ZN(n7482) );
  AND2_X1 U7442 ( .A1(n7897), .A2(n12003), .ZN(n7190) );
  NAND2_X2 U7443 ( .A1(n8964), .A2(n8963), .ZN(n11998) );
  NAND2_X1 U7444 ( .A1(n8567), .A2(n8566), .ZN(n8570) );
  XNOR2_X1 U7445 ( .A(n7193), .B(n11507), .ZN(n15748) );
  NAND2_X1 U7446 ( .A1(n7761), .A2(n15642), .ZN(n7760) );
  AND2_X1 U7447 ( .A1(n7568), .A2(n15506), .ZN(n15511) );
  OAI21_X1 U7448 ( .B1(n7193), .B2(n11533), .A(n7192), .ZN(n11681) );
  NAND2_X1 U7449 ( .A1(n11492), .A2(n11491), .ZN(n7193) );
  AND2_X1 U7450 ( .A1(n15640), .A2(n15639), .ZN(n15643) );
  INV_X2 U7451 ( .A(n15721), .ZN(n15947) );
  NAND2_X1 U7452 ( .A1(n11836), .A2(n11489), .ZN(n11555) );
  INV_X1 U7453 ( .A(n11837), .ZN(n11834) );
  NAND2_X2 U7454 ( .A1(n9048), .A2(n9047), .ZN(n11405) );
  OR2_X1 U7455 ( .A1(n11532), .A2(n11531), .ZN(n7192) );
  AND2_X1 U7456 ( .A1(n10177), .A2(n10178), .ZN(n12233) );
  NOR2_X1 U7457 ( .A1(n9869), .A2(n14616), .ZN(n9870) );
  NAND2_X1 U7458 ( .A1(n9024), .A2(n9023), .ZN(n11336) );
  NAND2_X1 U7459 ( .A1(n8463), .A2(n8064), .ZN(n8063) );
  NAND2_X1 U7460 ( .A1(n11611), .A2(n11488), .ZN(n11838) );
  NAND2_X1 U7461 ( .A1(n9732), .A2(n8217), .ZN(n7476) );
  NAND2_X1 U7462 ( .A1(n11099), .A2(n11235), .ZN(n11227) );
  NAND2_X1 U7463 ( .A1(n10157), .A2(n10162), .ZN(n10306) );
  NAND2_X1 U7464 ( .A1(n9002), .A2(n9001), .ZN(n11383) );
  INV_X2 U7465 ( .A(n13565), .ZN(n13635) );
  AND2_X2 U7466 ( .A1(n12892), .A2(n15660), .ZN(n15667) );
  AND2_X1 U7467 ( .A1(n10341), .A2(n10340), .ZN(n8159) );
  XNOR2_X1 U7468 ( .A(n14072), .B(n11569), .ZN(n11377) );
  INV_X2 U7469 ( .A(n13103), .ZN(n13041) );
  NAND2_X1 U7470 ( .A1(n9018), .A2(n9026), .ZN(n9040) );
  AND3_X1 U7471 ( .A1(n8331), .A2(n8330), .A3(n8329), .ZN(n12132) );
  NOR2_X1 U7472 ( .A1(n9616), .A2(n9602), .ZN(n9603) );
  BUF_X2 U7473 ( .A(n10396), .Z(n7394) );
  INV_X1 U7474 ( .A(n11397), .ZN(n11569) );
  CLKBUF_X1 U7475 ( .A(n11397), .Z(n7436) );
  INV_X4 U7476 ( .A(n10550), .ZN(n10554) );
  CLKBUF_X2 U7477 ( .A(n8381), .Z(n8766) );
  OR2_X1 U7478 ( .A1(n8326), .A2(n8325), .ZN(n8294) );
  BUF_X4 U7479 ( .A(n10533), .Z(n7478) );
  NAND2_X1 U7480 ( .A1(n7178), .A2(n9709), .ZN(n9710) );
  NOR2_X1 U7481 ( .A1(n15468), .A2(n15467), .ZN(n15472) );
  INV_X1 U7482 ( .A(n9192), .ZN(n10533) );
  CLKBUF_X2 U7483 ( .A(n9000), .Z(n9195) );
  AND4_X1 U7484 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9054), .ZN(n11429)
         );
  CLKBUF_X2 U7485 ( .A(n10344), .Z(n14194) );
  AND3_X1 U7486 ( .A1(n8397), .A2(n8396), .A3(n8395), .ZN(n11443) );
  AND2_X1 U7487 ( .A1(n8977), .A2(n10806), .ZN(n9000) );
  AND2_X1 U7488 ( .A1(n7180), .A2(n7179), .ZN(n7178) );
  NAND2_X1 U7489 ( .A1(n7445), .A2(n7442), .ZN(n13784) );
  INV_X2 U7490 ( .A(n11820), .ZN(n11900) );
  INV_X2 U7491 ( .A(n10140), .ZN(n10112) );
  BUF_X2 U7492 ( .A(n7237), .Z(n9232) );
  OR2_X1 U7493 ( .A1(n9757), .A2(n10807), .ZN(n7180) );
  NAND4_X2 U7494 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(n14743)
         );
  NAND2_X1 U7495 ( .A1(n7433), .A2(n8933), .ZN(n10770) );
  AND2_X2 U7496 ( .A1(n10940), .A2(n10714), .ZN(n10680) );
  OR3_X2 U7497 ( .A1(n12906), .A2(n15228), .A3(n15231), .ZN(n10714) );
  OR2_X1 U7498 ( .A1(n9890), .A2(n8846), .ZN(n7179) );
  OR2_X1 U7499 ( .A1(n9750), .A2(n9701), .ZN(n9702) );
  NAND2_X1 U7500 ( .A1(n13777), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8259) );
  CLKBUF_X3 U7501 ( .A(n10872), .Z(n7207) );
  NAND2_X1 U7502 ( .A1(n7626), .A2(n7625), .ZN(n7433) );
  INV_X1 U7503 ( .A(n10939), .ZN(n15236) );
  NAND2_X1 U7504 ( .A1(n8256), .A2(n8255), .ZN(n13777) );
  XNOR2_X1 U7505 ( .A(n10092), .B(n10091), .ZN(n15231) );
  XNOR2_X1 U7506 ( .A(n10086), .B(n10085), .ZN(n12906) );
  INV_X1 U7507 ( .A(n9420), .ZN(n15339) );
  OR2_X1 U7508 ( .A1(n8758), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U7509 ( .A1(n9552), .A2(n15220), .ZN(n9723) );
  NOR2_X1 U7510 ( .A1(n9800), .A2(n9799), .ZN(n9798) );
  OAI21_X1 U7511 ( .B1(n10090), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10086) );
  INV_X1 U7512 ( .A(n9553), .ZN(n15220) );
  OR2_X1 U7513 ( .A1(n14562), .A2(n14563), .ZN(n8932) );
  NAND2_X1 U7514 ( .A1(n8933), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U7515 ( .A1(n7466), .A2(n7465), .ZN(n8919) );
  OR2_X1 U7516 ( .A1(n9417), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n9418) );
  XNOR2_X1 U7517 ( .A(n9902), .B(P1_IR_REG_20__SCAN_IN), .ZN(n10719) );
  NAND2_X1 U7518 ( .A1(n10090), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10092) );
  NAND2_X1 U7519 ( .A1(n8273), .A2(n8272), .ZN(n13789) );
  XOR2_X1 U7520 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(n15450), .Z(n15452) );
  NOR2_X1 U7521 ( .A1(n9763), .A2(n9676), .ZN(n9675) );
  NAND2_X2 U7522 ( .A1(n10801), .A2(P2_U3088), .ZN(n14578) );
  OAI21_X1 U7523 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(n15447), .A(n15446), .ZN(
        n15450) );
  INV_X1 U7524 ( .A(n8801), .ZN(n8254) );
  AOI21_X1 U7525 ( .B1(n8662), .B2(n8052), .A(n7337), .ZN(n8050) );
  BUF_X2 U7526 ( .A(n11062), .Z(n7498) );
  NAND2_X1 U7527 ( .A1(n7995), .A2(n7902), .ZN(n7177) );
  INV_X1 U7528 ( .A(n8052), .ZN(n8051) );
  AND4_X1 U7529 ( .A1(n8912), .A2(n8911), .A3(n8910), .A4(n9487), .ZN(n8913)
         );
  AND4_X1 U7530 ( .A1(n7294), .A2(n7896), .A3(n9905), .A4(n9912), .ZN(n7214)
         );
  AND2_X1 U7531 ( .A1(n7678), .A2(n7676), .ZN(n8850) );
  AND2_X1 U7532 ( .A1(n8975), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8364) );
  AND2_X1 U7533 ( .A1(n9538), .A2(n10088), .ZN(n8219) );
  NAND2_X1 U7534 ( .A1(n8916), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7625) );
  AND2_X2 U7535 ( .A1(n8987), .A2(n8907), .ZN(n8944) );
  AND4_X1 U7536 ( .A1(n8243), .A2(n8242), .A3(n8241), .A4(n8347), .ZN(n8244)
         );
  AND2_X1 U7537 ( .A1(n7387), .A2(n9927), .ZN(n7896) );
  AND2_X1 U7538 ( .A1(n7578), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n15436) );
  AND4_X1 U7539 ( .A1(n9640), .A2(n9638), .A3(n9651), .A4(n9634), .ZN(n9532)
         );
  AND4_X1 U7540 ( .A1(n9225), .A2(n9498), .A3(n9484), .A4(n9491), .ZN(n8910)
         );
  NAND3_X1 U7541 ( .A1(n7346), .A2(n7345), .A3(n9533), .ZN(n9692) );
  INV_X1 U7542 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9640) );
  NOR2_X1 U7543 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8905) );
  INV_X1 U7544 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9484) );
  INV_X1 U7545 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9638) );
  INV_X1 U7546 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9409) );
  INV_X1 U7547 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8274) );
  NOR2_X1 U7548 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9529) );
  NOR2_X1 U7549 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8246) );
  INV_X4 U7550 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7551 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9912) );
  INV_X1 U7552 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9911) );
  NOR2_X1 U7553 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n9905) );
  INV_X1 U7554 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9415) );
  INV_X1 U7555 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10091) );
  INV_X1 U7556 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10085) );
  CLKBUF_X1 U7557 ( .A(P2_IR_REG_8__SCAN_IN), .Z(n7469) );
  NOR2_X1 U7558 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7622) );
  NOR2_X1 U7559 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7623) );
  NOR2_X1 U7560 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7624) );
  NOR2_X1 U7561 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n9622) );
  NOR2_X1 U7562 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9636) );
  INV_X1 U7563 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10805) );
  INV_X1 U7564 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9651) );
  NOR2_X1 U7565 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n8243) );
  NOR2_X1 U7566 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8242) );
  NOR2_X1 U7567 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8241) );
  INV_X4 U7568 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X2 U7569 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8987) );
  MUX2_X1 U7570 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n7175), .S(n16001), .Z(
        P1_U3557) );
  MUX2_X1 U7571 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n7175), .S(n16005), .Z(
        P1_U3525) );
  NAND2_X1 U7572 ( .A1(n7413), .A2(n7414), .ZN(n7175) );
  NAND2_X2 U7573 ( .A1(n15223), .A2(n15227), .ZN(n9715) );
  INV_X1 U7574 ( .A(n9710), .ZN(n15670) );
  NAND2_X1 U7575 ( .A1(n11838), .A2(n11837), .ZN(n11836) );
  XNOR2_X2 U7576 ( .A(n7516), .B(n15686), .ZN(n11837) );
  NAND2_X1 U7577 ( .A1(n11502), .A2(n11612), .ZN(n11611) );
  OR2_X1 U7578 ( .A1(n12669), .A2(n11087), .ZN(n11094) );
  NAND2_X1 U7579 ( .A1(n7866), .A2(n7868), .ZN(n12317) );
  AND2_X1 U7580 ( .A1(n14568), .A2(n14573), .ZN(n9003) );
  OR2_X2 U7581 ( .A1(n12696), .A2(n12697), .ZN(n7772) );
  NAND2_X1 U7582 ( .A1(n15602), .A2(n7574), .ZN(n15490) );
  NOR2_X2 U7583 ( .A1(n15473), .A2(n15474), .ZN(n15604) );
  OAI222_X1 U7584 ( .A1(P1_U3086), .A2(n12729), .B1(n15233), .B2(n12728), .C1(
        n12727), .C2(n15224), .ZN(P1_U3334) );
  NAND2_X1 U7585 ( .A1(n14684), .A2(n7276), .ZN(n14601) );
  NOR2_X1 U7586 ( .A1(n10960), .A2(n10672), .ZN(n10999) );
  INV_X1 U7587 ( .A(n12729), .ZN(n7968) );
  NAND2_X1 U7588 ( .A1(n10441), .A2(n7194), .ZN(n7275) );
  AND2_X1 U7589 ( .A1(n10440), .A2(n7195), .ZN(n7194) );
  INV_X1 U7590 ( .A(n10445), .ZN(n7195) );
  AND2_X1 U7591 ( .A1(n7502), .A2(n8181), .ZN(n7196) );
  AND2_X1 U7592 ( .A1(n7501), .A2(n7275), .ZN(n7197) );
  INV_X1 U7593 ( .A(n12503), .ZN(n7198) );
  NAND2_X1 U7594 ( .A1(n9418), .A2(n9419), .ZN(n11087) );
  AOI211_X1 U7595 ( .C1(n11967), .C2(n11966), .A(n11965), .B(n15947), .ZN(
        n11968) );
  NAND2_X1 U7596 ( .A1(n9410), .A2(n9409), .ZN(n9497) );
  NAND3_X1 U7597 ( .A1(n9413), .A2(n9497), .A3(n9412), .ZN(n12792) );
  NAND2_X1 U7598 ( .A1(n11094), .A2(n12792), .ZN(n11096) );
  INV_X1 U7599 ( .A(n8233), .ZN(n12492) );
  XNOR2_X1 U7600 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8357) );
  NAND2_X2 U7601 ( .A1(n8708), .A2(n8707), .ZN(n13647) );
  NAND2_X1 U7602 ( .A1(n9416), .A2(n7202), .ZN(n7199) );
  AND2_X1 U7603 ( .A1(n7199), .A2(n7200), .ZN(n9419) );
  OR2_X1 U7604 ( .A1(n7201), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7200) );
  INV_X1 U7605 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7201) );
  AND2_X1 U7606 ( .A1(n9415), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U7607 ( .A1(n8977), .A2(n10801), .ZN(n9192) );
  OAI211_X2 U7608 ( .C1(n9192), .C2(n10807), .A(n8991), .B(n8990), .ZN(n11397)
         );
  AND3_X2 U7609 ( .A1(n8908), .A2(n8944), .A3(n9134), .ZN(n7203) );
  AND3_X1 U7610 ( .A1(n8908), .A2(n8944), .A3(n9134), .ZN(n7205) );
  NAND2_X1 U7611 ( .A1(n9226), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7204) );
  NAND2_X1 U7612 ( .A1(n9226), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U7613 ( .A1(n7740), .A2(n7738), .ZN(n12230) );
  AND2_X1 U7614 ( .A1(n9414), .A2(n7895), .ZN(n9410) );
  AND4_X2 U7615 ( .A1(n9561), .A2(n9560), .A3(n9559), .A4(n9558), .ZN(n14887)
         );
  NAND2_X1 U7616 ( .A1(n11684), .A2(n11683), .ZN(n11703) );
  NAND2_X4 U7617 ( .A1(n15215), .A2(n9553), .ZN(n9898) );
  INV_X1 U7618 ( .A(n7203), .ZN(n9193) );
  NAND2_X1 U7619 ( .A1(n10345), .A2(n7164), .ZN(n10346) );
  NAND2_X2 U7620 ( .A1(n9715), .A2(n10806), .ZN(n9757) );
  NAND2_X1 U7621 ( .A1(n10338), .A2(n10339), .ZN(n10353) );
  NAND4_X2 U7622 ( .A1(n9036), .A2(n9035), .A3(n9034), .A4(n9033), .ZN(n14191)
         );
  OR2_X1 U7623 ( .A1(n9398), .A2(n11474), .ZN(n9036) );
  OAI222_X1 U7624 ( .A1(P1_U3086), .A2(n15223), .B1(n15233), .B2(n15222), .C1(
        n15221), .C2(n15235), .ZN(P1_U3327) );
  OAI21_X2 U7625 ( .B1(n10383), .B2(n10382), .A(n10381), .ZN(n10390) );
  INV_X2 U7626 ( .A(n12492), .ZN(n7208) );
  INV_X8 U7627 ( .A(n7208), .ZN(n7209) );
  OR2_X1 U7628 ( .A1(n14444), .A2(n9391), .ZN(n9463) );
  OAI21_X1 U7629 ( .B1(n9206), .B2(n9207), .A(n8077), .ZN(n9222) );
  NAND2_X1 U7630 ( .A1(n7437), .A2(n8077), .ZN(n7668) );
  INV_X1 U7631 ( .A(n9191), .ZN(n7437) );
  NAND2_X1 U7632 ( .A1(n9191), .A2(n7670), .ZN(n7669) );
  NOR2_X1 U7633 ( .A1(n8079), .A2(n7671), .ZN(n7670) );
  INV_X1 U7634 ( .A(n8897), .ZN(n7671) );
  INV_X1 U7635 ( .A(n9148), .ZN(n8889) );
  NOR2_X1 U7636 ( .A1(n8142), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n8141) );
  AND2_X1 U7637 ( .A1(n8566), .A2(n8544), .ZN(n8545) );
  NAND2_X1 U7638 ( .A1(n8342), .A2(n8341), .ZN(n8345) );
  NAND2_X1 U7639 ( .A1(n8058), .A2(n8057), .ZN(n8342) );
  AND2_X1 U7640 ( .A1(n8061), .A2(n8296), .ZN(n8057) );
  INV_X1 U7641 ( .A(n8339), .ZN(n8061) );
  INV_X1 U7642 ( .A(n14274), .ZN(n7851) );
  INV_X1 U7643 ( .A(n8003), .ZN(n8002) );
  NAND2_X1 U7644 ( .A1(n9665), .A2(n9664), .ZN(n12364) );
  OAI21_X1 U7645 ( .B1(n9958), .B2(n9957), .A(n9956), .ZN(n9962) );
  AND2_X1 U7646 ( .A1(n9951), .A2(n7477), .ZN(n9958) );
  NAND2_X1 U7647 ( .A1(n7987), .A2(n9973), .ZN(n7986) );
  NAND2_X1 U7648 ( .A1(n7350), .A2(n7349), .ZN(n10001) );
  NAND2_X1 U7649 ( .A1(n8178), .A2(n8180), .ZN(n8177) );
  INV_X1 U7650 ( .A(n10496), .ZN(n8178) );
  AND2_X1 U7651 ( .A1(n10495), .A2(n10496), .ZN(n8179) );
  NAND2_X1 U7652 ( .A1(n10040), .A2(n10037), .ZN(n7961) );
  AND2_X1 U7653 ( .A1(n10039), .A2(n7963), .ZN(n7962) );
  INV_X1 U7654 ( .A(n10037), .ZN(n7963) );
  NAND2_X1 U7655 ( .A1(n7705), .A2(n7706), .ZN(n7704) );
  INV_X1 U7656 ( .A(n13180), .ZN(n7705) );
  NAND2_X1 U7657 ( .A1(n7729), .A2(n11723), .ZN(n7728) );
  INV_X1 U7658 ( .A(n13784), .ZN(n8261) );
  AND2_X1 U7659 ( .A1(n13753), .A2(n13590), .ZN(n10301) );
  OR2_X1 U7660 ( .A1(n13582), .A2(n13590), .ZN(n7406) );
  NAND2_X1 U7661 ( .A1(n8152), .A2(n8150), .ZN(n13555) );
  NOR2_X1 U7662 ( .A1(n13552), .A2(n8151), .ZN(n8150) );
  NOR2_X1 U7663 ( .A1(n14466), .A2(n14469), .ZN(n7637) );
  OR2_X1 U7664 ( .A1(n9332), .A2(n14091), .ZN(n9348) );
  NAND2_X1 U7665 ( .A1(n14402), .A2(n9238), .ZN(n14390) );
  INV_X1 U7666 ( .A(n7827), .ZN(n7826) );
  OAI21_X1 U7667 ( .B1(n7830), .B2(n7828), .A(n12434), .ZN(n7827) );
  AOI21_X1 U7668 ( .B1(n9130), .B2(n9131), .A(n7280), .ZN(n8014) );
  INV_X1 U7669 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U7670 ( .A1(n14664), .A2(n12987), .ZN(n12997) );
  NOR2_X1 U7671 ( .A1(n15009), .A2(n15031), .ZN(n7935) );
  NOR2_X1 U7672 ( .A1(n7918), .A2(n7817), .ZN(n7816) );
  INV_X1 U7673 ( .A(n12864), .ZN(n7817) );
  NOR2_X1 U7674 ( .A1(n12631), .A2(n8109), .ZN(n8106) );
  NAND2_X1 U7675 ( .A1(n7818), .A2(n11534), .ZN(n11678) );
  INV_X1 U7676 ( .A(n11528), .ZN(n7818) );
  AOI21_X1 U7677 ( .B1(n7238), .B2(n7914), .A(n7912), .ZN(n7911) );
  NAND2_X1 U7678 ( .A1(n9523), .A2(n9522), .ZN(n9889) );
  OAI21_X1 U7679 ( .B1(n9360), .B2(n9359), .A(n9358), .ZN(n9376) );
  NAND2_X1 U7680 ( .A1(n9271), .A2(n9270), .ZN(n9286) );
  OAI21_X1 U7681 ( .B1(n9241), .B2(n7682), .A(n7681), .ZN(n9271) );
  INV_X1 U7682 ( .A(n7683), .ZN(n7682) );
  NOR2_X1 U7683 ( .A1(n9239), .A2(SI_19_), .ZN(n7687) );
  INV_X1 U7684 ( .A(n8901), .ZN(n8899) );
  NAND2_X1 U7685 ( .A1(n9191), .A2(n8897), .ZN(n9206) );
  AOI21_X1 U7686 ( .B1(n9147), .B2(n8090), .A(n7297), .ZN(n8088) );
  INV_X1 U7687 ( .A(n8891), .ZN(n8093) );
  NAND2_X1 U7688 ( .A1(n8886), .A2(n8885), .ZN(n9148) );
  NAND2_X1 U7689 ( .A1(n7665), .A2(n7664), .ZN(n7663) );
  NAND2_X1 U7690 ( .A1(n8068), .A2(n7654), .ZN(n9064) );
  OAI21_X1 U7691 ( .B1(n8863), .B2(n10831), .A(n7689), .ZN(n7688) );
  NAND2_X1 U7692 ( .A1(n8863), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U7693 ( .A1(n7688), .A2(SI_5_), .ZN(n8866) );
  OAI22_X1 U7694 ( .A1(n15482), .A2(n15481), .B1(P3_ADDR_REG_6__SCAN_IN), .B2(
        n15480), .ZN(n15486) );
  BUF_X1 U7695 ( .A(n8417), .Z(n8403) );
  INV_X1 U7696 ( .A(n13066), .ZN(n7698) );
  NAND2_X1 U7697 ( .A1(n13113), .A2(n13059), .ZN(n13062) );
  NAND2_X1 U7698 ( .A1(n10147), .A2(n10146), .ZN(n10148) );
  NAND2_X1 U7699 ( .A1(n7507), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7947) );
  NAND2_X1 U7700 ( .A1(n7946), .A2(n7945), .ZN(n12155) );
  INV_X1 U7701 ( .A(n11755), .ZN(n7945) );
  XNOR2_X1 U7702 ( .A(n7508), .B(n15642), .ZN(n15634) );
  NAND2_X1 U7703 ( .A1(n13311), .A2(n13310), .ZN(n7767) );
  NAND2_X1 U7704 ( .A1(n13311), .A2(n7770), .ZN(n7769) );
  NOR2_X1 U7705 ( .A1(n7771), .A2(n13320), .ZN(n7770) );
  INV_X1 U7706 ( .A(n13607), .ZN(n13574) );
  NAND2_X1 U7707 ( .A1(n13594), .A2(n13593), .ZN(n13596) );
  INV_X1 U7708 ( .A(n10142), .ZN(n8693) );
  AOI21_X1 U7709 ( .B1(n8799), .B2(n13996), .A(n7456), .ZN(n8807) );
  AND3_X2 U7710 ( .A1(n7756), .A2(n7754), .A3(n8298), .ZN(n8252) );
  NOR2_X1 U7711 ( .A1(n8749), .A2(n7755), .ZN(n7754) );
  NAND2_X1 U7712 ( .A1(n8252), .A2(n8251), .ZN(n8795) );
  AOI21_X1 U7713 ( .B1(n8040), .B2(n8038), .A(n8037), .ZN(n8036) );
  INV_X1 U7714 ( .A(n8040), .ZN(n8039) );
  INV_X1 U7715 ( .A(n8545), .ZN(n8037) );
  INV_X1 U7716 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U7717 ( .A1(n8294), .A2(n8059), .ZN(n8058) );
  NOR2_X1 U7718 ( .A1(n8295), .A2(n8060), .ZN(n8059) );
  INV_X1 U7719 ( .A(n8293), .ZN(n8060) );
  XNOR2_X1 U7720 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8310) );
  XNOR2_X1 U7721 ( .A(n8328), .B(P3_IR_REG_7__SCAN_IN), .ZN(n15617) );
  OAI21_X1 U7722 ( .B1(n7864), .B2(n7861), .A(n7860), .ZN(n7859) );
  NOR2_X1 U7723 ( .A1(n7865), .A2(n7863), .ZN(n7861) );
  NAND2_X1 U7724 ( .A1(n7864), .A2(n14070), .ZN(n7860) );
  NAND2_X1 U7725 ( .A1(n7425), .A2(n7424), .ZN(n7608) );
  INV_X1 U7726 ( .A(n15273), .ZN(n7424) );
  NAND2_X1 U7727 ( .A1(n7608), .A2(n7607), .ZN(n7606) );
  NAND2_X1 U7728 ( .A1(n15270), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7607) );
  OR2_X1 U7729 ( .A1(n15287), .A2(n15286), .ZN(n7609) );
  OR2_X1 U7730 ( .A1(n14524), .A2(n14262), .ZN(n7652) );
  NAND2_X1 U7731 ( .A1(n14343), .A2(n9453), .ZN(n7845) );
  INV_X1 U7732 ( .A(n8010), .ZN(n8007) );
  CLKBUF_X1 U7733 ( .A(n14390), .Z(n7397) );
  NOR2_X1 U7734 ( .A1(n12671), .A2(n8021), .ZN(n8020) );
  INV_X1 U7735 ( .A(n9205), .ZN(n8021) );
  NAND2_X1 U7736 ( .A1(n9244), .A2(n9243), .ZN(n14392) );
  NAND2_X1 U7737 ( .A1(n14423), .A2(n9421), .ZN(n15964) );
  OR2_X1 U7738 ( .A1(n9493), .A2(n14584), .ZN(n9512) );
  INV_X1 U7739 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9491) );
  INV_X1 U7740 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U7741 ( .A1(n12983), .A2(n14694), .ZN(n14613) );
  NAND2_X1 U7742 ( .A1(n14620), .A2(n14622), .ZN(n14621) );
  OAI21_X1 U7743 ( .B1(n10793), .B2(n8189), .A(n8187), .ZN(n12204) );
  NAND2_X1 U7744 ( .A1(n8195), .A2(n8194), .ZN(n8189) );
  OR2_X1 U7745 ( .A1(n8191), .A2(n8188), .ZN(n8187) );
  INV_X1 U7746 ( .A(n8194), .ZN(n8188) );
  NAND2_X1 U7747 ( .A1(n7343), .A2(n10685), .ZN(n8214) );
  NAND2_X1 U7748 ( .A1(n14621), .A2(n10684), .ZN(n7343) );
  XNOR2_X1 U7749 ( .A(n9903), .B(n14855), .ZN(n10067) );
  NAND2_X1 U7750 ( .A1(n10101), .A2(n10070), .ZN(n10078) );
  AND4_X1 U7751 ( .A1(n9579), .A2(n9578), .A3(n9577), .A4(n9576), .ZN(n14888)
         );
  AND2_X1 U7752 ( .A1(n9609), .A2(n9608), .ZN(n15000) );
  OR2_X1 U7753 ( .A1(n9809), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9734) );
  NOR2_X1 U7754 ( .A1(n15396), .A2(n7536), .ZN(n14834) );
  NAND2_X1 U7755 ( .A1(n9601), .A2(n9600), .ZN(n14988) );
  NAND2_X1 U7756 ( .A1(n9813), .A2(n9812), .ZN(n15077) );
  INV_X1 U7757 ( .A(n9715), .ZN(n10872) );
  NAND2_X1 U7758 ( .A1(n9715), .A2(n10801), .ZN(n9890) );
  AND2_X1 U7759 ( .A1(n7903), .A2(n7995), .ZN(n9543) );
  OAI21_X1 U7760 ( .B1(n7688), .B2(SI_5_), .A(n8866), .ZN(n9041) );
  NOR2_X1 U7761 ( .A1(n9731), .A2(n9730), .ZN(n10993) );
  AOI21_X1 U7762 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n15519), .A(n15518), .ZN(
        n15531) );
  NOR2_X1 U7763 ( .A1(n15517), .A2(n15516), .ZN(n15518) );
  INV_X1 U7764 ( .A(n13698), .ZN(n13198) );
  AND2_X1 U7765 ( .A1(P3_U3897), .A2(n12903), .ZN(n15638) );
  OAI22_X1 U7766 ( .A1(n13072), .A2(n13627), .B1(n13427), .B2(n10630), .ZN(
        n10631) );
  OAI21_X1 U7767 ( .B1(n8763), .B2(n8762), .A(n8771), .ZN(n13443) );
  AOI21_X1 U7768 ( .B1(n7849), .B2(n7848), .A(n7847), .ZN(n7846) );
  NAND2_X1 U7769 ( .A1(n15533), .A2(n15532), .ZN(n15536) );
  INV_X1 U7770 ( .A(n10413), .ZN(n8161) );
  NAND2_X1 U7771 ( .A1(n10428), .A2(n10429), .ZN(n7393) );
  INV_X1 U7772 ( .A(n10428), .ZN(n7391) );
  OAI21_X1 U7773 ( .B1(n9962), .B2(n9961), .A(n9960), .ZN(n9964) );
  OR2_X1 U7774 ( .A1(n7987), .A2(n9973), .ZN(n7985) );
  INV_X1 U7775 ( .A(n7986), .ZN(n7357) );
  NAND2_X1 U7776 ( .A1(n7991), .A2(n9977), .ZN(n7990) );
  AND2_X1 U7777 ( .A1(n7989), .A2(n7356), .ZN(n7351) );
  INV_X1 U7778 ( .A(n9981), .ZN(n9984) );
  INV_X1 U7779 ( .A(n9989), .ZN(n7376) );
  INV_X1 U7780 ( .A(n10476), .ZN(n7459) );
  OAI21_X1 U7781 ( .B1(n10475), .B2(n10554), .A(n10474), .ZN(n10476) );
  INV_X1 U7782 ( .A(n10479), .ZN(n8173) );
  INV_X1 U7783 ( .A(n10480), .ZN(n8174) );
  NAND2_X1 U7784 ( .A1(n7977), .A2(n10004), .ZN(n7976) );
  NAND2_X1 U7785 ( .A1(n10010), .A2(n7972), .ZN(n7971) );
  INV_X1 U7786 ( .A(n10009), .ZN(n7972) );
  NAND2_X1 U7787 ( .A1(n10492), .A2(n10491), .ZN(n10497) );
  OAI21_X1 U7788 ( .B1(n10497), .B2(n8179), .A(n7517), .ZN(n10503) );
  AND2_X1 U7789 ( .A1(n8177), .A2(n7518), .ZN(n7517) );
  INV_X1 U7790 ( .A(n10502), .ZN(n7518) );
  NAND2_X1 U7791 ( .A1(n8179), .A2(n8177), .ZN(n8176) );
  NOR2_X1 U7792 ( .A1(n9599), .A2(n7288), .ZN(n7964) );
  NAND2_X1 U7793 ( .A1(n10020), .A2(n10018), .ZN(n7983) );
  OR2_X1 U7794 ( .A1(n10020), .A2(n10018), .ZN(n7982) );
  NAND2_X1 U7795 ( .A1(n10942), .A2(n7969), .ZN(n9944) );
  INV_X1 U7796 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8551) );
  AOI21_X1 U7797 ( .B1(n10522), .B2(n10521), .A(n10523), .ZN(n7472) );
  NAND2_X1 U7798 ( .A1(n8169), .A2(n10526), .ZN(n8163) );
  NAND2_X1 U7799 ( .A1(n10573), .A2(n10553), .ZN(n10576) );
  INV_X1 U7800 ( .A(n7637), .ZN(n7636) );
  AOI21_X1 U7801 ( .B1(n7683), .B2(n7684), .A(n9267), .ZN(n7681) );
  INV_X1 U7802 ( .A(n8097), .ZN(n7660) );
  AOI21_X1 U7803 ( .B1(n8097), .B2(n8098), .A(n8095), .ZN(n8094) );
  INV_X1 U7804 ( .A(n9132), .ZN(n8095) );
  NOR2_X1 U7805 ( .A1(n8942), .A2(n8100), .ZN(n8099) );
  INV_X1 U7806 ( .A(n8880), .ZN(n8100) );
  NAND2_X1 U7807 ( .A1(n7797), .A2(n8856), .ZN(n7796) );
  INV_X1 U7808 ( .A(n8993), .ZN(n8856) );
  NAND2_X1 U7809 ( .A1(n13067), .A2(n13505), .ZN(n7708) );
  AND2_X1 U7810 ( .A1(n10145), .A2(n10144), .ZN(n10318) );
  INV_X1 U7811 ( .A(n11173), .ZN(n7944) );
  AND2_X1 U7812 ( .A1(n12337), .A2(n12336), .ZN(n12688) );
  INV_X1 U7813 ( .A(n10217), .ZN(n8129) );
  NOR2_X1 U7814 ( .A1(n12540), .A2(n13213), .ZN(n7748) );
  AND2_X1 U7815 ( .A1(n8149), .A2(n10194), .ZN(n8148) );
  NAND2_X1 U7816 ( .A1(n12290), .A2(n8776), .ZN(n12387) );
  NAND2_X1 U7817 ( .A1(n12217), .A2(n15762), .ZN(n10177) );
  OR2_X1 U7818 ( .A1(n13647), .A2(n13068), .ZN(n10154) );
  NAND2_X1 U7819 ( .A1(n13555), .A2(n10245), .ZN(n13540) );
  INV_X1 U7820 ( .A(n10276), .ZN(n11040) );
  INV_X1 U7821 ( .A(n8033), .ZN(n8032) );
  OAI21_X1 U7822 ( .B1(n8691), .B2(n8034), .A(n8720), .ZN(n8033) );
  INV_X1 U7823 ( .A(n8704), .ZN(n8034) );
  INV_X1 U7824 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8251) );
  AND2_X1 U7825 ( .A1(n8244), .A2(n7264), .ZN(n7756) );
  INV_X1 U7826 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8156) );
  INV_X1 U7827 ( .A(n7894), .ZN(n7892) );
  NOR2_X1 U7828 ( .A1(n14512), .A2(n14557), .ZN(n7643) );
  NOR2_X1 U7829 ( .A1(n14500), .A2(n7642), .ZN(n7641) );
  INV_X1 U7830 ( .A(n7643), .ZN(n7642) );
  AND2_X1 U7831 ( .A1(n7833), .A2(n7251), .ZN(n7832) );
  AND2_X1 U7832 ( .A1(n11794), .A2(n7631), .ZN(n7630) );
  INV_X1 U7833 ( .A(n15918), .ZN(n7631) );
  INV_X1 U7834 ( .A(n11285), .ZN(n7999) );
  OAI22_X1 U7835 ( .A1(n7979), .A2(n7978), .B1(n10045), .B2(n7980), .ZN(n10048) );
  AOI21_X1 U7836 ( .B1(n7960), .B2(n7958), .A(n7449), .ZN(n7978) );
  NOR2_X1 U7837 ( .A1(n14821), .A2(n7533), .ZN(n14825) );
  AND2_X1 U7838 ( .A1(n14822), .A2(n14823), .ZN(n7533) );
  NAND2_X1 U7839 ( .A1(n7597), .A2(n7595), .ZN(n14852) );
  NOR2_X1 U7840 ( .A1(n15114), .A2(n7596), .ZN(n7595) );
  NAND2_X1 U7841 ( .A1(n7599), .A2(n14724), .ZN(n7596) );
  OR2_X1 U7842 ( .A1(n7244), .A2(n7172), .ZN(n7909) );
  INV_X1 U7843 ( .A(n7789), .ZN(n7787) );
  NAND2_X1 U7844 ( .A1(n15141), .A2(n14958), .ZN(n7795) );
  NAND2_X1 U7845 ( .A1(n7591), .A2(n14732), .ZN(n10034) );
  INV_X1 U7846 ( .A(n15154), .ZN(n7590) );
  AND2_X1 U7847 ( .A1(n7586), .A2(n15880), .ZN(n7585) );
  NAND2_X1 U7848 ( .A1(n10939), .A2(n12729), .ZN(n11511) );
  NAND2_X1 U7849 ( .A1(n7598), .A2(n14904), .ZN(n7808) );
  AND2_X1 U7850 ( .A1(n14886), .A2(n14868), .ZN(n14869) );
  NAND2_X1 U7851 ( .A1(n7915), .A2(n12878), .ZN(n7914) );
  INV_X1 U7852 ( .A(n12876), .ZN(n7915) );
  INV_X1 U7853 ( .A(n12878), .ZN(n7913) );
  NOR2_X1 U7854 ( .A1(n15081), .A2(n7917), .ZN(n7916) );
  INV_X1 U7855 ( .A(n12875), .ZN(n7917) );
  OR2_X1 U7856 ( .A1(n12877), .A2(n12876), .ZN(n7919) );
  NAND2_X1 U7857 ( .A1(n15236), .A2(n14849), .ZN(n10942) );
  AND2_X1 U7858 ( .A1(n10698), .A2(n10697), .ZN(n10700) );
  OAI21_X1 U7859 ( .B1(n9342), .B2(n9341), .A(n9343), .ZN(n9360) );
  INV_X1 U7860 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9927) );
  AND2_X1 U7861 ( .A1(n9915), .A2(n7308), .ZN(n7994) );
  NOR2_X1 U7862 ( .A1(n9914), .A2(n9913), .ZN(n9915) );
  INV_X1 U7863 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7386) );
  NOR2_X1 U7864 ( .A1(n7675), .A2(n7673), .ZN(n7672) );
  NOR2_X1 U7865 ( .A1(n7674), .A2(n8897), .ZN(n7673) );
  INV_X1 U7866 ( .A(n9176), .ZN(n7658) );
  INV_X1 U7867 ( .A(n8088), .ZN(n7656) );
  NAND2_X1 U7868 ( .A1(n8887), .A2(SI_13_), .ZN(n8890) );
  AOI21_X1 U7869 ( .B1(n8085), .B2(n8087), .A(n8084), .ZN(n8083) );
  INV_X1 U7870 ( .A(n8875), .ZN(n8084) );
  NAND2_X1 U7871 ( .A1(n7796), .A2(n8857), .ZN(n9015) );
  INV_X1 U7872 ( .A(n7796), .ZN(n7475) );
  NOR2_X1 U7873 ( .A1(n7704), .A2(n7220), .ZN(n7695) );
  INV_X1 U7874 ( .A(n7704), .ZN(n7697) );
  NOR2_X1 U7875 ( .A1(n13180), .A2(n7241), .ZN(n7703) );
  NOR2_X1 U7876 ( .A1(n13070), .A2(n13486), .ZN(n7702) );
  NOR2_X1 U7877 ( .A1(n7255), .A2(n7218), .ZN(n7709) );
  NOR2_X1 U7878 ( .A1(n7716), .A2(n7291), .ZN(n7715) );
  INV_X1 U7879 ( .A(n13044), .ZN(n7716) );
  NOR2_X1 U7880 ( .A1(n12805), .A2(n7723), .ZN(n7722) );
  INV_X1 U7881 ( .A(n12779), .ZN(n7723) );
  NAND2_X1 U7882 ( .A1(n7720), .A2(n7722), .ZN(n7719) );
  INV_X1 U7883 ( .A(n12774), .ZN(n7720) );
  OAI211_X1 U7884 ( .C1(n11724), .C2(n7726), .A(n7725), .B(n11905), .ZN(n12062) );
  OR2_X1 U7885 ( .A1(n7707), .A2(n13122), .ZN(n7706) );
  INV_X1 U7886 ( .A(n7708), .ZN(n7707) );
  NAND2_X1 U7887 ( .A1(n7711), .A2(n13205), .ZN(n7693) );
  NOR2_X1 U7888 ( .A1(n8056), .A2(n10317), .ZN(n10320) );
  NAND2_X1 U7889 ( .A1(n7758), .A2(n7757), .ZN(n11140) );
  OR2_X1 U7890 ( .A1(n11062), .A2(n15682), .ZN(n7758) );
  NAND2_X1 U7891 ( .A1(n7498), .A2(n15682), .ZN(n7757) );
  NAND2_X1 U7892 ( .A1(n11188), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n13237) );
  NAND2_X1 U7893 ( .A1(n11765), .A2(n11766), .ZN(n12166) );
  NAND2_X1 U7894 ( .A1(n12176), .A2(n7315), .ZN(n7759) );
  NAND2_X1 U7895 ( .A1(n7763), .A2(n15642), .ZN(n7762) );
  INV_X1 U7896 ( .A(n12175), .ZN(n7763) );
  NAND2_X1 U7897 ( .A1(n12155), .A2(n12154), .ZN(n7508) );
  XNOR2_X1 U7898 ( .A(n12688), .B(n7941), .ZN(n12338) );
  NOR2_X1 U7899 ( .A1(n12338), .A2(n12329), .ZN(n12689) );
  AND2_X1 U7900 ( .A1(n13314), .A2(n13313), .ZN(n13345) );
  INV_X1 U7901 ( .A(n7733), .ZN(n7730) );
  AOI21_X1 U7902 ( .B1(n13387), .B2(n13386), .A(n13385), .ZN(n13408) );
  NOR2_X1 U7903 ( .A1(n13388), .A2(n13389), .ZN(n13406) );
  INV_X1 U7904 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8276) );
  INV_X1 U7905 ( .A(n13382), .ZN(n7939) );
  NAND2_X1 U7906 ( .A1(n13532), .A2(n8661), .ZN(n13514) );
  AND2_X1 U7907 ( .A1(n8783), .A2(n10254), .ZN(n8155) );
  AND2_X1 U7908 ( .A1(n8628), .A2(n13971), .ZN(n8642) );
  NAND2_X1 U7909 ( .A1(n13587), .A2(n8599), .ZN(n13573) );
  NAND2_X1 U7910 ( .A1(n13605), .A2(n7741), .ZN(n13587) );
  NOR2_X1 U7911 ( .A1(n13593), .A2(n7742), .ZN(n7741) );
  INV_X1 U7912 ( .A(n8583), .ZN(n7742) );
  NAND2_X1 U7913 ( .A1(n13605), .A2(n8583), .ZN(n13585) );
  AND2_X1 U7914 ( .A1(n10229), .A2(n10232), .ZN(n13612) );
  INV_X1 U7915 ( .A(n13209), .ZN(n13626) );
  NAND2_X1 U7916 ( .A1(n12816), .A2(n7269), .ZN(n13621) );
  AND2_X1 U7917 ( .A1(n10225), .A2(n10224), .ZN(n13631) );
  NAND2_X1 U7918 ( .A1(n12818), .A2(n12817), .ZN(n12816) );
  AND2_X1 U7919 ( .A1(n12768), .A2(n10216), .ZN(n8132) );
  NAND2_X1 U7920 ( .A1(n12542), .A2(n10202), .ZN(n12663) );
  AND2_X1 U7921 ( .A1(n12734), .A2(n10205), .ZN(n12773) );
  OAI21_X1 U7922 ( .B1(n12387), .B2(n8147), .A(n8145), .ZN(n12542) );
  INV_X1 U7923 ( .A(n8146), .ZN(n8145) );
  OAI21_X1 U7924 ( .B1(n8148), .B2(n8147), .A(n12717), .ZN(n8146) );
  INV_X1 U7925 ( .A(n10197), .ZN(n8147) );
  AND4_X1 U7926 ( .A1(n8338), .A2(n8337), .A3(n8336), .A4(n8335), .ZN(n12573)
         );
  AND4_X1 U7927 ( .A1(n8476), .A2(n8475), .A3(n8474), .A4(n8473), .ZN(n12804)
         );
  AND2_X1 U7928 ( .A1(n10202), .A2(n12778), .ZN(n12717) );
  NAND2_X1 U7929 ( .A1(n13215), .A2(n15857), .ZN(n10194) );
  NAND2_X1 U7930 ( .A1(n7411), .A2(n8148), .ZN(n12455) );
  AND3_X1 U7931 ( .A1(n8303), .A2(n8302), .A3(n8301), .ZN(n12469) );
  CLKBUF_X1 U7932 ( .A(n12387), .Z(n7411) );
  INV_X1 U7933 ( .A(n8138), .ZN(n8137) );
  OAI21_X1 U7934 ( .B1(n12215), .B2(n8139), .A(n12124), .ZN(n8138) );
  NAND2_X1 U7935 ( .A1(n8775), .A2(n10177), .ZN(n12216) );
  NAND2_X1 U7936 ( .A1(n12216), .A2(n12215), .ZN(n12214) );
  NOR2_X1 U7937 ( .A1(n12233), .A2(n7739), .ZN(n7738) );
  INV_X1 U7938 ( .A(n8416), .ZN(n7739) );
  NAND2_X1 U7939 ( .A1(n11739), .A2(n10162), .ZN(n8772) );
  AND3_X1 U7940 ( .A1(n8378), .A2(n8379), .A3(n8377), .ZN(n11365) );
  OR2_X1 U7941 ( .A1(n7486), .A2(SI_2_), .ZN(n8379) );
  NAND2_X1 U7942 ( .A1(n8739), .A2(n8738), .ZN(n10626) );
  XNOR2_X1 U7943 ( .A(n13463), .B(n13473), .ZN(n13454) );
  INV_X1 U7944 ( .A(n10259), .ZN(n8123) );
  AND2_X2 U7945 ( .A1(n10265), .A2(n10273), .ZN(n13482) );
  AND3_X1 U7946 ( .A1(n8646), .A2(n8645), .A3(n8644), .ZN(n13560) );
  NAND2_X1 U7947 ( .A1(n8660), .A2(n8781), .ZN(n13532) );
  NAND2_X1 U7948 ( .A1(n8832), .A2(n8791), .ZN(n13556) );
  NAND2_X1 U7949 ( .A1(n8152), .A2(n10300), .ZN(n13553) );
  NOR2_X1 U7950 ( .A1(n8835), .A2(n8834), .ZN(n11217) );
  NAND2_X1 U7951 ( .A1(n11307), .A2(n11040), .ZN(n13627) );
  INV_X1 U7952 ( .A(n13224), .ZN(n11738) );
  NAND2_X1 U7953 ( .A1(n8770), .A2(n11040), .ZN(n13629) );
  NOR2_X2 U7954 ( .A1(n8272), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n8256) );
  INV_X1 U7955 ( .A(n13777), .ZN(n7444) );
  NOR2_X1 U7956 ( .A1(P3_IR_REG_29__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7443) );
  NAND2_X1 U7957 ( .A1(n8737), .A2(n8736), .ZN(n10109) );
  NAND2_X1 U7958 ( .A1(n8252), .A2(n8140), .ZN(n8144) );
  INV_X1 U7959 ( .A(n8142), .ZN(n8140) );
  INV_X1 U7960 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8751) );
  INV_X1 U7961 ( .A(n8756), .ZN(n8752) );
  NAND2_X1 U7962 ( .A1(n7468), .A2(n12504), .ZN(n8621) );
  NAND2_X1 U7963 ( .A1(n8620), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U7964 ( .A1(n8601), .A2(n8600), .ZN(n8604) );
  AND2_X1 U7965 ( .A1(n8584), .A2(n8568), .ZN(n8569) );
  AOI21_X1 U7966 ( .B1(n8042), .B2(n8525), .A(n8041), .ZN(n8040) );
  INV_X1 U7967 ( .A(n8542), .ZN(n8041) );
  AND2_X1 U7968 ( .A1(n8043), .A2(n8045), .ZN(n8042) );
  INV_X1 U7969 ( .A(n8528), .ZN(n8043) );
  OR2_X1 U7970 ( .A1(n8526), .A2(n8525), .ZN(n8044) );
  NAND2_X1 U7971 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n8046), .ZN(n8045) );
  AND2_X1 U7972 ( .A1(n8482), .A2(n7317), .ZN(n8062) );
  OR2_X1 U7973 ( .A1(n8346), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U7974 ( .A1(n8291), .A2(n8290), .ZN(n8326) );
  INV_X1 U7975 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8429) );
  NAND2_X1 U7976 ( .A1(n7780), .A2(n7779), .ZN(n7956) );
  INV_X1 U7977 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7779) );
  INV_X1 U7978 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7780) );
  OR2_X1 U7979 ( .A1(n14011), .A2(n14010), .ZN(n7881) );
  AOI21_X1 U7980 ( .B1(n7879), .B2(n14137), .A(n7878), .ZN(n7877) );
  INV_X1 U7981 ( .A(n14014), .ZN(n7878) );
  OR2_X1 U7982 ( .A1(n14020), .A2(n14019), .ZN(n14021) );
  INV_X1 U7983 ( .A(n9232), .ZN(n10532) );
  NAND2_X1 U7984 ( .A1(n7169), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9056) );
  AND2_X1 U7985 ( .A1(n14199), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7618) );
  OR2_X1 U7986 ( .A1(n14213), .A2(n14212), .ZN(n7617) );
  INV_X1 U7987 ( .A(n14221), .ZN(n7605) );
  OR2_X1 U7988 ( .A1(n14235), .A2(n14234), .ZN(n7615) );
  AND2_X1 U7989 ( .A1(n7615), .A2(n7614), .ZN(n11270) );
  NAND2_X1 U7990 ( .A1(n11267), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7614) );
  NAND2_X1 U7991 ( .A1(n11270), .A2(n11269), .ZN(n11923) );
  AND2_X1 U7992 ( .A1(n15373), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7621) );
  AND2_X1 U7993 ( .A1(n12838), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7619) );
  NAND2_X1 U7994 ( .A1(n7609), .A2(n15301), .ZN(n15303) );
  NOR2_X1 U7995 ( .A1(n7648), .A2(n7653), .ZN(n7647) );
  NAND2_X1 U7996 ( .A1(n7649), .A2(n14283), .ZN(n7648) );
  INV_X1 U7997 ( .A(n7652), .ZN(n7649) );
  NOR2_X1 U7998 ( .A1(n7652), .A2(n14444), .ZN(n7646) );
  NAND2_X1 U7999 ( .A1(n9463), .A2(n9392), .ZN(n14274) );
  NAND2_X1 U8000 ( .A1(n14286), .A2(n14289), .ZN(n7852) );
  NOR3_X1 U8001 ( .A1(n14361), .A2(n14323), .A3(n7634), .ZN(n7633) );
  OAI21_X1 U8002 ( .B1(n14321), .B2(n9339), .A(n9340), .ZN(n14307) );
  AND2_X1 U8003 ( .A1(n9348), .A2(n9333), .ZN(n14324) );
  AOI21_X1 U8004 ( .B1(n7843), .B2(n7841), .A(n7840), .ZN(n7839) );
  INV_X1 U8005 ( .A(n7843), .ZN(n7842) );
  INV_X1 U8006 ( .A(n9453), .ZN(n7841) );
  AOI21_X1 U8007 ( .B1(n8006), .B2(n8004), .A(n7298), .ZN(n8003) );
  INV_X1 U8008 ( .A(n7242), .ZN(n8004) );
  XNOR2_X1 U8009 ( .A(n14540), .B(n14172), .ZN(n14357) );
  NAND2_X1 U8010 ( .A1(n14356), .A2(n14357), .ZN(n14355) );
  AND2_X1 U8011 ( .A1(n9450), .A2(n9449), .ZN(n14379) );
  NAND2_X1 U8012 ( .A1(n14386), .A2(n7423), .ZN(n9450) );
  OR2_X1 U8013 ( .A1(n14392), .A2(n9448), .ZN(n7423) );
  NOR2_X1 U8014 ( .A1(n14392), .A2(n14403), .ZN(n14391) );
  NOR2_X1 U8015 ( .A1(n8019), .A2(n14420), .ZN(n8016) );
  NAND2_X1 U8016 ( .A1(n9204), .A2(n12592), .ZN(n12590) );
  AOI21_X1 U8017 ( .B1(n7826), .B2(n7828), .A(n7284), .ZN(n7824) );
  OR2_X1 U8018 ( .A1(n12655), .A2(n12524), .ZN(n12444) );
  AOI21_X1 U8019 ( .B1(n8014), .B2(n8012), .A(n7258), .ZN(n8011) );
  NAND2_X1 U8020 ( .A1(n9438), .A2(n9437), .ZN(n12528) );
  NAND2_X1 U8021 ( .A1(n8015), .A2(n11974), .ZN(n11973) );
  INV_X1 U8022 ( .A(n7251), .ZN(n7835) );
  OR2_X1 U8023 ( .A1(n7821), .A2(n7820), .ZN(n7819) );
  INV_X1 U8024 ( .A(n11667), .ZN(n7820) );
  NAND2_X1 U8025 ( .A1(n9431), .A2(n9430), .ZN(n11635) );
  NAND2_X1 U8026 ( .A1(n11285), .A2(n11286), .ZN(n15697) );
  NAND2_X1 U8027 ( .A1(n9467), .A2(n9466), .ZN(n15797) );
  NAND2_X1 U8028 ( .A1(n10937), .A2(n7478), .ZN(n8951) );
  OR2_X1 U8029 ( .A1(n10832), .A2(n9192), .ZN(n9048) );
  NOR2_X1 U8030 ( .A1(n15241), .A2(n9510), .ZN(n9516) );
  NOR2_X1 U8031 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n8027) );
  NAND2_X1 U8032 ( .A1(n9483), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U8033 ( .A1(n9485), .A2(n9484), .ZN(n9490) );
  XNOR2_X1 U8034 ( .A(n9499), .B(n9498), .ZN(n10756) );
  CLKBUF_X1 U8035 ( .A(n9224), .Z(n8920) );
  INV_X1 U8036 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8907) );
  CLKBUF_X1 U8037 ( .A(n8987), .Z(n8997) );
  OR2_X1 U8038 ( .A1(n10791), .A2(n10738), .ZN(n10739) );
  AND2_X1 U8039 ( .A1(n12998), .A2(n12996), .ZN(n14665) );
  NAND2_X1 U8040 ( .A1(n12204), .A2(n12203), .ZN(n12257) );
  AND2_X1 U8041 ( .A1(n8206), .A2(n12963), .ZN(n8205) );
  NOR2_X1 U8042 ( .A1(n12561), .A2(n7565), .ZN(n7564) );
  INV_X1 U8043 ( .A(n8213), .ZN(n7565) );
  NAND2_X1 U8044 ( .A1(n12938), .A2(n7344), .ZN(n8224) );
  INV_X1 U8045 ( .A(n12937), .ZN(n7344) );
  NAND2_X1 U8046 ( .A1(n7299), .A2(n12952), .ZN(n7545) );
  OR2_X1 U8047 ( .A1(n16007), .A2(n8212), .ZN(n8211) );
  AND2_X1 U8048 ( .A1(n8215), .A2(n7334), .ZN(n7560) );
  AND2_X1 U8049 ( .A1(n8199), .A2(n13006), .ZN(n8198) );
  NAND2_X1 U8050 ( .A1(n7379), .A2(n10055), .ZN(n7378) );
  AND2_X1 U8051 ( .A1(n10061), .A2(n10060), .ZN(n10101) );
  NAND2_X1 U8052 ( .A1(n10059), .A2(n10081), .ZN(n10060) );
  NOR2_X1 U8053 ( .A1(n10095), .A2(n12759), .ZN(n10061) );
  INV_X1 U8054 ( .A(n10102), .ZN(n7448) );
  INV_X1 U8055 ( .A(n10105), .ZN(n7500) );
  OR2_X1 U8056 ( .A1(n9734), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9768) );
  OR2_X1 U8057 ( .A1(n10869), .A2(n10870), .ZN(n7528) );
  OR2_X1 U8058 ( .A1(n10971), .A2(n10972), .ZN(n7532) );
  AND2_X1 U8059 ( .A1(n7532), .A2(n7531), .ZN(n11458) );
  NAND2_X1 U8060 ( .A1(n11457), .A2(n11456), .ZN(n7531) );
  OR2_X1 U8061 ( .A1(n11458), .A2(n11459), .ZN(n7530) );
  XNOR2_X1 U8062 ( .A(n14825), .B(n15424), .ZN(n15421) );
  NAND2_X1 U8063 ( .A1(n15421), .A2(n16000), .ZN(n15420) );
  NAND2_X1 U8064 ( .A1(n14831), .A2(n15404), .ZN(n7535) );
  AND2_X1 U8065 ( .A1(n10720), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11494) );
  AND2_X1 U8066 ( .A1(n15114), .A2(n14904), .ZN(n7474) );
  NOR2_X1 U8067 ( .A1(n8234), .A2(n7811), .ZN(n7807) );
  NAND2_X1 U8068 ( .A1(n14899), .A2(n14900), .ZN(n14898) );
  NOR2_X1 U8069 ( .A1(n7592), .A2(n15135), .ZN(n14932) );
  AOI21_X1 U8070 ( .B1(n7789), .B2(n7791), .A(n12871), .ZN(n7786) );
  OR2_X1 U8071 ( .A1(n14964), .A2(n7787), .ZN(n7785) );
  NAND2_X1 U8072 ( .A1(n7792), .A2(n7795), .ZN(n7789) );
  NAND2_X1 U8073 ( .A1(n14939), .A2(n7249), .ZN(n7792) );
  NAND2_X1 U8074 ( .A1(n10034), .A2(n12884), .ZN(n14965) );
  NOR2_X1 U8075 ( .A1(n10028), .A2(n7799), .ZN(n7798) );
  INV_X1 U8076 ( .A(n7801), .ZN(n7799) );
  NAND2_X1 U8077 ( .A1(n15010), .A2(n14995), .ZN(n7804) );
  NOR2_X1 U8078 ( .A1(n14990), .A2(n7935), .ZN(n7934) );
  NAND2_X1 U8079 ( .A1(n7928), .A2(n12883), .ZN(n7927) );
  NAND2_X1 U8080 ( .A1(n7931), .A2(n7928), .ZN(n7936) );
  INV_X1 U8081 ( .A(n7935), .ZN(n7933) );
  NAND2_X1 U8082 ( .A1(n15027), .A2(n7928), .ZN(n7920) );
  NAND2_X1 U8083 ( .A1(n15018), .A2(n15001), .ZN(n7930) );
  NAND2_X1 U8084 ( .A1(n7932), .A2(n15026), .ZN(n7931) );
  INV_X1 U8085 ( .A(n15027), .ZN(n7932) );
  NOR2_X1 U8086 ( .A1(n15039), .A2(n8115), .ZN(n8114) );
  INV_X1 U8087 ( .A(n12866), .ZN(n8115) );
  NAND2_X1 U8088 ( .A1(n10657), .A2(n12485), .ZN(n11509) );
  AOI21_X1 U8089 ( .B1(n7813), .B2(n7816), .A(n7281), .ZN(n7812) );
  INV_X1 U8090 ( .A(n8106), .ZN(n7813) );
  INV_X1 U8091 ( .A(n7816), .ZN(n7814) );
  NAND2_X1 U8092 ( .A1(n12626), .A2(n8110), .ZN(n8109) );
  INV_X1 U8093 ( .A(n12406), .ZN(n8111) );
  OR2_X1 U8094 ( .A1(n12407), .A2(n8112), .ZN(n8107) );
  NAND2_X1 U8095 ( .A1(n8107), .A2(n8106), .ZN(n12865) );
  NAND2_X1 U8096 ( .A1(n12420), .A2(n12421), .ZN(n12407) );
  AND4_X1 U8097 ( .A1(n9660), .A2(n9659), .A3(n9658), .A4(n9657), .ZN(n12423)
         );
  OR2_X1 U8098 ( .A1(n13009), .A2(n10941), .ZN(n11508) );
  NAND2_X1 U8099 ( .A1(n12086), .A2(n12085), .ZN(n12087) );
  NAND2_X1 U8100 ( .A1(n12087), .A2(n12096), .ZN(n12354) );
  AND2_X1 U8101 ( .A1(n11854), .A2(n11859), .ZN(n7898) );
  NAND2_X1 U8102 ( .A1(n7901), .A2(n7900), .ZN(n7899) );
  NAND2_X1 U8103 ( .A1(n11678), .A2(n11677), .ZN(n11679) );
  OAI21_X1 U8104 ( .B1(n10832), .B2(n9757), .A(n9736), .ZN(n11543) );
  AND2_X1 U8105 ( .A1(n10874), .A2(n10985), .ZN(n15075) );
  INV_X1 U8106 ( .A(n15993), .ZN(n15747) );
  CLKBUF_X1 U8107 ( .A(n11509), .Z(n15731) );
  NOR2_X1 U8108 ( .A1(n15656), .A2(n15236), .ZN(n15912) );
  AND2_X1 U8109 ( .A1(n10714), .A2(n10846), .ZN(n11497) );
  XNOR2_X1 U8110 ( .A(n9889), .B(n9888), .ZN(n14567) );
  INV_X1 U8111 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U8112 ( .A1(n7384), .A2(n9927), .ZN(n10090) );
  NAND2_X1 U8113 ( .A1(n9289), .A2(n9288), .ZN(n9305) );
  NAND2_X1 U8114 ( .A1(n7680), .A2(n7683), .ZN(n9268) );
  NAND2_X1 U8115 ( .A1(n8896), .A2(n8895), .ZN(n9191) );
  INV_X1 U8116 ( .A(n9189), .ZN(n8895) );
  NOR2_X1 U8117 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n9530) );
  OAI21_X1 U8118 ( .B1(n8889), .B2(n8089), .A(n8088), .ZN(n9175) );
  AND2_X1 U8119 ( .A1(n9117), .A2(n9116), .ZN(n10933) );
  OR2_X1 U8120 ( .A1(n8876), .A2(SI_9_), .ZN(n7665) );
  NAND2_X1 U8121 ( .A1(n9078), .A2(n9077), .ZN(n9080) );
  NAND2_X1 U8122 ( .A1(n9064), .A2(n8869), .ZN(n9078) );
  INV_X1 U8123 ( .A(n8086), .ZN(n8085) );
  OAI21_X1 U8124 ( .B1(n9077), .B2(n8087), .A(n9094), .ZN(n8086) );
  INV_X1 U8125 ( .A(n8872), .ZN(n8087) );
  AND2_X1 U8126 ( .A1(n9042), .A2(n9026), .ZN(n8860) );
  NOR2_X1 U8127 ( .A1(n8864), .A2(n9041), .ZN(n8865) );
  OAI21_X1 U8128 ( .B1(n15604), .B2(n15603), .A(n7575), .ZN(n7574) );
  INV_X1 U8129 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7575) );
  NOR2_X1 U8130 ( .A1(n15489), .A2(n15488), .ZN(n15495) );
  OAI21_X1 U8131 ( .B1(n15504), .B2(n15505), .A(n7569), .ZN(n7568) );
  INV_X1 U8132 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7569) );
  OAI21_X1 U8133 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15542), .A(n15541), .ZN(
        n15548) );
  OAI21_X1 U8134 ( .B1(n15554), .B2(n15553), .A(n7567), .ZN(n7566) );
  INV_X1 U8135 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7567) );
  AND4_X1 U8136 ( .A1(n8441), .A2(n8440), .A3(n8439), .A4(n8438), .ZN(n12236)
         );
  OR2_X1 U8137 ( .A1(n10140), .A2(SI_3_), .ZN(n8397) );
  INV_X1 U8138 ( .A(n13487), .ZN(n13515) );
  AND4_X1 U8139 ( .A1(n8616), .A2(n8615), .A3(n8614), .A4(n8613), .ZN(n13590)
         );
  INV_X1 U8140 ( .A(n13082), .ZN(n13211) );
  AND2_X1 U8141 ( .A1(n11180), .A2(n11191), .ZN(n7492) );
  NAND2_X1 U8142 ( .A1(n7947), .A2(n7253), .ZN(n7946) );
  OR2_X1 U8143 ( .A1(n12160), .A2(n12159), .ZN(n12337) );
  INV_X1 U8144 ( .A(n7769), .ZN(n7768) );
  AOI21_X1 U8145 ( .B1(n13320), .B2(n7767), .A(n7766), .ZN(n13331) );
  OR2_X1 U8146 ( .A1(n13992), .A2(n8693), .ZN(n8695) );
  AND2_X1 U8147 ( .A1(n8533), .A2(n8532), .ZN(n13698) );
  AND3_X1 U8148 ( .A1(n8351), .A2(n8350), .A3(n8349), .ZN(n15871) );
  OAI211_X1 U8149 ( .C1(n8693), .C2(n10811), .A(n8317), .B(n8316), .ZN(n15841)
         );
  NOR2_X1 U8150 ( .A1(n13436), .A2(n10636), .ZN(n10643) );
  OR2_X1 U8151 ( .A1(n13443), .A2(n8792), .ZN(n7421) );
  NAND2_X1 U8152 ( .A1(n8625), .A2(n8624), .ZN(n13746) );
  AND2_X1 U8153 ( .A1(n8555), .A2(n8554), .ZN(n13768) );
  OR2_X1 U8154 ( .A1(n15895), .A2(n15886), .ZN(n13767) );
  AOI21_X1 U8155 ( .B1(n8807), .B2(n8803), .A(n7289), .ZN(n13773) );
  AND2_X1 U8156 ( .A1(n11200), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13772) );
  INV_X1 U8157 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8269) );
  NAND2_X1 U8158 ( .A1(n8272), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8270) );
  MUX2_X1 U8159 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8271), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n8273) );
  OAI21_X1 U8160 ( .B1(n8547), .B2(n7731), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8607) );
  NAND2_X1 U8161 ( .A1(n7733), .A2(n7732), .ZN(n7731) );
  NAND2_X1 U8162 ( .A1(n9363), .A2(n9362), .ZN(n14448) );
  NOR2_X1 U8163 ( .A1(n12648), .A2(n12649), .ZN(n12747) );
  NAND2_X1 U8164 ( .A1(n7870), .A2(n7254), .ZN(n7869) );
  NAND2_X1 U8165 ( .A1(n11385), .A2(n7888), .ZN(n11110) );
  NAND2_X1 U8166 ( .A1(n7859), .A2(n7862), .ZN(n7858) );
  OR2_X1 U8167 ( .A1(n7864), .A2(n7863), .ZN(n7862) );
  AOI21_X1 U8168 ( .B1(n7228), .B2(n7859), .A(n14163), .ZN(n7857) );
  NAND2_X1 U8169 ( .A1(n7419), .A2(n7418), .ZN(n7417) );
  INV_X1 U8170 ( .A(n14037), .ZN(n7418) );
  INV_X1 U8171 ( .A(n14036), .ZN(n7419) );
  XNOR2_X1 U8172 ( .A(n11098), .B(n11377), .ZN(n11235) );
  NOR2_X1 U8173 ( .A1(n11406), .A2(n11407), .ZN(n11423) );
  NAND2_X1 U8174 ( .A1(n7884), .A2(n7883), .ZN(n11406) );
  NAND3_X1 U8175 ( .A1(n7886), .A2(n11385), .A3(n7248), .ZN(n7883) );
  AND2_X1 U8176 ( .A1(n11108), .A2(n11092), .ZN(n14095) );
  INV_X1 U8177 ( .A(n12792), .ZN(n10621) );
  AND2_X1 U8178 ( .A1(n7617), .A2(n7616), .ZN(n10769) );
  NAND2_X1 U8179 ( .A1(n14210), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7616) );
  OR2_X1 U8180 ( .A1(n14254), .A2(n14253), .ZN(n14439) );
  NOR2_X1 U8181 ( .A1(n14276), .A2(n7652), .ZN(n14254) );
  NAND2_X1 U8182 ( .A1(n7845), .A2(n9454), .ZN(n14331) );
  NAND2_X1 U8183 ( .A1(n8008), .A2(n8010), .ZN(n14371) );
  NAND2_X1 U8184 ( .A1(n8009), .A2(n7242), .ZN(n8008) );
  INV_X1 U8185 ( .A(n7397), .ZN(n8009) );
  OR2_X1 U8186 ( .A1(n10857), .A2(n9192), .ZN(n9102) );
  NAND2_X1 U8187 ( .A1(n9397), .A2(n9396), .ZN(n14262) );
  AND2_X1 U8188 ( .A1(n15970), .A2(n15959), .ZN(n14510) );
  NAND2_X1 U8189 ( .A1(n9479), .A2(n7853), .ZN(n9517) );
  NAND2_X1 U8190 ( .A1(n14264), .A2(n9478), .ZN(n7691) );
  AND2_X1 U8191 ( .A1(n14266), .A2(n15964), .ZN(n7692) );
  INV_X1 U8192 ( .A(n14376), .ZN(n14545) );
  OR2_X1 U8193 ( .A1(n10925), .A2(n9192), .ZN(n8964) );
  OAI21_X1 U8194 ( .B1(n9512), .B2(P2_D_REG_0__SCAN_IN), .A(n9511), .ZN(n15249) );
  INV_X1 U8195 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10924) );
  INV_X1 U8196 ( .A(n12364), .ZN(n15880) );
  NAND2_X1 U8197 ( .A1(n8209), .A2(n12956), .ZN(n14630) );
  NAND2_X1 U8198 ( .A1(n14706), .A2(n14705), .ZN(n8209) );
  NAND2_X1 U8199 ( .A1(n8102), .A2(n9613), .ZN(n15170) );
  NOR2_X1 U8200 ( .A1(n7219), .A2(n16022), .ZN(n7547) );
  NAND2_X1 U8201 ( .A1(n7550), .A2(n7553), .ZN(n7549) );
  NAND2_X1 U8202 ( .A1(n14595), .A2(n13029), .ZN(n7553) );
  NAND2_X1 U8203 ( .A1(n9825), .A2(n9824), .ZN(n16026) );
  NAND2_X1 U8204 ( .A1(n14636), .A2(n12976), .ZN(n14697) );
  AND2_X1 U8205 ( .A1(n15237), .A2(n9715), .ZN(n14959) );
  AND4_X1 U8206 ( .A1(n9671), .A2(n9670), .A3(n9669), .A4(n9668), .ZN(n12362)
         );
  NAND2_X1 U8207 ( .A1(n10988), .A2(n10989), .ZN(n10987) );
  NAND2_X1 U8208 ( .A1(n14790), .A2(n14789), .ZN(n14788) );
  OAI22_X1 U8209 ( .A1(n14845), .A2(n15397), .B1(n14846), .B2(n15413), .ZN(
        n7540) );
  NAND2_X1 U8210 ( .A1(n9674), .A2(n9673), .ZN(n12273) );
  AOI21_X1 U8211 ( .B1(n7207), .B2(n10993), .A(n8218), .ZN(n8217) );
  NAND2_X1 U8212 ( .A1(n10804), .A2(n7170), .ZN(n9732) );
  AND2_X1 U8213 ( .A1(n9715), .A2(n7582), .ZN(n8218) );
  INV_X1 U8214 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10923) );
  NAND2_X1 U8215 ( .A1(n7577), .A2(n7576), .ZN(n15437) );
  NAND2_X1 U8216 ( .A1(n15432), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n7576) );
  INV_X1 U8217 ( .A(n15436), .ZN(n7577) );
  INV_X1 U8218 ( .A(n7571), .ZN(n15535) );
  NAND2_X1 U8219 ( .A1(n15580), .A2(n7570), .ZN(n15581) );
  OAI21_X1 U8220 ( .B1(n15579), .B2(n15578), .A(n15299), .ZN(n7570) );
  NOR2_X1 U8221 ( .A1(n15581), .A2(n15582), .ZN(n15584) );
  OR2_X1 U8222 ( .A1(n11094), .A2(n11292), .ZN(n8238) );
  NAND2_X1 U8223 ( .A1(n7236), .A2(n8182), .ZN(n8181) );
  MUX2_X1 U8224 ( .A(n10660), .B(n9710), .S(n10054), .Z(n9954) );
  NAND2_X1 U8225 ( .A1(n8162), .A2(n8161), .ZN(n8160) );
  INV_X1 U8226 ( .A(n10412), .ZN(n8162) );
  NAND2_X1 U8227 ( .A1(n7391), .A2(n7390), .ZN(n7389) );
  INV_X1 U8228 ( .A(n10429), .ZN(n7390) );
  NAND2_X1 U8229 ( .A1(n7369), .A2(n7368), .ZN(n9970) );
  OR2_X1 U8230 ( .A1(n9965), .A2(n7957), .ZN(n7370) );
  OR2_X1 U8231 ( .A1(n7991), .A2(n9977), .ZN(n7989) );
  NAND2_X1 U8232 ( .A1(n9975), .A2(n7355), .ZN(n7356) );
  NAND2_X1 U8233 ( .A1(n7984), .A2(n7353), .ZN(n7352) );
  NAND2_X1 U8234 ( .A1(n7354), .A2(n7286), .ZN(n7353) );
  NAND2_X1 U8235 ( .A1(n7355), .A2(n7986), .ZN(n7354) );
  INV_X1 U8236 ( .A(n10451), .ZN(n7520) );
  NAND2_X1 U8237 ( .A1(n9986), .A2(n9985), .ZN(n9988) );
  AND2_X1 U8238 ( .A1(n7992), .A2(n7374), .ZN(n7373) );
  NAND2_X1 U8239 ( .A1(n9991), .A2(n7993), .ZN(n7992) );
  NAND2_X1 U8240 ( .A1(n9987), .A2(n7376), .ZN(n7374) );
  NAND2_X1 U8241 ( .A1(n7372), .A2(n7371), .ZN(n9995) );
  AOI21_X1 U8242 ( .B1(n7373), .B2(n7375), .A(n7212), .ZN(n7371) );
  NAND2_X1 U8243 ( .A1(n9988), .A2(n7373), .ZN(n7372) );
  NOR2_X1 U8244 ( .A1(n9987), .A2(n7376), .ZN(n7375) );
  NAND2_X1 U8245 ( .A1(n8174), .A2(n8173), .ZN(n8172) );
  OAI21_X1 U8246 ( .B1(n10473), .B2(n10472), .A(n7293), .ZN(n8171) );
  NAND2_X1 U8247 ( .A1(n7348), .A2(n7347), .ZN(n10003) );
  INV_X1 U8248 ( .A(n10002), .ZN(n7347) );
  NAND2_X1 U8249 ( .A1(n10005), .A2(n7975), .ZN(n7974) );
  INV_X1 U8250 ( .A(n10004), .ZN(n7975) );
  NAND2_X1 U8251 ( .A1(n7360), .A2(n7973), .ZN(n10014) );
  NAND2_X1 U8252 ( .A1(n10011), .A2(n10009), .ZN(n7973) );
  NAND2_X1 U8253 ( .A1(n7243), .A2(n8184), .ZN(n8183) );
  OR2_X1 U8254 ( .A1(n10512), .A2(n10511), .ZN(n8239) );
  OAI21_X1 U8255 ( .B1(n10026), .B2(n7211), .A(n7363), .ZN(n7366) );
  NOR2_X1 U8256 ( .A1(n7364), .A2(n7367), .ZN(n7363) );
  NOR2_X1 U8257 ( .A1(n7211), .A2(n10025), .ZN(n7364) );
  INV_X1 U8258 ( .A(n7956), .ZN(n8375) );
  NOR2_X1 U8259 ( .A1(n8674), .A2(n8053), .ZN(n8052) );
  INV_X1 U8260 ( .A(n8665), .ZN(n8053) );
  AOI21_X1 U8261 ( .B1(n7962), .B2(n7961), .A(n7959), .ZN(n7958) );
  INV_X1 U8262 ( .A(n10041), .ZN(n7449) );
  OAI21_X1 U8263 ( .B1(n10038), .B2(n7962), .A(n7292), .ZN(n10043) );
  NAND2_X1 U8264 ( .A1(n9944), .A2(n10719), .ZN(n7967) );
  NOR2_X1 U8265 ( .A1(n15105), .A2(n9939), .ZN(n7599) );
  OR2_X1 U8266 ( .A1(n15231), .A2(P1_B_REG_SCAN_IN), .ZN(n10696) );
  INV_X1 U8267 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U8268 ( .A1(n8078), .A2(n8080), .B1(n9207), .B2(n8077), .ZN(n8076)
         );
  NOR2_X1 U8269 ( .A1(n9164), .A2(n8091), .ZN(n8090) );
  INV_X1 U8270 ( .A(n8890), .ZN(n8091) );
  OAI21_X1 U8271 ( .B1(n10801), .B2(n7462), .A(n7461), .ZN(n8867) );
  NAND2_X1 U8272 ( .A1(n10801), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7461) );
  NOR2_X1 U8273 ( .A1(n8073), .A2(n8072), .ZN(n8069) );
  INV_X1 U8274 ( .A(n8860), .ZN(n8073) );
  INV_X1 U8275 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15447) );
  AND3_X1 U8276 ( .A1(n10156), .A2(n13104), .A3(n13454), .ZN(n10299) );
  AND2_X1 U8277 ( .A1(n13233), .A2(n7781), .ZN(n11770) );
  NAND2_X1 U8278 ( .A1(n11769), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7781) );
  NAND2_X1 U8279 ( .A1(n13314), .A2(n7952), .ZN(n7951) );
  NOR2_X1 U8280 ( .A1(n7953), .A2(n13320), .ZN(n7952) );
  AOI21_X1 U8281 ( .B1(n13314), .B2(n13313), .A(n13346), .ZN(n7954) );
  AOI21_X1 U8282 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n13365), .A(n13361), .ZN(
        n13394) );
  INV_X1 U8283 ( .A(n13399), .ZN(n7778) );
  INV_X1 U8284 ( .A(n10181), .ZN(n8139) );
  NOR2_X1 U8285 ( .A1(n8139), .A2(n8136), .ZN(n8135) );
  INV_X1 U8286 ( .A(n10177), .ZN(n8136) );
  NAND2_X1 U8287 ( .A1(n8766), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8322) );
  INV_X1 U8288 ( .A(n12074), .ZN(n12069) );
  NAND2_X1 U8289 ( .A1(n13222), .A2(n15678), .ZN(n10160) );
  INV_X1 U8290 ( .A(n8126), .ZN(n8125) );
  OAI21_X1 U8291 ( .B1(n13482), .B2(n8127), .A(n10154), .ZN(n8126) );
  NOR2_X1 U8292 ( .A1(n10301), .A2(n8154), .ZN(n8153) );
  INV_X1 U8293 ( .A(n10235), .ZN(n8154) );
  NAND2_X1 U8294 ( .A1(n8251), .A2(n8143), .ZN(n8142) );
  INV_X1 U8295 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8143) );
  NOR2_X1 U8296 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n8250) );
  INV_X1 U8297 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8249) );
  INV_X1 U8298 ( .A(n8042), .ZN(n8038) );
  INV_X1 U8299 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8245) );
  OR2_X1 U8300 ( .A1(n8444), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U8301 ( .A1(n12851), .A2(n12850), .ZN(n7894) );
  OR2_X1 U8302 ( .A1(n7198), .A2(n15339), .ZN(n10537) );
  NOR2_X1 U8303 ( .A1(n10576), .A2(n10558), .ZN(n8167) );
  OR2_X1 U8304 ( .A1(n15325), .A2(n15324), .ZN(n15327) );
  INV_X1 U8305 ( .A(n9455), .ZN(n7840) );
  OR2_X1 U8306 ( .A1(n9312), .A2(n9311), .ZN(n9332) );
  AND2_X1 U8307 ( .A1(n9455), .A2(n9320), .ZN(n10607) );
  AND2_X1 U8308 ( .A1(n8001), .A2(n7690), .ZN(n7480) );
  INV_X1 U8309 ( .A(n14357), .ZN(n7690) );
  NAND2_X1 U8310 ( .A1(n8003), .A2(n8005), .ZN(n8001) );
  NAND2_X1 U8311 ( .A1(n8929), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9214) );
  INV_X1 U8312 ( .A(n9212), .ZN(n8929) );
  NOR2_X1 U8313 ( .A1(n9169), .A2(n12651), .ZN(n7388) );
  INV_X1 U8314 ( .A(n7829), .ZN(n7828) );
  NOR2_X1 U8315 ( .A1(n9441), .A2(n7831), .ZN(n7830) );
  INV_X1 U8316 ( .A(n9439), .ZN(n7831) );
  OR2_X1 U8317 ( .A1(n12655), .A2(n12642), .ZN(n7829) );
  INV_X1 U8318 ( .A(n9131), .ZN(n8012) );
  AND2_X1 U8319 ( .A1(n11656), .A2(n9432), .ZN(n7821) );
  INV_X1 U8320 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9103) );
  AND2_X1 U8321 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n9032) );
  NOR2_X1 U8322 ( .A1(n11473), .A2(n11470), .ZN(n11026) );
  NOR2_X1 U8323 ( .A1(n7636), .A2(n7265), .ZN(n14322) );
  NAND2_X1 U8324 ( .A1(n12597), .A2(n12863), .ZN(n12678) );
  NAND2_X1 U8325 ( .A1(n15708), .A2(n15695), .ZN(n15694) );
  OR2_X1 U8326 ( .A1(n9028), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9045) );
  AND2_X1 U8327 ( .A1(n7555), .A2(n7558), .ZN(n7554) );
  NAND2_X1 U8328 ( .A1(n14595), .A2(n7556), .ZN(n7555) );
  NAND2_X1 U8329 ( .A1(n12191), .A2(n12192), .ZN(n8194) );
  AND2_X1 U8330 ( .A1(n12193), .A2(n8192), .ZN(n8191) );
  NAND2_X1 U8331 ( .A1(n8193), .A2(n8195), .ZN(n8192) );
  INV_X1 U8332 ( .A(n10739), .ZN(n8193) );
  NOR2_X1 U8333 ( .A1(n8208), .A2(n8204), .ZN(n8203) );
  INV_X1 U8334 ( .A(n14629), .ZN(n8208) );
  INV_X1 U8335 ( .A(n14705), .ZN(n8204) );
  NAND2_X1 U8336 ( .A1(n14629), .A2(n8207), .ZN(n8206) );
  INV_X1 U8337 ( .A(n12956), .ZN(n8207) );
  INV_X1 U8338 ( .A(n12729), .ZN(n9945) );
  INV_X1 U8339 ( .A(n9850), .ZN(n9575) );
  NOR2_X1 U8340 ( .A1(n8201), .A2(n8197), .ZN(n8196) );
  INV_X1 U8341 ( .A(n14665), .ZN(n8197) );
  INV_X1 U8342 ( .A(n14656), .ZN(n8201) );
  NAND2_X1 U8343 ( .A1(n14656), .A2(n8200), .ZN(n8199) );
  INV_X1 U8344 ( .A(n12998), .ZN(n8200) );
  NAND2_X1 U8345 ( .A1(n15161), .A2(n14733), .ZN(n7938) );
  INV_X1 U8346 ( .A(n7938), .ZN(n7924) );
  AOI21_X1 U8347 ( .B1(n12097), .B2(n12353), .A(n7259), .ZN(n8104) );
  AND2_X1 U8348 ( .A1(n7232), .A2(n11541), .ZN(n11867) );
  NOR2_X1 U8349 ( .A1(n11531), .A2(n11559), .ZN(n11541) );
  AND2_X1 U8350 ( .A1(n12485), .A2(n12404), .ZN(n10715) );
  NAND2_X1 U8351 ( .A1(n11541), .A2(n7216), .ZN(n11715) );
  NAND2_X1 U8352 ( .A1(n9379), .A2(n9378), .ZN(n9395) );
  NAND2_X1 U8353 ( .A1(n9308), .A2(n9307), .ZN(n9323) );
  AOI21_X1 U8354 ( .B1(n9240), .B2(n7686), .A(n7329), .ZN(n7683) );
  INV_X1 U8355 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U8356 ( .A1(n8894), .A2(SI_16_), .ZN(n8897) );
  AOI21_X1 U8357 ( .B1(n8099), .B2(n8879), .A(n7290), .ZN(n8097) );
  INV_X1 U8358 ( .A(n8099), .ZN(n8098) );
  INV_X1 U8359 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7346) );
  OAI21_X1 U8360 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n15510), .A(n15509), .ZN(
        n15517) );
  AOI22_X1 U8361 ( .A1(n15531), .A2(n15530), .B1(P1_ADDR_REG_11__SCAN_IN), 
        .B2(n15529), .ZN(n15539) );
  OAI21_X1 U8362 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15571), .A(n15570), .ZN(
        n15574) );
  XNOR2_X1 U8363 ( .A(n11443), .B(n13041), .ZN(n11722) );
  NAND2_X1 U8364 ( .A1(n12775), .A2(n12774), .ZN(n7724) );
  INV_X1 U8365 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13961) );
  INV_X1 U8366 ( .A(n7728), .ZN(n7727) );
  NAND2_X1 U8367 ( .A1(n7724), .A2(n7722), .ZN(n12809) );
  INV_X1 U8368 ( .A(n10318), .ZN(n10147) );
  AND4_X2 U8369 ( .A1(n8309), .A2(n8308), .A3(n8307), .A4(n8306), .ZN(n12247)
         );
  OR2_X1 U8370 ( .A1(n11117), .A2(n11116), .ZN(n11119) );
  OR2_X1 U8371 ( .A1(n11121), .A2(n11748), .ZN(n11123) );
  OAI21_X1 U8372 ( .B1(n7165), .B2(n11116), .A(n7494), .ZN(n11036) );
  NAND2_X1 U8373 ( .A1(n13789), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U8374 ( .A1(n11139), .A2(n11140), .ZN(n11138) );
  XNOR2_X1 U8375 ( .A(n11770), .B(n15617), .ZN(n15622) );
  NOR2_X1 U8376 ( .A1(n15622), .A2(n15822), .ZN(n15621) );
  AOI21_X1 U8377 ( .B1(n12169), .B2(n12168), .A(n12167), .ZN(n15639) );
  AND2_X1 U8378 ( .A1(n7765), .A2(n7764), .ZN(n12182) );
  AND2_X1 U8379 ( .A1(n12176), .A2(n12175), .ZN(n12177) );
  NAND2_X1 U8380 ( .A1(n12171), .A2(n12172), .ZN(n12331) );
  AOI21_X1 U8381 ( .B1(n12702), .B2(n7941), .A(n12701), .ZN(n12707) );
  INV_X1 U8382 ( .A(n7482), .ZN(n12695) );
  OR2_X1 U8383 ( .A1(n12689), .A2(n12690), .ZN(n7948) );
  AND2_X1 U8384 ( .A1(n13249), .A2(n13253), .ZN(n13279) );
  XNOR2_X1 U8385 ( .A(n13272), .B(n13280), .ZN(n13263) );
  NOR2_X1 U8386 ( .A1(n13262), .A2(n13263), .ZN(n13273) );
  NOR2_X1 U8387 ( .A1(n13341), .A2(n7497), .ZN(n7496) );
  INV_X1 U8388 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n7497) );
  NOR2_X1 U8389 ( .A1(n13370), .A2(n13369), .ZN(n13385) );
  XNOR2_X1 U8390 ( .A(n13394), .B(n13395), .ZN(n13362) );
  NOR2_X1 U8391 ( .A1(n13362), .A2(n13363), .ZN(n13396) );
  NAND2_X1 U8392 ( .A1(n13397), .A2(n7778), .ZN(n7776) );
  INV_X1 U8393 ( .A(n7776), .ZN(n7774) );
  OR2_X1 U8394 ( .A1(n13362), .A2(n7777), .ZN(n7775) );
  NAND2_X1 U8395 ( .A1(n7778), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7777) );
  AND4_X1 U8396 ( .A1(n10130), .A2(n10129), .A3(n10128), .A4(n10127), .ZN(
        n10630) );
  NOR2_X1 U8397 ( .A1(n13104), .A2(n7753), .ZN(n7752) );
  INV_X1 U8398 ( .A(n8732), .ZN(n7753) );
  OAI21_X1 U8399 ( .B1(n7404), .B2(n8781), .A(n7296), .ZN(n7403) );
  NAND2_X1 U8400 ( .A1(n13972), .A2(n8655), .ZN(n8668) );
  INV_X1 U8401 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n13972) );
  INV_X1 U8402 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n13971) );
  OR2_X1 U8403 ( .A1(n8593), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8611) );
  INV_X1 U8404 ( .A(n13612), .ZN(n8582) );
  INV_X1 U8405 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13960) );
  AND2_X1 U8406 ( .A1(n8556), .A2(n13961), .ZN(n8576) );
  NAND2_X1 U8407 ( .A1(n8576), .A2(n13960), .ZN(n8593) );
  AOI21_X1 U8408 ( .B1(n8132), .B2(n8130), .A(n8129), .ZN(n8128) );
  INV_X1 U8409 ( .A(n8132), .ZN(n8131) );
  INV_X1 U8410 ( .A(n8778), .ZN(n8130) );
  INV_X1 U8411 ( .A(n12817), .ZN(n12822) );
  OR2_X1 U8412 ( .A1(n8456), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8471) );
  INV_X1 U8413 ( .A(n12773), .ZN(n7749) );
  INV_X1 U8414 ( .A(n7454), .ZN(n12391) );
  NOR2_X1 U8415 ( .A1(n8437), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8318) );
  INV_X1 U8416 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n13857) );
  AND2_X1 U8417 ( .A1(n8318), .A2(n13857), .ZN(n8305) );
  OR2_X1 U8418 ( .A1(n8435), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8437) );
  CLKBUF_X1 U8419 ( .A(n11823), .Z(n11824) );
  AND2_X1 U8420 ( .A1(n12140), .A2(n12141), .ZN(n8400) );
  INV_X1 U8421 ( .A(n11818), .ZN(n8773) );
  NOR2_X1 U8422 ( .A1(n11220), .A2(n15886), .ZN(n11314) );
  NOR2_X1 U8423 ( .A1(n8120), .A2(n8118), .ZN(n8117) );
  INV_X1 U8424 ( .A(n13629), .ZN(n13606) );
  NAND2_X1 U8425 ( .A1(n13530), .A2(n8647), .ZN(n13542) );
  NAND2_X1 U8426 ( .A1(n7743), .A2(n8633), .ZN(n13543) );
  AND2_X1 U8427 ( .A1(n8501), .A2(n8500), .ZN(n8509) );
  NAND2_X1 U8428 ( .A1(n7740), .A2(n8416), .ZN(n12232) );
  NAND2_X1 U8429 ( .A1(n13772), .A2(n11201), .ZN(n11220) );
  INV_X1 U8430 ( .A(n13556), .ZN(n15764) );
  CLKBUF_X1 U8431 ( .A(n8399), .Z(n7398) );
  NAND2_X1 U8432 ( .A1(n12119), .A2(n11900), .ZN(n15886) );
  INV_X1 U8433 ( .A(n8807), .ZN(n10860) );
  NAND2_X1 U8434 ( .A1(n10111), .A2(n10110), .ZN(n10117) );
  NAND2_X1 U8435 ( .A1(n8031), .A2(n8029), .ZN(n8735) );
  AOI21_X1 U8436 ( .B1(n8032), .B2(n8034), .A(n8030), .ZN(n8029) );
  INV_X1 U8437 ( .A(n8722), .ZN(n8030) );
  XNOR2_X1 U8438 ( .A(n8823), .B(n8822), .ZN(n11200) );
  OAI21_X1 U8439 ( .B1(n8821), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8823) );
  AND2_X1 U8440 ( .A1(n8649), .A2(n8636), .ZN(n8637) );
  OR2_X1 U8441 ( .A1(n8750), .A2(n8749), .ZN(n8756) );
  AND2_X1 U8442 ( .A1(n7250), .A2(n7736), .ZN(n7733) );
  INV_X1 U8443 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7736) );
  INV_X1 U8444 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7732) );
  AND2_X1 U8445 ( .A1(n8600), .A2(n8586), .ZN(n8587) );
  NOR2_X1 U8446 ( .A1(n8547), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8552) );
  INV_X1 U8447 ( .A(n8547), .ZN(n7734) );
  OR2_X1 U8448 ( .A1(n8750), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U8449 ( .A1(n7756), .A2(n8299), .ZN(n8750) );
  AND2_X1 U8450 ( .A1(n8299), .A2(n8244), .ZN(n8485) );
  NOR2_X1 U8451 ( .A1(n8478), .A2(n8065), .ZN(n8064) );
  INV_X1 U8452 ( .A(n8462), .ZN(n8065) );
  INV_X1 U8453 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n8480) );
  AND2_X1 U8454 ( .A1(n8493), .A2(n8481), .ZN(n8482) );
  NOR2_X1 U8455 ( .A1(n8327), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8312) );
  AND2_X1 U8456 ( .A1(n8288), .A2(n8287), .ZN(n8425) );
  BUF_X1 U8457 ( .A(n8298), .Z(n8299) );
  INV_X1 U8458 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8549) );
  INV_X1 U8459 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8158) );
  INV_X1 U8460 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n8157) );
  AND2_X1 U8461 ( .A1(n8282), .A2(n8281), .ZN(n8388) );
  NAND2_X1 U8462 ( .A1(n7956), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U8463 ( .A1(n8364), .A2(n8357), .ZN(n8356) );
  NAND2_X1 U8464 ( .A1(n11101), .A2(n7889), .ZN(n7888) );
  INV_X1 U8465 ( .A(n11103), .ZN(n7889) );
  OR2_X1 U8466 ( .A1(n14138), .A2(n14137), .ZN(n7882) );
  INV_X1 U8467 ( .A(n14070), .ZN(n7863) );
  XNOR2_X1 U8468 ( .A(n14073), .B(n14072), .ZN(n7864) );
  NAND2_X1 U8469 ( .A1(n7877), .A2(n7316), .ZN(n7875) );
  INV_X1 U8470 ( .A(n7875), .ZN(n7874) );
  OAI21_X1 U8471 ( .B1(n12648), .B2(n7891), .A(n7890), .ZN(n12854) );
  NAND2_X1 U8472 ( .A1(n7893), .A2(n7894), .ZN(n7890) );
  OR2_X1 U8473 ( .A1(n12649), .A2(n7892), .ZN(n7891) );
  NAND2_X1 U8474 ( .A1(n12745), .A2(n12852), .ZN(n7893) );
  NAND2_X1 U8475 ( .A1(n12854), .A2(n12855), .ZN(n14003) );
  INV_X1 U8476 ( .A(n7881), .ZN(n7880) );
  NAND2_X1 U8477 ( .A1(n9245), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n9260) );
  INV_X1 U8478 ( .A(n9246), .ZN(n9245) );
  OR2_X1 U8479 ( .A1(n9155), .A2(n12497), .ZN(n9169) );
  OR2_X1 U8480 ( .A1(n9274), .A2(n14131), .ZN(n9294) );
  INV_X1 U8481 ( .A(n11977), .ZN(n14153) );
  INV_X1 U8482 ( .A(n7388), .ZN(n9182) );
  AND2_X1 U8483 ( .A1(n9354), .A2(n9353), .ZN(n14000) );
  NAND4_X1 U8484 ( .A1(n8974), .A2(n8973), .A3(n8972), .A4(n8971), .ZN(n10344)
         );
  NAND2_X1 U8485 ( .A1(n7237), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U8486 ( .A1(n7422), .A2(n7325), .ZN(n7425) );
  OR2_X1 U8487 ( .A1(n11924), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7613) );
  AND2_X1 U8488 ( .A1(n12026), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7620) );
  AND2_X1 U8489 ( .A1(n15303), .A2(n15304), .ZN(n15325) );
  NOR2_X1 U8490 ( .A1(n15328), .A2(n15329), .ZN(n15338) );
  INV_X1 U8491 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8275) );
  OR2_X1 U8492 ( .A1(n14276), .A2(n14262), .ZN(n14251) );
  NAND2_X1 U8493 ( .A1(n14295), .A2(n14283), .ZN(n14276) );
  INV_X1 U8494 ( .A(n14289), .ZN(n7848) );
  INV_X1 U8495 ( .A(n9463), .ZN(n7847) );
  NOR2_X1 U8496 ( .A1(n14332), .A2(n7844), .ZN(n7843) );
  INV_X1 U8497 ( .A(n9454), .ZN(n7844) );
  NAND2_X1 U8498 ( .A1(n14380), .A2(n14379), .ZN(n14378) );
  OR2_X1 U8499 ( .A1(n14392), .A2(n14174), .ZN(n8010) );
  OR2_X1 U8500 ( .A1(n9230), .A2(n9229), .ZN(n9246) );
  NAND2_X1 U8501 ( .A1(n7838), .A2(n14176), .ZN(n7837) );
  NAND2_X1 U8502 ( .A1(n12597), .A2(n7224), .ZN(n14403) );
  NAND2_X1 U8503 ( .A1(n12597), .A2(n7641), .ZN(n14427) );
  NAND2_X1 U8504 ( .A1(n7388), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U8505 ( .A1(n7825), .A2(n7829), .ZN(n12433) );
  NAND2_X1 U8506 ( .A1(n9440), .A2(n7830), .ZN(n7825) );
  NAND2_X1 U8507 ( .A1(n7630), .A2(n7270), .ZN(n12524) );
  NAND2_X1 U8508 ( .A1(n7836), .A2(n9436), .ZN(n12510) );
  AND2_X1 U8509 ( .A1(n7630), .A2(n7217), .ZN(n12523) );
  NAND2_X1 U8510 ( .A1(n8927), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9125) );
  INV_X1 U8511 ( .A(n9123), .ZN(n8927) );
  INV_X1 U8512 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8952) );
  OR2_X1 U8513 ( .A1(n9125), .A2(n8952), .ZN(n9141) );
  NAND2_X1 U8514 ( .A1(n11794), .A2(n9480), .ZN(n11979) );
  OR2_X1 U8515 ( .A1(n9104), .A2(n9103), .ZN(n9106) );
  INV_X1 U8516 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8965) );
  OR2_X1 U8517 ( .A1(n9106), .A2(n8965), .ZN(n9123) );
  NAND2_X1 U8518 ( .A1(n7822), .A2(n7821), .ZN(n11668) );
  NOR2_X1 U8519 ( .A1(n11998), .A2(n11663), .ZN(n11794) );
  INV_X1 U8520 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9085) );
  OR2_X1 U8521 ( .A1(n9086), .A2(n9085), .ZN(n9104) );
  NOR2_X1 U8522 ( .A1(n15804), .A2(n15831), .ZN(n11651) );
  OR2_X1 U8523 ( .A1(n11027), .A2(n15801), .ZN(n15804) );
  NAND2_X1 U8524 ( .A1(n11478), .A2(n9426), .ZN(n11029) );
  NAND2_X1 U8525 ( .A1(n11469), .A2(n9037), .ZN(n11025) );
  NAND2_X1 U8526 ( .A1(n7628), .A2(n11782), .ZN(n11470) );
  INV_X1 U8527 ( .A(n15694), .ZN(n7628) );
  CLKBUF_X1 U8528 ( .A(n8233), .Z(n14360) );
  NAND2_X1 U8529 ( .A1(n15699), .A2(n9424), .ZN(n11331) );
  NOR2_X1 U8530 ( .A1(n7436), .A2(n7629), .ZN(n15695) );
  NAND2_X1 U8531 ( .A1(n9258), .A2(n9257), .ZN(n14376) );
  AND2_X1 U8532 ( .A1(n10649), .A2(n10756), .ZN(n11084) );
  INV_X1 U8533 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9487) );
  OR2_X1 U8534 ( .A1(n9497), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9482) );
  OR2_X1 U8535 ( .A1(n9151), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9177) );
  OR2_X1 U8536 ( .A1(n9081), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9098) );
  OR2_X1 U8537 ( .A1(n9098), .A2(n7469), .ZN(n9099) );
  NOR2_X1 U8538 ( .A1(n9045), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9135) );
  INV_X1 U8539 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9772) );
  INV_X1 U8540 ( .A(n9574), .ZN(n9566) );
  INV_X1 U8541 ( .A(n7554), .ZN(n7552) );
  INV_X1 U8542 ( .A(n9858), .ZN(n9851) );
  INV_X1 U8543 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9676) );
  AND2_X1 U8544 ( .A1(n12973), .A2(n12971), .ZN(n8220) );
  OR2_X1 U8545 ( .A1(n12558), .A2(n12559), .ZN(n8213) );
  XNOR2_X1 U8546 ( .A(n10673), .B(n13025), .ZN(n10676) );
  NAND2_X1 U8547 ( .A1(n9826), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9836) );
  INV_X1 U8548 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9814) );
  OR2_X1 U8549 ( .A1(n9789), .A2(n9788), .ZN(n9815) );
  OR2_X1 U8550 ( .A1(n9768), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9633) );
  INV_X1 U8551 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15510) );
  AND2_X1 U8552 ( .A1(n15420), .A2(n14826), .ZN(n15410) );
  NAND2_X1 U8553 ( .A1(n9541), .A2(n9540), .ZN(n9903) );
  AND2_X1 U8554 ( .A1(n7909), .A2(n12885), .ZN(n7908) );
  OR2_X1 U8555 ( .A1(n15114), .A2(n15121), .ZN(n7594) );
  NAND2_X1 U8556 ( .A1(n14936), .A2(n14731), .ZN(n8074) );
  NAND2_X1 U8557 ( .A1(n7784), .A2(n7783), .ZN(n14912) );
  AOI21_X1 U8558 ( .B1(n7786), .B2(n7787), .A(n7229), .ZN(n7783) );
  NOR2_X1 U8559 ( .A1(n14981), .A2(n15141), .ZN(n7588) );
  INV_X1 U8560 ( .A(n14981), .ZN(n7589) );
  AOI21_X1 U8561 ( .B1(n7803), .B2(n7937), .A(n12869), .ZN(n7801) );
  INV_X1 U8562 ( .A(n7803), .ZN(n7802) );
  NAND2_X1 U8563 ( .A1(n7922), .A2(n7921), .ZN(n14968) );
  NAND2_X1 U8564 ( .A1(n7926), .A2(n7938), .ZN(n7921) );
  NAND2_X1 U8565 ( .A1(n15027), .A2(n7923), .ZN(n7922) );
  NOR2_X1 U8566 ( .A1(n7929), .A2(n7924), .ZN(n7923) );
  AND2_X1 U8567 ( .A1(n7260), .A2(n14990), .ZN(n7803) );
  NOR2_X1 U8568 ( .A1(n15170), .A2(n15017), .ZN(n14999) );
  NAND2_X1 U8569 ( .A1(n15040), .A2(n15018), .ZN(n15017) );
  NOR2_X1 U8570 ( .A1(n15062), .A2(n16026), .ZN(n15040) );
  NOR2_X1 U8571 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  NAND2_X1 U8572 ( .A1(n15074), .A2(n15189), .ZN(n15062) );
  NOR2_X1 U8573 ( .A1(n15070), .A2(n15077), .ZN(n15074) );
  OR2_X1 U8574 ( .A1(n9667), .A2(n9655), .ZN(n9800) );
  INV_X1 U8575 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9799) );
  AND4_X1 U8576 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n14649)
         );
  AND2_X1 U8577 ( .A1(n12095), .A2(n12094), .ZN(n12098) );
  NAND2_X1 U8578 ( .A1(n12098), .A2(n12097), .ZN(n12347) );
  AOI21_X1 U8579 ( .B1(n7898), .B2(n11860), .A(n7221), .ZN(n7897) );
  OR2_X1 U8580 ( .A1(n9773), .A2(n9772), .ZN(n9775) );
  INV_X1 U8581 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9761) );
  OR2_X1 U8582 ( .A1(n9775), .A2(n9761), .ZN(n9763) );
  OR2_X1 U8583 ( .A1(n11845), .A2(n14624), .ZN(n11559) );
  NOR2_X1 U8584 ( .A1(n10806), .A2(n10833), .ZN(n7582) );
  NAND2_X1 U8585 ( .A1(n11846), .A2(n15686), .ZN(n11845) );
  INV_X1 U8586 ( .A(n15731), .ZN(n15071) );
  OR2_X1 U8587 ( .A1(n10725), .A2(n10985), .ZN(n15042) );
  NOR2_X1 U8588 ( .A1(n15101), .A2(n15100), .ZN(n15102) );
  NAND2_X1 U8589 ( .A1(n7809), .A2(n7806), .ZN(n15106) );
  AND2_X1 U8590 ( .A1(n14871), .A2(n7808), .ZN(n7806) );
  AND2_X1 U8591 ( .A1(n7809), .A2(n7808), .ZN(n14872) );
  NAND2_X1 U8592 ( .A1(n7910), .A2(n7238), .ZN(n15056) );
  OR2_X1 U8593 ( .A1(n12877), .A2(n7914), .ZN(n7910) );
  NAND2_X1 U8594 ( .A1(n7919), .A2(n12875), .ZN(n15082) );
  NAND2_X1 U8595 ( .A1(n7919), .A2(n7916), .ZN(n15994) );
  INV_X1 U8596 ( .A(n15998), .ZN(n15953) );
  OR2_X1 U8597 ( .A1(n11508), .A2(n14849), .ZN(n15671) );
  INV_X1 U8598 ( .A(n15949), .ZN(n15990) );
  INV_X1 U8599 ( .A(n10700), .ZN(n10843) );
  XNOR2_X1 U8600 ( .A(n9376), .B(n9361), .ZN(n14579) );
  XNOR2_X1 U8601 ( .A(n9323), .B(n9321), .ZN(n14589) );
  NOR2_X1 U8602 ( .A1(n7384), .A2(n7383), .ZN(n7382) );
  OR2_X1 U8603 ( .A1(n9908), .A2(n7386), .ZN(n7385) );
  NOR2_X1 U8604 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7383) );
  INV_X1 U8605 ( .A(n7687), .ZN(n7685) );
  NAND2_X1 U8606 ( .A1(n7995), .A2(n7387), .ZN(n9907) );
  AND2_X1 U8607 ( .A1(n9223), .A2(n8902), .ZN(n12150) );
  NAND2_X1 U8608 ( .A1(n7460), .A2(n7655), .ZN(n9188) );
  AOI21_X1 U8609 ( .B1(n7657), .B2(n7656), .A(n7328), .ZN(n7655) );
  NAND2_X1 U8610 ( .A1(n9148), .A2(n7657), .ZN(n7460) );
  NAND2_X1 U8611 ( .A1(n9150), .A2(n8890), .ZN(n9165) );
  AND2_X1 U8612 ( .A1(n9782), .A2(n9642), .ZN(n11893) );
  XNOR2_X1 U8613 ( .A(n8943), .B(n8942), .ZN(n10937) );
  AND2_X1 U8614 ( .A1(n9019), .A2(n9018), .ZN(n10808) );
  NAND2_X1 U8615 ( .A1(n7797), .A2(n8857), .ZN(n8994) );
  NOR2_X1 U8616 ( .A1(n8852), .A2(n9713), .ZN(n8982) );
  NAND2_X1 U8617 ( .A1(n7346), .A2(n7345), .ZN(n9707) );
  INV_X1 U8618 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15432) );
  AOI22_X1 U8619 ( .A1(n15478), .A2(n15477), .B1(P1_ADDR_REG_5__SCAN_IN), .B2(
        n15476), .ZN(n15481) );
  NAND2_X1 U8620 ( .A1(n7573), .A2(n7572), .ZN(n7571) );
  NAND2_X1 U8621 ( .A1(n15527), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7572) );
  INV_X1 U8622 ( .A(n15526), .ZN(n7573) );
  AND4_X1 U8623 ( .A1(n8747), .A2(n8746), .A3(n8745), .A4(n8744), .ZN(n13072)
         );
  OAI211_X1 U8624 ( .C1(n7711), .C2(n7696), .A(n7694), .B(n7701), .ZN(n13102)
         );
  AOI21_X1 U8625 ( .B1(n7703), .B2(n7706), .A(n7702), .ZN(n7701) );
  NAND2_X1 U8626 ( .A1(n7697), .A2(n7698), .ZN(n7696) );
  AND4_X1 U8627 ( .A1(n8508), .A2(n8507), .A3(n8506), .A4(n8505), .ZN(n13082)
         );
  AND3_X1 U8628 ( .A1(n8632), .A2(n8631), .A3(n8630), .ZN(n13575) );
  AND4_X1 U8629 ( .A1(n10130), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n13108)
         );
  NAND2_X1 U8630 ( .A1(n7447), .A2(n7446), .ZN(n11367) );
  INV_X1 U8631 ( .A(n11306), .ZN(n7446) );
  AND2_X1 U8632 ( .A1(n8640), .A2(n8639), .ZN(n13120) );
  NAND2_X1 U8633 ( .A1(n7724), .A2(n12779), .ZN(n12781) );
  NAND2_X1 U8634 ( .A1(n7710), .A2(n7709), .ZN(n13121) );
  NOR2_X1 U8635 ( .A1(n8226), .A2(n7713), .ZN(n7712) );
  INV_X1 U8636 ( .A(n13129), .ZN(n7713) );
  AND2_X1 U8637 ( .A1(n7714), .A2(n7717), .ZN(n13130) );
  INV_X1 U8638 ( .A(n13608), .ZN(n13139) );
  NAND2_X1 U8639 ( .A1(n11724), .A2(n11723), .ZN(n11730) );
  NAND2_X1 U8640 ( .A1(n7737), .A2(n12473), .ZN(n12476) );
  CLKBUF_X1 U8641 ( .A(n8368), .Z(n11303) );
  INV_X1 U8642 ( .A(n7722), .ZN(n7721) );
  AND2_X1 U8643 ( .A1(n12808), .A2(n7719), .ZN(n7718) );
  OR2_X1 U8644 ( .A1(n11218), .A2(n11307), .ZN(n13174) );
  NAND2_X1 U8645 ( .A1(n11207), .A2(n11206), .ZN(n13190) );
  AND2_X1 U8646 ( .A1(n12062), .A2(n12061), .ZN(n12064) );
  NAND2_X1 U8647 ( .A1(n7710), .A2(n7241), .ZN(n7700) );
  INV_X1 U8648 ( .A(n13172), .ZN(n13195) );
  NAND2_X1 U8649 ( .A1(n13045), .A2(n13044), .ZN(n13188) );
  INV_X1 U8650 ( .A(n13178), .ZN(n13197) );
  XNOR2_X1 U8651 ( .A(n8753), .B(P3_IR_REG_22__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U8652 ( .A1(n7441), .A2(n7440), .ZN(n8049) );
  INV_X1 U8653 ( .A(n10153), .ZN(n7440) );
  INV_X1 U8654 ( .A(n13560), .ZN(n13206) );
  INV_X1 U8655 ( .A(n12804), .ZN(n13212) );
  INV_X1 U8656 ( .A(n12573), .ZN(n13214) );
  INV_X1 U8657 ( .A(n12236), .ZN(n13218) );
  INV_X1 U8658 ( .A(n8120), .ZN(n8119) );
  INV_X1 U8659 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11162) );
  NOR2_X1 U8660 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11046), .ZN(n11156) );
  NAND2_X1 U8661 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8358) );
  XNOR2_X1 U8662 ( .A(n11037), .B(n7409), .ZN(n11133) );
  OR2_X1 U8663 ( .A1(n11165), .A2(n15727), .ZN(n11167) );
  AOI21_X1 U8664 ( .B1(n13237), .B2(n11752), .A(n13238), .ZN(n13244) );
  INV_X1 U8665 ( .A(n7947), .ZN(n15610) );
  INV_X1 U8666 ( .A(n7508), .ZN(n12156) );
  XNOR2_X1 U8667 ( .A(n7482), .B(n12687), .ZN(n12328) );
  INV_X1 U8668 ( .A(n7948), .ZN(n12694) );
  XNOR2_X1 U8669 ( .A(n13279), .B(n13280), .ZN(n13250) );
  NOR2_X1 U8670 ( .A1(n13332), .A2(n13331), .ZN(n13335) );
  NOR2_X1 U8671 ( .A1(n13335), .A2(n13334), .ZN(n13361) );
  NOR2_X1 U8672 ( .A1(n13360), .A2(n13359), .ZN(n13381) );
  MUX2_X1 U8673 ( .A(n11057), .B(n13223), .S(n11044), .Z(n15641) );
  NOR2_X1 U8674 ( .A1(n13406), .A2(n7495), .ZN(n13391) );
  AND2_X1 U8675 ( .A1(n13388), .A2(n13389), .ZN(n7495) );
  NAND2_X1 U8676 ( .A1(n8681), .A2(n8680), .ZN(n13654) );
  NAND2_X1 U8677 ( .A1(n7746), .A2(n13532), .ZN(n13517) );
  NAND2_X1 U8678 ( .A1(n8782), .A2(n10254), .ZN(n13524) );
  NAND2_X1 U8679 ( .A1(n13596), .A2(n10235), .ZN(n13579) );
  NAND2_X1 U8680 ( .A1(n8610), .A2(n8609), .ZN(n13582) );
  AND2_X1 U8681 ( .A1(n8592), .A2(n8591), .ZN(n13599) );
  AND2_X1 U8682 ( .A1(n8575), .A2(n8574), .ZN(n13618) );
  NAND2_X1 U8683 ( .A1(n12816), .A2(n8541), .ZN(n13623) );
  NAND2_X1 U8684 ( .A1(n8133), .A2(n8132), .ZN(n12767) );
  AND2_X1 U8685 ( .A1(n8133), .A2(n10216), .ZN(n12769) );
  NAND2_X1 U8686 ( .A1(n12735), .A2(n8778), .ZN(n8133) );
  NAND2_X1 U8687 ( .A1(n12455), .A2(n10197), .ZN(n12543) );
  NAND2_X1 U8688 ( .A1(n7411), .A2(n10194), .ZN(n12453) );
  INV_X1 U8689 ( .A(n12469), .ZN(n15857) );
  NAND2_X1 U8690 ( .A1(n12214), .A2(n10181), .ZN(n12125) );
  AND3_X1 U8691 ( .A1(n8433), .A2(n8432), .A3(n8431), .ZN(n15762) );
  INV_X1 U8692 ( .A(n13637), .ZN(n13568) );
  NAND2_X1 U8693 ( .A1(n11314), .A2(n11821), .ZN(n13520) );
  OR2_X1 U8694 ( .A1(n11320), .A2(n11940), .ZN(n13637) );
  NAND2_X1 U8695 ( .A1(n11320), .A2(n13520), .ZN(n13565) );
  INV_X1 U8696 ( .A(n13520), .ZN(n13634) );
  AOI21_X1 U8697 ( .B1(n13780), .B2(n10142), .A(n10141), .ZN(n13705) );
  INV_X1 U8698 ( .A(n10131), .ZN(n13708) );
  AND2_X1 U8699 ( .A1(n13453), .A2(n13452), .ZN(n13711) );
  XNOR2_X1 U8700 ( .A(n13468), .B(n13467), .ZN(n13716) );
  NAND2_X1 U8701 ( .A1(n13480), .A2(n13482), .ZN(n8124) );
  NOR2_X1 U8702 ( .A1(n13501), .A2(n13500), .ZN(n13727) );
  NAND2_X1 U8703 ( .A1(n8654), .A2(n8653), .ZN(n13734) );
  INV_X1 U8704 ( .A(n13120), .ZN(n13740) );
  AND3_X1 U8705 ( .A1(n13564), .A2(n13563), .A3(n13562), .ZN(n13744) );
  INV_X1 U8706 ( .A(n13599), .ZN(n13757) );
  INV_X1 U8707 ( .A(n13618), .ZN(n13761) );
  INV_X1 U8708 ( .A(n8509), .ZN(n12833) );
  AND2_X1 U8709 ( .A1(n8806), .A2(n8805), .ZN(n13771) );
  OR2_X1 U8710 ( .A1(n8258), .A2(n8255), .ZN(n7445) );
  NOR2_X1 U8711 ( .A1(n7444), .A2(n7443), .ZN(n7442) );
  XNOR2_X1 U8712 ( .A(n8721), .B(n8719), .ZN(n12743) );
  NAND2_X1 U8713 ( .A1(n8705), .A2(n8704), .ZN(n8721) );
  INV_X1 U8714 ( .A(n8252), .ZN(n8793) );
  NAND2_X1 U8715 ( .A1(n8054), .A2(n8665), .ZN(n8675) );
  NAND2_X1 U8716 ( .A1(n8664), .A2(n8663), .ZN(n8054) );
  NAND2_X1 U8717 ( .A1(n8621), .A2(n8634), .ZN(n8622) );
  NAND2_X1 U8718 ( .A1(n8035), .A2(n8040), .ZN(n8546) );
  NAND2_X1 U8719 ( .A1(n8526), .A2(n8042), .ZN(n8035) );
  NAND2_X1 U8720 ( .A1(n8044), .A2(n8042), .ZN(n8543) );
  NAND2_X1 U8721 ( .A1(n8044), .A2(n8045), .ZN(n8529) );
  INV_X1 U8722 ( .A(SI_12_), .ZN(n13914) );
  NAND2_X1 U8723 ( .A1(n8463), .A2(n8462), .ZN(n8479) );
  XNOR2_X1 U8724 ( .A(n8347), .B(n8348), .ZN(n12335) );
  NAND2_X1 U8725 ( .A1(n8058), .A2(n8296), .ZN(n8340) );
  NAND2_X1 U8726 ( .A1(n8294), .A2(n8293), .ZN(n8311) );
  OR2_X1 U8727 ( .A1(n7956), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n8392) );
  NOR2_X1 U8728 ( .A1(n10649), .A2(n10648), .ZN(n10758) );
  NAND2_X1 U8729 ( .A1(n7416), .A2(n7865), .ZN(n14071) );
  INV_X1 U8730 ( .A(n14042), .ZN(n7416) );
  INV_X1 U8731 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n12651) );
  NAND2_X1 U8732 ( .A1(n7882), .A2(n7881), .ZN(n14064) );
  OAI21_X1 U8733 ( .B1(n14138), .B2(n7875), .A(n7871), .ZN(n14082) );
  AOI21_X1 U8734 ( .B1(n7874), .B2(n7873), .A(n7872), .ZN(n7871) );
  INV_X1 U8735 ( .A(n14117), .ZN(n7872) );
  INV_X1 U8736 ( .A(n7879), .ZN(n7873) );
  NOR2_X1 U8737 ( .A1(n11344), .A2(n11345), .ZN(n11411) );
  NAND2_X1 U8738 ( .A1(n11987), .A2(n11994), .ZN(n12048) );
  NAND2_X1 U8739 ( .A1(n7876), .A2(n7877), .ZN(n14119) );
  NAND2_X1 U8740 ( .A1(n14138), .A2(n7879), .ZN(n7876) );
  AND2_X1 U8741 ( .A1(n7867), .A2(n12282), .ZN(n7866) );
  AND2_X1 U8742 ( .A1(n7868), .A2(n7867), .ZN(n12283) );
  NAND2_X1 U8743 ( .A1(n11102), .A2(n11378), .ZN(n11385) );
  AOI21_X1 U8744 ( .B1(n11425), .B2(n11424), .A(n11423), .ZN(n11428) );
  NOR2_X1 U8745 ( .A1(n12747), .A2(n12746), .ZN(n12853) );
  INV_X1 U8746 ( .A(n14135), .ZN(n14159) );
  OR2_X1 U8747 ( .A1(n10615), .A2(n11390), .ZN(n10616) );
  OR2_X1 U8748 ( .A1(n14279), .A2(n9398), .ZN(n9390) );
  INV_X1 U8749 ( .A(n14000), .ZN(n14168) );
  NAND2_X1 U8750 ( .A1(n9338), .A2(n9337), .ZN(n14169) );
  NAND2_X1 U8751 ( .A1(n9232), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9013) );
  NAND2_X1 U8752 ( .A1(n9003), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8981) );
  INV_X1 U8753 ( .A(n7617), .ZN(n14211) );
  NOR2_X1 U8754 ( .A1(n10769), .A2(n10768), .ZN(n10777) );
  INV_X1 U8755 ( .A(n7608), .ZN(n15272) );
  INV_X1 U8756 ( .A(n7425), .ZN(n15274) );
  INV_X1 U8757 ( .A(n7606), .ZN(n14222) );
  INV_X1 U8758 ( .A(n7615), .ZN(n14233) );
  NOR2_X1 U8759 ( .A1(n10772), .A2(P2_U3088), .ZN(n15271) );
  NOR2_X1 U8760 ( .A1(n15284), .A2(n15285), .ZN(n15287) );
  INV_X1 U8761 ( .A(n7609), .ZN(n15300) );
  NAND2_X1 U8762 ( .A1(n7256), .A2(n15340), .ZN(n7610) );
  OAI21_X1 U8763 ( .B1(n15377), .B2(n8275), .A(n15348), .ZN(n7427) );
  NAND2_X1 U8764 ( .A1(n7651), .A2(n7650), .ZN(n14246) );
  NAND2_X1 U8765 ( .A1(n7645), .A2(n7653), .ZN(n7650) );
  OAI21_X1 U8766 ( .B1(n14275), .B2(n14274), .A(n14273), .ZN(n14442) );
  NAND2_X1 U8767 ( .A1(n14292), .A2(n7213), .ZN(n14273) );
  AND2_X1 U8768 ( .A1(n14292), .A2(n9373), .ZN(n14275) );
  NAND2_X1 U8769 ( .A1(n7852), .A2(n7849), .ZN(n14271) );
  NAND2_X1 U8770 ( .A1(n7852), .A2(n9462), .ZN(n14269) );
  NAND2_X1 U8771 ( .A1(n9291), .A2(n9290), .ZN(n14469) );
  NAND2_X1 U8772 ( .A1(n7397), .A2(n8006), .ZN(n8000) );
  NAND2_X1 U8773 ( .A1(n8017), .A2(n8018), .ZN(n14421) );
  AND2_X1 U8774 ( .A1(n12590), .A2(n9205), .ZN(n12677) );
  NAND2_X1 U8775 ( .A1(n9180), .A2(n9179), .ZN(n15960) );
  NAND2_X1 U8776 ( .A1(n9440), .A2(n9439), .ZN(n12373) );
  NAND2_X1 U8777 ( .A1(n11973), .A2(n9131), .ZN(n12508) );
  AOI21_X1 U8778 ( .B1(n11789), .B2(n9435), .A(n7835), .ZN(n11975) );
  NOR2_X1 U8779 ( .A1(n11656), .A2(n7998), .ZN(n7997) );
  INV_X1 U8780 ( .A(n9093), .ZN(n7998) );
  NAND2_X1 U8781 ( .A1(n7822), .A2(n9432), .ZN(n11646) );
  INV_X1 U8782 ( .A(n15717), .ZN(n15934) );
  AND2_X1 U8783 ( .A1(n15721), .A2(n15707), .ZN(n15917) );
  NAND2_X1 U8784 ( .A1(n9154), .A2(n9153), .ZN(n12537) );
  NAND2_X1 U8785 ( .A1(n10536), .A2(n10535), .ZN(n14524) );
  INV_X1 U8786 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7505) );
  NAND2_X1 U8787 ( .A1(n9273), .A2(n9272), .ZN(n14540) );
  AND3_X1 U8788 ( .A1(n14484), .A2(n14483), .A3(n14482), .ZN(n14543) );
  INV_X1 U8789 ( .A(n14392), .ZN(n14549) );
  NAND2_X1 U8790 ( .A1(n9210), .A2(n9209), .ZN(n14557) );
  NAND2_X1 U8791 ( .A1(n9139), .A2(n9138), .ZN(n15918) );
  NAND2_X1 U8792 ( .A1(n10933), .A2(n7478), .ZN(n9121) );
  INV_X2 U8793 ( .A(n15971), .ZN(n15973) );
  AND2_X1 U8794 ( .A1(n8027), .A2(n8026), .ZN(n8025) );
  INV_X1 U8795 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8026) );
  INV_X1 U8796 ( .A(n8935), .ZN(n14573) );
  XNOR2_X1 U8797 ( .A(n9492), .B(n9491), .ZN(n14584) );
  NAND2_X1 U8798 ( .A1(n9490), .A2(n9486), .ZN(n14586) );
  OR2_X1 U8799 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  XNOR2_X1 U8800 ( .A(n9488), .B(n9487), .ZN(n14590) );
  NAND2_X1 U8801 ( .A1(n14563), .A2(n9409), .ZN(n9412) );
  INV_X1 U8802 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n12153) );
  INV_X1 U8803 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11278) );
  INV_X1 U8804 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11152) );
  INV_X1 U8805 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10855) );
  INV_X1 U8806 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10850) );
  INV_X1 U8807 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10821) );
  INV_X1 U8808 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10825) );
  INV_X1 U8809 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10810) );
  NOR2_X1 U8810 ( .A1(n9022), .A2(n9021), .ZN(n14210) );
  MUX2_X1 U8811 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7600), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8989) );
  NAND2_X1 U8812 ( .A1(n10873), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10713) );
  NAND2_X1 U8813 ( .A1(n8190), .A2(n8195), .ZN(n12194) );
  NAND2_X1 U8814 ( .A1(n10793), .A2(n10739), .ZN(n8190) );
  NAND2_X1 U8815 ( .A1(n14684), .A2(n12925), .ZN(n14603) );
  NOR2_X1 U8816 ( .A1(n10962), .A2(n10961), .ZN(n10960) );
  NAND2_X1 U8817 ( .A1(n14678), .A2(n12971), .ZN(n14638) );
  NAND2_X1 U8818 ( .A1(n9590), .A2(n9589), .ZN(n15154) );
  NAND2_X1 U8819 ( .A1(n7563), .A2(n7279), .ZN(n14645) );
  NAND2_X1 U8820 ( .A1(n14655), .A2(n14656), .ZN(n14654) );
  NAND2_X1 U8821 ( .A1(n14668), .A2(n12998), .ZN(n14655) );
  NOR2_X1 U8822 ( .A1(n10724), .A2(n10723), .ZN(n16011) );
  NAND2_X1 U8823 ( .A1(n7562), .A2(n8215), .ZN(n10737) );
  NAND2_X1 U8824 ( .A1(n8210), .A2(n12945), .ZN(n16021) );
  NAND2_X1 U8825 ( .A1(n16006), .A2(n16007), .ZN(n8210) );
  AND2_X1 U8826 ( .A1(n8214), .A2(n8215), .ZN(n11575) );
  NAND2_X1 U8827 ( .A1(n12257), .A2(n12256), .ZN(n12361) );
  INV_X1 U8828 ( .A(n7563), .ZN(n12908) );
  NAND2_X1 U8829 ( .A1(n12557), .A2(n8213), .ZN(n12560) );
  INV_X1 U8830 ( .A(n7545), .ZN(n7544) );
  NAND2_X1 U8831 ( .A1(n7545), .A2(n7226), .ZN(n7542) );
  AND4_X1 U8832 ( .A1(n9743), .A2(n9742), .A3(n9741), .A4(n9740), .ZN(n11686)
         );
  NAND2_X1 U8833 ( .A1(n15975), .A2(n15976), .ZN(n15974) );
  NAND2_X1 U8834 ( .A1(n10052), .A2(n7378), .ZN(n7377) );
  AND2_X1 U8835 ( .A1(n10076), .A2(n7439), .ZN(n7453) );
  AND2_X1 U8836 ( .A1(n10057), .A2(n10077), .ZN(n7439) );
  NAND2_X1 U8837 ( .A1(n10057), .A2(n7500), .ZN(n7499) );
  OAI21_X1 U8838 ( .B1(n14945), .B2(n9722), .A(n9876), .ZN(n14958) );
  NAND2_X1 U8839 ( .A1(n9598), .A2(n9597), .ZN(n14984) );
  INV_X1 U8840 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10951) );
  INV_X1 U8841 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10953) );
  AND4_X1 U8842 ( .A1(n9691), .A2(n9690), .A3(n9689), .A4(n9688), .ZN(n11709)
         );
  CLKBUF_X1 U8843 ( .A(n10660), .Z(n14744) );
  NAND2_X1 U8844 ( .A1(n10987), .A2(n7277), .ZN(n14762) );
  NAND2_X1 U8845 ( .A1(n14788), .A2(n7322), .ZN(n10869) );
  INV_X1 U8846 ( .A(n7528), .ZN(n10897) );
  AND2_X1 U8847 ( .A1(n7528), .A2(n7527), .ZN(n10899) );
  NAND2_X1 U8848 ( .A1(n10903), .A2(n10898), .ZN(n7527) );
  INV_X1 U8849 ( .A(n7532), .ZN(n11455) );
  INV_X1 U8850 ( .A(n7530), .ZN(n11884) );
  AND2_X1 U8851 ( .A1(n7530), .A2(n7529), .ZN(n14808) );
  NAND2_X1 U8852 ( .A1(n11891), .A2(n11885), .ZN(n7529) );
  XNOR2_X1 U8853 ( .A(n9783), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14823) );
  NOR2_X1 U8854 ( .A1(n14832), .A2(n7534), .ZN(n15396) );
  NAND2_X1 U8855 ( .A1(n14898), .A2(n7810), .ZN(n14882) );
  NAND2_X1 U8856 ( .A1(n14913), .A2(n8231), .ZN(n14901) );
  NAND2_X1 U8857 ( .A1(n9848), .A2(n9847), .ZN(n14919) );
  NAND2_X1 U8858 ( .A1(n7788), .A2(n7789), .ZN(n14925) );
  NAND2_X1 U8859 ( .A1(n7785), .A2(n7786), .ZN(n14924) );
  NAND2_X1 U8860 ( .A1(n14964), .A2(n7790), .ZN(n7788) );
  AND2_X1 U8861 ( .A1(n7793), .A2(n7249), .ZN(n14940) );
  NAND2_X1 U8862 ( .A1(n14964), .A2(n14965), .ZN(n7793) );
  AND2_X1 U8863 ( .A1(n7804), .A2(n7260), .ZN(n14991) );
  AND2_X1 U8864 ( .A1(n7804), .A2(n7803), .ZN(n15162) );
  NAND2_X1 U8865 ( .A1(n7936), .A2(n7933), .ZN(n14979) );
  NAND2_X1 U8866 ( .A1(n7931), .A2(n7930), .ZN(n14996) );
  NAND2_X1 U8867 ( .A1(n8116), .A2(n12866), .ZN(n15038) );
  NAND2_X1 U8868 ( .A1(n9628), .A2(n9627), .ZN(n16008) );
  OR2_X1 U8869 ( .A1(n11572), .A2(n9757), .ZN(n9628) );
  INV_X1 U8870 ( .A(n12865), .ZN(n7815) );
  INV_X1 U8871 ( .A(n8109), .ZN(n8108) );
  AND2_X1 U8872 ( .A1(n15021), .A2(n15993), .ZN(n15083) );
  NAND2_X1 U8873 ( .A1(n12349), .A2(n15880), .ZN(n12350) );
  NAND2_X1 U8874 ( .A1(n12354), .A2(n12353), .ZN(n12405) );
  NAND2_X1 U8875 ( .A1(n7899), .A2(n7898), .ZN(n12005) );
  NAND2_X1 U8876 ( .A1(n7899), .A2(n11859), .ZN(n11862) );
  NAND2_X1 U8877 ( .A1(n8113), .A2(n11506), .ZN(n11524) );
  NAND2_X1 U8878 ( .A1(n15021), .A2(n12090), .ZN(n15069) );
  NAND2_X1 U8879 ( .A1(n11498), .A2(n11497), .ZN(n15660) );
  AND2_X1 U8880 ( .A1(n7214), .A2(n7906), .ZN(n7905) );
  AND2_X1 U8881 ( .A1(n8219), .A2(n7907), .ZN(n7906) );
  AND2_X1 U8882 ( .A1(n9536), .A2(n9544), .ZN(n7907) );
  NAND2_X1 U8883 ( .A1(n7380), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7438) );
  XNOR2_X1 U8884 ( .A(n10089), .B(n10088), .ZN(n15228) );
  XNOR2_X1 U8885 ( .A(n9581), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15237) );
  INV_X1 U8886 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n12151) );
  INV_X1 U8887 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11570) );
  INV_X1 U8888 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11550) );
  INV_X1 U8889 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11279) );
  INV_X1 U8890 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n11150) );
  INV_X1 U8891 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10935) );
  NAND2_X1 U8892 ( .A1(n7662), .A2(n8877), .ZN(n8961) );
  NAND2_X1 U8893 ( .A1(n7665), .A2(n8877), .ZN(n8959) );
  OAI21_X1 U8894 ( .B1(n9078), .B2(n8087), .A(n8085), .ZN(n9097) );
  INV_X1 U8895 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10851) );
  NAND2_X1 U8896 ( .A1(n7805), .A2(n9044), .ZN(n10832) );
  AOI21_X1 U8897 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(n15438), .A(n15606), .ZN(
        n15440) );
  XNOR2_X1 U8898 ( .A(n15490), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15485) );
  OAI21_X1 U8899 ( .B1(n15502), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n15501), .ZN(
        n15504) );
  NAND2_X1 U8900 ( .A1(n15504), .A2(n15505), .ZN(n15506) );
  NOR2_X1 U8901 ( .A1(n15512), .A2(n15511), .ZN(n15513) );
  NAND2_X1 U8902 ( .A1(n15554), .A2(n15553), .ZN(n15555) );
  NOR2_X1 U8903 ( .A1(n15562), .A2(n15561), .ZN(n15563) );
  NAND2_X1 U8904 ( .A1(n15567), .A2(n15566), .ZN(n15579) );
  NOR2_X1 U8905 ( .A1(n15585), .A2(n15584), .ZN(n15594) );
  AND2_X1 U8906 ( .A1(n10650), .A2(n13772), .ZN(P3_U3897) );
  INV_X1 U8907 ( .A(n7946), .ZN(n11756) );
  OR2_X1 U8908 ( .A1(n7230), .A2(n7768), .ZN(n13312) );
  XNOR2_X1 U8909 ( .A(n7401), .B(n13409), .ZN(n13426) );
  NOR2_X1 U8910 ( .A1(n7319), .A2(n7488), .ZN(n7487) );
  INV_X1 U8911 ( .A(n7421), .ZN(n8843) );
  NOR2_X1 U8912 ( .A1(n15894), .A2(n8844), .ZN(n7488) );
  OAI22_X1 U8913 ( .A1(n13437), .A2(n13767), .B1(n15898), .B2(n10644), .ZN(
        n10645) );
  OAI21_X1 U8914 ( .B1(n7421), .B2(n15895), .A(n7420), .ZN(n8831) );
  NAND2_X1 U8915 ( .A1(n15895), .A2(n8830), .ZN(n7420) );
  INV_X1 U8916 ( .A(n7857), .ZN(n7856) );
  NAND2_X1 U8917 ( .A1(n7428), .A2(n7426), .ZN(P2_U3233) );
  NAND2_X1 U8918 ( .A1(n7611), .A2(n15251), .ZN(n7428) );
  NOR2_X1 U8919 ( .A1(n7610), .A2(n7427), .ZN(n7426) );
  XNOR2_X1 U8920 ( .A(n7612), .B(n7338), .ZN(n7611) );
  OR2_X1 U8921 ( .A1(n15970), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7854) );
  NOR2_X1 U8922 ( .A1(n7318), .A2(n7504), .ZN(n7503) );
  NAND2_X1 U8923 ( .A1(n9517), .A2(n15973), .ZN(n7506) );
  NOR2_X1 U8924 ( .A1(n15973), .A2(n7505), .ZN(n7504) );
  NOR2_X1 U8925 ( .A1(n10714), .A2(n10713), .ZN(P1_U4016) );
  NAND2_X1 U8926 ( .A1(n7549), .A2(n16010), .ZN(n7548) );
  AOI21_X1 U8927 ( .B1(n15381), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n14851), .ZN(
        n7538) );
  NAND2_X1 U8928 ( .A1(n7540), .A2(n12404), .ZN(n7539) );
  NAND2_X1 U8929 ( .A1(n14850), .A2(n14849), .ZN(n7537) );
  XNOR2_X1 U8930 ( .A(n7581), .B(n7579), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8931 ( .A(n15601), .B(n7580), .ZN(n7579) );
  AOI21_X1 U8932 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15596), .A(n15595), .ZN(
        n7581) );
  XNOR2_X1 U8933 ( .A(n7340), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7580) );
  INV_X2 U8934 ( .A(n9949), .ZN(n10054) );
  OAI21_X2 U8935 ( .B1(n9944), .B2(n9945), .A(n7967), .ZN(n9949) );
  INV_X2 U8936 ( .A(n10375), .ZN(n10396) );
  AND2_X1 U8937 ( .A1(n7966), .A2(n10029), .ZN(n7211) );
  AND2_X1 U8938 ( .A1(n9990), .A2(n9992), .ZN(n7212) );
  NAND2_X1 U8939 ( .A1(n9797), .A2(n9796), .ZN(n12915) );
  INV_X1 U8940 ( .A(n12915), .ZN(n7584) );
  INV_X1 U8941 ( .A(n15055), .ZN(n7912) );
  INV_X1 U8942 ( .A(n12624), .ZN(n8112) );
  AND2_X1 U8943 ( .A1(n14274), .A2(n9373), .ZN(n7213) );
  AND2_X1 U8944 ( .A1(n8176), .A2(n10502), .ZN(n7215) );
  INV_X1 U8945 ( .A(n8382), .ZN(n8470) );
  INV_X2 U8946 ( .A(n8470), .ZN(n8434) );
  NAND2_X1 U8947 ( .A1(n9550), .A2(n9549), .ZN(n15105) );
  AND2_X1 U8948 ( .A1(n11682), .A2(n11705), .ZN(n7216) );
  XNOR2_X1 U8949 ( .A(n15170), .B(n8101), .ZN(n14995) );
  INV_X1 U8950 ( .A(n14995), .ZN(n7937) );
  AND2_X1 U8951 ( .A1(n9480), .A2(n7632), .ZN(n7217) );
  NAND2_X1 U8952 ( .A1(n9331), .A2(n9330), .ZN(n14323) );
  INV_X1 U8953 ( .A(n14500), .ZN(n7838) );
  AND3_X1 U8954 ( .A1(n13065), .A2(n13528), .A3(n13515), .ZN(n7218) );
  AND2_X1 U8955 ( .A1(n7550), .A2(n7287), .ZN(n7219) );
  OR2_X1 U8956 ( .A1(n13066), .A2(n13205), .ZN(n7220) );
  INV_X1 U8957 ( .A(n9976), .ZN(n7355) );
  AND2_X1 U8958 ( .A1(n12213), .A2(n14738), .ZN(n7221) );
  NOR2_X1 U8959 ( .A1(n14361), .A2(n7636), .ZN(n7635) );
  AND4_X1 U8960 ( .A1(n13513), .A2(n7745), .A3(n10316), .A4(n13542), .ZN(n7222) );
  AND2_X1 U8961 ( .A1(n7591), .A2(n7590), .ZN(n7223) );
  AND2_X1 U8962 ( .A1(n7641), .A2(n7640), .ZN(n7224) );
  AND2_X1 U8963 ( .A1(n7585), .A2(n7584), .ZN(n7225) );
  INV_X1 U8964 ( .A(n9147), .ZN(n8888) );
  NAND2_X1 U8965 ( .A1(n12952), .A2(n12945), .ZN(n7226) );
  NAND2_X1 U8966 ( .A1(n8063), .A2(n7317), .ZN(n7227) );
  NAND2_X1 U8967 ( .A1(n7864), .A2(n7865), .ZN(n7228) );
  AND2_X1 U8968 ( .A1(n14936), .A2(n7794), .ZN(n7229) );
  AND2_X1 U8969 ( .A1(n7767), .A2(n13320), .ZN(n7230) );
  NAND2_X1 U8970 ( .A1(n12909), .A2(n12910), .ZN(n7231) );
  AND2_X1 U8971 ( .A1(n7216), .A2(n7583), .ZN(n7232) );
  INV_X1 U8972 ( .A(n10056), .ZN(n7379) );
  NAND2_X1 U8973 ( .A1(n7734), .A2(n7250), .ZN(n8572) );
  AND2_X1 U8974 ( .A1(n9843), .A2(n9842), .ZN(n16018) );
  AND2_X1 U8975 ( .A1(n12865), .A2(n12864), .ZN(n7233) );
  INV_X1 U8976 ( .A(n16022), .ZN(n16010) );
  AND2_X1 U8977 ( .A1(n7585), .A2(n12349), .ZN(n7234) );
  NAND2_X1 U8978 ( .A1(n9612), .A2(n9901), .ZN(n12404) );
  INV_X1 U8979 ( .A(n8781), .ZN(n7745) );
  INV_X2 U8980 ( .A(n12999), .ZN(n13024) );
  XOR2_X1 U8981 ( .A(n14540), .B(n14072), .Z(n7235) );
  NAND2_X2 U8982 ( .A1(n8951), .A2(n8950), .ZN(n12279) );
  AND2_X1 U8983 ( .A1(n10398), .A2(n10397), .ZN(n7236) );
  INV_X2 U8984 ( .A(n8850), .ZN(n10806) );
  NAND2_X1 U8985 ( .A1(n8124), .A2(n10273), .ZN(n13467) );
  OR2_X1 U8986 ( .A1(n7916), .A2(n7913), .ZN(n7238) );
  INV_X1 U8987 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9537) );
  INV_X1 U8988 ( .A(n15114), .ZN(n7598) );
  AND2_X1 U8989 ( .A1(n7606), .A2(n7605), .ZN(n7239) );
  OR2_X1 U8990 ( .A1(n14361), .A2(n14469), .ZN(n7240) );
  AND2_X1 U8991 ( .A1(n7708), .A2(n7709), .ZN(n7241) );
  NAND2_X1 U8992 ( .A1(n14392), .A2(n14174), .ZN(n7242) );
  NAND2_X1 U8993 ( .A1(n7937), .A2(n7930), .ZN(n7929) );
  NAND2_X1 U8994 ( .A1(n10528), .A2(n10527), .ZN(n10578) );
  INV_X1 U8995 ( .A(n12669), .ZN(n11390) );
  AND2_X1 U8996 ( .A1(n10505), .A2(n10504), .ZN(n7243) );
  INV_X1 U8997 ( .A(n8090), .ZN(n8089) );
  AND2_X1 U8998 ( .A1(n14914), .A2(n8074), .ZN(n7244) );
  INV_X1 U8999 ( .A(n15135), .ZN(n14936) );
  NAND2_X1 U9000 ( .A1(n9857), .A2(n9856), .ZN(n15135) );
  INV_X1 U9001 ( .A(n9207), .ZN(n8081) );
  AND2_X1 U9002 ( .A1(n11297), .A2(n11298), .ZN(n7245) );
  OR2_X1 U9003 ( .A1(n10078), .A2(n10077), .ZN(n7246) );
  OR2_X1 U9004 ( .A1(n14981), .A2(n15154), .ZN(n7247) );
  INV_X1 U9005 ( .A(n10578), .ZN(n7653) );
  INV_X1 U9006 ( .A(n14595), .ZN(n7557) );
  NAND2_X1 U9007 ( .A1(n11404), .A2(n11403), .ZN(n7248) );
  OR2_X1 U9008 ( .A1(n14959), .A2(n14732), .ZN(n7249) );
  AND2_X1 U9009 ( .A1(n8551), .A2(n7735), .ZN(n7250) );
  NAND2_X1 U9010 ( .A1(n12043), .A2(n12038), .ZN(n7251) );
  INV_X1 U9011 ( .A(n10273), .ZN(n8127) );
  NAND2_X1 U9012 ( .A1(n15974), .A2(n8224), .ZN(n16006) );
  NAND2_X1 U9013 ( .A1(n9572), .A2(n9571), .ZN(n15121) );
  INV_X1 U9014 ( .A(n15121), .ZN(n14724) );
  NAND2_X1 U9015 ( .A1(n9381), .A2(n9380), .ZN(n14444) );
  INV_X1 U9016 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8914) );
  AND2_X1 U9017 ( .A1(n8000), .A2(n8003), .ZN(n7252) );
  INV_X1 U9018 ( .A(n11129), .ZN(n7493) );
  INV_X1 U9019 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9544) );
  INV_X1 U9020 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9904) );
  OR2_X1 U9021 ( .A1(n15617), .A2(n11753), .ZN(n7253) );
  AND2_X1 U9022 ( .A1(n12045), .A2(n12037), .ZN(n7254) );
  AND2_X1 U9023 ( .A1(n13146), .A2(n13064), .ZN(n7255) );
  INV_X1 U9024 ( .A(n14959), .ZN(n7591) );
  INV_X1 U9025 ( .A(n15081), .ZN(n7918) );
  INV_X1 U9026 ( .A(n11447), .ZN(n8118) );
  OR2_X1 U9027 ( .A1(n15364), .A2(n15347), .ZN(n7256) );
  NAND2_X1 U9028 ( .A1(n9197), .A2(n9196), .ZN(n14512) );
  INV_X1 U9029 ( .A(n10029), .ZN(n7965) );
  NAND2_X1 U9030 ( .A1(n12997), .A2(n14665), .ZN(n14668) );
  AND2_X1 U9031 ( .A1(n9345), .A2(n9344), .ZN(n14531) );
  INV_X1 U9032 ( .A(n14531), .ZN(n7634) );
  AND2_X1 U9033 ( .A1(n7545), .A2(n15976), .ZN(n7257) );
  AND2_X1 U9034 ( .A1(n15918), .A2(n14182), .ZN(n7258) );
  AND2_X1 U9035 ( .A1(n15900), .A2(n14736), .ZN(n7259) );
  OR2_X1 U9036 ( .A1(n15170), .A2(n15031), .ZN(n7260) );
  AND2_X1 U9037 ( .A1(n7870), .A2(n11994), .ZN(n7261) );
  AND2_X1 U9038 ( .A1(n8608), .A2(n11129), .ZN(n7262) );
  INV_X1 U9039 ( .A(n7592), .ZN(n14944) );
  NAND2_X1 U9040 ( .A1(n9868), .A2(n9867), .ZN(n15141) );
  INV_X1 U9041 ( .A(n11860), .ZN(n7900) );
  INV_X4 U9042 ( .A(n10806), .ZN(n10801) );
  NOR2_X1 U9043 ( .A1(n14376), .A2(n14173), .ZN(n7263) );
  AND2_X1 U9044 ( .A1(n8245), .A2(n8156), .ZN(n7264) );
  OR2_X1 U9045 ( .A1(n14361), .A2(n14323), .ZN(n7265) );
  NAND2_X1 U9046 ( .A1(n7385), .A2(n7382), .ZN(n10939) );
  AOI21_X1 U9047 ( .B1(n8089), .B2(n8088), .A(n7658), .ZN(n7657) );
  INV_X1 U9048 ( .A(n8079), .ZN(n8078) );
  INV_X1 U9049 ( .A(n10042), .ZN(n7959) );
  AND2_X1 U9050 ( .A1(n14500), .A2(n14008), .ZN(n7266) );
  AND2_X1 U9051 ( .A1(n13311), .A2(n13310), .ZN(n7267) );
  INV_X1 U9052 ( .A(n7635), .ZN(n7639) );
  AND2_X1 U9053 ( .A1(n10000), .A2(n9999), .ZN(n7268) );
  INV_X1 U9054 ( .A(n7593), .ZN(n14957) );
  NAND2_X1 U9055 ( .A1(n7223), .A2(n7589), .ZN(n7593) );
  AND2_X1 U9056 ( .A1(n8564), .A2(n8541), .ZN(n7269) );
  AND2_X1 U9057 ( .A1(n7217), .A2(n15941), .ZN(n7270) );
  AND2_X1 U9058 ( .A1(n7845), .A2(n7843), .ZN(n7271) );
  INV_X1 U9059 ( .A(n7791), .ZN(n7790) );
  NAND2_X1 U9060 ( .A1(n14965), .A2(n7795), .ZN(n7791) );
  OR2_X1 U9061 ( .A1(n10457), .A2(n10458), .ZN(n7272) );
  AND2_X1 U9062 ( .A1(n8648), .A2(n8633), .ZN(n7273) );
  AND2_X1 U9063 ( .A1(n12929), .A2(n12925), .ZN(n7276) );
  OR2_X1 U9064 ( .A1(n10881), .A2(n10863), .ZN(n7277) );
  INV_X1 U9065 ( .A(n7811), .ZN(n7810) );
  OR2_X1 U9066 ( .A1(n7236), .A2(n8182), .ZN(n7278) );
  INV_X1 U9067 ( .A(n8019), .ZN(n8018) );
  NOR2_X1 U9068 ( .A1(n8020), .A2(n9220), .ZN(n8019) );
  AND2_X1 U9069 ( .A1(n7231), .A2(n14646), .ZN(n7279) );
  AND2_X1 U9070 ( .A1(n10234), .A2(n10235), .ZN(n13593) );
  INV_X1 U9071 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7387) );
  NOR2_X1 U9072 ( .A1(n15918), .A2(n14182), .ZN(n7280) );
  NOR2_X1 U9073 ( .A1(n15077), .A2(n15058), .ZN(n7281) );
  NOR2_X1 U9074 ( .A1(n14405), .A2(n9447), .ZN(n7282) );
  NOR2_X1 U9075 ( .A1(n15900), .A2(n14736), .ZN(n7283) );
  NOR2_X1 U9076 ( .A1(n15960), .A2(n9442), .ZN(n7284) );
  NOR2_X1 U9077 ( .A1(n14444), .A2(n14166), .ZN(n7285) );
  OR2_X1 U9078 ( .A1(n7358), .A2(n7357), .ZN(n7286) );
  INV_X1 U9079 ( .A(n9939), .ZN(n15099) );
  NAND2_X1 U9080 ( .A1(n9881), .A2(n9880), .ZN(n9939) );
  OR2_X1 U9081 ( .A1(n7552), .A2(n13029), .ZN(n7287) );
  AND2_X1 U9082 ( .A1(n10027), .A2(n7965), .ZN(n7288) );
  INV_X1 U9083 ( .A(n9978), .ZN(n7991) );
  AND2_X1 U9084 ( .A1(n7456), .A2(n12507), .ZN(n7289) );
  AND2_X1 U9085 ( .A1(n8882), .A2(n13912), .ZN(n7290) );
  AND2_X1 U9086 ( .A1(n13186), .A2(n13209), .ZN(n7291) );
  AND2_X1 U9087 ( .A1(n7959), .A2(n7961), .ZN(n7292) );
  INV_X1 U9088 ( .A(n15018), .ZN(n15175) );
  AND2_X1 U9089 ( .A1(n9834), .A2(n9833), .ZN(n15018) );
  INV_X1 U9090 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10831) );
  INV_X1 U9091 ( .A(n7404), .ZN(n7746) );
  NAND2_X1 U9092 ( .A1(n10479), .A2(n10480), .ZN(n7293) );
  AND3_X1 U9093 ( .A1(n10091), .A2(n9911), .A3(n10085), .ZN(n7294) );
  AND2_X1 U9094 ( .A1(n8022), .A2(n12592), .ZN(n7295) );
  NAND2_X1 U9095 ( .A1(n13657), .A2(n13204), .ZN(n7296) );
  AND2_X1 U9096 ( .A1(n13499), .A2(n10271), .ZN(n13513) );
  INV_X1 U9097 ( .A(n13513), .ZN(n7747) );
  NAND2_X1 U9098 ( .A1(n7995), .A2(n7994), .ZN(n9926) );
  INV_X1 U9099 ( .A(n9926), .ZN(n7384) );
  AND2_X1 U9100 ( .A1(n8093), .A2(n8092), .ZN(n7297) );
  AND2_X1 U9101 ( .A1(n14376), .A2(n14173), .ZN(n7298) );
  NAND2_X1 U9102 ( .A1(n10791), .A2(n10738), .ZN(n8195) );
  NAND2_X1 U9103 ( .A1(n16020), .A2(n8211), .ZN(n7299) );
  INV_X1 U9104 ( .A(n9975), .ZN(n7358) );
  INV_X1 U9105 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8916) );
  INV_X1 U9106 ( .A(n7926), .ZN(n7925) );
  NAND2_X1 U9107 ( .A1(n7927), .A2(n7934), .ZN(n7926) );
  INV_X1 U9108 ( .A(n10005), .ZN(n7977) );
  OR2_X1 U9109 ( .A1(n13395), .A2(n13380), .ZN(n7300) );
  NOR2_X1 U9110 ( .A1(n13396), .A2(n13397), .ZN(n7301) );
  INV_X1 U9111 ( .A(n10495), .ZN(n8180) );
  OR2_X1 U9112 ( .A1(n10518), .A2(n7332), .ZN(n7302) );
  INV_X1 U9113 ( .A(n7412), .ZN(n8075) );
  NAND2_X1 U9114 ( .A1(n10287), .A2(n10284), .ZN(n10635) );
  AND2_X1 U9115 ( .A1(n12473), .A2(n12474), .ZN(n7303) );
  AND2_X1 U9116 ( .A1(n11506), .A2(n11525), .ZN(n7304) );
  AND2_X1 U9117 ( .A1(n7246), .A2(n10103), .ZN(n7305) );
  INV_X1 U9118 ( .A(n12945), .ZN(n8212) );
  AND2_X1 U9119 ( .A1(n10684), .A2(n8216), .ZN(n7306) );
  OR2_X1 U9120 ( .A1(n8169), .A2(n10526), .ZN(n7307) );
  INV_X1 U9121 ( .A(n15105), .ZN(n14868) );
  AND2_X1 U9122 ( .A1(n9610), .A2(n7387), .ZN(n7308) );
  AND2_X1 U9123 ( .A1(n8075), .A2(n8074), .ZN(n7309) );
  INV_X1 U9124 ( .A(n8958), .ZN(n7664) );
  AND2_X1 U9125 ( .A1(n10047), .A2(n10046), .ZN(n7310) );
  OR2_X1 U9126 ( .A1(n7243), .A2(n8184), .ZN(n7311) );
  NAND2_X1 U9127 ( .A1(n12278), .A2(n12277), .ZN(n7312) );
  INV_X1 U9128 ( .A(n12921), .ZN(n15926) );
  NAND2_X1 U9129 ( .A1(n9645), .A2(n9644), .ZN(n12921) );
  AND2_X1 U9130 ( .A1(n7858), .A2(n14102), .ZN(n7313) );
  NAND2_X1 U9131 ( .A1(n10045), .A2(n7980), .ZN(n7314) );
  INV_X1 U9132 ( .A(n9974), .ZN(n7987) );
  INV_X1 U9133 ( .A(n7850), .ZN(n7849) );
  NAND2_X1 U9134 ( .A1(n7851), .A2(n9462), .ZN(n7850) );
  INV_X1 U9135 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7462) );
  INV_X1 U9136 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10088) );
  INV_X1 U9137 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7735) );
  INV_X1 U9138 ( .A(n12687), .ZN(n7941) );
  NAND2_X1 U9139 ( .A1(n12557), .A2(n7564), .ZN(n7563) );
  INV_X1 U9140 ( .A(n12452), .ZN(n8149) );
  INV_X1 U9141 ( .A(n14041), .ZN(n7865) );
  NAND2_X1 U9142 ( .A1(n8485), .A2(n8245), .ZN(n8487) );
  INV_X1 U9143 ( .A(n14731), .ZN(n7794) );
  AND3_X2 U9144 ( .A1(n9532), .A2(n9636), .A3(n9531), .ZN(n9621) );
  INV_X1 U9145 ( .A(n7498), .ZN(n7409) );
  INV_X1 U9146 ( .A(n9004), .ZN(n9088) );
  NAND2_X1 U9147 ( .A1(n12407), .A2(n12406), .ZN(n12625) );
  AND2_X1 U9148 ( .A1(n12175), .A2(n12178), .ZN(n7315) );
  INV_X1 U9149 ( .A(n10300), .ZN(n8151) );
  OR2_X1 U9150 ( .A1(n14016), .A2(n14015), .ZN(n7316) );
  INV_X1 U9151 ( .A(n14715), .ZN(n7556) );
  NAND2_X1 U9152 ( .A1(n9310), .A2(n9309), .ZN(n14466) );
  INV_X1 U9153 ( .A(n14466), .ZN(n7638) );
  NAND2_X1 U9154 ( .A1(n8480), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7317) );
  INV_X1 U9155 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9634) );
  AND2_X1 U9156 ( .A1(n14262), .A2(n14558), .ZN(n7318) );
  INV_X1 U9157 ( .A(n8077), .ZN(n7674) );
  NOR2_X1 U9158 ( .A1(n8080), .A2(n13898), .ZN(n8077) );
  NOR2_X1 U9159 ( .A1(n13446), .A2(n13694), .ZN(n7319) );
  AND2_X1 U9160 ( .A1(n7800), .A2(n7801), .ZN(n7320) );
  AND2_X1 U9161 ( .A1(n7882), .A2(n7879), .ZN(n7321) );
  INV_X1 U9162 ( .A(n8006), .ZN(n8005) );
  NOR2_X1 U9163 ( .A1(n7263), .A2(n8007), .ZN(n8006) );
  NAND2_X1 U9164 ( .A1(n12597), .A2(n7643), .ZN(n7644) );
  OR2_X1 U9165 ( .A1(n10889), .A2(n10868), .ZN(n7322) );
  AND2_X1 U9166 ( .A1(n8107), .A2(n8108), .ZN(n7323) );
  OR2_X1 U9167 ( .A1(n7815), .A2(n7814), .ZN(n7324) );
  INV_X1 U9168 ( .A(n7929), .ZN(n7928) );
  NAND2_X1 U9169 ( .A1(n11263), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7325) );
  AND2_X1 U9170 ( .A1(n7563), .A2(n7231), .ZN(n7326) );
  AND2_X1 U9171 ( .A1(n7920), .A2(n7925), .ZN(n7327) );
  INV_X1 U9172 ( .A(SI_18_), .ZN(n13898) );
  AND2_X1 U9173 ( .A1(n8893), .A2(n13821), .ZN(n7328) );
  AND2_X1 U9174 ( .A1(n9256), .A2(SI_20_), .ZN(n7329) );
  AND2_X1 U9175 ( .A1(n10501), .A2(n10500), .ZN(n7330) );
  OR2_X1 U9176 ( .A1(n8547), .A2(n7730), .ZN(n7331) );
  INV_X1 U9177 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11419) );
  AND2_X1 U9178 ( .A1(n10515), .A2(n10514), .ZN(n7332) );
  INV_X1 U9179 ( .A(n7686), .ZN(n7684) );
  NOR2_X1 U9180 ( .A1(n9254), .A2(n7687), .ZN(n7686) );
  XNOR2_X1 U9181 ( .A(n9239), .B(SI_19_), .ZN(n9240) );
  INV_X1 U9182 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8255) );
  INV_X1 U9183 ( .A(n15031), .ZN(n8101) );
  INV_X1 U9184 ( .A(SI_14_), .ZN(n8092) );
  INV_X1 U9185 ( .A(n14405), .ZN(n7640) );
  INV_X1 U9186 ( .A(n14163), .ZN(n14102) );
  NAND2_X1 U9187 ( .A1(n11987), .A2(n7261), .ZN(n7868) );
  AND2_X1 U9188 ( .A1(n11541), .A2(n11682), .ZN(n7333) );
  AND2_X2 U9189 ( .A1(n9516), .A2(n9513), .ZN(n15970) );
  OAI22_X1 U9190 ( .A1(n11792), .A2(n11793), .B1(n12043), .B2(n14184), .ZN(
        n11972) );
  INV_X1 U9191 ( .A(n11972), .ZN(n8015) );
  NAND2_X1 U9192 ( .A1(n9654), .A2(n9653), .ZN(n15900) );
  INV_X1 U9193 ( .A(n15900), .ZN(n7586) );
  NAND2_X1 U9194 ( .A1(n7996), .A2(n9093), .ZN(n11655) );
  NAND2_X1 U9195 ( .A1(n10690), .A2(n10691), .ZN(n7334) );
  AND2_X1 U9196 ( .A1(n7868), .A2(n7869), .ZN(n7335) );
  NAND2_X1 U9197 ( .A1(n7225), .A2(n12349), .ZN(n7587) );
  AND2_X1 U9198 ( .A1(n15358), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7336) );
  INV_X1 U9199 ( .A(n8226), .ZN(n7717) );
  INV_X1 U9200 ( .A(n11858), .ZN(n7583) );
  XNOR2_X1 U9201 ( .A(n7438), .B(n9538), .ZN(n15227) );
  INV_X1 U9202 ( .A(n12279), .ZN(n7632) );
  INV_X1 U9203 ( .A(n7885), .ZN(n11345) );
  NAND2_X1 U9204 ( .A1(n7886), .A2(n11385), .ZN(n7885) );
  AND2_X1 U9205 ( .A1(n8676), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7337) );
  INV_X1 U9206 ( .A(n13395), .ZN(n13386) );
  NOR2_X1 U9207 ( .A1(n8999), .A2(n8944), .ZN(n14199) );
  INV_X1 U9208 ( .A(n14199), .ZN(n7464) );
  XOR2_X1 U9209 ( .A(n9420), .B(P2_REG1_REG_19__SCAN_IN), .Z(n7338) );
  AND2_X1 U9210 ( .A1(n8915), .A2(n8025), .ZN(n14562) );
  NAND2_X1 U9211 ( .A1(n7943), .A2(n11053), .ZN(n7339) );
  XOR2_X1 U9212 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n7340) );
  INV_X1 U9213 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U9214 ( .A1(n7342), .A2(n7341), .ZN(n10961) );
  OR2_X1 U9215 ( .A1(n10927), .A2(n13025), .ZN(n7341) );
  NAND2_X1 U9216 ( .A1(n10926), .A2(n10927), .ZN(n7342) );
  NAND2_X1 U9217 ( .A1(n7559), .A2(n10736), .ZN(n10793) );
  NAND2_X4 U9218 ( .A1(n10680), .A2(n15063), .ZN(n13023) );
  NOR2_X1 U9219 ( .A1(n11001), .A2(n8225), .ZN(n14620) );
  NAND2_X1 U9220 ( .A1(n12997), .A2(n8196), .ZN(n7541) );
  NAND2_X2 U9221 ( .A1(n14613), .A2(n14614), .ZN(n14664) );
  AND2_X1 U9222 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9707), .ZN(n9729) );
  INV_X2 U9223 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7345) );
  OR2_X2 U9224 ( .A1(n14677), .A2(n14676), .ZN(n14678) );
  INV_X1 U9225 ( .A(n10001), .ZN(n7348) );
  NAND2_X1 U9226 ( .A1(n9998), .A2(n9997), .ZN(n7349) );
  NAND2_X1 U9227 ( .A1(n9994), .A2(n9993), .ZN(n7350) );
  NAND2_X1 U9228 ( .A1(n7352), .A2(n7351), .ZN(n7988) );
  NAND2_X1 U9229 ( .A1(n10808), .A2(n7170), .ZN(n9695) );
  NAND2_X1 U9230 ( .A1(n10823), .A2(n7170), .ZN(n9748) );
  NAND2_X1 U9231 ( .A1(n10835), .A2(n7170), .ZN(n9685) );
  NAND2_X1 U9232 ( .A1(n10848), .A2(n7170), .ZN(n9771) );
  NAND2_X1 U9233 ( .A1(n10933), .A2(n7170), .ZN(n9665) );
  NAND2_X1 U9234 ( .A1(n11149), .A2(n7170), .ZN(n9797) );
  NAND2_X1 U9235 ( .A1(n10937), .A2(n7170), .ZN(n9654) );
  NAND2_X1 U9236 ( .A1(n11277), .A2(n7170), .ZN(n9645) );
  NAND2_X1 U9237 ( .A1(n11548), .A2(n7170), .ZN(n9813) );
  NAND2_X1 U9238 ( .A1(n11418), .A2(n7170), .ZN(n9786) );
  NAND2_X1 U9239 ( .A1(n11933), .A2(n7170), .ZN(n9825) );
  NAND2_X1 U9240 ( .A1(n12150), .A2(n7170), .ZN(n9834) );
  NAND2_X1 U9241 ( .A1(n12402), .A2(n7170), .ZN(n8102) );
  NAND2_X1 U9242 ( .A1(n12483), .A2(n7170), .ZN(n9601) );
  NAND2_X1 U9243 ( .A1(n12668), .A2(n7170), .ZN(n9590) );
  NAND2_X1 U9244 ( .A1(n12758), .A2(n7170), .ZN(n9868) );
  NAND2_X1 U9245 ( .A1(n14589), .A2(n7170), .ZN(n9857) );
  NAND2_X1 U9246 ( .A1(n12905), .A2(n7170), .ZN(n9848) );
  NAND2_X1 U9247 ( .A1(n14582), .A2(n7170), .ZN(n9572) );
  NAND2_X1 U9248 ( .A1(n14579), .A2(n7170), .ZN(n9564) );
  NAND2_X1 U9249 ( .A1(n14574), .A2(n7170), .ZN(n9550) );
  NAND2_X1 U9250 ( .A1(n14571), .A2(n7170), .ZN(n9881) );
  NAND2_X1 U9251 ( .A1(n14567), .A2(n7170), .ZN(n9892) );
  NAND2_X1 U9252 ( .A1(n14561), .A2(n7170), .ZN(n9541) );
  OAI211_X1 U9253 ( .C1(n10007), .C2(n10008), .A(n7361), .B(n7971), .ZN(n7360)
         );
  NAND2_X1 U9254 ( .A1(n7362), .A2(n10006), .ZN(n7361) );
  NAND2_X1 U9255 ( .A1(n10007), .A2(n10008), .ZN(n7362) );
  NAND3_X1 U9256 ( .A1(n7366), .A2(n10033), .A3(n7365), .ZN(n10036) );
  NAND3_X1 U9257 ( .A1(n10022), .A2(n7964), .A3(n10021), .ZN(n7365) );
  INV_X1 U9258 ( .A(n7964), .ZN(n7367) );
  NAND2_X1 U9259 ( .A1(n9965), .A2(n7957), .ZN(n7368) );
  NAND3_X1 U9260 ( .A1(n7370), .A2(n9964), .A3(n9963), .ZN(n7369) );
  OAI22_X1 U9261 ( .A1(n7377), .A2(n7310), .B1(n7379), .B2(n10055), .ZN(n10076) );
  NAND4_X1 U9262 ( .A1(n7214), .A2(n9621), .A3(n7381), .A4(n10088), .ZN(n7380)
         );
  NAND2_X1 U9263 ( .A1(n7995), .A2(n7214), .ZN(n10087) );
  AND2_X4 U9264 ( .A1(n9621), .A2(n7381), .ZN(n7995) );
  NOR2_X2 U9265 ( .A1(n9692), .A2(n9535), .ZN(n7381) );
  NAND2_X1 U9266 ( .A1(n7988), .A2(n7990), .ZN(n9981) );
  NAND2_X1 U9267 ( .A1(n10036), .A2(n10035), .ZN(n10038) );
  NOR2_X1 U9268 ( .A1(n7453), .A2(n7452), .ZN(n7451) );
  OAI21_X1 U9269 ( .B1(n7268), .B2(n7515), .A(n7976), .ZN(n10007) );
  OR2_X1 U9270 ( .A1(n9953), .A2(n9952), .ZN(n7477) );
  INV_X1 U9271 ( .A(n9382), .ZN(n9383) );
  NAND2_X1 U9272 ( .A1(n9292), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U9273 ( .A1(n8928), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9155) );
  NOR2_X1 U9274 ( .A1(n12835), .A2(n15969), .ZN(n15284) );
  INV_X1 U9275 ( .A(n11262), .ZN(n7422) );
  NOR2_X1 U9276 ( .A1(n15367), .A2(n7621), .ZN(n11928) );
  NAND2_X1 U9277 ( .A1(n11923), .A2(n7613), .ZN(n15369) );
  NOR2_X1 U9278 ( .A1(n12834), .A2(n7619), .ZN(n15283) );
  NOR2_X1 U9279 ( .A1(n15353), .A2(n7336), .ZN(n12618) );
  NAND2_X1 U9280 ( .A1(n10441), .A2(n10440), .ZN(n10446) );
  NAND2_X1 U9281 ( .A1(n7521), .A2(n7519), .ZN(n10457) );
  NAND2_X1 U9282 ( .A1(n10469), .A2(n10468), .ZN(n10473) );
  NAND2_X1 U9283 ( .A1(n8185), .A2(n8186), .ZN(n10522) );
  OAI21_X1 U9284 ( .B1(n7525), .B2(n7524), .A(n8183), .ZN(n10512) );
  NAND2_X1 U9285 ( .A1(n7392), .A2(n7389), .ZN(n10436) );
  OAI21_X1 U9286 ( .B1(n8159), .B2(n10351), .A(n7470), .ZN(n7458) );
  NAND3_X1 U9287 ( .A1(n10425), .A2(n10424), .A3(n7393), .ZN(n7392) );
  NAND2_X1 U9288 ( .A1(n7510), .A2(n7509), .ZN(n7797) );
  AOI21_X1 U9289 ( .B1(n10457), .B2(n10458), .A(n8232), .ZN(n7473) );
  INV_X1 U9290 ( .A(n10335), .ZN(n10345) );
  AND2_X1 U9291 ( .A1(n10336), .A2(n10337), .ZN(n10354) );
  AOI21_X1 U9292 ( .B1(n10446), .B2(n10445), .A(n10444), .ZN(n10447) );
  NAND2_X1 U9293 ( .A1(n10591), .A2(n10588), .ZN(n10589) );
  OAI21_X1 U9294 ( .B1(n8171), .B2(n8170), .A(n8172), .ZN(n10487) );
  NAND2_X1 U9295 ( .A1(n10412), .A2(n10413), .ZN(n7490) );
  INV_X1 U9296 ( .A(n10591), .ZN(n7395) );
  AOI21_X1 U9297 ( .B1(n10473), .B2(n10472), .A(n7459), .ZN(n8170) );
  NAND2_X1 U9298 ( .A1(n8159), .A2(n10351), .ZN(n7396) );
  CLKBUF_X2 U9299 ( .A(n10335), .Z(n10375) );
  NAND3_X1 U9300 ( .A1(n7458), .A2(n10352), .A3(n7396), .ZN(n7435) );
  NAND2_X1 U9301 ( .A1(n9204), .A2(n7295), .ZN(n8017) );
  NAND2_X1 U9302 ( .A1(n9237), .A2(n14411), .ZN(n14402) );
  INV_X1 U9303 ( .A(n8014), .ZN(n8013) );
  OAI21_X1 U9304 ( .B1(n14390), .B2(n8002), .A(n7480), .ZN(n7479) );
  OAI22_X1 U9305 ( .A1(n12381), .A2(n12380), .B1(n12655), .B2(n14180), .ZN(
        n12440) );
  INV_X1 U9306 ( .A(SI_2_), .ZN(n7509) );
  NAND2_X1 U9307 ( .A1(n14686), .A2(n14685), .ZN(n14684) );
  NOR2_X1 U9308 ( .A1(n7692), .A2(n7691), .ZN(n7853) );
  OAI21_X1 U9309 ( .B1(n11972), .B2(n8013), .A(n8011), .ZN(n12522) );
  NAND2_X1 U9310 ( .A1(n9080), .A2(n8872), .ZN(n9095) );
  NAND2_X1 U9311 ( .A1(n8853), .A2(n8982), .ZN(n8986) );
  NAND2_X1 U9312 ( .A1(n7506), .A2(n7503), .ZN(P2_U3496) );
  OR2_X2 U9313 ( .A1(n13403), .A2(n15636), .ZN(n7481) );
  NAND2_X1 U9314 ( .A1(n7948), .A2(n12704), .ZN(n13261) );
  NAND2_X1 U9315 ( .A1(n11135), .A2(n11136), .ZN(n11134) );
  AOI21_X1 U9316 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n11769), .A(n13244), .ZN(
        n11753) );
  NOR2_X1 U9317 ( .A1(n13274), .A2(n13273), .ZN(n13278) );
  NOR2_X1 U9318 ( .A1(n11187), .A2(n11186), .ZN(n13240) );
  AOI21_X1 U9319 ( .B1(n11170), .B2(n11053), .A(n11054), .ZN(n11184) );
  NOR2_X1 U9320 ( .A1(n13347), .A2(n13348), .ZN(n13351) );
  NAND2_X1 U9321 ( .A1(n7399), .A2(n7300), .ZN(n7940) );
  XNOR2_X1 U9322 ( .A(n13380), .B(n13395), .ZN(n13360) );
  NAND2_X1 U9323 ( .A1(n12073), .A2(n12074), .ZN(n7740) );
  NAND2_X2 U9324 ( .A1(n7407), .A2(n8455), .ZN(n12540) );
  OAI21_X2 U9325 ( .B1(n8660), .B2(n7404), .A(n7744), .ZN(n13502) );
  NAND2_X1 U9326 ( .A1(n12730), .A2(n8510), .ZN(n12764) );
  NAND2_X1 U9327 ( .A1(n8718), .A2(n8717), .ZN(n13455) );
  NAND2_X1 U9328 ( .A1(n7940), .A2(n7939), .ZN(n7400) );
  INV_X1 U9329 ( .A(n13381), .ZN(n7399) );
  OAI22_X1 U9330 ( .A1(n13502), .A2(n8687), .B1(n13654), .B2(n13487), .ZN(
        n13481) );
  NAND3_X1 U9331 ( .A1(n7943), .A2(n11053), .A3(P3_REG2_REG_3__SCAN_IN), .ZN(
        n11170) );
  INV_X1 U9332 ( .A(n7400), .ZN(n13405) );
  NAND2_X1 U9333 ( .A1(n7400), .A2(n13404), .ZN(n7401) );
  NOR2_X1 U9334 ( .A1(n13351), .A2(n13350), .ZN(n13358) );
  NOR2_X1 U9335 ( .A1(n13358), .A2(n7496), .ZN(n13380) );
  INV_X1 U9336 ( .A(n15014), .ZN(n7402) );
  NAND2_X1 U9337 ( .A1(n8113), .A2(n7304), .ZN(n11527) );
  OAI21_X1 U9338 ( .B1(n10963), .B2(n13023), .A(n10659), .ZN(n10926) );
  XNOR2_X1 U9339 ( .A(n7457), .B(n7557), .ZN(n14600) );
  OAI21_X1 U9340 ( .B1(n15103), .B2(n15953), .A(n15102), .ZN(n7415) );
  INV_X1 U9341 ( .A(n7415), .ZN(n7414) );
  NAND2_X1 U9342 ( .A1(n8638), .A2(n8637), .ZN(n8650) );
  NAND2_X1 U9343 ( .A1(n8588), .A2(n8587), .ZN(n8601) );
  NAND2_X1 U9344 ( .A1(n8389), .A2(n8388), .ZN(n8391) );
  NAND2_X1 U9345 ( .A1(n8426), .A2(n8425), .ZN(n8428) );
  NAND2_X1 U9346 ( .A1(n8286), .A2(n8285), .ZN(n8426) );
  NAND2_X1 U9347 ( .A1(n7405), .A2(n10278), .ZN(n10263) );
  NAND2_X1 U9348 ( .A1(n13470), .A2(n13454), .ZN(n7405) );
  NAND2_X1 U9349 ( .A1(n8585), .A2(n8584), .ZN(n8588) );
  INV_X1 U9350 ( .A(n8055), .ZN(n8677) );
  NAND2_X1 U9351 ( .A1(n13217), .A2(n15818), .ZN(n10186) );
  INV_X1 U9352 ( .A(n12123), .ZN(n7410) );
  NAND2_X1 U9353 ( .A1(n8332), .A2(n12294), .ZN(n7454) );
  NAND2_X1 U9354 ( .A1(n13621), .A2(n8565), .ZN(n13602) );
  NAND2_X1 U9355 ( .A1(n12764), .A2(n12763), .ZN(n12762) );
  NAND2_X1 U9356 ( .A1(n11823), .A2(n8400), .ZN(n12142) );
  OAI21_X2 U9357 ( .B1(n13573), .B2(n8617), .A(n7406), .ZN(n13558) );
  NAND2_X1 U9358 ( .A1(n7410), .A2(n8451), .ZN(n12297) );
  NAND2_X1 U9359 ( .A1(n8380), .A2(n11818), .ZN(n11823) );
  NAND2_X1 U9360 ( .A1(n12230), .A2(n8450), .ZN(n12120) );
  NAND2_X1 U9361 ( .A1(n12731), .A2(n12806), .ZN(n12730) );
  NAND2_X1 U9362 ( .A1(n13221), .A2(n15723), .ZN(n10159) );
  NAND2_X1 U9363 ( .A1(n12120), .A2(n8454), .ZN(n12457) );
  NAND2_X1 U9364 ( .A1(n12142), .A2(n8401), .ZN(n12073) );
  NAND2_X1 U9365 ( .A1(n12762), .A2(n8523), .ZN(n12818) );
  NAND2_X1 U9366 ( .A1(n12457), .A2(n7408), .ZN(n7407) );
  OR2_X2 U9367 ( .A1(n13455), .A2(n13454), .ZN(n13457) );
  AND2_X1 U9368 ( .A1(n12456), .A2(n12452), .ZN(n7408) );
  INV_X1 U9369 ( .A(n12297), .ZN(n7455) );
  NAND2_X1 U9370 ( .A1(n8469), .A2(n15887), .ZN(n7751) );
  NOR2_X1 U9371 ( .A1(n10140), .A2(n10819), .ZN(n7484) );
  NAND2_X1 U9372 ( .A1(n13529), .A2(n13530), .ZN(n8660) );
  INV_X1 U9373 ( .A(n11301), .ZN(n11941) );
  NAND2_X1 U9374 ( .A1(n15613), .A2(n11764), .ZN(n11765) );
  NOR2_X1 U9375 ( .A1(n13319), .A2(n13318), .ZN(n13336) );
  NOR2_X1 U9376 ( .A1(n13257), .A2(n13256), .ZN(n13259) );
  AOI211_X2 U9377 ( .C1(n13416), .C2(n15638), .A(n13415), .B(n13414), .ZN(
        n13425) );
  NAND2_X1 U9378 ( .A1(n13497), .A2(n8785), .ZN(n13496) );
  NAND2_X1 U9379 ( .A1(n7455), .A2(n8452), .ZN(n12294) );
  NAND2_X1 U9380 ( .A1(n12229), .A2(n12233), .ZN(n8775) );
  NAND2_X1 U9381 ( .A1(n12823), .A2(n12822), .ZN(n12821) );
  NAND2_X1 U9382 ( .A1(n13296), .A2(n13297), .ZN(n13298) );
  XNOR2_X1 U9383 ( .A(n10152), .B(n13412), .ZN(n7441) );
  OAI21_X1 U9384 ( .B1(n14954), .B2(n14965), .A(n12884), .ZN(n14943) );
  NAND2_X1 U9385 ( .A1(n14863), .A2(n9879), .ZN(n14866) );
  NAND2_X1 U9386 ( .A1(n15095), .A2(n15993), .ZN(n7413) );
  NAND2_X1 U9387 ( .A1(n12490), .A2(n12489), .ZN(n12647) );
  NAND2_X1 U9388 ( .A1(n12412), .A2(n12411), .ZN(n12628) );
  INV_X1 U9389 ( .A(n12047), .ZN(n7870) );
  XNOR2_X1 U9390 ( .A(n15283), .B(n15289), .ZN(n12835) );
  NOR2_X1 U9391 ( .A1(n15354), .A2(n15355), .ZN(n15353) );
  NOR2_X1 U9392 ( .A1(n12618), .A2(n12619), .ZN(n12834) );
  NOR2_X1 U9393 ( .A1(n11928), .A2(n11927), .ZN(n12021) );
  NAND2_X1 U9394 ( .A1(n12024), .A2(n12023), .ZN(n12614) );
  NOR2_X1 U9395 ( .A1(n14197), .A2(n14196), .ZN(n14195) );
  NOR2_X1 U9396 ( .A1(n15369), .A2(n15370), .ZN(n15367) );
  NAND2_X1 U9397 ( .A1(n9423), .A2(n10593), .ZN(n15699) );
  NOR2_X1 U9398 ( .A1(n12021), .A2(n7620), .ZN(n12024) );
  NOR2_X1 U9399 ( .A1(n14195), .A2(n7618), .ZN(n14213) );
  AOI21_X2 U9400 ( .B1(n14272), .B2(n14271), .A(n14270), .ZN(n14446) );
  NAND2_X2 U9401 ( .A1(n9460), .A2(n9459), .ZN(n14286) );
  NAND2_X1 U9402 ( .A1(n7429), .A2(n15337), .ZN(n7612) );
  INV_X1 U9403 ( .A(n15338), .ZN(n7429) );
  INV_X1 U9404 ( .A(n13602), .ZN(n7430) );
  XNOR2_X1 U9405 ( .A(n7431), .B(n10635), .ZN(n10633) );
  NAND2_X1 U9406 ( .A1(n10627), .A2(n10628), .ZN(n7431) );
  NAND2_X1 U9407 ( .A1(n12660), .A2(n8492), .ZN(n12731) );
  CLKBUF_X1 U9408 ( .A(n11941), .Z(n7432) );
  OAI21_X1 U9409 ( .B1(n10618), .B2(n10619), .A(n10617), .ZN(n10625) );
  INV_X1 U9410 ( .A(n7473), .ZN(n7434) );
  NAND2_X1 U9411 ( .A1(n7434), .A2(n7272), .ZN(n10464) );
  NAND2_X1 U9412 ( .A1(n7435), .A2(n10357), .ZN(n10363) );
  NAND2_X1 U9413 ( .A1(n7501), .A2(n7275), .ZN(n10452) );
  OAI21_X1 U9414 ( .B1(n7629), .B2(n10583), .A(n9421), .ZN(n10342) );
  NAND2_X1 U9415 ( .A1(n9116), .A2(n8880), .ZN(n8943) );
  OAI22_X1 U9416 ( .A1(n10378), .A2(n10377), .B1(n10380), .B2(n10379), .ZN(
        n10383) );
  OAI21_X1 U9417 ( .B1(n10522), .B2(n10521), .A(n7307), .ZN(n7471) );
  INV_X2 U9418 ( .A(n7476), .ZN(n15686) );
  NAND2_X1 U9419 ( .A1(n13615), .A2(n10232), .ZN(n13594) );
  NAND2_X1 U9420 ( .A1(n8780), .A2(n10249), .ZN(n13527) );
  OAI21_X1 U9421 ( .B1(n8048), .B2(n10324), .A(n10328), .ZN(n8047) );
  INV_X1 U9422 ( .A(n8620), .ZN(n7468) );
  NAND2_X1 U9423 ( .A1(n8570), .A2(n8569), .ZN(n8585) );
  NAND4_X1 U9424 ( .A1(n8247), .A2(n8246), .A3(n7735), .A4(n8551), .ZN(n8749)
         );
  NAND3_X1 U9425 ( .A1(n7751), .A2(n7750), .A3(n7749), .ZN(n12660) );
  NOR2_X1 U9426 ( .A1(n7954), .A2(n7950), .ZN(n13347) );
  AOI21_X1 U9427 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n11185), .A(n11184), .ZN(
        n11187) );
  INV_X1 U9428 ( .A(n10593), .ZN(n15698) );
  INV_X1 U9429 ( .A(n12588), .ZN(n9204) );
  NAND2_X1 U9430 ( .A1(n11632), .A2(n11633), .ZN(n7996) );
  NAND2_X1 U9431 ( .A1(n7479), .A2(n9282), .ZN(n14347) );
  NAND2_X1 U9432 ( .A1(n12291), .A2(n12299), .ZN(n12290) );
  AND4_X2 U9433 ( .A1(n8372), .A2(n8371), .A3(n8370), .A4(n8369), .ZN(n8399)
         );
  NAND2_X1 U9434 ( .A1(n7475), .A2(n8857), .ZN(n8996) );
  NAND2_X1 U9435 ( .A1(n8134), .A2(n8137), .ZN(n12127) );
  NAND2_X1 U9436 ( .A1(n7483), .A2(n8359), .ZN(n11301) );
  INV_X2 U9437 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U9438 ( .A1(n8752), .A2(n8751), .ZN(n8758) );
  NAND2_X1 U9439 ( .A1(n12471), .A2(n12470), .ZN(n7737) );
  INV_X1 U9440 ( .A(n11305), .ZN(n7447) );
  OAI21_X1 U9441 ( .B1(n12775), .B2(n7721), .A(n7718), .ZN(n13040) );
  NAND2_X4 U9442 ( .A1(n11299), .A2(n7245), .ZN(n13103) );
  NAND2_X1 U9443 ( .A1(n7700), .A2(n7706), .ZN(n13179) );
  INV_X1 U9444 ( .A(n13063), .ZN(n7711) );
  INV_X1 U9445 ( .A(n7456), .ZN(n8825) );
  NAND2_X1 U9446 ( .A1(n8802), .A2(n8801), .ZN(n7456) );
  NAND2_X1 U9447 ( .A1(n7499), .A2(n7305), .ZN(n7452) );
  AOI21_X1 U9448 ( .B1(n8877), .B2(n8958), .A(n7660), .ZN(n7659) );
  NAND2_X1 U9449 ( .A1(n14712), .A2(n14715), .ZN(n7457) );
  NAND2_X1 U9450 ( .A1(n7541), .A2(n8198), .ZN(n14713) );
  NAND2_X1 U9451 ( .A1(n8202), .A2(n8205), .ZN(n14677) );
  NOR2_X1 U9452 ( .A1(n10999), .A2(n11000), .ZN(n11001) );
  NAND2_X1 U9453 ( .A1(n11967), .A2(n12792), .ZN(n10334) );
  INV_X1 U9454 ( .A(n10104), .ZN(n7450) );
  NAND2_X1 U9455 ( .A1(n7451), .A2(n7450), .ZN(P1_U3242) );
  NAND2_X1 U9456 ( .A1(n7454), .A2(n8453), .ZN(n12456) );
  NAND2_X1 U9457 ( .A1(n12064), .A2(n12063), .ZN(n12105) );
  NAND2_X1 U9458 ( .A1(n7714), .A2(n7712), .ZN(n13128) );
  NAND2_X1 U9459 ( .A1(n8214), .A2(n11576), .ZN(n7562) );
  NAND2_X1 U9460 ( .A1(n7995), .A2(n7308), .ZN(n9909) );
  AOI21_X1 U9461 ( .B1(n12361), .B2(n12360), .A(n12359), .ZN(n12367) );
  NAND2_X1 U9462 ( .A1(n11679), .A2(n11685), .ZN(n11699) );
  OAI22_X1 U9463 ( .A1(n14912), .A2(n14914), .B1(n14926), .B2(n15128), .ZN(
        n14899) );
  NAND2_X1 U9464 ( .A1(n11553), .A2(n11552), .ZN(n8113) );
  NAND2_X1 U9465 ( .A1(n15036), .A2(n12867), .ZN(n15014) );
  NAND2_X1 U9466 ( .A1(n15053), .A2(n7912), .ZN(n8116) );
  NAND2_X1 U9467 ( .A1(n7237), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8978) );
  NOR2_X2 U9468 ( .A1(n11087), .A2(n9420), .ZN(n11967) );
  NAND2_X1 U9469 ( .A1(n10368), .A2(n10367), .ZN(n10378) );
  NAND4_X1 U9470 ( .A1(n8276), .A2(n7677), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U9471 ( .A1(n9078), .A2(n8085), .ZN(n8082) );
  OAI21_X1 U9472 ( .B1(n7661), .B2(n7665), .A(n7659), .ZN(n8096) );
  AOI21_X1 U9473 ( .B1(n9000), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n7463), .ZN(
        n9001) );
  NOR2_X1 U9474 ( .A1(n8977), .A2(n7464), .ZN(n7463) );
  NAND2_X1 U9475 ( .A1(n8914), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7465) );
  INV_X1 U9476 ( .A(n7467), .ZN(n7466) );
  AOI21_X1 U9477 ( .B1(n8918), .B2(P2_IR_REG_31__SCAN_IN), .A(n8914), .ZN(
        n7467) );
  NAND2_X1 U9478 ( .A1(n8786), .A2(n13104), .ZN(n10106) );
  NAND2_X1 U9479 ( .A1(n10327), .A2(n8049), .ZN(n8048) );
  NAND2_X1 U9480 ( .A1(n8356), .A2(n8277), .ZN(n8374) );
  NAND3_X1 U9481 ( .A1(n8634), .A2(n12484), .A3(n8621), .ZN(n8635) );
  NAND2_X1 U9482 ( .A1(n8028), .A2(n8280), .ZN(n8389) );
  AOI21_X1 U9483 ( .B1(n8125), .B2(n8127), .A(n8123), .ZN(n8122) );
  OAI21_X2 U9484 ( .B1(n8688), .B2(n14591), .A(n8689), .ZN(n8692) );
  NAND2_X1 U9485 ( .A1(n7502), .A2(n8181), .ZN(n10406) );
  NAND2_X1 U9486 ( .A1(n10406), .A2(n10407), .ZN(n10405) );
  NAND2_X1 U9487 ( .A1(n10349), .A2(n10350), .ZN(n7470) );
  OAI21_X1 U9488 ( .B1(n7471), .B2(n7472), .A(n8163), .ZN(n8168) );
  NAND2_X1 U9489 ( .A1(n7489), .A2(n8160), .ZN(n10420) );
  INV_X1 U9490 ( .A(n10399), .ZN(n8182) );
  INV_X1 U9491 ( .A(n8855), .ZN(n7510) );
  CLKBUF_X2 U9492 ( .A(n10334), .Z(n9421) );
  NAND4_X4 U9493 ( .A1(n8978), .A2(n8979), .A3(n8981), .A4(n8980), .ZN(n10348)
         );
  XNOR2_X2 U9494 ( .A(n9545), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9553) );
  INV_X1 U9495 ( .A(n7995), .ZN(n9625) );
  NAND2_X1 U9496 ( .A1(n7905), .A2(n7995), .ZN(n15210) );
  OAI211_X1 U9497 ( .C1(n10076), .C2(n10075), .A(n10074), .B(n10073), .ZN(
        n10104) );
  NAND2_X1 U9498 ( .A1(n13453), .A2(n10260), .ZN(n8786) );
  NAND2_X1 U9499 ( .A1(n8047), .A2(n10333), .ZN(P3_U3296) );
  NAND2_X1 U9500 ( .A1(n8782), .A2(n8155), .ZN(n13497) );
  NAND2_X2 U9501 ( .A1(n12663), .A2(n12773), .ZN(n12735) );
  INV_X1 U9502 ( .A(n11365), .ZN(n15678) );
  AND2_X1 U9503 ( .A1(n8996), .A2(n8995), .ZN(n10804) );
  NAND2_X1 U9504 ( .A1(n8915), .A2(n8914), .ZN(n8917) );
  OAI22_X1 U9505 ( .A1(n14330), .A2(n10607), .B1(n14466), .B2(n14170), .ZN(
        n14321) );
  NAND2_X1 U9506 ( .A1(n7772), .A2(n12703), .ZN(n13249) );
  NAND3_X1 U9507 ( .A1(n13401), .A2(n13402), .A3(n7481), .ZN(P3_U3200) );
  OAI21_X1 U9508 ( .B1(n13231), .B2(n13230), .A(n13229), .ZN(n13233) );
  XNOR2_X2 U9509 ( .A(n8394), .B(n8393), .ZN(n11173) );
  OAI21_X2 U9510 ( .B1(n10633), .B2(n13625), .A(n10632), .ZN(n13436) );
  NAND2_X2 U9511 ( .A1(n13484), .A2(n8703), .ZN(n13469) );
  NOR2_X1 U9512 ( .A1(n7262), .A2(n7484), .ZN(n7483) );
  NAND3_X1 U9513 ( .A1(n10513), .A2(n8239), .A3(n7302), .ZN(n8185) );
  NAND3_X1 U9514 ( .A1(n10409), .A2(n7485), .A3(n7490), .ZN(n7489) );
  NAND2_X1 U9515 ( .A1(n7196), .A2(n10408), .ZN(n7485) );
  NAND2_X1 U9516 ( .A1(n8917), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7627) );
  OAI21_X1 U9517 ( .B1(n8843), .B2(n15892), .A(n7487), .ZN(P3_U3487) );
  OAI21_X2 U9518 ( .B1(n8977), .B2(P2_IR_REG_0__SCAN_IN), .A(n7491), .ZN(
        n11292) );
  NAND2_X1 U9519 ( .A1(n8977), .A2(n14593), .ZN(n7491) );
  NAND3_X1 U9520 ( .A1(n10342), .A2(n10343), .A3(n8237), .ZN(n10347) );
  NAND2_X1 U9521 ( .A1(n10518), .A2(n7332), .ZN(n8186) );
  NOR2_X2 U9522 ( .A1(n10334), .A2(n12669), .ZN(n10335) );
  NAND2_X1 U9523 ( .A1(n12331), .A2(n12332), .ZN(n12333) );
  XNOR2_X1 U9524 ( .A(n13336), .B(n13320), .ZN(n13323) );
  NOR2_X1 U9525 ( .A1(n13298), .A2(n13299), .ZN(n13318) );
  NAND2_X2 U9526 ( .A1(n8919), .A2(n8917), .ZN(n14580) );
  INV_X1 U9527 ( .A(n15611), .ZN(n7507) );
  OAI22_X2 U9528 ( .A1(n14057), .A2(n14055), .B1(n14027), .B2(n14026), .ZN(
        n14110) );
  INV_X1 U9529 ( .A(n9188), .ZN(n8896) );
  INV_X1 U9530 ( .A(n8070), .ZN(n7654) );
  INV_X2 U9531 ( .A(n10806), .ZN(n8863) );
  NAND2_X1 U9532 ( .A1(n7197), .A2(n7520), .ZN(n7519) );
  INV_X1 U9533 ( .A(n10450), .ZN(n7522) );
  INV_X1 U9534 ( .A(n10447), .ZN(n7501) );
  NAND3_X1 U9535 ( .A1(n10395), .A2(n10394), .A3(n7278), .ZN(n7502) );
  NAND2_X1 U9536 ( .A1(n7203), .A2(n8913), .ZN(n8918) );
  NAND2_X1 U9537 ( .A1(n8017), .A2(n8016), .ZN(n14418) );
  NAND2_X1 U9538 ( .A1(n15693), .A2(n15698), .ZN(n15692) );
  NOR2_X1 U9539 ( .A1(n15633), .A2(n12157), .ZN(n12160) );
  NAND2_X1 U9540 ( .A1(n8986), .A2(n8854), .ZN(n8855) );
  NAND2_X2 U9541 ( .A1(n9015), .A2(n8859), .ZN(n9018) );
  INV_X1 U9542 ( .A(n7663), .ZN(n7662) );
  NAND2_X1 U9543 ( .A1(n7523), .A2(n7522), .ZN(n7521) );
  NAND3_X1 U9544 ( .A1(n7512), .A2(n7511), .A3(n7985), .ZN(n7984) );
  NAND2_X1 U9545 ( .A1(n9968), .A2(n9967), .ZN(n7511) );
  NAND2_X1 U9546 ( .A1(n9972), .A2(n9971), .ZN(n7512) );
  NAND3_X1 U9547 ( .A1(n7514), .A2(n7513), .A3(n7982), .ZN(n7981) );
  NAND2_X1 U9548 ( .A1(n10017), .A2(n10016), .ZN(n7513) );
  NAND2_X1 U9549 ( .A1(n10013), .A2(n10012), .ZN(n7514) );
  NAND2_X1 U9550 ( .A1(n10003), .A2(n7974), .ZN(n7515) );
  NAND2_X1 U9551 ( .A1(n10043), .A2(n7314), .ZN(n7979) );
  NAND2_X1 U9552 ( .A1(n10452), .A2(n10451), .ZN(n7523) );
  NAND2_X1 U9553 ( .A1(n10354), .A2(n10353), .ZN(n10352) );
  NAND2_X1 U9554 ( .A1(n10503), .A2(n7311), .ZN(n7525) );
  NAND2_X1 U9555 ( .A1(n7627), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U9556 ( .A1(n10436), .A2(n10437), .ZN(n10435) );
  NAND2_X1 U9557 ( .A1(n10420), .A2(n10421), .ZN(n10419) );
  OR2_X1 U9558 ( .A1(n14832), .A2(n7536), .ZN(n15398) );
  INV_X1 U9559 ( .A(n7535), .ZN(n7536) );
  NAND2_X1 U9560 ( .A1(n7535), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7534) );
  MUX2_X1 U9561 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10863), .S(n10993), .Z(
        n10989) );
  NAND3_X1 U9562 ( .A1(n7539), .A2(n7538), .A3(n7537), .ZN(P1_U3262) );
  OAI211_X1 U9563 ( .C1(n14712), .C2(n7548), .A(n13033), .B(n7546), .ZN(
        P1_U3220) );
  NAND2_X1 U9564 ( .A1(n14712), .A2(n7547), .ZN(n7546) );
  OAI22_X1 U9565 ( .A1(n7552), .A2(n7551), .B1(n13029), .B2(n7554), .ZN(n7550)
         );
  NOR2_X1 U9566 ( .A1(n14595), .A2(n13029), .ZN(n7551) );
  NAND2_X1 U9567 ( .A1(n13022), .A2(n13021), .ZN(n7558) );
  NAND2_X1 U9568 ( .A1(n7562), .A2(n7560), .ZN(n7559) );
  OR2_X1 U9569 ( .A1(n7562), .A2(n7561), .ZN(n11574) );
  INV_X1 U9570 ( .A(n8215), .ZN(n7561) );
  NAND3_X1 U9571 ( .A1(n15063), .A2(n10680), .A3(n10660), .ZN(n10665) );
  INV_X1 U9572 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7578) );
  NAND2_X1 U9573 ( .A1(n11867), .A2(n12213), .ZN(n12013) );
  NAND3_X1 U9574 ( .A1(n7225), .A2(n15926), .A3(n12349), .ZN(n12636) );
  INV_X1 U9575 ( .A(n7587), .ZN(n12427) );
  NAND2_X1 U9576 ( .A1(n7223), .A2(n7588), .ZN(n7592) );
  NOR2_X1 U9577 ( .A1(n7594), .A2(n14915), .ZN(n14886) );
  INV_X1 U9578 ( .A(n14915), .ZN(n7597) );
  OR2_X1 U9579 ( .A1(n15121), .A2(n14915), .ZN(n14902) );
  NAND2_X1 U9580 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7600) );
  NAND2_X1 U9581 ( .A1(n9193), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U9582 ( .A1(n9045), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U9583 ( .A1(n8920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9208) );
  MUX2_X1 U9584 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7601), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9029) );
  NAND2_X1 U9585 ( .A1(n9028), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7601) );
  NAND2_X1 U9586 ( .A1(n8922), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U9587 ( .A1(n9081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U9588 ( .A1(n9497), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9499) );
  MUX2_X1 U9589 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7602), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9137) );
  NAND2_X1 U9590 ( .A1(n9136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9591 ( .A1(n9482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U9592 ( .A1(n9099), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U9593 ( .A1(n9177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9166) );
  MUX2_X1 U9594 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7603), .S(n7469), .Z(n9100)
         );
  NAND2_X1 U9595 ( .A1(n9098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7603) );
  MUX2_X1 U9596 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7604), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9152) );
  NAND2_X1 U9597 ( .A1(n9151), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7604) );
  OAI21_X1 U9598 ( .B1(n9177), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U9599 ( .A1(n9118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U9600 ( .A1(n9490), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9492) );
  OAI21_X1 U9601 ( .B1(n9118), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U9602 ( .A1(n7217), .A2(n11794), .ZN(n12509) );
  NAND2_X1 U9603 ( .A1(n7637), .A2(n7633), .ZN(n14309) );
  INV_X1 U9604 ( .A(n7644), .ZN(n14426) );
  NAND2_X1 U9605 ( .A1(n14295), .A2(n7646), .ZN(n7645) );
  NAND2_X1 U9606 ( .A1(n14295), .A2(n7647), .ZN(n7651) );
  INV_X1 U9607 ( .A(n8877), .ZN(n7661) );
  NAND2_X1 U9608 ( .A1(n7663), .A2(n8877), .ZN(n9115) );
  NAND3_X1 U9609 ( .A1(n7669), .A2(n7667), .A3(n7668), .ZN(n9223) );
  NAND2_X1 U9610 ( .A1(n7666), .A2(n7669), .ZN(n8900) );
  AND2_X1 U9611 ( .A1(n7668), .A2(n7672), .ZN(n7666) );
  AND2_X1 U9612 ( .A1(n7672), .A2(n8899), .ZN(n7667) );
  INV_X1 U9613 ( .A(n8076), .ZN(n7675) );
  INV_X1 U9614 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7679) );
  INV_X1 U9615 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7677) );
  NAND4_X1 U9616 ( .A1(n8275), .A2(n8274), .A3(n7679), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7678) );
  OAI21_X1 U9617 ( .B1(n9241), .B2(n9240), .A(n7685), .ZN(n9255) );
  NAND2_X1 U9618 ( .A1(n9241), .A2(n7686), .ZN(n7680) );
  NAND2_X1 U9619 ( .A1(n13162), .A2(n7695), .ZN(n7694) );
  OAI211_X1 U9620 ( .C1(n13063), .C2(n13162), .A(n7693), .B(n7698), .ZN(n7710)
         );
  NAND2_X1 U9621 ( .A1(n13162), .A2(n13541), .ZN(n7699) );
  AND2_X1 U9622 ( .A1(n7699), .A2(n7711), .ZN(n13144) );
  NAND2_X1 U9623 ( .A1(n13045), .A2(n7715), .ZN(n7714) );
  INV_X1 U9624 ( .A(n11729), .ZN(n7729) );
  NAND2_X1 U9625 ( .A1(n7728), .A2(n11902), .ZN(n7725) );
  INV_X1 U9626 ( .A(n11902), .ZN(n7726) );
  NAND2_X1 U9627 ( .A1(n11903), .A2(n11902), .ZN(n11904) );
  NAND2_X1 U9628 ( .A1(n11724), .A2(n7727), .ZN(n11903) );
  NAND2_X1 U9629 ( .A1(n7737), .A2(n7303), .ZN(n12576) );
  XNOR2_X1 U9630 ( .A(n11365), .B(n13041), .ZN(n11434) );
  NOR2_X2 U9631 ( .A1(n8410), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8298) );
  NAND4_X1 U9632 ( .A1(n8376), .A2(n8157), .A3(n8158), .A4(n8240), .ZN(n8410)
         );
  INV_X1 U9633 ( .A(n7748), .ZN(n7750) );
  NAND2_X1 U9634 ( .A1(n7750), .A2(n7751), .ZN(n12658) );
  NAND2_X1 U9635 ( .A1(n13457), .A2(n8732), .ZN(n8761) );
  NAND3_X1 U9636 ( .A1(n8250), .A2(n8248), .A3(n8249), .ZN(n7755) );
  NAND2_X1 U9637 ( .A1(n11123), .A2(n11061), .ZN(n11139) );
  XNOR2_X2 U9638 ( .A(n7955), .B(n8376), .ZN(n11062) );
  NAND2_X1 U9639 ( .A1(n11138), .A2(n11063), .ZN(n11064) );
  INV_X1 U9640 ( .A(n12176), .ZN(n7761) );
  NAND3_X1 U9641 ( .A1(n7760), .A2(n7762), .A3(n7759), .ZN(n15630) );
  NAND4_X1 U9642 ( .A1(n7760), .A2(n7762), .A3(n7759), .A4(
        P3_REG1_REG_9__SCAN_IN), .ZN(n7765) );
  INV_X1 U9643 ( .A(n7765), .ZN(n15629) );
  INV_X1 U9644 ( .A(n12179), .ZN(n7764) );
  NAND2_X1 U9645 ( .A1(n7769), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7766) );
  INV_X1 U9646 ( .A(n13310), .ZN(n7771) );
  NAND2_X1 U9647 ( .A1(n7775), .A2(n7776), .ZN(n13419) );
  NAND2_X1 U9648 ( .A1(n12087), .A2(n8104), .ZN(n7782) );
  NAND2_X1 U9649 ( .A1(n14964), .A2(n7786), .ZN(n7784) );
  NAND2_X1 U9650 ( .A1(n7800), .A2(n7798), .ZN(n14969) );
  OR2_X2 U9651 ( .A1(n15010), .A2(n7802), .ZN(n7800) );
  NAND3_X1 U9652 ( .A1(n9043), .A2(n9041), .A3(n9042), .ZN(n7805) );
  NAND2_X1 U9653 ( .A1(n14898), .A2(n7807), .ZN(n7809) );
  INV_X1 U9654 ( .A(n7809), .ZN(n14881) );
  NOR2_X1 U9655 ( .A1(n14724), .A2(n14888), .ZN(n7811) );
  NAND3_X1 U9656 ( .A1(n7526), .A2(n14580), .A3(n15257), .ZN(n8990) );
  INV_X1 U9657 ( .A(n11656), .ZN(n9111) );
  NAND2_X1 U9658 ( .A1(n9440), .A2(n7826), .ZN(n7823) );
  NAND2_X1 U9659 ( .A1(n7823), .A2(n7824), .ZN(n12593) );
  NOR2_X1 U9660 ( .A1(n11974), .A2(n7832), .ZN(n7834) );
  INV_X1 U9661 ( .A(n9435), .ZN(n7833) );
  OAI21_X1 U9662 ( .B1(n11789), .B2(n7835), .A(n7834), .ZN(n7836) );
  NAND2_X1 U9663 ( .A1(n12510), .A2(n12511), .ZN(n9438) );
  AOI21_X2 U9664 ( .B1(n14417), .B2(n7837), .A(n7266), .ZN(n14410) );
  OAI21_X2 U9665 ( .B1(n14343), .B2(n7842), .A(n7839), .ZN(n14317) );
  OAI21_X1 U9666 ( .B1(n14286), .B2(n7850), .A(n7846), .ZN(n9465) );
  AND2_X1 U9667 ( .A1(n9479), .A2(n9478), .ZN(n14268) );
  NAND2_X1 U9668 ( .A1(n9444), .A2(n9443), .ZN(n12672) );
  XNOR2_X2 U9669 ( .A(n11104), .B(n11336), .ZN(n11324) );
  AND2_X1 U9670 ( .A1(n9009), .A2(n9424), .ZN(n10593) );
  XNOR2_X2 U9671 ( .A(n8358), .B(P3_IR_REG_1__SCAN_IN), .ZN(n11129) );
  NAND2_X4 U9672 ( .A1(n11096), .A2(n11095), .ZN(n14072) );
  NAND2_X1 U9673 ( .A1(n14042), .A2(n7313), .ZN(n7855) );
  OAI211_X1 U9674 ( .C1(n14042), .C2(n7856), .A(n7855), .B(n14079), .ZN(
        P2_U3192) );
  AND2_X1 U9675 ( .A1(n7869), .A2(n7312), .ZN(n7867) );
  NAND2_X1 U9676 ( .A1(n11344), .A2(n7248), .ZN(n7884) );
  NOR2_X1 U9677 ( .A1(n11109), .A2(n7887), .ZN(n7886) );
  INV_X1 U9678 ( .A(n7888), .ZN(n7887) );
  XNOR2_X2 U9679 ( .A(n9417), .B(n7895), .ZN(n12669) );
  INV_X2 U9680 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7895) );
  OR2_X2 U9681 ( .A1(n9414), .A2(n14563), .ZN(n9417) );
  AND2_X2 U9682 ( .A1(n9408), .A2(n9407), .ZN(n9414) );
  INV_X1 U9683 ( .A(n11861), .ZN(n7901) );
  AND2_X1 U9684 ( .A1(n7214), .A2(n8219), .ZN(n7902) );
  AND2_X1 U9685 ( .A1(n7214), .A2(n7904), .ZN(n7903) );
  AND2_X1 U9686 ( .A1(n8219), .A2(n9536), .ZN(n7904) );
  INV_X1 U9687 ( .A(n7940), .ZN(n13383) );
  INV_X1 U9688 ( .A(n11051), .ZN(n7942) );
  NAND2_X1 U9689 ( .A1(n7942), .A2(n7944), .ZN(n7943) );
  NAND2_X1 U9690 ( .A1(n7339), .A2(n11168), .ZN(n11169) );
  OR2_X1 U9691 ( .A1(n7954), .A2(n7949), .ZN(n13316) );
  INV_X1 U9692 ( .A(n7951), .ZN(n7949) );
  NAND2_X1 U9693 ( .A1(n7951), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7950) );
  INV_X1 U9694 ( .A(n13313), .ZN(n7953) );
  INV_X1 U9695 ( .A(n9966), .ZN(n7957) );
  NAND2_X1 U9696 ( .A1(n10038), .A2(n7961), .ZN(n7960) );
  INV_X1 U9697 ( .A(n10027), .ZN(n7966) );
  OAI21_X2 U9698 ( .B1(n9901), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U9699 ( .A1(n12404), .A2(n10939), .ZN(n7969) );
  INV_X1 U9700 ( .A(n12404), .ZN(n14849) );
  INV_X1 U9701 ( .A(n10044), .ZN(n7980) );
  NAND2_X1 U9702 ( .A1(n7981), .A2(n7983), .ZN(n10023) );
  INV_X1 U9703 ( .A(n9990), .ZN(n7993) );
  NAND2_X1 U9704 ( .A1(n7996), .A2(n7997), .ZN(n15848) );
  NAND2_X1 U9705 ( .A1(n11241), .A2(n7999), .ZN(n11283) );
  XNOR2_X2 U9706 ( .A(n11397), .B(n10348), .ZN(n11285) );
  INV_X1 U9707 ( .A(n9220), .ZN(n8022) );
  NAND2_X1 U9708 ( .A1(n8023), .A2(n8024), .ZN(n9405) );
  NAND2_X1 U9709 ( .A1(n14290), .A2(n7213), .ZN(n8023) );
  OR2_X1 U9710 ( .A1(n14290), .A2(n14289), .ZN(n14292) );
  NAND2_X1 U9711 ( .A1(n8915), .A2(n8027), .ZN(n8933) );
  NAND2_X1 U9712 ( .A1(n8374), .A2(n8279), .ZN(n8028) );
  INV_X1 U9713 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8975) );
  NAND2_X1 U9714 ( .A1(n8635), .A2(n8634), .ZN(n8638) );
  NAND2_X1 U9715 ( .A1(n8692), .A2(n8032), .ZN(n8031) );
  NAND2_X1 U9716 ( .A1(n8692), .A2(n8691), .ZN(n8705) );
  OAI21_X2 U9717 ( .B1(n8526), .B2(n8039), .A(n8036), .ZN(n8567) );
  NAND4_X1 U9718 ( .A1(n10285), .A2(n10298), .A3(n10299), .A4(n7222), .ZN(
        n8056) );
  AND2_X2 U9719 ( .A1(n8748), .A2(n10266), .ZN(n13104) );
  NAND2_X1 U9720 ( .A1(n8063), .A2(n8062), .ZN(n8494) );
  OAI21_X1 U9721 ( .B1(n9018), .B2(n8067), .A(n8066), .ZN(n9062) );
  AOI21_X1 U9722 ( .B1(n8865), .B2(n8073), .A(n8072), .ZN(n8066) );
  INV_X1 U9723 ( .A(n8865), .ZN(n8067) );
  NAND2_X1 U9724 ( .A1(n9018), .A2(n8069), .ZN(n8068) );
  OAI21_X1 U9725 ( .B1(n8865), .B2(n8072), .A(n9061), .ZN(n8070) );
  NAND2_X1 U9726 ( .A1(n8071), .A2(n8865), .ZN(n9044) );
  NAND2_X1 U9727 ( .A1(n9018), .A2(n8860), .ZN(n8071) );
  INV_X1 U9728 ( .A(n8866), .ZN(n8072) );
  OAI21_X1 U9729 ( .B1(n8081), .B2(n8080), .A(n13898), .ZN(n8079) );
  NOR2_X1 U9730 ( .A1(n8898), .A2(SI_17_), .ZN(n8080) );
  NAND2_X1 U9731 ( .A1(n8082), .A2(n8083), .ZN(n8876) );
  NAND2_X1 U9732 ( .A1(n8889), .A2(n8888), .ZN(n9150) );
  NAND2_X1 U9733 ( .A1(n9115), .A2(n9114), .ZN(n9116) );
  OAI21_X1 U9734 ( .B1(n9115), .B2(n8098), .A(n8097), .ZN(n9133) );
  NAND2_X1 U9735 ( .A1(n8096), .A2(n8094), .ZN(n8886) );
  INV_X1 U9736 ( .A(n12353), .ZN(n8105) );
  NAND2_X2 U9737 ( .A1(n14969), .A2(n12870), .ZN(n14964) );
  NAND2_X1 U9738 ( .A1(n12624), .A2(n8111), .ZN(n8110) );
  NAND2_X1 U9739 ( .A1(n8116), .A2(n8114), .ZN(n15036) );
  NAND2_X1 U9740 ( .A1(n8117), .A2(n8363), .ZN(n11739) );
  NAND2_X1 U9741 ( .A1(n8363), .A2(n8119), .ZN(n13224) );
  NAND3_X1 U9742 ( .A1(n8361), .A2(n8360), .A3(n8362), .ZN(n8120) );
  NAND2_X1 U9743 ( .A1(n8121), .A2(n8122), .ZN(n13451) );
  NAND2_X1 U9744 ( .A1(n13480), .A2(n8125), .ZN(n8121) );
  OAI21_X2 U9745 ( .B1(n12735), .B2(n8131), .A(n8128), .ZN(n12823) );
  NAND2_X1 U9746 ( .A1(n8775), .A2(n8135), .ZN(n8134) );
  INV_X1 U9747 ( .A(n10582), .ZN(n8165) );
  NAND2_X1 U9748 ( .A1(n8166), .A2(n8165), .ZN(n8164) );
  NAND2_X1 U9749 ( .A1(n8168), .A2(n8167), .ZN(n8166) );
  INV_X1 U9750 ( .A(n10524), .ZN(n8169) );
  NAND2_X1 U9751 ( .A1(n10497), .A2(n8177), .ZN(n8175) );
  INV_X1 U9752 ( .A(n10506), .ZN(n8184) );
  NAND2_X1 U9753 ( .A1(n14706), .A2(n8203), .ZN(n8202) );
  NAND2_X1 U9754 ( .A1(n14621), .A2(n7306), .ZN(n8215) );
  INV_X1 U9755 ( .A(n10685), .ZN(n8216) );
  INV_X1 U9756 ( .A(n10660), .ZN(n9711) );
  OAI21_X1 U9757 ( .B1(n11502), .B2(n11621), .A(n11501), .ZN(n11835) );
  OAI22_X2 U9758 ( .A1(n14127), .A2(n14125), .B1(n7235), .B2(n14023), .ZN(
        n14024) );
  NAND2_X1 U9759 ( .A1(n13412), .A2(n11787), .ZN(n11298) );
  INV_X1 U9760 ( .A(n13412), .ZN(n10151) );
  NAND4_X2 U9761 ( .A1(n9014), .A2(n9013), .A3(n9012), .A4(n9011), .ZN(n14192)
         );
  NAND2_X1 U9762 ( .A1(n10626), .A2(n13459), .ZN(n10628) );
  INV_X1 U9763 ( .A(n10626), .ZN(n13446) );
  OR2_X1 U9764 ( .A1(n10626), .A2(n13072), .ZN(n8748) );
  AOI21_X2 U9765 ( .B1(n12672), .B2(n12671), .A(n9445), .ZN(n14417) );
  OAI21_X1 U9766 ( .B1(n8495), .B2(n11279), .A(n8511), .ZN(n8496) );
  NAND2_X1 U9767 ( .A1(n8494), .A2(n8493), .ZN(n8495) );
  INV_X1 U9768 ( .A(n10014), .ZN(n10017) );
  AOI21_X2 U9769 ( .B1(n10297), .B2(n10319), .A(n10318), .ZN(n10326) );
  NAND2_X2 U9770 ( .A1(n9553), .A2(n9552), .ZN(n9722) );
  NAND2_X1 U9771 ( .A1(n11504), .A2(n11503), .ZN(n11552) );
  CLKBUF_X1 U9772 ( .A(n12120), .Z(n12296) );
  NAND2_X1 U9773 ( .A1(n8774), .A2(n8773), .ZN(n11816) );
  INV_X1 U9774 ( .A(n11819), .ZN(n8774) );
  NAND2_X1 U9775 ( .A1(n9411), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9413) );
  CLKBUF_X1 U9776 ( .A(n11736), .Z(n11826) );
  NAND2_X1 U9777 ( .A1(n11393), .A2(n9420), .ZN(n15717) );
  INV_X1 U9778 ( .A(n10363), .ZN(n10366) );
  INV_X1 U9779 ( .A(n11511), .ZN(n10657) );
  OR2_X1 U9780 ( .A1(n11572), .A2(n9192), .ZN(n9197) );
  OAI21_X1 U9781 ( .B1(n8850), .B2(n8846), .A(n8845), .ZN(n8848) );
  NAND2_X1 U9782 ( .A1(n8850), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U9783 ( .A1(n10634), .A2(n10287), .ZN(n10150) );
  NAND2_X1 U9784 ( .A1(n8403), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8320) );
  INV_X2 U9785 ( .A(n9157), .ZN(n9398) );
  OAI22_X1 U9786 ( .A1(n7516), .A2(n13024), .B1(n15686), .B2(n7171), .ZN(
        n10673) );
  AND4_X4 U9787 ( .A1(n8320), .A2(n8322), .A3(n8321), .A4(n8323), .ZN(n12302)
         );
  NAND4_X1 U9788 ( .A1(n9008), .A2(n9007), .A3(n9006), .A4(n9005), .ZN(n14193)
         );
  NOR2_X2 U9789 ( .A1(n14568), .A2(n8935), .ZN(n9004) );
  INV_X1 U9790 ( .A(n8260), .ZN(n13036) );
  AND2_X1 U9791 ( .A1(n13435), .A2(n15891), .ZN(n10636) );
  AND2_X2 U9792 ( .A1(n14568), .A2(n8935), .ZN(n9157) );
  OAI222_X1 U9793 ( .A1(P3_U3151), .A2(n7165), .B1(n13993), .B2(n13788), .C1(
        n13888), .C2(n13787), .ZN(P3_U3268) );
  AND2_X1 U9794 ( .A1(n11058), .A2(n7206), .ZN(n13422) );
  NAND3_X1 U9795 ( .A1(n10080), .A2(n10081), .A3(n10079), .ZN(n10099) );
  INV_X1 U9796 ( .A(n9552), .ZN(n15215) );
  AND2_X4 U9797 ( .A1(n10651), .A2(n10714), .ZN(n12999) );
  AND3_X1 U9798 ( .A1(n8229), .A2(n12887), .A3(n9899), .ZN(n8221) );
  INV_X1 U9799 ( .A(n15894), .ZN(n15892) );
  AND2_X2 U9800 ( .A1(n8829), .A2(n8828), .ZN(n15895) );
  AND4_X1 U9801 ( .A1(n9877), .A2(n14914), .A3(n12871), .A4(n14942), .ZN(n8222) );
  OR2_X1 U9802 ( .A1(n8668), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8223) );
  AND2_X1 U9803 ( .A1(n10679), .A2(n10678), .ZN(n8225) );
  AND2_X1 U9804 ( .A1(n13046), .A2(n13626), .ZN(n8226) );
  OR2_X1 U9805 ( .A1(n13446), .A2(n13767), .ZN(n8227) );
  AND2_X1 U9806 ( .A1(n9616), .A2(n9602), .ZN(n8228) );
  AND4_X1 U9807 ( .A1(n9879), .A2(n8234), .A3(n9878), .A4(n8222), .ZN(n8229)
         );
  OR2_X1 U9808 ( .A1(n14868), .A2(n14887), .ZN(n8230) );
  OR2_X1 U9809 ( .A1(n15128), .A2(n14730), .ZN(n8231) );
  INV_X1 U9810 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8846) );
  INV_X1 U9811 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8262) );
  INV_X1 U9812 ( .A(n10216), .ZN(n8777) );
  AND2_X1 U9813 ( .A1(n10456), .A2(n10455), .ZN(n8232) );
  OR2_X2 U9814 ( .A1(n11088), .A2(n7198), .ZN(n8233) );
  XOR2_X2 U9815 ( .A(n15114), .B(n14904), .Z(n8234) );
  OR2_X1 U9816 ( .A1(n13713), .A2(n13712), .ZN(P3_U3454) );
  OR2_X1 U9817 ( .A1(n13466), .A2(n13465), .ZN(P3_U3206) );
  OR2_X1 U9818 ( .A1(n11292), .A2(n11390), .ZN(n8237) );
  INV_X1 U9819 ( .A(n13552), .ZN(n8779) );
  NAND2_X1 U9820 ( .A1(n11392), .A2(n15714), .ZN(n15721) );
  INV_X1 U9821 ( .A(n11854), .ZN(n11863) );
  INV_X2 U9822 ( .A(n15667), .ZN(n15021) );
  INV_X1 U9823 ( .A(n10364), .ZN(n10365) );
  INV_X1 U9824 ( .A(n9982), .ZN(n9983) );
  INV_X1 U9825 ( .A(n10461), .ZN(n10462) );
  INV_X1 U9826 ( .A(n10015), .ZN(n10016) );
  AND2_X1 U9827 ( .A1(n14953), .A2(n10032), .ZN(n10033) );
  INV_X1 U9828 ( .A(n10039), .ZN(n10040) );
  INV_X1 U9829 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8248) );
  INV_X1 U9830 ( .A(n13542), .ZN(n8648) );
  NAND2_X1 U9831 ( .A1(n10317), .A2(n10145), .ZN(n10146) );
  INV_X1 U9832 ( .A(n13631), .ZN(n8564) );
  AND2_X1 U9833 ( .A1(n10560), .A2(n10559), .ZN(n10558) );
  OR2_X1 U9834 ( .A1(n10683), .A2(n10682), .ZN(n10684) );
  XNOR2_X1 U9835 ( .A(n9900), .B(n14849), .ZN(n9922) );
  NOR2_X1 U9836 ( .A1(n10143), .A2(n10296), .ZN(n10149) );
  NAND2_X1 U9837 ( .A1(n10330), .A2(n11820), .ZN(n10276) );
  INV_X1 U9838 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8240) );
  INV_X1 U9839 ( .A(n9294), .ZN(n9292) );
  INV_X1 U9840 ( .A(n9141), .ZN(n8928) );
  XNOR2_X1 U9841 ( .A(n11473), .B(n14191), .ZN(n11479) );
  INV_X1 U9842 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8945) );
  INV_X1 U9843 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9655) );
  OR2_X1 U9844 ( .A1(n12932), .A2(n12931), .ZN(n12933) );
  OR2_X1 U9845 ( .A1(n15121), .A2(n14888), .ZN(n12885) );
  NAND2_X1 U9846 ( .A1(n9711), .A2(n9710), .ZN(n11488) );
  INV_X1 U9847 ( .A(n9253), .ZN(n9256) );
  INV_X1 U9848 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9533) );
  NOR2_X1 U9849 ( .A1(n8534), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8556) );
  NOR2_X1 U9850 ( .A1(n8471), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8503) );
  OR2_X1 U9851 ( .A1(n8517), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8534) );
  NOR2_X1 U9852 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n8223), .ZN(n8697) );
  INV_X1 U9853 ( .A(n7747), .ZN(n8783) );
  INV_X1 U9854 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U9855 ( .A1(n10306), .A2(n11737), .ZN(n11736) );
  INV_X1 U9856 ( .A(n12487), .ZN(n12488) );
  AND2_X1 U9857 ( .A1(n9364), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9382) );
  NAND2_X1 U9858 ( .A1(n9259), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9274) );
  OR2_X1 U9859 ( .A1(n9214), .A2(n8930), .ZN(n9230) );
  XNOR2_X1 U9860 ( .A(n14512), .B(n9203), .ZN(n12592) );
  XNOR2_X1 U9861 ( .A(n15960), .B(n14179), .ZN(n12434) );
  INV_X1 U9862 ( .A(n14604), .ZN(n12929) );
  INV_X1 U9863 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9737) );
  INV_X1 U9864 ( .A(n12917), .ZN(n12918) );
  AND2_X1 U9866 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n9566), .ZN(n9554) );
  OR2_X1 U9867 ( .A1(n9591), .A2(n14698), .ZN(n9869) );
  OR2_X1 U9868 ( .A1(n9836), .A2(n9835), .ZN(n9838) );
  AND2_X1 U9869 ( .A1(n14988), .A2(n14733), .ZN(n12869) );
  INV_X1 U9870 ( .A(n16008), .ZN(n15189) );
  INV_X1 U9871 ( .A(SI_15_), .ZN(n13821) );
  OR2_X1 U9872 ( .A1(n11011), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n15462) );
  OR2_X1 U9873 ( .A1(n8333), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8456) );
  NOR2_X1 U9874 ( .A1(n8611), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8628) );
  INV_X1 U9875 ( .A(n13486), .ZN(n13068) );
  NAND2_X1 U9876 ( .A1(n10326), .A2(n10325), .ZN(n10327) );
  INV_X1 U9877 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15476) );
  AND2_X1 U9878 ( .A1(n11043), .A2(n11072), .ZN(n11058) );
  INV_X1 U9879 ( .A(n10631), .ZN(n10632) );
  INV_X1 U9880 ( .A(n13472), .ZN(n13505) );
  AND2_X1 U9881 ( .A1(n8642), .A2(n8641), .ZN(n8655) );
  INV_X1 U9882 ( .A(n13588), .ZN(n13628) );
  INV_X1 U9883 ( .A(n13627), .ZN(n13609) );
  OR2_X1 U9884 ( .A1(n8838), .A2(n12119), .ZN(n8832) );
  INV_X1 U9885 ( .A(n13771), .ZN(n11315) );
  AND2_X1 U9886 ( .A1(n10151), .A2(n11787), .ZN(n11821) );
  AND2_X1 U9887 ( .A1(n8820), .A2(n10153), .ZN(n13625) );
  INV_X1 U9888 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8822) );
  AND2_X1 U9889 ( .A1(n8618), .A2(n8602), .ZN(n8603) );
  INV_X1 U9890 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8313) );
  OR2_X1 U9891 ( .A1(n11355), .A2(n11343), .ZN(n11344) );
  INV_X1 U9892 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n12497) );
  INV_X1 U9893 ( .A(n14095), .ZN(n14157) );
  AND2_X1 U9894 ( .A1(n10621), .A2(n11390), .ZN(n11106) );
  AND2_X1 U9895 ( .A1(n9383), .A2(n9366), .ZN(n14296) );
  OR2_X1 U9896 ( .A1(n9199), .A2(n9198), .ZN(n9212) );
  OR2_X1 U9897 ( .A1(n11919), .A2(n11920), .ZN(n12028) );
  OR2_X1 U9898 ( .A1(n15365), .A2(n15366), .ZN(n15362) );
  OR2_X1 U9899 ( .A1(n15351), .A2(n15352), .ZN(n15349) );
  AND2_X1 U9900 ( .A1(n15311), .A2(n15310), .ZN(n15320) );
  INV_X1 U9901 ( .A(n14183), .ZN(n12280) );
  INV_X1 U9902 ( .A(n14188), .ZN(n11595) );
  INV_X1 U9903 ( .A(n15917), .ZN(n15940) );
  INV_X1 U9904 ( .A(n15797), .ZN(n15702) );
  OR2_X1 U9905 ( .A1(n9136), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U9906 ( .A1(n12916), .A2(n12918), .ZN(n12919) );
  AND3_X1 U9907 ( .A1(n10714), .A2(n10873), .A3(n10928), .ZN(n10720) );
  OR2_X1 U9908 ( .A1(n9838), .A2(n9614), .ZN(n9616) );
  INV_X1 U9909 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15451) );
  INV_X1 U9910 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15480) );
  INV_X1 U9911 ( .A(n12871), .ZN(n14929) );
  NAND2_X1 U9912 ( .A1(n15021), .A2(n11512), .ZN(n15078) );
  INV_X1 U9913 ( .A(n12887), .ZN(n12872) );
  INV_X1 U9914 ( .A(n15075), .ZN(n15041) );
  INV_X1 U9915 ( .A(n12003), .ZN(n12008) );
  AND2_X1 U9916 ( .A1(n10657), .A2(n10716), .ZN(n15949) );
  OR2_X1 U9917 ( .A1(n12404), .A2(n10719), .ZN(n15656) );
  XNOR2_X1 U9918 ( .A(n8898), .B(SI_17_), .ZN(n9207) );
  XNOR2_X1 U9919 ( .A(n8891), .B(SI_14_), .ZN(n9164) );
  AOI22_X1 U9920 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n11011), .B1(n15463), .B2(
        n15462), .ZN(n15478) );
  OAI21_X1 U9921 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n15498), .A(n15497), .ZN(
        n15507) );
  INV_X1 U9922 ( .A(n13174), .ZN(n13191) );
  AND2_X1 U9923 ( .A1(n11308), .A2(n11307), .ZN(n13172) );
  INV_X1 U9924 ( .A(n13200), .ZN(n13168) );
  INV_X1 U9925 ( .A(n12113), .ZN(n10328) );
  AND4_X1 U9926 ( .A1(n8673), .A2(n8672), .A3(n8671), .A4(n8670), .ZN(n13528)
         );
  AND3_X1 U9927 ( .A1(n8659), .A2(n8658), .A3(n8657), .ZN(n13541) );
  INV_X1 U9928 ( .A(n15641), .ZN(n15618) );
  INV_X1 U9929 ( .A(n13512), .ZN(n13639) );
  INV_X1 U9930 ( .A(n15886), .ZN(n15872) );
  AND3_X1 U9931 ( .A1(n8837), .A2(n8836), .A3(n8835), .ZN(n11318) );
  OR2_X1 U9932 ( .A1(n13556), .A2(n15873), .ZN(n15891) );
  AND2_X1 U9933 ( .A1(n11821), .A2(n12119), .ZN(n15873) );
  INV_X1 U9934 ( .A(n13625), .ZN(n13604) );
  INV_X1 U9935 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8606) );
  AND2_X1 U9936 ( .A1(n8462), .A2(n8343), .ZN(n8344) );
  OR2_X1 U9937 ( .A1(n9496), .A2(n14584), .ZN(n10649) );
  INV_X1 U9938 ( .A(n14092), .ZN(n14155) );
  INV_X1 U9939 ( .A(n12754), .ZN(n10617) );
  AND2_X1 U9940 ( .A1(n10772), .A2(n14575), .ZN(n10767) );
  AND2_X1 U9941 ( .A1(n10772), .A2(n10771), .ZN(n15374) );
  INV_X1 U9942 ( .A(n15364), .ZN(n15333) );
  INV_X1 U9943 ( .A(n10607), .ZN(n14332) );
  AND2_X1 U9944 ( .A1(n15721), .A2(n15713), .ZN(n15807) );
  NAND2_X1 U9945 ( .A1(n15250), .A2(n11090), .ZN(n15714) );
  INV_X1 U9946 ( .A(n15964), .ZN(n15834) );
  INV_X1 U9947 ( .A(n9421), .ZN(n15758) );
  AND2_X1 U9948 ( .A1(n15973), .A2(n15959), .ZN(n14558) );
  INV_X1 U9949 ( .A(n16016), .ZN(n15980) );
  AND2_X1 U9950 ( .A1(n9816), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9826) );
  INV_X1 U9951 ( .A(n16031), .ZN(n14721) );
  AND2_X1 U9952 ( .A1(n10929), .A2(n15949), .ZN(n16027) );
  AND2_X1 U9953 ( .A1(n9588), .A2(n9587), .ZN(n14972) );
  NAND2_X1 U9954 ( .A1(n9893), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9718) );
  OR2_X1 U9955 ( .A1(n15383), .A2(n10985), .ZN(n14812) );
  INV_X1 U9956 ( .A(n14824), .ZN(n15424) );
  INV_X1 U9957 ( .A(n14812), .ZN(n15423) );
  INV_X1 U9958 ( .A(n12362), .ZN(n12565) );
  INV_X1 U9959 ( .A(n15086), .ZN(n15049) );
  INV_X1 U9960 ( .A(n15078), .ZN(n15066) );
  AND2_X1 U9961 ( .A1(n10712), .A2(n10844), .ZN(n11493) );
  AND2_X1 U9962 ( .A1(n15030), .A2(n15029), .ZN(n15182) );
  NAND2_X1 U9963 ( .A1(n10943), .A2(n10942), .ZN(n15993) );
  NAND2_X1 U9964 ( .A1(n15671), .A2(n15773), .ZN(n15998) );
  INV_X1 U9965 ( .A(n11493), .ZN(n11879) );
  INV_X1 U9966 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9536) );
  AND2_X1 U9967 ( .A1(n11073), .A2(n11072), .ZN(n15246) );
  NAND2_X1 U9968 ( .A1(n11221), .A2(n11314), .ZN(n13178) );
  NAND2_X1 U9969 ( .A1(n11214), .A2(n11213), .ZN(n13200) );
  NAND4_X1 U9970 ( .A1(n8731), .A2(n8730), .A3(n8729), .A4(n8728), .ZN(n13473)
         );
  INV_X1 U9971 ( .A(n13575), .ZN(n13207) );
  INV_X1 U9972 ( .A(n15638), .ZN(n13390) );
  INV_X1 U9973 ( .A(n15246), .ZN(n15651) );
  INV_X1 U9974 ( .A(n13422), .ZN(n15631) );
  OR2_X1 U9975 ( .A1(n11057), .A2(n11056), .ZN(n15636) );
  AND2_X1 U9976 ( .A1(n13611), .A2(n13610), .ZN(n13686) );
  AND2_X1 U9977 ( .A1(n12662), .A2(n12661), .ZN(n12796) );
  INV_X1 U9978 ( .A(n12467), .ZN(n13571) );
  NAND2_X1 U9979 ( .A1(n15894), .A2(n15872), .ZN(n13694) );
  AND3_X2 U9980 ( .A1(n8842), .A2(n11318), .A3(n8841), .ZN(n15894) );
  OR2_X1 U9981 ( .A1(n15895), .A2(n15858), .ZN(n13749) );
  AND2_X1 U9982 ( .A1(n15876), .A2(n15875), .ZN(n15878) );
  NAND2_X1 U9983 ( .A1(n10860), .A2(n13772), .ZN(n10861) );
  INV_X1 U9984 ( .A(SI_26_), .ZN(n13812) );
  OR2_X1 U9985 ( .A1(n8489), .A2(n8488), .ZN(n13252) );
  INV_X1 U9986 ( .A(SI_11_), .ZN(n13912) );
  INV_X1 U9987 ( .A(n12117), .ZN(n13995) );
  INV_X1 U9988 ( .A(n14512), .ZN(n12863) );
  AND2_X1 U9989 ( .A1(n11091), .A2(n15714), .ZN(n14135) );
  NAND2_X1 U9990 ( .A1(n11085), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14092) );
  NAND2_X1 U9991 ( .A1(n9372), .A2(n9371), .ZN(n14167) );
  NAND2_X1 U9992 ( .A1(n10767), .A2(n14580), .ZN(n15368) );
  NAND2_X1 U9993 ( .A1(n10767), .A2(n10759), .ZN(n15364) );
  INV_X1 U9994 ( .A(n15271), .ZN(n15377) );
  AND2_X1 U9995 ( .A1(n12439), .A2(n12438), .ZN(n15967) );
  INV_X1 U9996 ( .A(n15807), .ZN(n14369) );
  INV_X1 U9997 ( .A(n15970), .ZN(n15968) );
  INV_X1 U9998 ( .A(n14510), .ZN(n14498) );
  INV_X1 U9999 ( .A(n14323), .ZN(n14535) );
  AND2_X1 U10000 ( .A1(n15967), .A2(n15966), .ZN(n15972) );
  NAND2_X1 U10001 ( .A1(n9516), .A2(n15249), .ZN(n15971) );
  OR2_X1 U10002 ( .A1(n15247), .A2(n15244), .ZN(n15245) );
  AND2_X1 U10003 ( .A1(n11084), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15250) );
  INV_X1 U10004 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12504) );
  INV_X1 U10005 ( .A(n12839), .ZN(n15289) );
  INV_X1 U10006 ( .A(n15141), .ZN(n14949) );
  INV_X1 U10007 ( .A(n12198), .ZN(n12213) );
  INV_X1 U10008 ( .A(n14919), .ZN(n15128) );
  INV_X1 U10009 ( .A(n14988), .ZN(n15161) );
  OR2_X1 U10010 ( .A1(n10724), .A2(n10717), .ZN(n16022) );
  NAND2_X1 U10011 ( .A1(n10722), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16031) );
  NAND2_X1 U10012 ( .A1(n9866), .A2(n9865), .ZN(n14731) );
  INV_X1 U10013 ( .A(n16018), .ZN(n15001) );
  INV_X1 U10014 ( .A(n12423), .ZN(n14736) );
  OR2_X1 U10015 ( .A1(n15383), .A2(n15379), .ZN(n15397) );
  OR2_X1 U10016 ( .A1(n15383), .A2(n10891), .ZN(n15413) );
  INV_X1 U10017 ( .A(n15381), .ZN(n15430) );
  NAND2_X1 U10018 ( .A1(n15021), .A2(n12404), .ZN(n15086) );
  INV_X1 U10019 ( .A(n15034), .ZN(n12432) );
  AND2_X2 U10020 ( .A1(n11880), .A2(n11493), .ZN(n16001) );
  INV_X1 U10021 ( .A(n16005), .ZN(n16002) );
  AND2_X2 U10022 ( .A1(n11880), .A2(n11879), .ZN(n16005) );
  INV_X1 U10023 ( .A(n10713), .ZN(n10846) );
  INV_X1 U10024 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11936) );
  INV_X1 U10025 ( .A(n11893), .ZN(n14811) );
  INV_X1 U10026 ( .A(n15212), .ZN(n15224) );
  AND2_X1 U10027 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10758), .ZN(P2_U3947) );
  NAND2_X1 U10028 ( .A1(n9515), .A2(n9514), .ZN(P2_U3528) );
  NOR2_X1 U10029 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), 
        .ZN(n8247) );
  INV_X1 U10030 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8253) );
  INV_X1 U10031 ( .A(n8256), .ZN(n8257) );
  NAND2_X1 U10032 ( .A1(n8257), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8258) );
  XNOR2_X2 U10033 ( .A(n8259), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8260) );
  AND2_X2 U10034 ( .A1(n13784), .A2(n8260), .ZN(n8382) );
  NAND2_X1 U10035 ( .A1(n8434), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8268) );
  AND2_X2 U10036 ( .A1(n8261), .A2(n13036), .ZN(n8381) );
  NAND2_X1 U10037 ( .A1(n8766), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8267) );
  NOR2_X1 U10038 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8419) );
  NAND2_X1 U10039 ( .A1(n8419), .A2(n8418), .ZN(n8435) );
  NAND2_X1 U10040 ( .A1(n8305), .A2(n8262), .ZN(n8333) );
  OR2_X1 U10041 ( .A1(n8305), .A2(n8262), .ZN(n8263) );
  NAND2_X1 U10042 ( .A1(n8333), .A2(n8263), .ZN(n12479) );
  NAND2_X1 U10043 ( .A1(n8383), .A2(n12479), .ZN(n8266) );
  AND2_X2 U10044 ( .A1(n13784), .A2(n13036), .ZN(n8417) );
  CLKBUF_X1 U10045 ( .A(n8417), .Z(n8264) );
  NAND2_X1 U10046 ( .A1(n8264), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8265) );
  AND4_X2 U10047 ( .A1(n8268), .A2(n8267), .A3(n8266), .A4(n8265), .ZN(n12580)
         );
  INV_X1 U10048 ( .A(n12580), .ZN(n13215) );
  XNOR2_X2 U10049 ( .A(n8270), .B(n8269), .ZN(n12903) );
  NAND2_X1 U10050 ( .A1(n8801), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8271) );
  AND2_X4 U10051 ( .A1(n11042), .A2(n10806), .ZN(n10142) );
  INV_X1 U10052 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10803) );
  NAND2_X1 U10053 ( .A1(n10803), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U10054 ( .A1(n10805), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8280) );
  INV_X1 U10055 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10833) );
  NAND2_X1 U10056 ( .A1(n10833), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8278) );
  NAND2_X1 U10057 ( .A1(n8280), .A2(n8278), .ZN(n8373) );
  INV_X1 U10058 ( .A(n8373), .ZN(n8279) );
  NAND2_X1 U10059 ( .A1(n10810), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8282) );
  INV_X1 U10060 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10829) );
  NAND2_X1 U10061 ( .A1(n10829), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U10062 ( .A1(n8391), .A2(n8282), .ZN(n8409) );
  NAND2_X1 U10063 ( .A1(n10825), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8285) );
  INV_X1 U10064 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10827) );
  NAND2_X1 U10065 ( .A1(n10827), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10066 ( .A1(n8285), .A2(n8283), .ZN(n8408) );
  INV_X1 U10067 ( .A(n8408), .ZN(n8284) );
  NAND2_X1 U10068 ( .A1(n8409), .A2(n8284), .ZN(n8286) );
  NAND2_X1 U10069 ( .A1(n10821), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8288) );
  NAND2_X1 U10070 ( .A1(n10831), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U10071 ( .A1(n8428), .A2(n8288), .ZN(n8443) );
  NAND2_X1 U10072 ( .A1(n7462), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U10073 ( .A1(n8443), .A2(n8289), .ZN(n8291) );
  NAND2_X1 U10074 ( .A1(n10953), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10075 ( .A1(n10851), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U10076 ( .A1(n10850), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8292) );
  NAND2_X1 U10077 ( .A1(n8293), .A2(n8292), .ZN(n8325) );
  INV_X1 U10078 ( .A(n8310), .ZN(n8295) );
  NAND2_X1 U10079 ( .A1(n10855), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10080 ( .A1(n10923), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10081 ( .A1(n10924), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U10082 ( .A1(n8341), .A2(n8297), .ZN(n8339) );
  XNOR2_X1 U10083 ( .A(n8340), .B(n8339), .ZN(n10841) );
  NAND2_X1 U10084 ( .A1(n10142), .A2(n10841), .ZN(n8303) );
  INV_X1 U10085 ( .A(SI_9_), .ZN(n13827) );
  NAND2_X1 U10086 ( .A1(n10112), .A2(n13827), .ZN(n8302) );
  INV_X4 U10087 ( .A(n11042), .ZN(n8608) );
  NAND2_X1 U10088 ( .A1(n8299), .A2(n8429), .ZN(n8444) );
  NAND2_X1 U10089 ( .A1(n8312), .A2(n8313), .ZN(n8346) );
  NAND2_X1 U10090 ( .A1(n8346), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8300) );
  XNOR2_X1 U10091 ( .A(n8300), .B(P3_IR_REG_9__SCAN_IN), .ZN(n12178) );
  INV_X1 U10092 ( .A(n12178), .ZN(n15642) );
  NAND2_X1 U10093 ( .A1(n8608), .A2(n15642), .ZN(n8301) );
  NAND2_X1 U10094 ( .A1(n13215), .A2(n12469), .ZN(n8453) );
  NAND2_X1 U10095 ( .A1(n12580), .A2(n12469), .ZN(n10193) );
  NAND2_X1 U10096 ( .A1(n10193), .A2(n10194), .ZN(n12394) );
  BUF_X4 U10097 ( .A(n8381), .Z(n10125) );
  NAND2_X1 U10098 ( .A1(n10125), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U10099 ( .A1(n8434), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8308) );
  NOR2_X1 U10100 ( .A1(n8318), .A2(n13857), .ZN(n8304) );
  OR2_X1 U10101 ( .A1(n8305), .A2(n8304), .ZN(n12307) );
  NAND2_X1 U10102 ( .A1(n8383), .A2(n12307), .ZN(n8307) );
  NAND2_X1 U10103 ( .A1(n8264), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8306) );
  XNOR2_X1 U10104 ( .A(n8311), .B(n8310), .ZN(n10811) );
  NAND2_X1 U10105 ( .A1(n10112), .A2(SI_8_), .ZN(n8317) );
  OR2_X1 U10106 ( .A1(n8312), .A2(n8549), .ZN(n8314) );
  MUX2_X1 U10107 ( .A(n8314), .B(P3_IR_REG_31__SCAN_IN), .S(n8313), .Z(n8315)
         );
  NAND2_X1 U10108 ( .A1(n8315), .A2(n8346), .ZN(n12174) );
  INV_X1 U10109 ( .A(n12174), .ZN(n12168) );
  NAND2_X1 U10110 ( .A1(n8608), .A2(n12168), .ZN(n8316) );
  INV_X1 U10111 ( .A(n15841), .ZN(n12250) );
  NAND2_X1 U10112 ( .A1(n12247), .A2(n12250), .ZN(n12389) );
  AND2_X1 U10113 ( .A1(n12394), .A2(n12389), .ZN(n8332) );
  NAND2_X1 U10114 ( .A1(n12247), .A2(n15841), .ZN(n10188) );
  NAND2_X1 U10115 ( .A1(n13216), .A2(n12250), .ZN(n10189) );
  AND2_X2 U10116 ( .A1(n10188), .A2(n10189), .ZN(n12299) );
  NAND2_X1 U10117 ( .A1(n8382), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8323) );
  AND2_X1 U10118 ( .A1(n8437), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8319) );
  OR2_X1 U10119 ( .A1(n8319), .A2(n8318), .ZN(n12131) );
  NAND2_X1 U10120 ( .A1(n8383), .A2(n12131), .ZN(n8321) );
  INV_X1 U10121 ( .A(n12302), .ZN(n13217) );
  INV_X1 U10122 ( .A(SI_7_), .ZN(n8324) );
  NAND2_X1 U10123 ( .A1(n10112), .A2(n8324), .ZN(n8331) );
  XNOR2_X1 U10124 ( .A(n8326), .B(n8325), .ZN(n10842) );
  NAND2_X1 U10125 ( .A1(n10142), .A2(n10842), .ZN(n8330) );
  NAND2_X1 U10126 ( .A1(n8327), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8328) );
  INV_X1 U10127 ( .A(n15617), .ZN(n11757) );
  NAND2_X1 U10128 ( .A1(n8608), .A2(n11757), .ZN(n8329) );
  NAND2_X1 U10129 ( .A1(n13217), .A2(n12132), .ZN(n8451) );
  NAND2_X1 U10130 ( .A1(n12302), .A2(n12132), .ZN(n10185) );
  INV_X1 U10131 ( .A(n12132), .ZN(n15818) );
  NAND2_X1 U10132 ( .A1(n8434), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U10133 ( .A1(n10125), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10134 ( .A1(n8333), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U10135 ( .A1(n8456), .A2(n8334), .ZN(n12571) );
  NAND2_X1 U10136 ( .A1(n8765), .A2(n12571), .ZN(n8336) );
  NAND2_X1 U10137 ( .A1(n10126), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U10138 ( .A1(n10935), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U10139 ( .A1(n10951), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8343) );
  OAI21_X1 U10140 ( .B1(n8345), .B2(n8344), .A(n8463), .ZN(n10838) );
  NAND2_X1 U10141 ( .A1(n10142), .A2(n10838), .ZN(n8351) );
  INV_X1 U10142 ( .A(SI_10_), .ZN(n13915) );
  NAND2_X1 U10143 ( .A1(n10112), .A2(n13915), .ZN(n8350) );
  NAND2_X1 U10144 ( .A1(n8464), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10145 ( .A1(n8608), .A2(n12335), .ZN(n8349) );
  NAND2_X1 U10146 ( .A1(n12573), .A2(n15871), .ZN(n10197) );
  INV_X1 U10147 ( .A(n15871), .ZN(n12579) );
  NAND2_X1 U10148 ( .A1(n13214), .A2(n12579), .ZN(n10198) );
  NAND2_X1 U10149 ( .A1(n10197), .A2(n10198), .ZN(n12452) );
  NAND2_X1 U10150 ( .A1(n8383), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8355) );
  NAND2_X1 U10151 ( .A1(n8381), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10152 ( .A1(n8417), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10153 ( .A1(n8382), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8352) );
  INV_X1 U10154 ( .A(SI_1_), .ZN(n10819) );
  OAI21_X1 U10155 ( .B1(n8357), .B2(n8364), .A(n8356), .ZN(n10818) );
  NAND2_X1 U10156 ( .A1(n10142), .A2(n10818), .ZN(n8359) );
  NAND2_X1 U10157 ( .A1(n8368), .A2(n11301), .ZN(n10162) );
  NAND2_X1 U10158 ( .A1(n8383), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U10159 ( .A1(n8381), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10160 ( .A1(n8417), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U10161 ( .A1(n8382), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8360) );
  INV_X1 U10162 ( .A(n8364), .ZN(n8366) );
  INV_X1 U10163 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U10164 ( .A1(n8851), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8365) );
  AND2_X1 U10165 ( .A1(n8366), .A2(n8365), .ZN(n8367) );
  NAND2_X1 U10166 ( .A1(n8863), .A2(SI_0_), .ZN(n8976) );
  OAI21_X1 U10167 ( .B1(n10801), .B2(n8367), .A(n8976), .ZN(n13999) );
  MUX2_X1 U10168 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13999), .S(n11042), .Z(n11447) );
  NAND2_X1 U10169 ( .A1(n13224), .A2(n11447), .ZN(n11737) );
  NAND2_X1 U10170 ( .A1(n11303), .A2(n7432), .ZN(n11825) );
  NAND2_X1 U10171 ( .A1(n11736), .A2(n11825), .ZN(n8380) );
  NAND2_X1 U10172 ( .A1(n8383), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U10173 ( .A1(n8381), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U10174 ( .A1(n8264), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10175 ( .A1(n8382), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8369) );
  INV_X1 U10176 ( .A(n8399), .ZN(n13222) );
  XNOR2_X1 U10177 ( .A(n8374), .B(n8373), .ZN(n10813) );
  NAND2_X1 U10178 ( .A1(n10142), .A2(n10813), .ZN(n8378) );
  NAND2_X1 U10179 ( .A1(n8608), .A2(n7498), .ZN(n8377) );
  NAND2_X1 U10180 ( .A1(n8399), .A2(n11365), .ZN(n10165) );
  NAND2_X1 U10181 ( .A1(n8381), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10182 ( .A1(n8382), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10183 ( .A1(n8417), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8385) );
  INV_X1 U10184 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n13944) );
  NAND2_X1 U10185 ( .A1(n8383), .A2(n13944), .ZN(n8384) );
  AND4_X2 U10186 ( .A1(n8387), .A2(n8386), .A3(n8385), .A4(n8384), .ZN(n8398)
         );
  OR2_X1 U10187 ( .A1(n8389), .A2(n8388), .ZN(n8390) );
  AND2_X1 U10188 ( .A1(n8391), .A2(n8390), .ZN(n10814) );
  NAND2_X1 U10189 ( .A1(n10142), .A2(n10814), .ZN(n8396) );
  NAND2_X1 U10190 ( .A1(n8392), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8394) );
  INV_X1 U10191 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U10192 ( .A1(n8608), .A2(n11173), .ZN(n8395) );
  NAND2_X1 U10193 ( .A1(n8398), .A2(n11443), .ZN(n10166) );
  INV_X1 U10194 ( .A(n11443), .ZN(n15723) );
  NAND2_X1 U10195 ( .A1(n10166), .A2(n10159), .ZN(n12140) );
  NAND2_X1 U10196 ( .A1(n8399), .A2(n15678), .ZN(n12141) );
  NAND2_X1 U10197 ( .A1(n13221), .A2(n11443), .ZN(n8401) );
  NAND2_X1 U10198 ( .A1(n8766), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8407) );
  AND2_X1 U10199 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8402) );
  OR2_X1 U10200 ( .A1(n8402), .A2(n8419), .ZN(n12081) );
  NAND2_X1 U10201 ( .A1(n8383), .A2(n12081), .ZN(n8406) );
  NAND2_X1 U10202 ( .A1(n8434), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U10203 ( .A1(n8403), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8404) );
  NAND4_X1 U10204 ( .A1(n8407), .A2(n8406), .A3(n8405), .A4(n8404), .ZN(n13220) );
  XNOR2_X1 U10205 ( .A(n8409), .B(n8408), .ZN(n10839) );
  NAND2_X1 U10206 ( .A1(n10142), .A2(n10839), .ZN(n8415) );
  INV_X1 U10207 ( .A(n8298), .ZN(n8413) );
  NAND2_X1 U10208 ( .A1(n8410), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8411) );
  MUX2_X1 U10209 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8411), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8412) );
  NAND2_X1 U10210 ( .A1(n8413), .A2(n8412), .ZN(n11185) );
  NAND2_X1 U10211 ( .A1(n8608), .A2(n11185), .ZN(n8414) );
  OAI211_X1 U10212 ( .C1(n7486), .C2(SI_4_), .A(n8415), .B(n8414), .ZN(n15737)
         );
  XNOR2_X1 U10213 ( .A(n13220), .B(n15737), .ZN(n12074) );
  INV_X1 U10214 ( .A(n15737), .ZN(n12082) );
  NAND2_X1 U10215 ( .A1(n13220), .A2(n12082), .ZN(n8416) );
  NAND2_X1 U10216 ( .A1(n10125), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U10217 ( .A1(n8403), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8423) );
  OR2_X1 U10218 ( .A1(n8419), .A2(n8418), .ZN(n8420) );
  NAND2_X1 U10219 ( .A1(n8435), .A2(n8420), .ZN(n12239) );
  NAND2_X1 U10220 ( .A1(n8383), .A2(n12239), .ZN(n8422) );
  NAND2_X1 U10221 ( .A1(n8434), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8421) );
  AND4_X2 U10222 ( .A1(n8424), .A2(n8423), .A3(n8422), .A4(n8421), .ZN(n12217)
         );
  NAND2_X1 U10223 ( .A1(n10112), .A2(n13836), .ZN(n8433) );
  OR2_X1 U10224 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  AND2_X1 U10225 ( .A1(n8428), .A2(n8427), .ZN(n10815) );
  NAND2_X1 U10226 ( .A1(n10142), .A2(n10815), .ZN(n8432) );
  OR2_X1 U10227 ( .A1(n8299), .A2(n8549), .ZN(n8430) );
  XNOR2_X1 U10228 ( .A(n8430), .B(n8429), .ZN(n11759) );
  NAND2_X1 U10229 ( .A1(n8608), .A2(n11759), .ZN(n8431) );
  INV_X1 U10230 ( .A(n12217), .ZN(n13219) );
  INV_X1 U10231 ( .A(n15762), .ZN(n8449) );
  NAND2_X1 U10232 ( .A1(n13219), .A2(n8449), .ZN(n10178) );
  NAND2_X1 U10233 ( .A1(n10125), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U10234 ( .A1(n8434), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U10235 ( .A1(n8435), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U10236 ( .A1(n8437), .A2(n8436), .ZN(n12225) );
  NAND2_X1 U10237 ( .A1(n8383), .A2(n12225), .ZN(n8439) );
  NAND2_X1 U10238 ( .A1(n8403), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8438) );
  INV_X1 U10239 ( .A(SI_6_), .ZN(n13923) );
  XNOR2_X1 U10240 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8442) );
  XNOR2_X1 U10241 ( .A(n8443), .B(n8442), .ZN(n10816) );
  NAND2_X1 U10242 ( .A1(n10142), .A2(n10816), .ZN(n8447) );
  NAND2_X1 U10243 ( .A1(n8444), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8445) );
  XNOR2_X1 U10244 ( .A(n8445), .B(P3_IR_REG_6__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U10245 ( .A1(n8608), .A2(n13236), .ZN(n8446) );
  OAI211_X1 U10246 ( .C1(n7486), .C2(n13923), .A(n8447), .B(n8446), .ZN(n15781) );
  NAND2_X1 U10247 ( .A1(n12236), .A2(n15781), .ZN(n10181) );
  INV_X1 U10248 ( .A(n15781), .ZN(n8448) );
  NAND2_X1 U10249 ( .A1(n13218), .A2(n8448), .ZN(n10182) );
  NAND2_X1 U10250 ( .A1(n10181), .A2(n10182), .ZN(n12218) );
  NAND2_X1 U10251 ( .A1(n12217), .A2(n8449), .ZN(n12219) );
  AND2_X1 U10252 ( .A1(n12218), .A2(n12219), .ZN(n8450) );
  NAND2_X1 U10253 ( .A1(n13218), .A2(n15781), .ZN(n12121) );
  AND2_X1 U10254 ( .A1(n12121), .A2(n8451), .ZN(n12295) );
  INV_X1 U10255 ( .A(n12299), .ZN(n8452) );
  AND2_X1 U10256 ( .A1(n12295), .A2(n8452), .ZN(n12293) );
  AND2_X1 U10257 ( .A1(n12293), .A2(n8453), .ZN(n8454) );
  NAND2_X1 U10258 ( .A1(n13214), .A2(n15871), .ZN(n8455) );
  NAND2_X1 U10259 ( .A1(n10125), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8461) );
  NAND2_X1 U10260 ( .A1(n8456), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10261 ( .A1(n8471), .A2(n8457), .ZN(n12719) );
  NAND2_X1 U10262 ( .A1(n8765), .A2(n12719), .ZN(n8460) );
  NAND2_X1 U10263 ( .A1(n8434), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8459) );
  NAND2_X1 U10264 ( .A1(n10126), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8458) );
  NAND4_X1 U10265 ( .A1(n8461), .A2(n8460), .A3(n8459), .A4(n8458), .ZN(n13213) );
  NAND2_X1 U10266 ( .A1(n12540), .A2(n13213), .ZN(n8469) );
  XNOR2_X1 U10267 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8477) );
  XNOR2_X1 U10268 ( .A(n8479), .B(n8477), .ZN(n10828) );
  NAND2_X1 U10269 ( .A1(n10142), .A2(n10828), .ZN(n8468) );
  OAI21_X1 U10270 ( .B1(n8464), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8466) );
  INV_X1 U10271 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8465) );
  XNOR2_X1 U10272 ( .A(n8466), .B(n8465), .ZN(n12687) );
  NAND2_X1 U10273 ( .A1(n8608), .A2(n12687), .ZN(n8467) );
  OAI211_X1 U10274 ( .C1(n7486), .C2(SI_11_), .A(n8468), .B(n8467), .ZN(n15887) );
  NAND2_X1 U10275 ( .A1(n8434), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10276 ( .A1(n10125), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8475) );
  AND2_X1 U10277 ( .A1(n8471), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8472) );
  OR2_X1 U10278 ( .A1(n8472), .A2(n8503), .ZN(n12783) );
  NAND2_X1 U10279 ( .A1(n8765), .A2(n12783), .ZN(n8474) );
  NAND2_X1 U10280 ( .A1(n10126), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8473) );
  INV_X1 U10281 ( .A(n8477), .ZN(n8478) );
  NAND2_X1 U10282 ( .A1(n11150), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U10283 ( .A1(n11152), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8481) );
  INV_X1 U10284 ( .A(n8482), .ZN(n8483) );
  NAND2_X1 U10285 ( .A1(n7227), .A2(n8483), .ZN(n8484) );
  AND2_X1 U10286 ( .A1(n8494), .A2(n8484), .ZN(n10858) );
  NAND2_X1 U10287 ( .A1(n10858), .A2(n10142), .ZN(n8491) );
  NOR2_X1 U10288 ( .A1(n8485), .A2(n8549), .ZN(n8486) );
  MUX2_X1 U10289 ( .A(n8549), .B(n8486), .S(P3_IR_REG_12__SCAN_IN), .Z(n8489)
         );
  INV_X1 U10290 ( .A(n8487), .ZN(n8488) );
  INV_X1 U10291 ( .A(n13252), .ZN(n12698) );
  AOI22_X1 U10292 ( .A1(n10112), .A2(SI_12_), .B1(n8608), .B2(n12698), .ZN(
        n8490) );
  NAND2_X1 U10293 ( .A1(n8491), .A2(n8490), .ZN(n12788) );
  NAND2_X1 U10294 ( .A1(n12804), .A2(n12788), .ZN(n12734) );
  INV_X1 U10295 ( .A(n12788), .ZN(n12803) );
  NAND2_X1 U10296 ( .A1(n12803), .A2(n13212), .ZN(n10205) );
  NAND2_X1 U10297 ( .A1(n13212), .A2(n12788), .ZN(n8492) );
  NAND2_X1 U10298 ( .A1(n8496), .A2(n11278), .ZN(n8497) );
  NAND2_X1 U10299 ( .A1(n8512), .A2(n8497), .ZN(n10921) );
  NAND2_X1 U10300 ( .A1(n10921), .A2(n10142), .ZN(n8501) );
  INV_X1 U10301 ( .A(SI_13_), .ZN(n13880) );
  NAND2_X1 U10302 ( .A1(n8487), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8498) );
  MUX2_X1 U10303 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8498), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8499) );
  NAND2_X1 U10304 ( .A1(n8499), .A2(n8750), .ZN(n13294) );
  AOI22_X1 U10305 ( .A1(n10112), .A2(n13880), .B1(n8608), .B2(n13294), .ZN(
        n8500) );
  NAND2_X1 U10306 ( .A1(n8434), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10307 ( .A1(n10125), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8507) );
  INV_X1 U10308 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U10309 ( .A1(n8503), .A2(n8502), .ZN(n8517) );
  OR2_X1 U10310 ( .A1(n8503), .A2(n8502), .ZN(n8504) );
  NAND2_X1 U10311 ( .A1(n8517), .A2(n8504), .ZN(n12813) );
  NAND2_X1 U10312 ( .A1(n8765), .A2(n12813), .ZN(n8506) );
  NAND2_X1 U10313 ( .A1(n10126), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U10314 ( .A1(n8509), .A2(n13082), .ZN(n10210) );
  NAND2_X1 U10315 ( .A1(n12833), .A2(n13211), .ZN(n10216) );
  NAND2_X1 U10316 ( .A1(n10210), .A2(n10216), .ZN(n12806) );
  NAND2_X1 U10317 ( .A1(n8509), .A2(n13211), .ZN(n8510) );
  NAND2_X2 U10318 ( .A1(n8512), .A2(n8511), .ZN(n8526) );
  XNOR2_X1 U10319 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8524) );
  XNOR2_X1 U10320 ( .A(n8526), .B(n8524), .ZN(n10932) );
  NAND2_X1 U10321 ( .A1(n10932), .A2(n10142), .ZN(n8516) );
  NAND2_X1 U10322 ( .A1(n8750), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8514) );
  INV_X1 U10323 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8513) );
  XNOR2_X1 U10324 ( .A(n8514), .B(n8513), .ZN(n13305) );
  AOI22_X1 U10325 ( .A1(n10112), .A2(n8092), .B1(n8608), .B2(n13305), .ZN(
        n8515) );
  NAND2_X1 U10326 ( .A1(n8516), .A2(n8515), .ZN(n13702) );
  NAND2_X1 U10327 ( .A1(n10125), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U10328 ( .A1(n8517), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10329 ( .A1(n8534), .A2(n8518), .ZN(n13079) );
  NAND2_X1 U10330 ( .A1(n8765), .A2(n13079), .ZN(n8521) );
  NAND2_X1 U10331 ( .A1(n8558), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U10332 ( .A1(n10126), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8519) );
  NAND4_X1 U10333 ( .A1(n8522), .A2(n8521), .A3(n8520), .A4(n8519), .ZN(n13210) );
  OR2_X1 U10334 ( .A1(n13702), .A2(n13210), .ZN(n10217) );
  NAND2_X1 U10335 ( .A1(n13702), .A2(n13210), .ZN(n10211) );
  NAND2_X1 U10336 ( .A1(n10217), .A2(n10211), .ZN(n12763) );
  INV_X1 U10337 ( .A(n13702), .ZN(n13084) );
  NAND2_X1 U10338 ( .A1(n13084), .A2(n13210), .ZN(n8523) );
  INV_X1 U10339 ( .A(n8524), .ZN(n8525) );
  NAND2_X1 U10340 ( .A1(n11550), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8542) );
  INV_X1 U10341 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U10342 ( .A1(n11549), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U10343 ( .A1(n8542), .A2(n8527), .ZN(n8528) );
  NAND2_X1 U10344 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  AND2_X1 U10345 ( .A1(n8543), .A2(n8530), .ZN(n10955) );
  NAND2_X1 U10346 ( .A1(n10955), .A2(n10142), .ZN(n8533) );
  NAND2_X1 U10347 ( .A1(n8547), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8531) );
  XNOR2_X1 U10348 ( .A(n8531), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U10349 ( .A1(n10112), .A2(SI_15_), .B1(n8608), .B2(n13346), .ZN(
        n8532) );
  NAND2_X1 U10350 ( .A1(n10125), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8540) );
  INV_X1 U10351 ( .A(n8556), .ZN(n8536) );
  NAND2_X1 U10352 ( .A1(n8534), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U10353 ( .A1(n8536), .A2(n8535), .ZN(n13189) );
  NAND2_X1 U10354 ( .A1(n8765), .A2(n13189), .ZN(n8539) );
  INV_X1 U10355 ( .A(n8470), .ZN(n8558) );
  NAND2_X1 U10356 ( .A1(n8558), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10357 ( .A1(n10126), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8537) );
  NAND4_X1 U10358 ( .A1(n8540), .A2(n8539), .A3(n8538), .A4(n8537), .ZN(n13209) );
  NAND2_X1 U10359 ( .A1(n13698), .A2(n13209), .ZN(n10213) );
  NAND2_X1 U10360 ( .A1(n13198), .A2(n13626), .ZN(n10219) );
  NAND2_X1 U10361 ( .A1(n10213), .A2(n10219), .ZN(n12817) );
  NAND2_X1 U10362 ( .A1(n13198), .A2(n13209), .ZN(n8541) );
  NAND2_X1 U10363 ( .A1(n11570), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8566) );
  INV_X1 U10364 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11573) );
  NAND2_X1 U10365 ( .A1(n11573), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8544) );
  OAI21_X1 U10366 ( .B1(n8546), .B2(n8545), .A(n8567), .ZN(n11024) );
  OR2_X1 U10367 ( .A1(n11024), .A2(n8693), .ZN(n8555) );
  NOR2_X1 U10368 ( .A1(n8552), .A2(n8549), .ZN(n8548) );
  MUX2_X1 U10369 ( .A(n8549), .B(n8548), .S(P3_IR_REG_16__SCAN_IN), .Z(n8550)
         );
  INV_X1 U10370 ( .A(n8550), .ZN(n8553) );
  NAND2_X1 U10371 ( .A1(n8553), .A2(n8572), .ZN(n13365) );
  INV_X1 U10372 ( .A(n13365), .ZN(n13341) );
  AOI22_X1 U10373 ( .A1(n10112), .A2(SI_16_), .B1(n8608), .B2(n13341), .ZN(
        n8554) );
  NAND2_X1 U10374 ( .A1(n10125), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8562) );
  NOR2_X1 U10375 ( .A1(n8556), .A2(n13961), .ZN(n8557) );
  OR2_X1 U10376 ( .A1(n8576), .A2(n8557), .ZN(n13633) );
  NAND2_X1 U10377 ( .A1(n8765), .A2(n13633), .ZN(n8561) );
  NAND2_X1 U10378 ( .A1(n8558), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U10379 ( .A1(n10126), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8559) );
  NAND4_X1 U10380 ( .A1(n8562), .A2(n8561), .A3(n8560), .A4(n8559), .ZN(n13608) );
  NAND2_X1 U10381 ( .A1(n13768), .A2(n13608), .ZN(n10225) );
  INV_X1 U10382 ( .A(n13768), .ZN(n8563) );
  NAND2_X1 U10383 ( .A1(n8563), .A2(n13139), .ZN(n10224) );
  NAND2_X1 U10384 ( .A1(n13768), .A2(n13139), .ZN(n8565) );
  NAND2_X1 U10385 ( .A1(n11936), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8584) );
  INV_X1 U10386 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11935) );
  NAND2_X1 U10387 ( .A1(n11935), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8568) );
  OAI21_X1 U10388 ( .B1(n8570), .B2(n8569), .A(n8585), .ZN(n11148) );
  OR2_X1 U10389 ( .A1(n11148), .A2(n8693), .ZN(n8575) );
  NAND2_X1 U10390 ( .A1(n8572), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8571) );
  MUX2_X1 U10391 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8571), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8573) );
  AND2_X1 U10392 ( .A1(n8573), .A2(n7331), .ZN(n13395) );
  AOI22_X1 U10393 ( .A1(n10112), .A2(SI_17_), .B1(n8608), .B2(n13395), .ZN(
        n8574) );
  NAND2_X1 U10394 ( .A1(n10125), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8581) );
  OR2_X1 U10395 ( .A1(n8576), .A2(n13960), .ZN(n8577) );
  NAND2_X1 U10396 ( .A1(n8593), .A2(n8577), .ZN(n13616) );
  NAND2_X1 U10397 ( .A1(n8765), .A2(n13616), .ZN(n8580) );
  NAND2_X1 U10398 ( .A1(n8558), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U10399 ( .A1(n10126), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8578) );
  NAND4_X1 U10400 ( .A1(n8581), .A2(n8580), .A3(n8579), .A4(n8578), .ZN(n13588) );
  NAND2_X1 U10401 ( .A1(n13618), .A2(n13588), .ZN(n10229) );
  NAND2_X1 U10402 ( .A1(n13761), .A2(n13628), .ZN(n10232) );
  NAND2_X1 U10403 ( .A1(n13761), .A2(n13588), .ZN(n8583) );
  NAND2_X1 U10404 ( .A1(n12151), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U10405 ( .A1(n12153), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8586) );
  OR2_X1 U10406 ( .A1(n8588), .A2(n8587), .ZN(n8589) );
  AND2_X1 U10407 ( .A1(n8601), .A2(n8589), .ZN(n11363) );
  NAND2_X1 U10408 ( .A1(n11363), .A2(n10142), .ZN(n8592) );
  NAND2_X1 U10409 ( .A1(n7331), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8590) );
  XNOR2_X1 U10410 ( .A(n8590), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13407) );
  AOI22_X1 U10411 ( .A1(n10112), .A2(SI_18_), .B1(n8608), .B2(n13407), .ZN(
        n8591) );
  NAND2_X1 U10412 ( .A1(n10125), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U10413 ( .A1(n8593), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U10414 ( .A1(n8611), .A2(n8594), .ZN(n13597) );
  NAND2_X1 U10415 ( .A1(n8765), .A2(n13597), .ZN(n8597) );
  NAND2_X1 U10416 ( .A1(n8558), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U10417 ( .A1(n10126), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8595) );
  NAND4_X1 U10418 ( .A1(n8598), .A2(n8597), .A3(n8596), .A4(n8595), .ZN(n13607) );
  NAND2_X1 U10419 ( .A1(n13599), .A2(n13607), .ZN(n10234) );
  NAND2_X1 U10420 ( .A1(n13757), .A2(n13574), .ZN(n10235) );
  NAND2_X1 U10421 ( .A1(n13599), .A2(n13574), .ZN(n8599) );
  INV_X1 U10422 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12403) );
  NAND2_X1 U10423 ( .A1(n12403), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8618) );
  INV_X1 U10424 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12900) );
  NAND2_X1 U10425 ( .A1(n12900), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8602) );
  OR2_X1 U10426 ( .A1(n8604), .A2(n8603), .ZN(n8605) );
  NAND2_X1 U10427 ( .A1(n8619), .A2(n8605), .ZN(n11360) );
  NAND2_X1 U10428 ( .A1(n11360), .A2(n10142), .ZN(n8610) );
  INV_X1 U10429 ( .A(SI_19_), .ZN(n11359) );
  XNOR2_X2 U10430 ( .A(n8607), .B(n8606), .ZN(n13412) );
  AOI22_X1 U10431 ( .A1(n10112), .A2(n11359), .B1(n8608), .B2(n13412), .ZN(
        n8609) );
  NAND2_X1 U10432 ( .A1(n8558), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U10433 ( .A1(n8766), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8615) );
  AND2_X1 U10434 ( .A1(n8611), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8612) );
  OR2_X1 U10435 ( .A1(n8612), .A2(n8628), .ZN(n13580) );
  NAND2_X1 U10436 ( .A1(n8765), .A2(n13580), .ZN(n8614) );
  NAND2_X1 U10437 ( .A1(n10126), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8613) );
  AND2_X1 U10438 ( .A1(n13582), .A2(n13590), .ZN(n8617) );
  NAND2_X1 U10439 ( .A1(n8622), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8623) );
  AND2_X1 U10440 ( .A1(n8635), .A2(n8623), .ZN(n11786) );
  NAND2_X1 U10441 ( .A1(n11786), .A2(n10142), .ZN(n8625) );
  NAND2_X1 U10442 ( .A1(n10112), .A2(SI_20_), .ZN(n8624) );
  NAND2_X1 U10443 ( .A1(n10125), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U10444 ( .A1(n10126), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8626) );
  AND2_X1 U10445 ( .A1(n8627), .A2(n8626), .ZN(n8632) );
  NOR2_X1 U10446 ( .A1(n8628), .A2(n13971), .ZN(n8629) );
  OR2_X1 U10447 ( .A1(n8642), .A2(n8629), .ZN(n13567) );
  NAND2_X1 U10448 ( .A1(n13567), .A2(n8765), .ZN(n8631) );
  NAND2_X1 U10449 ( .A1(n8558), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8630) );
  OR2_X1 U10450 ( .A1(n13746), .A2(n13575), .ZN(n10246) );
  NAND2_X1 U10451 ( .A1(n13746), .A2(n13575), .ZN(n10245) );
  NAND2_X1 U10452 ( .A1(n10246), .A2(n10245), .ZN(n13552) );
  NAND2_X1 U10453 ( .A1(n13746), .A2(n13207), .ZN(n8633) );
  INV_X1 U10454 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12727) );
  NAND2_X1 U10455 ( .A1(n12727), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8649) );
  INV_X1 U10456 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12670) );
  NAND2_X1 U10457 ( .A1(n12670), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8636) );
  OAI21_X1 U10458 ( .B1(n8638), .B2(n8637), .A(n8650), .ZN(n11901) );
  OR2_X1 U10459 ( .A1(n11901), .A2(n8693), .ZN(n8640) );
  NAND2_X1 U10460 ( .A1(n10112), .A2(SI_21_), .ZN(n8639) );
  INV_X1 U10461 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8641) );
  NOR2_X1 U10462 ( .A1(n8642), .A2(n8641), .ZN(n8643) );
  OR2_X1 U10463 ( .A1(n8655), .A2(n8643), .ZN(n13549) );
  NAND2_X1 U10464 ( .A1(n13549), .A2(n8765), .ZN(n8646) );
  AOI22_X1 U10465 ( .A1(n10125), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n8558), 
        .B2(P3_REG2_REG_21__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U10466 ( .A1(n10126), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U10467 ( .A1(n13120), .A2(n13560), .ZN(n13530) );
  NAND2_X1 U10468 ( .A1(n13740), .A2(n13206), .ZN(n8647) );
  NAND2_X2 U10469 ( .A1(n8650), .A2(n8649), .ZN(n8664) );
  INV_X1 U10470 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U10471 ( .A1(n8651), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8665) );
  INV_X1 U10472 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12794) );
  NAND2_X1 U10473 ( .A1(n12794), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U10474 ( .A1(n8665), .A2(n8652), .ZN(n8662) );
  XNOR2_X1 U10475 ( .A(n8664), .B(n8662), .ZN(n12116) );
  NAND2_X1 U10476 ( .A1(n12116), .A2(n10142), .ZN(n8654) );
  NAND2_X1 U10477 ( .A1(n10112), .A2(SI_22_), .ZN(n8653) );
  OR2_X1 U10478 ( .A1(n8655), .A2(n13972), .ZN(n8656) );
  NAND2_X1 U10479 ( .A1(n8656), .A2(n8668), .ZN(n13537) );
  NAND2_X1 U10480 ( .A1(n13537), .A2(n8765), .ZN(n8659) );
  AOI22_X1 U10481 ( .A1(n10125), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n8558), 
        .B2(P3_REG2_REG_22__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U10482 ( .A1(n10126), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8657) );
  OR2_X1 U10483 ( .A1(n13734), .A2(n13541), .ZN(n10253) );
  NAND2_X1 U10484 ( .A1(n13734), .A2(n13541), .ZN(n10254) );
  NAND2_X1 U10485 ( .A1(n10253), .A2(n10254), .ZN(n8781) );
  INV_X1 U10486 ( .A(n13541), .ZN(n13205) );
  OR2_X1 U10487 ( .A1(n13734), .A2(n13205), .ZN(n8661) );
  INV_X1 U10488 ( .A(n8662), .ZN(n8663) );
  INV_X1 U10489 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8676) );
  XNOR2_X1 U10490 ( .A(n8676), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n8674) );
  XNOR2_X1 U10491 ( .A(n8675), .B(n8674), .ZN(n12112) );
  NAND2_X1 U10492 ( .A1(n12112), .A2(n10142), .ZN(n8667) );
  NAND2_X1 U10493 ( .A1(n10112), .A2(SI_23_), .ZN(n8666) );
  NAND2_X2 U10494 ( .A1(n8667), .A2(n8666), .ZN(n13657) );
  NAND2_X1 U10495 ( .A1(n10125), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8673) );
  NAND2_X1 U10496 ( .A1(n8558), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U10497 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(n8668), .ZN(n8669) );
  NAND2_X1 U10498 ( .A1(n8669), .A2(n8223), .ZN(n13519) );
  NAND2_X1 U10499 ( .A1(n8765), .A2(n13519), .ZN(n8671) );
  NAND2_X1 U10500 ( .A1(n10126), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8670) );
  OR2_X2 U10501 ( .A1(n13657), .A2(n13528), .ZN(n13499) );
  NAND2_X1 U10502 ( .A1(n13657), .A2(n13528), .ZN(n10271) );
  INV_X1 U10503 ( .A(n13528), .ZN(n13204) );
  INV_X1 U10504 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n15234) );
  INV_X1 U10505 ( .A(n8677), .ZN(n8678) );
  NAND2_X1 U10506 ( .A1(n8678), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U10507 ( .A1(n8689), .A2(n8679), .ZN(n8688) );
  XNOR2_X1 U10508 ( .A(n8688), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n12505) );
  NAND2_X1 U10509 ( .A1(n12505), .A2(n10142), .ZN(n8681) );
  NAND2_X1 U10510 ( .A1(n10112), .A2(SI_24_), .ZN(n8680) );
  NAND2_X1 U10511 ( .A1(n10125), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8686) );
  NAND2_X1 U10512 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n8223), .ZN(n8682) );
  INV_X1 U10513 ( .A(n8697), .ZN(n8696) );
  NAND2_X1 U10514 ( .A1(n8682), .A2(n8696), .ZN(n13506) );
  NAND2_X1 U10515 ( .A1(n8765), .A2(n13506), .ZN(n8685) );
  NAND2_X1 U10516 ( .A1(n8558), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U10517 ( .A1(n10126), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8683) );
  NAND4_X1 U10518 ( .A1(n8686), .A2(n8685), .A3(n8684), .A4(n8683), .ZN(n13487) );
  AND2_X1 U10519 ( .A1(n13654), .A2(n13487), .ZN(n8687) );
  INV_X1 U10520 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n14591) );
  INV_X1 U10521 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12907) );
  NAND2_X1 U10522 ( .A1(n12907), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8704) );
  INV_X1 U10523 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14588) );
  NAND2_X1 U10524 ( .A1(n14588), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8690) );
  AND2_X1 U10525 ( .A1(n8704), .A2(n8690), .ZN(n8691) );
  OAI21_X1 U10526 ( .B1(n8692), .B2(n8691), .A(n8705), .ZN(n13992) );
  NAND2_X1 U10527 ( .A1(n10112), .A2(SI_25_), .ZN(n8694) );
  NAND2_X2 U10528 ( .A1(n8695), .A2(n8694), .ZN(n13493) );
  INV_X1 U10529 ( .A(n13493), .ZN(n13720) );
  NAND2_X1 U10530 ( .A1(n8766), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U10531 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(n8696), .ZN(n8698) );
  INV_X1 U10532 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n13957) );
  NAND2_X1 U10533 ( .A1(n8697), .A2(n13957), .ZN(n8709) );
  NAND2_X1 U10534 ( .A1(n8698), .A2(n8709), .ZN(n13492) );
  NAND2_X1 U10535 ( .A1(n8765), .A2(n13492), .ZN(n8701) );
  NAND2_X1 U10536 ( .A1(n8558), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8700) );
  NAND2_X1 U10537 ( .A1(n10126), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8699) );
  NAND4_X1 U10538 ( .A1(n8702), .A2(n8701), .A3(n8700), .A4(n8699), .ZN(n13472) );
  NAND2_X1 U10539 ( .A1(n13720), .A2(n13472), .ZN(n10265) );
  NAND2_X1 U10540 ( .A1(n13493), .A2(n13505), .ZN(n10273) );
  OR2_X2 U10541 ( .A1(n13481), .A2(n13482), .ZN(n13484) );
  NAND2_X1 U10542 ( .A1(n13493), .A2(n13472), .ZN(n8703) );
  INV_X1 U10543 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15230) );
  NAND2_X1 U10544 ( .A1(n15230), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8722) );
  INV_X1 U10545 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14583) );
  NAND2_X1 U10546 ( .A1(n14583), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U10547 ( .A1(n8722), .A2(n8706), .ZN(n8719) );
  NAND2_X1 U10548 ( .A1(n12743), .A2(n10142), .ZN(n8708) );
  NAND2_X1 U10549 ( .A1(n10112), .A2(SI_26_), .ZN(n8707) );
  NAND2_X1 U10550 ( .A1(n10125), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U10551 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n8709), .ZN(n8711) );
  INV_X1 U10552 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n13982) );
  INV_X1 U10553 ( .A(n8709), .ZN(n8710) );
  NAND2_X1 U10554 ( .A1(n13982), .A2(n8710), .ZN(n8726) );
  NAND2_X1 U10555 ( .A1(n8711), .A2(n8726), .ZN(n13477) );
  NAND2_X1 U10556 ( .A1(n8765), .A2(n13477), .ZN(n8714) );
  NAND2_X1 U10557 ( .A1(n8558), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U10558 ( .A1(n10126), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8712) );
  NAND4_X1 U10559 ( .A1(n8715), .A2(n8714), .A3(n8713), .A4(n8712), .ZN(n13486) );
  OR2_X1 U10560 ( .A1(n13647), .A2(n13486), .ZN(n8716) );
  NAND2_X1 U10561 ( .A1(n13469), .A2(n8716), .ZN(n8718) );
  NAND2_X1 U10562 ( .A1(n13647), .A2(n13486), .ZN(n8717) );
  INV_X1 U10563 ( .A(n8719), .ZN(n8720) );
  INV_X1 U10564 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15225) );
  NAND2_X1 U10565 ( .A1(n15225), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8736) );
  INV_X1 U10566 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14581) );
  NAND2_X1 U10567 ( .A1(n14581), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U10568 ( .A1(n8736), .A2(n8723), .ZN(n8733) );
  XNOR2_X1 U10569 ( .A(n8735), .B(n8733), .ZN(n13786) );
  NAND2_X1 U10570 ( .A1(n13786), .A2(n10142), .ZN(n8725) );
  NAND2_X1 U10571 ( .A1(n10112), .A2(SI_27_), .ZN(n8724) );
  NAND2_X2 U10572 ( .A1(n8725), .A2(n8724), .ZN(n13463) );
  NAND2_X1 U10573 ( .A1(n10125), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U10574 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n8726), .ZN(n8727) );
  NOR2_X1 U10575 ( .A1(n8726), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8740) );
  INV_X1 U10576 ( .A(n8740), .ZN(n8742) );
  NAND2_X1 U10577 ( .A1(n8727), .A2(n8742), .ZN(n13462) );
  NAND2_X1 U10578 ( .A1(n8765), .A2(n13462), .ZN(n8730) );
  NAND2_X1 U10579 ( .A1(n8558), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U10580 ( .A1(n10126), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8728) );
  OR2_X1 U10581 ( .A1(n13463), .A2(n13473), .ZN(n8732) );
  INV_X1 U10582 ( .A(n8733), .ZN(n8734) );
  NAND2_X1 U10583 ( .A1(n8735), .A2(n8734), .ZN(n8737) );
  INV_X1 U10584 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15221) );
  XNOR2_X1 U10585 ( .A(n15221), .B(P1_DATAO_REG_28__SCAN_IN), .ZN(n10107) );
  XNOR2_X1 U10586 ( .A(n10109), .B(n10107), .ZN(n12901) );
  NAND2_X1 U10587 ( .A1(n12901), .A2(n10142), .ZN(n8739) );
  NAND2_X1 U10588 ( .A1(n10112), .A2(SI_28_), .ZN(n8738) );
  NAND2_X1 U10589 ( .A1(n10125), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U10590 ( .A1(n10126), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8746) );
  INV_X1 U10591 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U10592 ( .A1(n8741), .A2(n8740), .ZN(n8764) );
  NAND2_X1 U10593 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(n8742), .ZN(n8743) );
  NAND2_X1 U10594 ( .A1(n8764), .A2(n8743), .ZN(n13444) );
  NAND2_X1 U10595 ( .A1(n8765), .A2(n13444), .ZN(n8745) );
  NAND2_X1 U10596 ( .A1(n8558), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U10597 ( .A1(n10626), .A2(n13072), .ZN(n10266) );
  NAND2_X1 U10598 ( .A1(n8761), .A2(n13104), .ZN(n8760) );
  NAND2_X1 U10599 ( .A1(n8821), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U10600 ( .A1(n10151), .A2(n10330), .ZN(n8820) );
  NAND2_X1 U10601 ( .A1(n8758), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8754) );
  MUX2_X1 U10602 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8754), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8755) );
  AND2_X2 U10603 ( .A1(n8755), .A2(n8821), .ZN(n11820) );
  NAND2_X1 U10604 ( .A1(n8756), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8757) );
  MUX2_X1 U10605 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8757), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8759) );
  NAND2_X1 U10606 ( .A1(n8759), .A2(n8758), .ZN(n11787) );
  INV_X1 U10607 ( .A(n11787), .ZN(n8819) );
  NAND2_X1 U10608 ( .A1(n11820), .A2(n8819), .ZN(n10153) );
  NAND2_X1 U10609 ( .A1(n8760), .A2(n13604), .ZN(n8763) );
  INV_X1 U10610 ( .A(n10627), .ZN(n8762) );
  INV_X1 U10611 ( .A(n8764), .ZN(n13430) );
  NAND2_X1 U10612 ( .A1(n8765), .A2(n13430), .ZN(n10130) );
  NAND2_X1 U10613 ( .A1(n8766), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U10614 ( .A1(n10126), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U10615 ( .A1(n8558), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8767) );
  INV_X1 U10616 ( .A(n13108), .ZN(n13203) );
  INV_X1 U10617 ( .A(n12903), .ZN(n11044) );
  INV_X1 U10618 ( .A(n7206), .ZN(n10329) );
  NAND2_X1 U10619 ( .A1(n11044), .A2(n10329), .ZN(n11056) );
  NAND2_X1 U10620 ( .A1(n11042), .A2(n11056), .ZN(n8770) );
  INV_X1 U10621 ( .A(n8770), .ZN(n11307) );
  AOI22_X1 U10622 ( .A1(n13203), .A2(n13606), .B1(n13609), .B2(n13473), .ZN(
        n8771) );
  NAND2_X1 U10623 ( .A1(n8772), .A2(n10157), .ZN(n11819) );
  NAND2_X1 U10624 ( .A1(n11816), .A2(n10165), .ZN(n12139) );
  INV_X1 U10625 ( .A(n12140), .ZN(n12138) );
  NAND2_X1 U10626 ( .A1(n12139), .A2(n12138), .ZN(n12137) );
  NAND2_X1 U10627 ( .A1(n12137), .A2(n10166), .ZN(n12070) );
  NAND2_X1 U10628 ( .A1(n12070), .A2(n12069), .ZN(n12072) );
  INV_X1 U10629 ( .A(n13220), .ZN(n12235) );
  NAND2_X1 U10630 ( .A1(n12235), .A2(n12082), .ZN(n10174) );
  NAND2_X1 U10631 ( .A1(n12072), .A2(n10174), .ZN(n12229) );
  INV_X1 U10632 ( .A(n12218), .ZN(n12215) );
  INV_X1 U10633 ( .A(n12123), .ZN(n12124) );
  NAND2_X1 U10634 ( .A1(n12127), .A2(n10185), .ZN(n12291) );
  INV_X1 U10635 ( .A(n10188), .ZN(n12385) );
  NOR2_X1 U10636 ( .A1(n12394), .A2(n12385), .ZN(n8776) );
  INV_X1 U10637 ( .A(n13213), .ZN(n12786) );
  INV_X1 U10638 ( .A(n15887), .ZN(n12776) );
  NAND2_X1 U10639 ( .A1(n12786), .A2(n12776), .ZN(n10202) );
  NAND2_X1 U10640 ( .A1(n13213), .A2(n15887), .ZN(n12778) );
  AND2_X1 U10641 ( .A1(n12734), .A2(n10210), .ZN(n8778) );
  INV_X1 U10642 ( .A(n12763), .ZN(n12768) );
  NAND2_X1 U10643 ( .A1(n12821), .A2(n10219), .ZN(n13632) );
  NAND2_X1 U10644 ( .A1(n13632), .A2(n13631), .ZN(n13630) );
  NAND2_X1 U10645 ( .A1(n13630), .A2(n10224), .ZN(n13613) );
  NAND2_X1 U10646 ( .A1(n13613), .A2(n13612), .ZN(n13615) );
  INV_X1 U10647 ( .A(n13582), .ZN(n13753) );
  INV_X1 U10648 ( .A(n13590), .ZN(n13208) );
  NAND2_X1 U10649 ( .A1(n13582), .A2(n13208), .ZN(n10300) );
  NAND2_X1 U10650 ( .A1(n13540), .A2(n13542), .ZN(n8780) );
  NAND2_X1 U10651 ( .A1(n13740), .A2(n13560), .ZN(n10249) );
  NAND2_X1 U10652 ( .A1(n13527), .A2(n7745), .ZN(n8782) );
  OR2_X1 U10653 ( .A1(n13654), .A2(n13515), .ZN(n10264) );
  NAND2_X1 U10654 ( .A1(n13654), .A2(n13515), .ZN(n10272) );
  NAND2_X1 U10655 ( .A1(n10264), .A2(n10272), .ZN(n13503) );
  INV_X1 U10656 ( .A(n13499), .ZN(n8784) );
  NOR2_X1 U10657 ( .A1(n13503), .A2(n8784), .ZN(n8785) );
  NAND2_X1 U10658 ( .A1(n13647), .A2(n13068), .ZN(n10259) );
  NAND2_X1 U10659 ( .A1(n13451), .A2(n13454), .ZN(n13453) );
  INV_X1 U10660 ( .A(n13473), .ZN(n13100) );
  NAND2_X1 U10661 ( .A1(n13463), .A2(n13100), .ZN(n10260) );
  OR2_X1 U10662 ( .A1(n8786), .A2(n13104), .ZN(n8787) );
  NAND2_X1 U10663 ( .A1(n10106), .A2(n8787), .ZN(n13448) );
  NAND2_X1 U10664 ( .A1(n11298), .A2(n8820), .ZN(n8838) );
  INV_X1 U10665 ( .A(n10330), .ZN(n12119) );
  NAND2_X1 U10666 ( .A1(n13412), .A2(n11900), .ZN(n8790) );
  AND2_X1 U10667 ( .A1(n11900), .A2(n11787), .ZN(n8840) );
  INV_X1 U10668 ( .A(n8840), .ZN(n8788) );
  XNOR2_X1 U10669 ( .A(n10330), .B(n8788), .ZN(n8789) );
  NAND2_X1 U10670 ( .A1(n8790), .A2(n8789), .ZN(n11208) );
  INV_X1 U10671 ( .A(n11298), .ZN(n10325) );
  NAND3_X1 U10672 ( .A1(n11208), .A2(n10325), .A3(n15886), .ZN(n8791) );
  AND2_X1 U10673 ( .A1(n13448), .A2(n15891), .ZN(n8792) );
  INV_X1 U10674 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U10675 ( .A1(n8793), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8794) );
  MUX2_X1 U10676 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8794), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8796) );
  NAND2_X1 U10677 ( .A1(n8796), .A2(n8795), .ZN(n12507) );
  XNOR2_X1 U10678 ( .A(n12507), .B(P3_B_REG_SCAN_IN), .ZN(n8799) );
  NAND2_X1 U10679 ( .A1(n8795), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8797) );
  MUX2_X1 U10680 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8797), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8798) );
  NAND2_X1 U10681 ( .A1(n8798), .A2(n8144), .ZN(n13996) );
  NAND2_X1 U10682 ( .A1(n8144), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8800) );
  MUX2_X1 U10683 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8800), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8802) );
  INV_X1 U10684 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8803) );
  INV_X1 U10685 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8804) );
  NAND2_X1 U10686 ( .A1(n8807), .A2(n8804), .ZN(n8806) );
  NAND2_X1 U10687 ( .A1(n7456), .A2(n13996), .ZN(n8805) );
  NAND2_X1 U10688 ( .A1(n13773), .A2(n13771), .ZN(n8837) );
  NOR2_X1 U10689 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n8811) );
  NOR4_X1 U10690 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8810) );
  NOR4_X1 U10691 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8809) );
  NOR4_X1 U10692 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8808) );
  NAND4_X1 U10693 ( .A1(n8811), .A2(n8810), .A3(n8809), .A4(n8808), .ZN(n8817)
         );
  NOR4_X1 U10694 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8815) );
  NOR4_X1 U10695 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8814) );
  NOR4_X1 U10696 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8813) );
  NOR4_X1 U10697 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n8812) );
  NAND4_X1 U10698 ( .A1(n8815), .A2(n8814), .A3(n8813), .A4(n8812), .ZN(n8816)
         );
  NOR2_X1 U10699 ( .A1(n8817), .A2(n8816), .ZN(n8818) );
  NOR2_X1 U10700 ( .A1(n10860), .A2(n8818), .ZN(n8834) );
  NOR2_X1 U10701 ( .A1(n8837), .A2(n8834), .ZN(n11219) );
  NAND2_X1 U10702 ( .A1(n11900), .A2(n8819), .ZN(n11295) );
  OR2_X1 U10703 ( .A1(n8820), .A2(n11295), .ZN(n11209) );
  NOR2_X1 U10704 ( .A1(n13996), .A2(n12507), .ZN(n8824) );
  NAND2_X1 U10705 ( .A1(n8825), .A2(n8824), .ZN(n11201) );
  NOR2_X1 U10706 ( .A1(n11298), .A2(n10276), .ZN(n11245) );
  INV_X1 U10707 ( .A(n11220), .ZN(n11213) );
  NAND2_X1 U10708 ( .A1(n11245), .A2(n11213), .ZN(n11215) );
  OAI21_X1 U10709 ( .B1(n11209), .B2(n11220), .A(n11215), .ZN(n8826) );
  NAND2_X1 U10710 ( .A1(n11219), .A2(n8826), .ZN(n8829) );
  INV_X1 U10711 ( .A(n13773), .ZN(n8827) );
  NAND2_X1 U10712 ( .A1(n8827), .A2(n11315), .ZN(n8835) );
  NAND3_X1 U10713 ( .A1(n11217), .A2(n11213), .A3(n11208), .ZN(n8828) );
  NAND2_X1 U10714 ( .A1(n8831), .A2(n8227), .ZN(P3_U3455) );
  INV_X1 U10715 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8844) );
  NAND2_X1 U10716 ( .A1(n8832), .A2(n10276), .ZN(n11316) );
  NAND2_X1 U10717 ( .A1(n11298), .A2(n11040), .ZN(n11317) );
  NAND2_X1 U10718 ( .A1(n11316), .A2(n11317), .ZN(n8833) );
  NAND2_X1 U10719 ( .A1(n8833), .A2(n13771), .ZN(n8842) );
  NOR2_X1 U10720 ( .A1(n8834), .A2(n11220), .ZN(n8836) );
  NAND2_X1 U10721 ( .A1(n8838), .A2(n11900), .ZN(n8839) );
  OAI211_X1 U10722 ( .C1(n10330), .C2(n8840), .A(n8839), .B(n11315), .ZN(n8841) );
  INV_X1 U10723 ( .A(n8848), .ZN(n8847) );
  NAND2_X1 U10724 ( .A1(n8847), .A2(n10819), .ZN(n8849) );
  NAND2_X1 U10725 ( .A1(n8848), .A2(SI_1_), .ZN(n8854) );
  NAND2_X1 U10726 ( .A1(n8849), .A2(n8854), .ZN(n8984) );
  INV_X1 U10727 ( .A(n8984), .ZN(n8853) );
  MUX2_X1 U10728 ( .A(n8851), .B(n8975), .S(n8850), .Z(n8852) );
  INV_X1 U10729 ( .A(SI_0_), .ZN(n9713) );
  NAND2_X1 U10730 ( .A1(n8855), .A2(SI_2_), .ZN(n8857) );
  MUX2_X1 U10731 ( .A(n10833), .B(n10805), .S(n8863), .Z(n8993) );
  MUX2_X1 U10732 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8863), .Z(n8858) );
  NAND2_X1 U10733 ( .A1(n8858), .A2(SI_3_), .ZN(n9026) );
  OAI21_X1 U10734 ( .B1(SI_3_), .B2(n8858), .A(n9026), .ZN(n9016) );
  INV_X1 U10735 ( .A(n9016), .ZN(n8859) );
  MUX2_X1 U10736 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8863), .Z(n8861) );
  NAND2_X1 U10737 ( .A1(n8861), .A2(SI_4_), .ZN(n9042) );
  INV_X1 U10738 ( .A(n8861), .ZN(n8862) );
  INV_X1 U10739 ( .A(SI_4_), .ZN(n10840) );
  NAND2_X1 U10740 ( .A1(n8862), .A2(n10840), .ZN(n9027) );
  INV_X1 U10741 ( .A(n9027), .ZN(n8864) );
  NAND2_X1 U10742 ( .A1(n8867), .A2(SI_6_), .ZN(n8869) );
  OAI21_X1 U10743 ( .B1(SI_6_), .B2(n8867), .A(n8869), .ZN(n8868) );
  INV_X1 U10744 ( .A(n8868), .ZN(n9061) );
  MUX2_X1 U10745 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10801), .Z(n8870) );
  NAND2_X1 U10746 ( .A1(n8870), .A2(SI_7_), .ZN(n8872) );
  OAI21_X1 U10747 ( .B1(n8870), .B2(SI_7_), .A(n8872), .ZN(n8871) );
  INV_X1 U10748 ( .A(n8871), .ZN(n9077) );
  MUX2_X1 U10749 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10801), .Z(n8873) );
  NAND2_X1 U10750 ( .A1(n8873), .A2(SI_8_), .ZN(n8875) );
  OAI21_X1 U10751 ( .B1(SI_8_), .B2(n8873), .A(n8875), .ZN(n8874) );
  INV_X1 U10752 ( .A(n8874), .ZN(n9094) );
  NAND2_X1 U10753 ( .A1(n8876), .A2(SI_9_), .ZN(n8877) );
  MUX2_X1 U10754 ( .A(n10923), .B(n10924), .S(n10801), .Z(n8958) );
  MUX2_X1 U10755 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10801), .Z(n8878) );
  NAND2_X1 U10756 ( .A1(n8878), .A2(SI_10_), .ZN(n8880) );
  OAI21_X1 U10757 ( .B1(SI_10_), .B2(n8878), .A(n8880), .ZN(n8879) );
  INV_X1 U10758 ( .A(n8879), .ZN(n9114) );
  MUX2_X1 U10759 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10801), .Z(n8881) );
  XNOR2_X1 U10760 ( .A(n8881), .B(SI_11_), .ZN(n8942) );
  INV_X1 U10761 ( .A(n8881), .ZN(n8882) );
  MUX2_X1 U10762 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n10801), .Z(n8883) );
  XNOR2_X1 U10763 ( .A(n8883), .B(n13914), .ZN(n9132) );
  INV_X1 U10764 ( .A(n8883), .ZN(n8884) );
  NAND2_X1 U10765 ( .A1(n8884), .A2(n13914), .ZN(n8885) );
  MUX2_X1 U10766 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10801), .Z(n8887) );
  OAI21_X1 U10767 ( .B1(SI_13_), .B2(n8887), .A(n8890), .ZN(n9147) );
  MUX2_X1 U10768 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10801), .Z(n8891) );
  MUX2_X1 U10769 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10801), .Z(n8892) );
  XNOR2_X1 U10770 ( .A(n8892), .B(n13821), .ZN(n9176) );
  INV_X1 U10771 ( .A(n8892), .ZN(n8893) );
  MUX2_X1 U10772 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n10801), .Z(n8894) );
  OAI21_X1 U10773 ( .B1(SI_16_), .B2(n8894), .A(n8897), .ZN(n9189) );
  MUX2_X1 U10774 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n10801), .Z(n8898) );
  MUX2_X1 U10775 ( .A(n12151), .B(n12153), .S(n10801), .Z(n8901) );
  NAND2_X1 U10776 ( .A1(n8900), .A2(n8901), .ZN(n8902) );
  NOR2_X1 U10777 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n8906) );
  AND4_X2 U10778 ( .A1(n8906), .A2(n8905), .A3(n8904), .A4(n8903), .ZN(n8908)
         );
  INV_X1 U10779 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8921) );
  INV_X1 U10780 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8909) );
  AND4_X1 U10781 ( .A1(n8921), .A2(n8909), .A3(n7895), .A4(n9409), .ZN(n8912)
         );
  NAND2_X1 U10782 ( .A1(n9415), .A2(n7201), .ZN(n9406) );
  INV_X1 U10783 ( .A(n9406), .ZN(n8911) );
  INV_X1 U10784 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U10785 ( .A1(n12150), .A2(n7478), .ZN(n8925) );
  NAND2_X1 U10786 ( .A1(n7205), .A2(n8909), .ZN(n9224) );
  NAND2_X1 U10787 ( .A1(n9208), .A2(n8921), .ZN(n8922) );
  XNOR2_X1 U10788 ( .A(n8923), .B(P2_IR_REG_18__SCAN_IN), .ZN(n15326) );
  AOI22_X1 U10789 ( .A1(n10534), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n10755), 
        .B2(n15326), .ZN(n8924) );
  NAND2_X1 U10790 ( .A1(n9032), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9069) );
  INV_X1 U10791 ( .A(n9069), .ZN(n8926) );
  NAND2_X1 U10792 ( .A1(n8926), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9086) );
  INV_X1 U10793 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9198) );
  INV_X1 U10794 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8930) );
  NAND2_X1 U10795 ( .A1(n9214), .A2(n8930), .ZN(n8931) );
  NAND2_X1 U10796 ( .A1(n9230), .A2(n8931), .ZN(n14140) );
  XNOR2_X2 U10797 ( .A(n8932), .B(P2_IR_REG_30__SCAN_IN), .ZN(n14568) );
  OR2_X1 U10798 ( .A1(n14140), .A2(n9398), .ZN(n8941) );
  INV_X1 U10799 ( .A(n7168), .ZN(n9473) );
  INV_X1 U10800 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U10801 ( .A1(n9232), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U10802 ( .A1(n10529), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8936) );
  OAI211_X1 U10803 ( .C1(n9473), .C2(n8938), .A(n8937), .B(n8936), .ZN(n8939)
         );
  INV_X1 U10804 ( .A(n8939), .ZN(n8940) );
  NAND2_X1 U10805 ( .A1(n8941), .A2(n8940), .ZN(n14176) );
  XNOR2_X1 U10806 ( .A(n14500), .B(n14176), .ZN(n14420) );
  NAND2_X1 U10807 ( .A1(n8944), .A2(n8945), .ZN(n9028) );
  INV_X1 U10808 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8946) );
  NAND2_X1 U10809 ( .A1(n9135), .A2(n8946), .ZN(n9081) );
  INV_X1 U10810 ( .A(n9099), .ZN(n8948) );
  INV_X1 U10811 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U10812 ( .A1(n8948), .A2(n8947), .ZN(n9118) );
  XNOR2_X1 U10813 ( .A(n8949), .B(P2_IR_REG_11__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U10814 ( .A1(n12026), .A2(n10755), .B1(n9195), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U10815 ( .A1(n9125), .A2(n8952), .ZN(n8953) );
  NAND2_X1 U10816 ( .A1(n9141), .A2(n8953), .ZN(n12284) );
  OR2_X1 U10817 ( .A1(n9398), .A2(n12284), .ZN(n8957) );
  NAND2_X1 U10818 ( .A1(n9232), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8956) );
  NAND2_X1 U10819 ( .A1(n7169), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U10820 ( .A1(n10529), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8954) );
  NAND4_X1 U10821 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n14183) );
  XNOR2_X1 U10822 ( .A(n12279), .B(n12280), .ZN(n11974) );
  INV_X1 U10823 ( .A(n11974), .ZN(n9130) );
  NAND2_X1 U10824 ( .A1(n8959), .A2(n8958), .ZN(n8960) );
  NAND2_X1 U10825 ( .A1(n8961), .A2(n8960), .ZN(n10925) );
  XNOR2_X1 U10826 ( .A(n8962), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U10827 ( .A1(n10755), .A2(n11924), .B1(n9195), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U10828 ( .A1(n9106), .A2(n8965), .ZN(n8966) );
  NAND2_X1 U10829 ( .A1(n9123), .A2(n8966), .ZN(n11991) );
  OR2_X1 U10830 ( .A1(n9398), .A2(n11991), .ZN(n8970) );
  NAND2_X1 U10831 ( .A1(n7169), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U10832 ( .A1(n10529), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8968) );
  NAND2_X1 U10833 ( .A1(n9232), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8967) );
  NAND4_X1 U10834 ( .A1(n8970), .A2(n8969), .A3(n8968), .A4(n8967), .ZN(n14185) );
  XNOR2_X1 U10835 ( .A(n11998), .B(n14185), .ZN(n10597) );
  INV_X1 U10836 ( .A(n10597), .ZN(n11669) );
  NAND2_X1 U10837 ( .A1(n9003), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U10838 ( .A1(n9157), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8972) );
  NAND2_X1 U10839 ( .A1(n9004), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8971) );
  INV_X1 U10840 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n15255) );
  XNOR2_X1 U10841 ( .A(n8976), .B(n8975), .ZN(n14593) );
  NAND2_X1 U10842 ( .A1(n14194), .A2(n7629), .ZN(n11241) );
  NAND2_X1 U10843 ( .A1(n9004), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8980) );
  NAND2_X1 U10844 ( .A1(n9157), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8979) );
  INV_X1 U10845 ( .A(n8982), .ZN(n8983) );
  NAND2_X1 U10846 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  NAND2_X1 U10847 ( .A1(n8986), .A2(n8985), .ZN(n10807) );
  NAND2_X1 U10848 ( .A1(n9000), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8991) );
  INV_X1 U10849 ( .A(n8997), .ZN(n8988) );
  NAND2_X1 U10850 ( .A1(n8989), .A2(n8988), .ZN(n10802) );
  INV_X1 U10851 ( .A(n10802), .ZN(n15257) );
  OR2_X1 U10852 ( .A1(n10348), .A2(n7436), .ZN(n8992) );
  NAND2_X1 U10853 ( .A1(n11283), .A2(n8992), .ZN(n15693) );
  NAND2_X1 U10854 ( .A1(n8994), .A2(n8993), .ZN(n8995) );
  NAND2_X1 U10855 ( .A1(n10804), .A2(n10533), .ZN(n9002) );
  NOR2_X1 U10856 ( .A1(n8997), .A2(n14563), .ZN(n8998) );
  MUX2_X1 U10857 ( .A(n14563), .B(n8998), .S(P2_IR_REG_2__SCAN_IN), .Z(n8999)
         );
  NAND2_X1 U10858 ( .A1(n7237), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U10859 ( .A1(n9003), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U10860 ( .A1(n9157), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U10861 ( .A1(n9004), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9005) );
  NAND2_X1 U10862 ( .A1(n15708), .A2(n14193), .ZN(n9009) );
  INV_X1 U10863 ( .A(n14193), .ZN(n11228) );
  NAND2_X1 U10864 ( .A1(n11383), .A2(n11228), .ZN(n9424) );
  NAND2_X1 U10865 ( .A1(n15708), .A2(n11228), .ZN(n9010) );
  NAND2_X1 U10866 ( .A1(n15692), .A2(n9010), .ZN(n11325) );
  OR2_X1 U10867 ( .A1(n9398), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U10868 ( .A1(n7168), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9012) );
  NAND2_X1 U10869 ( .A1(n9004), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9011) );
  INV_X1 U10870 ( .A(n9015), .ZN(n9017) );
  NAND2_X1 U10871 ( .A1(n9017), .A2(n9016), .ZN(n9019) );
  NAND2_X1 U10872 ( .A1(n10808), .A2(n10533), .ZN(n9024) );
  NOR2_X1 U10873 ( .A1(n8944), .A2(n14563), .ZN(n9020) );
  MUX2_X1 U10874 ( .A(n14563), .B(n9020), .S(P2_IR_REG_3__SCAN_IN), .Z(n9022)
         );
  INV_X1 U10875 ( .A(n9028), .ZN(n9021) );
  AOI22_X1 U10876 ( .A1(n9195), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n10755), 
        .B2(n14210), .ZN(n9023) );
  NAND2_X1 U10877 ( .A1(n11325), .A2(n11324), .ZN(n11327) );
  INV_X1 U10878 ( .A(n11336), .ZN(n11782) );
  NAND2_X1 U10879 ( .A1(n11782), .A2(n11104), .ZN(n9025) );
  NAND2_X1 U10880 ( .A1(n11327), .A2(n9025), .ZN(n11467) );
  NAND2_X1 U10881 ( .A1(n9042), .A2(n9027), .ZN(n9038) );
  XNOR2_X1 U10882 ( .A(n9040), .B(n9038), .ZN(n10823) );
  NAND2_X1 U10883 ( .A1(n10823), .A2(n7478), .ZN(n9031) );
  AND2_X1 U10884 ( .A1(n9029), .A2(n9045), .ZN(n10780) );
  AOI22_X1 U10885 ( .A1(n9195), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10755), 
        .B2(n10780), .ZN(n9030) );
  NAND2_X2 U10886 ( .A1(n9031), .A2(n9030), .ZN(n11473) );
  INV_X1 U10887 ( .A(n9032), .ZN(n9051) );
  OAI21_X1 U10888 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n9051), .ZN(n11474) );
  NAND2_X1 U10889 ( .A1(n9232), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U10890 ( .A1(n7168), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U10891 ( .A1(n9004), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9033) );
  INV_X1 U10892 ( .A(n11479), .ZN(n11466) );
  NAND2_X1 U10893 ( .A1(n11467), .A2(n11466), .ZN(n11469) );
  OR2_X1 U10894 ( .A1(n11473), .A2(n14191), .ZN(n9037) );
  INV_X1 U10895 ( .A(n9038), .ZN(n9039) );
  NAND2_X1 U10896 ( .A1(n9040), .A2(n9039), .ZN(n9043) );
  XNOR2_X1 U10897 ( .A(n9046), .B(P2_IR_REG_5__SCAN_IN), .ZN(n11263) );
  AOI22_X1 U10898 ( .A1(n9195), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10755), 
        .B2(n11263), .ZN(n9047) );
  NAND2_X1 U10899 ( .A1(n9232), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9057) );
  INV_X1 U10900 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U10901 ( .A1(n9051), .A2(n9050), .ZN(n9052) );
  NAND2_X1 U10902 ( .A1(n9069), .A2(n9052), .ZN(n11600) );
  OR2_X1 U10903 ( .A1(n9398), .A2(n11600), .ZN(n9055) );
  INV_X1 U10904 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9053) );
  OR2_X1 U10905 ( .A1(n9088), .A2(n9053), .ZN(n9054) );
  NAND2_X1 U10906 ( .A1(n11405), .A2(n14190), .ZN(n9058) );
  NAND2_X1 U10907 ( .A1(n11025), .A2(n9058), .ZN(n9060) );
  INV_X1 U10908 ( .A(n11405), .ZN(n11602) );
  NAND2_X1 U10909 ( .A1(n11602), .A2(n11429), .ZN(n9059) );
  NAND2_X1 U10910 ( .A1(n9060), .A2(n9059), .ZN(n15802) );
  OR2_X1 U10911 ( .A1(n9062), .A2(n9061), .ZN(n9063) );
  AND2_X1 U10912 ( .A1(n9064), .A2(n9063), .ZN(n10835) );
  NAND2_X1 U10913 ( .A1(n10835), .A2(n7478), .ZN(n9067) );
  OR2_X1 U10914 ( .A1(n9135), .A2(n14563), .ZN(n9065) );
  XNOR2_X1 U10915 ( .A(n9065), .B(P2_IR_REG_6__SCAN_IN), .ZN(n15270) );
  AOI22_X1 U10916 ( .A1(n10534), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10755), 
        .B2(n15270), .ZN(n9066) );
  NAND2_X1 U10917 ( .A1(n9067), .A2(n9066), .ZN(n15801) );
  INV_X1 U10918 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9068) );
  NAND2_X1 U10919 ( .A1(n9069), .A2(n9068), .ZN(n9070) );
  NAND2_X1 U10920 ( .A1(n9086), .A2(n9070), .ZN(n15799) );
  OR2_X1 U10921 ( .A1(n9398), .A2(n15799), .ZN(n9074) );
  NAND2_X1 U10922 ( .A1(n7168), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U10923 ( .A1(n9232), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U10924 ( .A1(n10529), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9071) );
  NAND4_X1 U10925 ( .A1(n9074), .A2(n9073), .A3(n9072), .A4(n9071), .ZN(n14189) );
  XNOR2_X1 U10926 ( .A(n15801), .B(n14189), .ZN(n15795) );
  INV_X1 U10927 ( .A(n15795), .ZN(n15803) );
  NAND2_X1 U10928 ( .A1(n15802), .A2(n15803), .ZN(n9076) );
  INV_X1 U10929 ( .A(n15801), .ZN(n15811) );
  INV_X1 U10930 ( .A(n14189), .ZN(n11803) );
  NAND2_X1 U10931 ( .A1(n15811), .A2(n11803), .ZN(n9075) );
  NAND2_X1 U10932 ( .A1(n9076), .A2(n9075), .ZN(n11632) );
  OR2_X1 U10933 ( .A1(n9078), .A2(n9077), .ZN(n9079) );
  AND2_X1 U10934 ( .A1(n9079), .A2(n9080), .ZN(n10848) );
  NAND2_X1 U10935 ( .A1(n10848), .A2(n7478), .ZN(n9084) );
  XNOR2_X1 U10936 ( .A(n9082), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14226) );
  AOI22_X1 U10937 ( .A1(n10534), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10755), 
        .B2(n14226), .ZN(n9083) );
  NAND2_X1 U10938 ( .A1(n9086), .A2(n9085), .ZN(n9087) );
  NAND2_X1 U10939 ( .A1(n9104), .A2(n9087), .ZN(n11809) );
  OR2_X1 U10940 ( .A1(n9398), .A2(n11809), .ZN(n9092) );
  NAND2_X1 U10941 ( .A1(n9232), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U10942 ( .A1(n7169), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9090) );
  NAND2_X1 U10943 ( .A1(n10529), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9089) );
  NAND4_X1 U10944 ( .A1(n9092), .A2(n9091), .A3(n9090), .A4(n9089), .ZN(n14188) );
  XNOR2_X1 U10945 ( .A(n15831), .B(n11595), .ZN(n11633) );
  OR2_X1 U10946 ( .A1(n15831), .A2(n14188), .ZN(n9093) );
  OR2_X1 U10947 ( .A1(n9095), .A2(n9094), .ZN(n9096) );
  NAND2_X1 U10948 ( .A1(n9097), .A2(n9096), .ZN(n10857) );
  NAND2_X1 U10949 ( .A1(n9100), .A2(n9099), .ZN(n14238) );
  INV_X1 U10950 ( .A(n14238), .ZN(n11267) );
  AOI22_X1 U10951 ( .A1(n10755), .A2(n11267), .B1(n9195), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U10952 ( .A1(n9102), .A2(n9101), .ZN(n11654) );
  NAND2_X1 U10953 ( .A1(n9104), .A2(n9103), .ZN(n9105) );
  NAND2_X1 U10954 ( .A1(n9106), .A2(n9105), .ZN(n11649) );
  OR2_X1 U10955 ( .A1(n9398), .A2(n11649), .ZN(n9110) );
  NAND2_X1 U10956 ( .A1(n9232), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U10957 ( .A1(n7169), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U10958 ( .A1(n10529), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9107) );
  NAND4_X1 U10959 ( .A1(n9110), .A2(n9109), .A3(n9108), .A4(n9107), .ZN(n14187) );
  XNOR2_X1 U10960 ( .A(n11654), .B(n14187), .ZN(n11656) );
  NAND2_X1 U10961 ( .A1(n11654), .A2(n14187), .ZN(n9112) );
  NAND2_X1 U10962 ( .A1(n15848), .A2(n9112), .ZN(n11660) );
  NAND2_X1 U10963 ( .A1(n11669), .A2(n11660), .ZN(n11662) );
  NAND2_X1 U10964 ( .A1(n11998), .A2(n14185), .ZN(n9113) );
  NAND2_X1 U10965 ( .A1(n11662), .A2(n9113), .ZN(n11792) );
  OR2_X1 U10966 ( .A1(n9115), .A2(n9114), .ZN(n9117) );
  XNOR2_X1 U10967 ( .A(n9119), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U10968 ( .A1(n15373), .A2(n10755), .B1(n9195), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n9120) );
  NAND2_X2 U10969 ( .A1(n9121), .A2(n9120), .ZN(n12043) );
  INV_X1 U10970 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9122) );
  NAND2_X1 U10971 ( .A1(n9123), .A2(n9122), .ZN(n9124) );
  NAND2_X1 U10972 ( .A1(n9125), .A2(n9124), .ZN(n12041) );
  OR2_X1 U10973 ( .A1(n9398), .A2(n12041), .ZN(n9129) );
  NAND2_X1 U10974 ( .A1(n9232), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U10975 ( .A1(n7168), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U10976 ( .A1(n10529), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9126) );
  NAND4_X1 U10977 ( .A1(n9129), .A2(n9128), .A3(n9127), .A4(n9126), .ZN(n14184) );
  XNOR2_X1 U10978 ( .A(n12043), .B(n14184), .ZN(n11793) );
  NAND2_X1 U10979 ( .A1(n12279), .A2(n14183), .ZN(n9131) );
  XNOR2_X1 U10980 ( .A(n9133), .B(n9132), .ZN(n11149) );
  NAND2_X1 U10981 ( .A1(n11149), .A2(n7478), .ZN(n9139) );
  NAND2_X1 U10982 ( .A1(n9135), .A2(n9134), .ZN(n9136) );
  AND2_X1 U10983 ( .A1(n9137), .A2(n9151), .ZN(n12615) );
  AOI22_X1 U10984 ( .A1(n10534), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10755), 
        .B2(n12615), .ZN(n9138) );
  INV_X1 U10985 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U10986 ( .A1(n9141), .A2(n9140), .ZN(n9142) );
  NAND2_X1 U10987 ( .A1(n9155), .A2(n9142), .ZN(n15915) );
  OR2_X1 U10988 ( .A1(n9398), .A2(n15915), .ZN(n9146) );
  NAND2_X1 U10989 ( .A1(n7169), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U10990 ( .A1(n10529), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U10991 ( .A1(n9232), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9143) );
  NAND4_X1 U10992 ( .A1(n9146), .A2(n9145), .A3(n9144), .A4(n9143), .ZN(n14182) );
  NAND2_X1 U10993 ( .A1(n9148), .A2(n9147), .ZN(n9149) );
  AND2_X1 U10994 ( .A1(n9150), .A2(n9149), .ZN(n11277) );
  NAND2_X1 U10995 ( .A1(n11277), .A2(n7478), .ZN(n9154) );
  NAND2_X1 U10996 ( .A1(n9152), .A2(n9177), .ZN(n12616) );
  INV_X1 U10997 ( .A(n12616), .ZN(n15358) );
  AOI22_X1 U10998 ( .A1(n10755), .A2(n15358), .B1(n9195), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n9153) );
  NAND2_X1 U10999 ( .A1(n9155), .A2(n12497), .ZN(n9156) );
  AND2_X1 U11000 ( .A1(n9169), .A2(n9156), .ZN(n15937) );
  NAND2_X1 U11001 ( .A1(n15937), .A2(n9157), .ZN(n9161) );
  NAND2_X1 U11002 ( .A1(n9232), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U11003 ( .A1(n7169), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U11004 ( .A1(n10529), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9158) );
  NAND4_X1 U11005 ( .A1(n9161), .A2(n9160), .A3(n9159), .A4(n9158), .ZN(n14181) );
  XNOR2_X1 U11006 ( .A(n12537), .B(n14181), .ZN(n12521) );
  INV_X1 U11007 ( .A(n12521), .ZN(n12527) );
  NAND2_X1 U11008 ( .A1(n12522), .A2(n12527), .ZN(n9163) );
  NAND2_X1 U11009 ( .A1(n12537), .A2(n14181), .ZN(n9162) );
  NAND2_X1 U11010 ( .A1(n9163), .A2(n9162), .ZN(n12381) );
  XNOR2_X1 U11011 ( .A(n9165), .B(n9164), .ZN(n11418) );
  NAND2_X1 U11012 ( .A1(n11418), .A2(n7478), .ZN(n9168) );
  XNOR2_X1 U11013 ( .A(n9166), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U11014 ( .A1(n10755), .A2(n12838), .B1(n9195), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U11015 ( .A1(n9169), .A2(n12651), .ZN(n9170) );
  NAND2_X1 U11016 ( .A1(n9182), .A2(n9170), .ZN(n12650) );
  NAND2_X1 U11017 ( .A1(n9232), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U11018 ( .A1(n7169), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9171) );
  AND2_X1 U11019 ( .A1(n9172), .A2(n9171), .ZN(n9174) );
  NAND2_X1 U11020 ( .A1(n10529), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9173) );
  OAI211_X1 U11021 ( .C1(n12650), .C2(n9398), .A(n9174), .B(n9173), .ZN(n14180) );
  XNOR2_X1 U11022 ( .A(n12655), .B(n14180), .ZN(n12380) );
  XNOR2_X1 U11023 ( .A(n9175), .B(n9176), .ZN(n11548) );
  NAND2_X1 U11024 ( .A1(n11548), .A2(n7478), .ZN(n9180) );
  XNOR2_X1 U11025 ( .A(n9178), .B(P2_IR_REG_15__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U11026 ( .A1(n12839), .A2(n10755), .B1(n9195), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n9179) );
  INV_X1 U11027 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9186) );
  INV_X1 U11028 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9181) );
  NAND2_X1 U11029 ( .A1(n9182), .A2(n9181), .ZN(n9183) );
  NAND2_X1 U11030 ( .A1(n9199), .A2(n9183), .ZN(n12750) );
  OR2_X1 U11031 ( .A1(n12750), .A2(n9398), .ZN(n9185) );
  AOI22_X1 U11032 ( .A1(n9232), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n7168), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n9184) );
  OAI211_X1 U11033 ( .C1(n9088), .C2(n9186), .A(n9185), .B(n9184), .ZN(n14179)
         );
  INV_X1 U11034 ( .A(n12434), .ZN(n12441) );
  NAND2_X1 U11035 ( .A1(n12440), .A2(n12441), .ZN(n12443) );
  OR2_X1 U11036 ( .A1(n15960), .A2(n14179), .ZN(n9187) );
  NAND2_X1 U11037 ( .A1(n12443), .A2(n9187), .ZN(n12588) );
  NAND2_X1 U11038 ( .A1(n9188), .A2(n9189), .ZN(n9190) );
  NAND2_X1 U11039 ( .A1(n9191), .A2(n9190), .ZN(n11572) );
  XNOR2_X1 U11040 ( .A(n9194), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15308) );
  AOI22_X1 U11041 ( .A1(n10534), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10755), 
        .B2(n15308), .ZN(n9196) );
  NAND2_X1 U11042 ( .A1(n9199), .A2(n9198), .ZN(n9200) );
  NAND2_X1 U11043 ( .A1(n9212), .A2(n9200), .ZN(n12857) );
  AOI22_X1 U11044 ( .A1(n9232), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n7169), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U11045 ( .A1(n10529), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9201) );
  OAI211_X1 U11046 ( .C1(n12857), .C2(n9398), .A(n9202), .B(n9201), .ZN(n14178) );
  INV_X1 U11047 ( .A(n14178), .ZN(n9203) );
  INV_X1 U11048 ( .A(n12592), .ZN(n12587) );
  NAND2_X1 U11049 ( .A1(n14512), .A2(n14178), .ZN(n9205) );
  XNOR2_X1 U11050 ( .A(n9206), .B(n9207), .ZN(n11933) );
  NAND2_X1 U11051 ( .A1(n11933), .A2(n7478), .ZN(n9210) );
  XNOR2_X1 U11052 ( .A(n9208), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15323) );
  AOI22_X1 U11053 ( .A1(n10534), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n10755), 
        .B2(n15323), .ZN(n9209) );
  INV_X1 U11054 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U11055 ( .A1(n9212), .A2(n9211), .ZN(n9213) );
  NAND2_X1 U11056 ( .A1(n9214), .A2(n9213), .ZN(n12681) );
  OR2_X1 U11057 ( .A1(n12681), .A2(n9398), .ZN(n9219) );
  INV_X1 U11058 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n15302) );
  NAND2_X1 U11059 ( .A1(n10529), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9216) );
  NAND2_X1 U11060 ( .A1(n7169), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9215) );
  OAI211_X1 U11061 ( .C1(n10532), .C2(n15302), .A(n9216), .B(n9215), .ZN(n9217) );
  INV_X1 U11062 ( .A(n9217), .ZN(n9218) );
  NAND2_X1 U11063 ( .A1(n9219), .A2(n9218), .ZN(n14177) );
  XNOR2_X1 U11064 ( .A(n14557), .B(n14177), .ZN(n12671) );
  INV_X1 U11065 ( .A(n12671), .ZN(n12676) );
  NOR2_X1 U11066 ( .A1(n14557), .A2(n14177), .ZN(n9220) );
  INV_X1 U11067 ( .A(n14176), .ZN(n14008) );
  NAND2_X1 U11068 ( .A1(n7838), .A2(n14008), .ZN(n9221) );
  NAND2_X1 U11069 ( .A1(n14418), .A2(n9221), .ZN(n14399) );
  INV_X1 U11070 ( .A(n14399), .ZN(n9237) );
  MUX2_X1 U11071 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n8863), .Z(n9239) );
  XNOR2_X1 U11072 ( .A(n9241), .B(n9240), .ZN(n12402) );
  NAND2_X1 U11073 ( .A1(n12402), .A2(n7478), .ZN(n9228) );
  NOR2_X2 U11074 ( .A1(n9224), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U11075 ( .A1(n9408), .A2(n9225), .ZN(n9226) );
  XNOR2_X2 U11076 ( .A(n7204), .B(n9415), .ZN(n9420) );
  AOI22_X1 U11077 ( .A1(n10534), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10755), 
        .B2(n15339), .ZN(n9227) );
  INV_X1 U11078 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U11079 ( .A1(n9230), .A2(n9229), .ZN(n9231) );
  NAND2_X1 U11080 ( .A1(n9246), .A2(n9231), .ZN(n14406) );
  INV_X1 U11081 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14407) );
  NAND2_X1 U11082 ( .A1(n9232), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U11083 ( .A1(n10529), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9233) );
  OAI211_X1 U11084 ( .C1(n9473), .C2(n14407), .A(n9234), .B(n9233), .ZN(n9235)
         );
  INV_X1 U11085 ( .A(n9235), .ZN(n9236) );
  OAI21_X1 U11086 ( .B1(n14406), .B2(n9398), .A(n9236), .ZN(n14175) );
  INV_X1 U11087 ( .A(n14175), .ZN(n9447) );
  XNOR2_X1 U11088 ( .A(n14405), .B(n9447), .ZN(n14411) );
  NAND2_X1 U11089 ( .A1(n14405), .A2(n14175), .ZN(n9238) );
  INV_X1 U11090 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12484) );
  MUX2_X1 U11091 ( .A(n12484), .B(n12504), .S(n10801), .Z(n9253) );
  XNOR2_X1 U11092 ( .A(n9253), .B(SI_20_), .ZN(n9242) );
  XNOR2_X1 U11093 ( .A(n9255), .B(n9242), .ZN(n12483) );
  NAND2_X1 U11094 ( .A1(n12483), .A2(n7478), .ZN(n9244) );
  NAND2_X1 U11095 ( .A1(n10534), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9243) );
  INV_X1 U11096 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n14120) );
  NAND2_X1 U11097 ( .A1(n9246), .A2(n14120), .ZN(n9247) );
  AND2_X1 U11098 ( .A1(n9260), .A2(n9247), .ZN(n14393) );
  NAND2_X1 U11099 ( .A1(n14393), .A2(n9157), .ZN(n9252) );
  INV_X1 U11100 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n14490) );
  NAND2_X1 U11101 ( .A1(n10529), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U11102 ( .A1(n7168), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9248) );
  OAI211_X1 U11103 ( .C1(n10532), .C2(n14490), .A(n9249), .B(n9248), .ZN(n9250) );
  INV_X1 U11104 ( .A(n9250), .ZN(n9251) );
  NAND2_X1 U11105 ( .A1(n9252), .A2(n9251), .ZN(n14174) );
  NOR2_X1 U11106 ( .A1(n9256), .A2(SI_20_), .ZN(n9254) );
  MUX2_X1 U11107 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10801), .Z(n9269) );
  XNOR2_X1 U11108 ( .A(n9269), .B(SI_21_), .ZN(n9267) );
  XNOR2_X1 U11109 ( .A(n9268), .B(n9267), .ZN(n12668) );
  NAND2_X1 U11110 ( .A1(n12668), .A2(n7478), .ZN(n9258) );
  NAND2_X1 U11111 ( .A1(n10534), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9257) );
  INV_X1 U11112 ( .A(n9260), .ZN(n9259) );
  INV_X1 U11113 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n14084) );
  NAND2_X1 U11114 ( .A1(n9260), .A2(n14084), .ZN(n9261) );
  NAND2_X1 U11115 ( .A1(n9274), .A2(n9261), .ZN(n14373) );
  OR2_X1 U11116 ( .A1(n14373), .A2(n9398), .ZN(n9266) );
  INV_X1 U11117 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14485) );
  NAND2_X1 U11118 ( .A1(n7169), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9263) );
  NAND2_X1 U11119 ( .A1(n10529), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9262) );
  OAI211_X1 U11120 ( .C1(n10532), .C2(n14485), .A(n9263), .B(n9262), .ZN(n9264) );
  INV_X1 U11121 ( .A(n9264), .ZN(n9265) );
  NAND2_X1 U11122 ( .A1(n9266), .A2(n9265), .ZN(n14173) );
  NAND2_X1 U11123 ( .A1(n9269), .A2(SI_21_), .ZN(n9270) );
  XNOR2_X1 U11124 ( .A(n9286), .B(SI_22_), .ZN(n9580) );
  MUX2_X1 U11125 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n8863), .Z(n9287) );
  XNOR2_X1 U11126 ( .A(n9580), .B(n9287), .ZN(n12791) );
  NAND2_X1 U11127 ( .A1(n12791), .A2(n7478), .ZN(n9273) );
  NAND2_X1 U11128 ( .A1(n10534), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9272) );
  INV_X1 U11129 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U11130 ( .A1(n9274), .A2(n14131), .ZN(n9275) );
  AND2_X1 U11131 ( .A1(n9294), .A2(n9275), .ZN(n14363) );
  NAND2_X1 U11132 ( .A1(n14363), .A2(n9157), .ZN(n9281) );
  INV_X1 U11133 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11134 ( .A1(n10529), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11135 ( .A1(n7168), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9276) );
  OAI211_X1 U11136 ( .C1(n10532), .C2(n9278), .A(n9277), .B(n9276), .ZN(n9279)
         );
  INV_X1 U11137 ( .A(n9279), .ZN(n9280) );
  NAND2_X1 U11138 ( .A1(n9281), .A2(n9280), .ZN(n14172) );
  NAND2_X1 U11139 ( .A1(n14540), .A2(n14172), .ZN(n9282) );
  INV_X1 U11140 ( .A(n9287), .ZN(n9284) );
  INV_X1 U11141 ( .A(SI_22_), .ZN(n9283) );
  NAND2_X1 U11142 ( .A1(n9284), .A2(n9283), .ZN(n9285) );
  NAND2_X1 U11143 ( .A1(n9286), .A2(n9285), .ZN(n9289) );
  NAND2_X1 U11144 ( .A1(n9287), .A2(SI_22_), .ZN(n9288) );
  MUX2_X1 U11145 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10801), .Z(n9306) );
  XNOR2_X1 U11146 ( .A(n9306), .B(SI_23_), .ZN(n9303) );
  XNOR2_X1 U11147 ( .A(n9305), .B(n9303), .ZN(n12758) );
  NAND2_X1 U11148 ( .A1(n12758), .A2(n7478), .ZN(n9291) );
  NAND2_X1 U11149 ( .A1(n10534), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9290) );
  INV_X1 U11150 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11151 ( .A1(n9294), .A2(n9293), .ZN(n9295) );
  NAND2_X1 U11152 ( .A1(n9312), .A2(n9295), .ZN(n14349) );
  OR2_X1 U11153 ( .A1(n14349), .A2(n9398), .ZN(n9301) );
  INV_X1 U11154 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U11155 ( .A1(n7168), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U11156 ( .A1(n10529), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9296) );
  OAI211_X1 U11157 ( .C1(n9298), .C2(n10532), .A(n9297), .B(n9296), .ZN(n9299)
         );
  INV_X1 U11158 ( .A(n9299), .ZN(n9300) );
  NAND2_X1 U11159 ( .A1(n9301), .A2(n9300), .ZN(n14171) );
  OR2_X1 U11160 ( .A1(n14469), .A2(n14171), .ZN(n10605) );
  NAND2_X1 U11161 ( .A1(n14347), .A2(n10605), .ZN(n9302) );
  NAND2_X1 U11162 ( .A1(n14469), .A2(n14171), .ZN(n10604) );
  NAND2_X1 U11163 ( .A1(n9302), .A2(n10604), .ZN(n14330) );
  INV_X1 U11164 ( .A(n9303), .ZN(n9304) );
  NAND2_X1 U11165 ( .A1(n9305), .A2(n9304), .ZN(n9308) );
  NAND2_X1 U11166 ( .A1(n9306), .A2(SI_23_), .ZN(n9307) );
  MUX2_X1 U11167 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10801), .Z(n9324) );
  XNOR2_X1 U11168 ( .A(n9324), .B(SI_24_), .ZN(n9321) );
  NAND2_X1 U11169 ( .A1(n14589), .A2(n7478), .ZN(n9310) );
  NAND2_X1 U11170 ( .A1(n10534), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9309) );
  INV_X1 U11171 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U11172 ( .A1(n9312), .A2(n9311), .ZN(n9313) );
  AND2_X1 U11173 ( .A1(n9332), .A2(n9313), .ZN(n14337) );
  NAND2_X1 U11174 ( .A1(n14337), .A2(n9157), .ZN(n9319) );
  INV_X1 U11175 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9316) );
  NAND2_X1 U11176 ( .A1(n7169), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U11177 ( .A1(n10529), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9314) );
  OAI211_X1 U11178 ( .C1(n9316), .C2(n10532), .A(n9315), .B(n9314), .ZN(n9317)
         );
  INV_X1 U11179 ( .A(n9317), .ZN(n9318) );
  NAND2_X1 U11180 ( .A1(n9319), .A2(n9318), .ZN(n14170) );
  INV_X1 U11181 ( .A(n14170), .ZN(n10517) );
  NAND2_X1 U11182 ( .A1(n14466), .A2(n10517), .ZN(n9455) );
  OR2_X1 U11183 ( .A1(n14466), .A2(n10517), .ZN(n9320) );
  INV_X1 U11184 ( .A(n9321), .ZN(n9322) );
  NAND2_X1 U11185 ( .A1(n9323), .A2(n9322), .ZN(n9326) );
  NAND2_X1 U11186 ( .A1(n9324), .A2(SI_24_), .ZN(n9325) );
  NAND2_X1 U11187 ( .A1(n9326), .A2(n9325), .ZN(n9342) );
  MUX2_X1 U11188 ( .A(n12907), .B(n14588), .S(n10801), .Z(n9327) );
  INV_X1 U11189 ( .A(SI_25_), .ZN(n13994) );
  NAND2_X1 U11190 ( .A1(n9327), .A2(n13994), .ZN(n9343) );
  INV_X1 U11191 ( .A(n9327), .ZN(n9328) );
  NAND2_X1 U11192 ( .A1(n9328), .A2(SI_25_), .ZN(n9329) );
  NAND2_X1 U11193 ( .A1(n9343), .A2(n9329), .ZN(n9341) );
  XNOR2_X1 U11194 ( .A(n9342), .B(n9341), .ZN(n12905) );
  NAND2_X1 U11195 ( .A1(n12905), .A2(n7478), .ZN(n9331) );
  NAND2_X1 U11196 ( .A1(n10534), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9330) );
  INV_X1 U11197 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n14091) );
  NAND2_X1 U11198 ( .A1(n9332), .A2(n14091), .ZN(n9333) );
  NAND2_X1 U11199 ( .A1(n14324), .A2(n9157), .ZN(n9338) );
  INV_X1 U11200 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14462) );
  NAND2_X1 U11201 ( .A1(n10529), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9335) );
  NAND2_X1 U11202 ( .A1(n7169), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9334) );
  OAI211_X1 U11203 ( .C1(n10532), .C2(n14462), .A(n9335), .B(n9334), .ZN(n9336) );
  INV_X1 U11204 ( .A(n9336), .ZN(n9337) );
  NOR2_X1 U11205 ( .A1(n14323), .A2(n14169), .ZN(n9339) );
  NAND2_X1 U11206 ( .A1(n14323), .A2(n14169), .ZN(n9340) );
  MUX2_X1 U11207 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10801), .Z(n9357) );
  XNOR2_X1 U11208 ( .A(n9357), .B(n13812), .ZN(n9356) );
  XNOR2_X1 U11209 ( .A(n9360), .B(n9356), .ZN(n14582) );
  NAND2_X1 U11210 ( .A1(n14582), .A2(n7478), .ZN(n9345) );
  NAND2_X1 U11211 ( .A1(n10534), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9344) );
  INV_X1 U11212 ( .A(n9348), .ZN(n9346) );
  NAND2_X1 U11213 ( .A1(n9346), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9365) );
  INV_X1 U11214 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9347) );
  NAND2_X1 U11215 ( .A1(n9348), .A2(n9347), .ZN(n9349) );
  NAND2_X1 U11216 ( .A1(n9365), .A2(n9349), .ZN(n14154) );
  OR2_X1 U11217 ( .A1(n14154), .A2(n9398), .ZN(n9354) );
  INV_X1 U11218 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14457) );
  NAND2_X1 U11219 ( .A1(n10529), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U11220 ( .A1(n7169), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9350) );
  OAI211_X1 U11221 ( .C1(n10532), .C2(n14457), .A(n9351), .B(n9350), .ZN(n9352) );
  INV_X1 U11222 ( .A(n9352), .ZN(n9353) );
  NOR2_X1 U11223 ( .A1(n14531), .A2(n14000), .ZN(n9355) );
  INV_X1 U11224 ( .A(n9356), .ZN(n9359) );
  NAND2_X1 U11225 ( .A1(n9357), .A2(SI_26_), .ZN(n9358) );
  MUX2_X1 U11226 ( .A(n15225), .B(n14581), .S(n10801), .Z(n9374) );
  INV_X1 U11227 ( .A(n9374), .ZN(n9377) );
  XNOR2_X1 U11228 ( .A(n9377), .B(SI_27_), .ZN(n9361) );
  NAND2_X1 U11229 ( .A1(n14579), .A2(n7478), .ZN(n9363) );
  NAND2_X1 U11230 ( .A1(n10534), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9362) );
  INV_X1 U11231 ( .A(n9365), .ZN(n9364) );
  INV_X1 U11232 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n14046) );
  NAND2_X1 U11233 ( .A1(n9365), .A2(n14046), .ZN(n9366) );
  NAND2_X1 U11234 ( .A1(n14296), .A2(n9157), .ZN(n9372) );
  INV_X1 U11235 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U11236 ( .A1(n10529), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U11237 ( .A1(n7168), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9367) );
  OAI211_X1 U11238 ( .C1(n10532), .C2(n9369), .A(n9368), .B(n9367), .ZN(n9370)
         );
  INV_X1 U11239 ( .A(n9370), .ZN(n9371) );
  XNOR2_X1 U11240 ( .A(n14448), .B(n14167), .ZN(n14289) );
  NAND2_X1 U11241 ( .A1(n14448), .A2(n14167), .ZN(n9373) );
  INV_X1 U11242 ( .A(SI_27_), .ZN(n13888) );
  NAND2_X1 U11243 ( .A1(n9374), .A2(n13888), .ZN(n9375) );
  NAND2_X1 U11244 ( .A1(n9376), .A2(n9375), .ZN(n9379) );
  NAND2_X1 U11245 ( .A1(n9377), .A2(SI_27_), .ZN(n9378) );
  MUX2_X1 U11246 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n8863), .Z(n9393) );
  XNOR2_X1 U11247 ( .A(n9393), .B(SI_28_), .ZN(n9394) );
  NAND2_X1 U11248 ( .A1(n14574), .A2(n7478), .ZN(n9381) );
  NAND2_X1 U11249 ( .A1(n10534), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9380) );
  NAND2_X1 U11250 ( .A1(n9382), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n14260) );
  INV_X1 U11251 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n14076) );
  NAND2_X1 U11252 ( .A1(n9383), .A2(n14076), .ZN(n9384) );
  NAND2_X1 U11253 ( .A1(n14260), .A2(n9384), .ZN(n14279) );
  INV_X1 U11254 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9387) );
  NAND2_X1 U11255 ( .A1(n10529), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U11256 ( .A1(n7168), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9385) );
  OAI211_X1 U11257 ( .C1(n10532), .C2(n9387), .A(n9386), .B(n9385), .ZN(n9388)
         );
  INV_X1 U11258 ( .A(n9388), .ZN(n9389) );
  NAND2_X1 U11259 ( .A1(n9390), .A2(n9389), .ZN(n14166) );
  INV_X1 U11260 ( .A(n14166), .ZN(n9391) );
  NAND2_X1 U11261 ( .A1(n14444), .A2(n9391), .ZN(n9392) );
  MUX2_X1 U11262 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n10801), .Z(n9520) );
  INV_X1 U11263 ( .A(SI_29_), .ZN(n13785) );
  XNOR2_X1 U11264 ( .A(n9520), .B(n13785), .ZN(n9518) );
  XNOR2_X1 U11265 ( .A(n9519), .B(n9518), .ZN(n14571) );
  NAND2_X1 U11266 ( .A1(n14571), .A2(n7478), .ZN(n9397) );
  NAND2_X1 U11267 ( .A1(n10534), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9396) );
  OR2_X1 U11268 ( .A1(n14260), .A2(n9398), .ZN(n9404) );
  INV_X1 U11269 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U11270 ( .A1(n7169), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9400) );
  NAND2_X1 U11271 ( .A1(n10529), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9399) );
  OAI211_X1 U11272 ( .C1(n10532), .C2(n9401), .A(n9400), .B(n9399), .ZN(n9402)
         );
  INV_X1 U11273 ( .A(n9402), .ZN(n9403) );
  NAND2_X1 U11274 ( .A1(n9404), .A2(n9403), .ZN(n14165) );
  XNOR2_X1 U11275 ( .A(n14262), .B(n14165), .ZN(n10609) );
  INV_X1 U11276 ( .A(n10609), .ZN(n9464) );
  XNOR2_X1 U11277 ( .A(n9405), .B(n9464), .ZN(n14266) );
  NOR2_X1 U11278 ( .A1(n9406), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n9407) );
  NOR2_X1 U11279 ( .A1(n9410), .A2(n14563), .ZN(n9411) );
  INV_X1 U11280 ( .A(n10537), .ZN(n11092) );
  NAND2_X1 U11281 ( .A1(n11106), .A2(n11092), .ZN(n10620) );
  NAND3_X1 U11282 ( .A1(n10620), .A2(n9420), .A3(n11096), .ZN(n14423) );
  INV_X1 U11283 ( .A(n14173), .ZN(n14017) );
  OR2_X1 U11284 ( .A1(n14376), .A2(n14017), .ZN(n9451) );
  NAND2_X1 U11285 ( .A1(n14376), .A2(n14017), .ZN(n9422) );
  NAND2_X1 U11286 ( .A1(n9451), .A2(n9422), .ZN(n14370) );
  INV_X1 U11287 ( .A(n14370), .ZN(n14380) );
  INV_X1 U11288 ( .A(n14174), .ZN(n9448) );
  INV_X1 U11289 ( .A(n11324), .ZN(n11330) );
  NOR2_X1 U11290 ( .A1(n14194), .A2(n11292), .ZN(n11286) );
  OR2_X1 U11291 ( .A1(n10348), .A2(n11569), .ZN(n15696) );
  NAND2_X1 U11292 ( .A1(n15697), .A2(n15696), .ZN(n9423) );
  NAND2_X1 U11293 ( .A1(n11330), .A2(n11331), .ZN(n11329) );
  NAND2_X1 U11294 ( .A1(n11336), .A2(n11104), .ZN(n9425) );
  NAND2_X1 U11295 ( .A1(n11329), .A2(n9425), .ZN(n11480) );
  NAND2_X1 U11296 ( .A1(n11480), .A2(n11479), .ZN(n11478) );
  INV_X1 U11297 ( .A(n14191), .ZN(n11341) );
  NAND2_X1 U11298 ( .A1(n11473), .A2(n11341), .ZN(n9426) );
  NAND2_X1 U11299 ( .A1(n11602), .A2(n14190), .ZN(n9427) );
  NAND2_X1 U11300 ( .A1(n11029), .A2(n9427), .ZN(n9429) );
  NAND2_X1 U11301 ( .A1(n11405), .A2(n11429), .ZN(n9428) );
  NAND2_X1 U11302 ( .A1(n9429), .A2(n9428), .ZN(n15794) );
  NAND2_X1 U11303 ( .A1(n15794), .A2(n15795), .ZN(n9431) );
  NAND2_X1 U11304 ( .A1(n15801), .A2(n11803), .ZN(n9430) );
  AND2_X1 U11305 ( .A1(n15831), .A2(n11595), .ZN(n9433) );
  OR2_X1 U11306 ( .A1(n15831), .A2(n11595), .ZN(n9432) );
  INV_X1 U11307 ( .A(n14187), .ZN(n11637) );
  NAND2_X1 U11308 ( .A1(n11654), .A2(n11637), .ZN(n11667) );
  INV_X1 U11309 ( .A(n14185), .ZN(n12044) );
  NAND2_X1 U11310 ( .A1(n11998), .A2(n12044), .ZN(n9434) );
  NAND2_X1 U11311 ( .A1(n11670), .A2(n9434), .ZN(n11789) );
  INV_X1 U11312 ( .A(n12043), .ZN(n9480) );
  NAND2_X1 U11313 ( .A1(n9480), .A2(n14184), .ZN(n9435) );
  INV_X1 U11314 ( .A(n14184), .ZN(n12038) );
  NAND2_X1 U11315 ( .A1(n12279), .A2(n12280), .ZN(n9436) );
  XNOR2_X1 U11316 ( .A(n15918), .B(n14182), .ZN(n12511) );
  INV_X1 U11317 ( .A(n14182), .ZN(n12312) );
  NAND2_X1 U11318 ( .A1(n15918), .A2(n12312), .ZN(n9437) );
  NAND2_X1 U11319 ( .A1(n12528), .A2(n12521), .ZN(n9440) );
  INV_X1 U11320 ( .A(n14181), .ZN(n12491) );
  NAND2_X1 U11321 ( .A1(n12537), .A2(n12491), .ZN(n9439) );
  INV_X1 U11322 ( .A(n14180), .ZN(n12642) );
  AND2_X1 U11323 ( .A1(n12655), .A2(n12642), .ZN(n9441) );
  INV_X1 U11324 ( .A(n14179), .ZN(n9442) );
  NAND2_X1 U11325 ( .A1(n12593), .A2(n12587), .ZN(n9444) );
  NAND2_X1 U11326 ( .A1(n12863), .A2(n14178), .ZN(n9443) );
  INV_X1 U11327 ( .A(n14177), .ZN(n10475) );
  NOR2_X1 U11328 ( .A1(n14557), .A2(n10475), .ZN(n9445) );
  NAND2_X1 U11329 ( .A1(n14405), .A2(n9447), .ZN(n9446) );
  NAND2_X1 U11330 ( .A1(n14392), .A2(n9448), .ZN(n9449) );
  NAND2_X1 U11331 ( .A1(n14378), .A2(n9451), .ZN(n14356) );
  INV_X1 U11332 ( .A(n14172), .ZN(n14022) );
  OR2_X1 U11333 ( .A1(n14540), .A2(n14022), .ZN(n9452) );
  INV_X1 U11334 ( .A(n14171), .ZN(n14056) );
  NAND2_X1 U11335 ( .A1(n14469), .A2(n14056), .ZN(n9453) );
  OR2_X1 U11336 ( .A1(n14469), .A2(n14056), .ZN(n9454) );
  INV_X1 U11337 ( .A(n14169), .ZN(n14147) );
  OR2_X1 U11338 ( .A1(n14323), .A2(n14147), .ZN(n9456) );
  NAND2_X1 U11339 ( .A1(n14317), .A2(n9456), .ZN(n9458) );
  NAND2_X1 U11340 ( .A1(n14323), .A2(n14147), .ZN(n9457) );
  XNOR2_X1 U11341 ( .A(n7634), .B(n14000), .ZN(n14303) );
  INV_X1 U11342 ( .A(n14303), .ZN(n14306) );
  NAND2_X1 U11343 ( .A1(n14302), .A2(n14306), .ZN(n9460) );
  OR2_X1 U11344 ( .A1(n14531), .A2(n14168), .ZN(n9459) );
  INV_X1 U11345 ( .A(n14167), .ZN(n9461) );
  NAND2_X1 U11346 ( .A1(n14448), .A2(n9461), .ZN(n9462) );
  XNOR2_X1 U11347 ( .A(n9465), .B(n9464), .ZN(n9468) );
  NAND2_X1 U11348 ( .A1(n10621), .A2(n15339), .ZN(n9467) );
  NAND2_X1 U11349 ( .A1(n7198), .A2(n11390), .ZN(n9466) );
  NAND2_X1 U11350 ( .A1(n9468), .A2(n15797), .ZN(n9479) );
  INV_X1 U11351 ( .A(n7526), .ZN(n9469) );
  AND2_X2 U11352 ( .A1(n11106), .A2(n9469), .ZN(n14152) );
  NAND2_X1 U11353 ( .A1(n11106), .A2(n7526), .ZN(n11977) );
  INV_X1 U11354 ( .A(P2_B_REG_SCAN_IN), .ZN(n9470) );
  NOR2_X1 U11355 ( .A1(n14580), .A2(n9470), .ZN(n9471) );
  NOR2_X1 U11356 ( .A1(n11977), .A2(n9471), .ZN(n14248) );
  INV_X1 U11357 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9472) );
  OR2_X1 U11358 ( .A1(n10532), .A2(n9472), .ZN(n9477) );
  INV_X1 U11359 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n14255) );
  OR2_X1 U11360 ( .A1(n9473), .A2(n14255), .ZN(n9476) );
  INV_X1 U11361 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9474) );
  OR2_X1 U11362 ( .A1(n9088), .A2(n9474), .ZN(n9475) );
  AND3_X1 U11363 ( .A1(n9477), .A2(n9476), .A3(n9475), .ZN(n10539) );
  INV_X1 U11364 ( .A(n10539), .ZN(n14164) );
  AOI22_X1 U11365 ( .A1(n14166), .A2(n14152), .B1(n14248), .B2(n14164), .ZN(
        n9478) );
  INV_X1 U11366 ( .A(n12537), .ZN(n15941) );
  NAND2_X1 U11367 ( .A1(n11026), .A2(n11602), .ZN(n11027) );
  INV_X1 U11368 ( .A(n11654), .ZN(n15852) );
  NAND2_X1 U11369 ( .A1(n11651), .A2(n15852), .ZN(n11663) );
  NAND2_X1 U11370 ( .A1(n14545), .A2(n14391), .ZN(n14372) );
  OR2_X1 U11371 ( .A1(n14540), .A2(n14372), .ZN(n14361) );
  NOR2_X2 U11372 ( .A1(n14309), .A2(n14448), .ZN(n14295) );
  INV_X1 U11373 ( .A(n14444), .ZN(n14283) );
  OR2_X2 U11374 ( .A1(n10621), .A2(n11390), .ZN(n11088) );
  INV_X2 U11375 ( .A(n8233), .ZN(n14308) );
  NAND2_X1 U11376 ( .A1(n14262), .A2(n14276), .ZN(n9481) );
  NAND3_X1 U11377 ( .A1(n14251), .A2(n14308), .A3(n9481), .ZN(n14264) );
  NAND2_X1 U11378 ( .A1(n9488), .A2(n9487), .ZN(n9483) );
  XNOR2_X1 U11379 ( .A(P2_B_REG_SCAN_IN), .B(n14590), .ZN(n9489) );
  AND2_X1 U11380 ( .A1(n14586), .A2(n9489), .ZN(n9493) );
  INV_X1 U11381 ( .A(n9512), .ZN(n15244) );
  INV_X1 U11382 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15243) );
  AOI22_X1 U11383 ( .A1(n15244), .A2(n15243), .B1(n14584), .B2(n14586), .ZN(
        n11081) );
  INV_X1 U11384 ( .A(n14586), .ZN(n9495) );
  INV_X1 U11385 ( .A(n14590), .ZN(n9494) );
  NAND2_X1 U11386 ( .A1(n9495), .A2(n9494), .ZN(n9496) );
  INV_X1 U11387 ( .A(n15250), .ZN(n15247) );
  OR2_X1 U11388 ( .A1(n11081), .A2(n15247), .ZN(n15241) );
  NOR4_X1 U11389 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9503) );
  NOR4_X1 U11390 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9502) );
  NOR4_X1 U11391 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9501) );
  NOR4_X1 U11392 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9500) );
  NAND4_X1 U11393 ( .A1(n9503), .A2(n9502), .A3(n9501), .A4(n9500), .ZN(n9509)
         );
  NOR2_X1 U11394 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9507) );
  NOR4_X1 U11395 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9506) );
  NOR4_X1 U11396 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9505) );
  NOR4_X1 U11397 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n9504) );
  NAND4_X1 U11398 ( .A1(n9507), .A2(n9506), .A3(n9505), .A4(n9504), .ZN(n9508)
         );
  OAI21_X1 U11399 ( .B1(n9509), .B2(n9508), .A(n15244), .ZN(n11080) );
  NAND2_X1 U11400 ( .A1(n11106), .A2(n10537), .ZN(n11388) );
  NAND2_X1 U11401 ( .A1(n14308), .A2(n15339), .ZN(n11089) );
  NAND3_X1 U11402 ( .A1(n11080), .A2(n11388), .A3(n11089), .ZN(n9510) );
  NAND2_X1 U11403 ( .A1(n14584), .A2(n14590), .ZN(n9511) );
  INV_X1 U11404 ( .A(n15249), .ZN(n9513) );
  NOR2_X2 U11405 ( .A1(n11088), .A2(n11092), .ZN(n15959) );
  NAND2_X1 U11406 ( .A1(n14262), .A2(n14510), .ZN(n9514) );
  NAND2_X1 U11407 ( .A1(n9519), .A2(n9518), .ZN(n9523) );
  INV_X1 U11408 ( .A(n9520), .ZN(n9521) );
  NAND2_X1 U11409 ( .A1(n9521), .A2(n13785), .ZN(n9522) );
  MUX2_X1 U11410 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8863), .Z(n9524) );
  XNOR2_X1 U11411 ( .A(n9524), .B(SI_30_), .ZN(n9887) );
  NAND2_X1 U11412 ( .A1(n9524), .A2(SI_30_), .ZN(n9525) );
  OAI21_X1 U11413 ( .B1(n9889), .B2(n9887), .A(n9525), .ZN(n9528) );
  MUX2_X1 U11414 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10801), .Z(n9526) );
  XNOR2_X1 U11415 ( .A(n9526), .B(SI_31_), .ZN(n9527) );
  XNOR2_X1 U11416 ( .A(n9528), .B(n9527), .ZN(n14561) );
  AND2_X1 U11417 ( .A1(n9530), .A2(n9529), .ZN(n9531) );
  NOR2_X1 U11418 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .ZN(n9534) );
  NAND2_X1 U11419 ( .A1(n9622), .A2(n9534), .ZN(n9535) );
  INV_X1 U11420 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9539) );
  OR2_X1 U11421 ( .A1(n7210), .A2(n9539), .ZN(n9540) );
  INV_X1 U11422 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9548) );
  NAND2_X1 U11423 ( .A1(n9893), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9547) );
  NAND2_X2 U11424 ( .A1(n15215), .A2(n15220), .ZN(n9750) );
  INV_X2 U11425 ( .A(n9750), .ZN(n9894) );
  NAND2_X1 U11426 ( .A1(n9894), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9546) );
  OAI211_X1 U11427 ( .C1(n9898), .C2(n9548), .A(n9547), .B(n9546), .ZN(n14855)
         );
  OR2_X1 U11428 ( .A1(n7210), .A2(n15221), .ZN(n9549) );
  NAND2_X1 U11429 ( .A1(n9894), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9561) );
  INV_X1 U11430 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9551) );
  OR2_X1 U11431 ( .A1(n9898), .A2(n9551), .ZN(n9560) );
  NAND2_X1 U11432 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9751) );
  NOR2_X1 U11433 ( .A1(n9751), .A2(n9737), .ZN(n9738) );
  NAND2_X1 U11434 ( .A1(n9738), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9773) );
  NAND2_X1 U11435 ( .A1(n9675), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9667) );
  NAND2_X1 U11436 ( .A1(n9798), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9789) );
  INV_X1 U11437 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9788) );
  INV_X1 U11438 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9835) );
  INV_X1 U11439 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9614) );
  INV_X1 U11440 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U11441 ( .A1(n9603), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9591) );
  INV_X1 U11442 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14698) );
  INV_X1 U11443 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14616) );
  NAND2_X1 U11444 ( .A1(n9870), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U11445 ( .A1(n9851), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9850) );
  NAND2_X1 U11446 ( .A1(n9575), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9574) );
  NAND2_X1 U11447 ( .A1(n9554), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n12889) );
  INV_X1 U11448 ( .A(n9554), .ZN(n9556) );
  INV_X1 U11449 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U11450 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  NAND2_X1 U11451 ( .A1(n12889), .A2(n9557), .ZN(n14873) );
  OR2_X1 U11452 ( .A1(n9722), .A2(n14873), .ZN(n9559) );
  INV_X1 U11453 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14874) );
  OR2_X1 U11454 ( .A1(n9882), .A2(n14874), .ZN(n9558) );
  NAND2_X1 U11455 ( .A1(n15105), .A2(n14887), .ZN(n9562) );
  INV_X1 U11456 ( .A(n14871), .ZN(n9879) );
  OR2_X1 U11457 ( .A1(n7210), .A2(n15225), .ZN(n9563) );
  NAND2_X1 U11458 ( .A1(n9894), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9570) );
  INV_X1 U11459 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9565) );
  OR2_X1 U11460 ( .A1(n9898), .A2(n9565), .ZN(n9569) );
  XNOR2_X1 U11461 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n9566), .ZN(n14889) );
  OR2_X1 U11462 ( .A1(n9722), .A2(n14889), .ZN(n9568) );
  INV_X1 U11463 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14893) );
  OR2_X1 U11464 ( .A1(n9882), .A2(n14893), .ZN(n9567) );
  AND4_X2 U11465 ( .A1(n9570), .A2(n9569), .A3(n9568), .A4(n9567), .ZN(n14904)
         );
  OR2_X1 U11466 ( .A1(n7210), .A2(n15230), .ZN(n9571) );
  NAND2_X1 U11467 ( .A1(n9894), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9579) );
  INV_X1 U11468 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9573) );
  OR2_X1 U11469 ( .A1(n9898), .A2(n9573), .ZN(n9578) );
  OAI21_X1 U11470 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n9575), .A(n9574), .ZN(
        n14718) );
  OR2_X1 U11471 ( .A1(n9722), .A2(n14718), .ZN(n9577) );
  INV_X1 U11472 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14908) );
  OR2_X1 U11473 ( .A1(n9882), .A2(n14908), .ZN(n9576) );
  XNOR2_X1 U11474 ( .A(n15121), .B(n14888), .ZN(n14900) );
  INV_X1 U11475 ( .A(n14900), .ZN(n9878) );
  OR2_X1 U11476 ( .A1(n9580), .A2(n10801), .ZN(n9581) );
  NAND2_X1 U11477 ( .A1(n9591), .A2(n14698), .ZN(n9582) );
  AND2_X1 U11478 ( .A1(n9869), .A2(n9582), .ZN(n14960) );
  NAND2_X1 U11479 ( .A1(n14960), .A2(n9860), .ZN(n9588) );
  INV_X1 U11480 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9585) );
  NAND2_X1 U11481 ( .A1(n9894), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U11482 ( .A1(n9893), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9583) );
  OAI211_X1 U11483 ( .C1(n9898), .C2(n9585), .A(n9584), .B(n9583), .ZN(n9586)
         );
  INV_X1 U11484 ( .A(n9586), .ZN(n9587) );
  NAND2_X1 U11485 ( .A1(n14959), .A2(n14972), .ZN(n12884) );
  INV_X1 U11486 ( .A(n14972), .ZN(n14732) );
  OR2_X1 U11487 ( .A1(n7210), .A2(n12727), .ZN(n9589) );
  OR2_X1 U11488 ( .A1(n9603), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9592) );
  AND2_X1 U11489 ( .A1(n9592), .A2(n9591), .ZN(n14971) );
  NAND2_X1 U11490 ( .A1(n14971), .A2(n9860), .ZN(n9598) );
  INV_X1 U11491 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U11492 ( .A1(n9894), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9594) );
  NAND2_X1 U11493 ( .A1(n9893), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9593) );
  OAI211_X1 U11494 ( .C1(n9898), .C2(n9595), .A(n9594), .B(n9593), .ZN(n9596)
         );
  INV_X1 U11495 ( .A(n9596), .ZN(n9597) );
  XNOR2_X1 U11496 ( .A(n15154), .B(n14984), .ZN(n10028) );
  INV_X1 U11497 ( .A(n10028), .ZN(n9599) );
  OR2_X1 U11498 ( .A1(n7210), .A2(n12484), .ZN(n9600) );
  NOR2_X1 U11499 ( .A1(n9603), .A2(n8228), .ZN(n14985) );
  NAND2_X1 U11500 ( .A1(n14985), .A2(n9860), .ZN(n9609) );
  INV_X1 U11501 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U11502 ( .A1(n9894), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9605) );
  NAND2_X1 U11503 ( .A1(n9893), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9604) );
  OAI211_X1 U11504 ( .C1(n9898), .C2(n9606), .A(n9605), .B(n9604), .ZN(n9607)
         );
  INV_X1 U11505 ( .A(n9607), .ZN(n9608) );
  XNOR2_X1 U11506 ( .A(n14988), .B(n15000), .ZN(n14990) );
  NAND2_X1 U11507 ( .A1(n9909), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9611) );
  MUX2_X1 U11508 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9611), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9612) );
  OR2_X2 U11509 ( .A1(n9909), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n9901) );
  AOI22_X1 U11510 ( .A1(n9832), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7207), 
        .B2(n14849), .ZN(n9613) );
  NAND2_X1 U11511 ( .A1(n9838), .A2(n9614), .ZN(n9615) );
  NAND2_X1 U11512 ( .A1(n9616), .A2(n9615), .ZN(n15004) );
  INV_X1 U11513 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14833) );
  NAND2_X1 U11514 ( .A1(n9894), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U11515 ( .A1(n9893), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9617) );
  OAI211_X1 U11516 ( .C1(n9898), .C2(n14833), .A(n9618), .B(n9617), .ZN(n9619)
         );
  INV_X1 U11517 ( .A(n9619), .ZN(n9620) );
  OAI21_X1 U11518 ( .B1(n15004), .B2(n9722), .A(n9620), .ZN(n15031) );
  INV_X1 U11519 ( .A(n9692), .ZN(n9730) );
  INV_X1 U11520 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9810) );
  NAND4_X1 U11521 ( .A1(n9621), .A2(n9730), .A3(n9622), .A4(n9810), .ZN(n9623)
         );
  NAND2_X1 U11522 ( .A1(n9623), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9624) );
  MUX2_X1 U11523 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9624), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9626) );
  NAND2_X1 U11524 ( .A1(n9626), .A2(n9625), .ZN(n14827) );
  INV_X1 U11525 ( .A(n14827), .ZN(n15418) );
  AOI22_X1 U11526 ( .A1(n9832), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7207), 
        .B2(n15418), .ZN(n9627) );
  NOR2_X1 U11527 ( .A1(n9816), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9629) );
  OR2_X1 U11528 ( .A1(n9826), .A2(n9629), .ZN(n16015) );
  AOI22_X1 U11529 ( .A1(n9721), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9893), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U11530 ( .A1(n9894), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9630) );
  OAI211_X1 U11531 ( .C1(n16015), .C2(n9722), .A(n9631), .B(n9630), .ZN(n15977) );
  XNOR2_X1 U11532 ( .A(n16008), .B(n15977), .ZN(n15055) );
  NOR2_X1 U11533 ( .A1(n9692), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9744) );
  INV_X1 U11534 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U11535 ( .A1(n9744), .A2(n9632), .ZN(n9809) );
  NAND2_X1 U11536 ( .A1(n9633), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U11537 ( .A1(n9758), .A2(n9634), .ZN(n9635) );
  NAND2_X1 U11538 ( .A1(n9635), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9672) );
  OR2_X1 U11539 ( .A1(n9636), .A2(n9537), .ZN(n9637) );
  NAND2_X1 U11540 ( .A1(n9672), .A2(n9637), .ZN(n9652) );
  OAI21_X1 U11541 ( .B1(n9652), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9795) );
  NAND2_X1 U11542 ( .A1(n9795), .A2(n9638), .ZN(n9639) );
  NAND2_X1 U11543 ( .A1(n9639), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9641) );
  NAND2_X1 U11544 ( .A1(n9641), .A2(n9640), .ZN(n9782) );
  OR2_X1 U11545 ( .A1(n9641), .A2(n9640), .ZN(n9642) );
  NOR2_X1 U11546 ( .A1(n7210), .A2(n11279), .ZN(n9643) );
  AOI21_X1 U11547 ( .B1(n11893), .B2(n7207), .A(n9643), .ZN(n9644) );
  NAND2_X1 U11548 ( .A1(n9894), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9650) );
  OR2_X1 U11549 ( .A1(n9898), .A2(n15931), .ZN(n9649) );
  OR2_X1 U11550 ( .A1(n9798), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9646) );
  NAND2_X1 U11551 ( .A1(n9789), .A2(n9646), .ZN(n14687) );
  OR2_X1 U11552 ( .A1(n9722), .A2(n14687), .ZN(n9648) );
  INV_X1 U11553 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11894) );
  OR2_X1 U11554 ( .A1(n9882), .A2(n11894), .ZN(n9647) );
  XNOR2_X1 U11555 ( .A(n12921), .B(n14649), .ZN(n12624) );
  XNOR2_X1 U11556 ( .A(n9651), .B(n9652), .ZN(n10977) );
  AOI22_X1 U11557 ( .A1(n9832), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10977), 
        .B2(n7207), .ZN(n9653) );
  NAND2_X1 U11558 ( .A1(n9894), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9660) );
  INV_X1 U11559 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11456) );
  OR2_X1 U11560 ( .A1(n9898), .A2(n11456), .ZN(n9659) );
  NAND2_X1 U11561 ( .A1(n9667), .A2(n9655), .ZN(n9656) );
  NAND2_X1 U11562 ( .A1(n9800), .A2(n9656), .ZN(n12567) );
  OR2_X1 U11563 ( .A1(n9722), .A2(n12567), .ZN(n9658) );
  INV_X1 U11564 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11451) );
  OR2_X1 U11565 ( .A1(n9882), .A2(n11451), .ZN(n9657) );
  XNOR2_X1 U11566 ( .A(n15900), .B(n12423), .ZN(n12355) );
  INV_X1 U11567 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U11568 ( .A1(n9672), .A2(n9661), .ZN(n9662) );
  NAND2_X1 U11569 ( .A1(n9662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9663) );
  XNOR2_X1 U11570 ( .A(n9663), .B(P1_IR_REG_10__SCAN_IN), .ZN(n14799) );
  AOI22_X1 U11571 ( .A1(n7207), .A2(n14799), .B1(n9832), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U11572 ( .A1(n9894), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9671) );
  INV_X1 U11573 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10970) );
  OR2_X1 U11574 ( .A1(n9898), .A2(n10970), .ZN(n9670) );
  OR2_X1 U11575 ( .A1(n9675), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U11576 ( .A1(n9667), .A2(n9666), .ZN(n12368) );
  OR2_X1 U11577 ( .A1(n9722), .A2(n12368), .ZN(n9669) );
  INV_X1 U11578 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12091) );
  OR2_X1 U11579 ( .A1(n9882), .A2(n12091), .ZN(n9668) );
  XNOR2_X1 U11580 ( .A(n12364), .B(n12362), .ZN(n12096) );
  OR2_X1 U11581 ( .A1(n10925), .A2(n9757), .ZN(n9674) );
  XNOR2_X1 U11582 ( .A(n9672), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U11583 ( .A1(n9832), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7207), .B2(
        n10922), .ZN(n9673) );
  NAND2_X1 U11584 ( .A1(n9894), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9682) );
  INV_X1 U11585 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10969) );
  OR2_X1 U11586 ( .A1(n9898), .A2(n10969), .ZN(n9681) );
  INV_X1 U11587 ( .A(n9675), .ZN(n9678) );
  NAND2_X1 U11588 ( .A1(n9763), .A2(n9676), .ZN(n9677) );
  NAND2_X1 U11589 ( .A1(n9678), .A2(n9677), .ZN(n12271) );
  OR2_X1 U11590 ( .A1(n9722), .A2(n12271), .ZN(n9680) );
  INV_X1 U11591 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n12012) );
  OR2_X1 U11592 ( .A1(n9882), .A2(n12012), .ZN(n9679) );
  NAND4_X1 U11593 ( .A1(n9682), .A2(n9681), .A3(n9680), .A4(n9679), .ZN(n14737) );
  XNOR2_X1 U11594 ( .A(n12273), .B(n14737), .ZN(n12003) );
  NAND2_X1 U11595 ( .A1(n9734), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9683) );
  XNOR2_X1 U11596 ( .A(n9683), .B(P1_IR_REG_6__SCAN_IN), .ZN(n14772) );
  AOI22_X1 U11597 ( .A1(n9832), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7207), .B2(
        n14772), .ZN(n9684) );
  NAND2_X1 U11598 ( .A1(n9685), .A2(n9684), .ZN(n11694) );
  NAND2_X1 U11599 ( .A1(n9721), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9691) );
  INV_X1 U11600 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11691) );
  OR2_X1 U11601 ( .A1(n9882), .A2(n11691), .ZN(n9690) );
  OR2_X1 U11602 ( .A1(n9738), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U11603 ( .A1(n9773), .A2(n9686), .ZN(n11690) );
  OR2_X1 U11604 ( .A1(n9722), .A2(n11690), .ZN(n9689) );
  INV_X1 U11605 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9687) );
  OR2_X1 U11606 ( .A1(n9750), .A2(n9687), .ZN(n9688) );
  XNOR2_X1 U11607 ( .A(n11694), .B(n11709), .ZN(n11685) );
  NAND2_X1 U11608 ( .A1(n9692), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9693) );
  XNOR2_X1 U11609 ( .A(n9693), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14760) );
  AOI22_X1 U11610 ( .A1(n9832), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n7207), .B2(
        n14760), .ZN(n9694) );
  NAND2_X1 U11611 ( .A1(n9695), .A2(n9694), .ZN(n14624) );
  NAND2_X1 U11612 ( .A1(n9721), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9700) );
  OR2_X1 U11613 ( .A1(n9722), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9699) );
  INV_X1 U11614 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10884) );
  OR2_X1 U11615 ( .A1(n9723), .A2(n10884), .ZN(n9698) );
  INV_X1 U11616 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9696) );
  OR2_X1 U11617 ( .A1(n9750), .A2(n9696), .ZN(n9697) );
  XNOR2_X1 U11618 ( .A(n14624), .B(n14742), .ZN(n11554) );
  OR2_X1 U11619 ( .A1(n9898), .A2(n15676), .ZN(n9705) );
  INV_X1 U11620 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10880) );
  OR2_X1 U11621 ( .A1(n9723), .A2(n10880), .ZN(n9704) );
  INV_X1 U11622 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11616) );
  OR2_X1 U11623 ( .A1(n9722), .A2(n11616), .ZN(n9703) );
  INV_X1 U11624 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9701) );
  NAND4_X2 U11625 ( .A1(n9705), .A2(n9704), .A3(n9703), .A4(n9702), .ZN(n10660) );
  NAND2_X1 U11626 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9706) );
  MUX2_X1 U11627 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9706), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9708) );
  NAND2_X1 U11628 ( .A1(n9708), .A2(n9707), .ZN(n10879) );
  OR2_X1 U11629 ( .A1(n9715), .A2(n10879), .ZN(n9709) );
  NAND2_X1 U11630 ( .A1(n10660), .A2(n15670), .ZN(n9712) );
  AND2_X2 U11631 ( .A1(n9712), .A2(n11488), .ZN(n11502) );
  NOR2_X1 U11632 ( .A1(n10801), .A2(n9713), .ZN(n9714) );
  XNOR2_X1 U11633 ( .A(n9714), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15238) );
  MUX2_X1 U11634 ( .A(n7345), .B(n15238), .S(n9715), .Z(n11617) );
  NAND2_X1 U11635 ( .A1(n9860), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9720) );
  INV_X1 U11636 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10652) );
  OR2_X1 U11637 ( .A1(n9898), .A2(n10652), .ZN(n9719) );
  INV_X1 U11638 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9716) );
  OR2_X1 U11639 ( .A1(n9750), .A2(n9716), .ZN(n9717) );
  NAND4_X2 U11640 ( .A1(n9720), .A2(n9719), .A3(n9718), .A4(n9717), .ZN(n14746) );
  NOR2_X1 U11641 ( .A1(n14746), .A2(n11617), .ZN(n11612) );
  AOI21_X1 U11642 ( .B1(n11617), .B2(n14746), .A(n11612), .ZN(n10945) );
  NAND2_X1 U11643 ( .A1(n9721), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9728) );
  INV_X1 U11644 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11847) );
  OR2_X1 U11645 ( .A1(n9722), .A2(n11847), .ZN(n9727) );
  INV_X1 U11646 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10882) );
  OR2_X1 U11647 ( .A1(n9723), .A2(n10882), .ZN(n9726) );
  INV_X1 U11648 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9724) );
  OR2_X1 U11649 ( .A1(n9750), .A2(n9724), .ZN(n9725) );
  MUX2_X1 U11650 ( .A(n9537), .B(n9729), .S(P1_IR_REG_2__SCAN_IN), .Z(n9731)
         );
  NAND4_X1 U11651 ( .A1(n11554), .A2(n11502), .A3(n10945), .A4(n11837), .ZN(
        n9756) );
  NAND2_X1 U11652 ( .A1(n9809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9733) );
  MUX2_X1 U11653 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9733), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9735) );
  AND2_X1 U11654 ( .A1(n9735), .A2(n9734), .ZN(n10914) );
  AOI22_X1 U11655 ( .A1(n9832), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7207), .B2(
        n10914), .ZN(n9736) );
  NAND2_X1 U11656 ( .A1(n9894), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9743) );
  INV_X1 U11657 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10866) );
  OR2_X1 U11658 ( .A1(n9898), .A2(n10866), .ZN(n9742) );
  AND2_X1 U11659 ( .A1(n9751), .A2(n9737), .ZN(n9739) );
  OR2_X1 U11660 ( .A1(n9739), .A2(n9738), .ZN(n11544) );
  OR2_X1 U11661 ( .A1(n9722), .A2(n11544), .ZN(n9741) );
  INV_X1 U11662 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10887) );
  OR2_X1 U11663 ( .A1(n9882), .A2(n10887), .ZN(n9740) );
  XNOR2_X1 U11664 ( .A(n11543), .B(n11686), .ZN(n11534) );
  OR2_X1 U11665 ( .A1(n9744), .A2(n9537), .ZN(n9745) );
  MUX2_X1 U11666 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9745), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9746) );
  AND2_X1 U11667 ( .A1(n9746), .A2(n9809), .ZN(n10885) );
  AOI22_X1 U11668 ( .A1(n9832), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n7207), .B2(
        n10885), .ZN(n9747) );
  NAND2_X1 U11669 ( .A1(n9748), .A2(n9747), .ZN(n11531) );
  NAND2_X1 U11670 ( .A1(n9721), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9755) );
  INV_X1 U11671 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9749) );
  OR2_X1 U11672 ( .A1(n9750), .A2(n9749), .ZN(n9754) );
  OAI21_X1 U11673 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9751), .ZN(n11515) );
  OR2_X1 U11674 ( .A1(n9722), .A2(n11515), .ZN(n9753) );
  INV_X1 U11675 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11517) );
  OR2_X1 U11676 ( .A1(n9882), .A2(n11517), .ZN(n9752) );
  NAND4_X1 U11677 ( .A1(n9755), .A2(n9754), .A3(n9753), .A4(n9752), .ZN(n14741) );
  OR2_X1 U11678 ( .A1(n11531), .A2(n14741), .ZN(n11525) );
  NAND2_X1 U11679 ( .A1(n11531), .A2(n14741), .ZN(n11526) );
  AND2_X1 U11680 ( .A1(n11525), .A2(n11526), .ZN(n11507) );
  NOR4_X1 U11681 ( .A1(n11685), .A2(n9756), .A3(n11534), .A4(n11507), .ZN(
        n9780) );
  OR2_X1 U11682 ( .A1(n10857), .A2(n9757), .ZN(n9760) );
  XNOR2_X1 U11683 ( .A(n9758), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U11684 ( .A1(n9832), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7207), .B2(
        n10890), .ZN(n9759) );
  NAND2_X1 U11685 ( .A1(n9760), .A2(n9759), .ZN(n12198) );
  NAND2_X1 U11686 ( .A1(n9894), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9767) );
  INV_X1 U11687 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10898) );
  OR2_X1 U11688 ( .A1(n9898), .A2(n10898), .ZN(n9766) );
  NAND2_X1 U11689 ( .A1(n9775), .A2(n9761), .ZN(n9762) );
  NAND2_X1 U11690 ( .A1(n9763), .A2(n9762), .ZN(n12206) );
  OR2_X1 U11691 ( .A1(n9722), .A2(n12206), .ZN(n9765) );
  INV_X1 U11692 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11869) );
  OR2_X1 U11693 ( .A1(n9882), .A2(n11869), .ZN(n9764) );
  NAND4_X1 U11694 ( .A1(n9767), .A2(n9766), .A3(n9765), .A4(n9764), .ZN(n14738) );
  XNOR2_X1 U11695 ( .A(n12198), .B(n14738), .ZN(n11854) );
  NAND2_X1 U11696 ( .A1(n9768), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9769) );
  XNOR2_X1 U11697 ( .A(n9769), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14784) );
  AOI22_X1 U11698 ( .A1(n9832), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7207), .B2(
        n14784), .ZN(n9770) );
  NAND2_X1 U11699 ( .A1(n9771), .A2(n9770), .ZN(n11858) );
  NAND2_X1 U11700 ( .A1(n9894), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9779) );
  INV_X1 U11701 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10868) );
  OR2_X1 U11702 ( .A1(n9898), .A2(n10868), .ZN(n9778) );
  NAND2_X1 U11703 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  NAND2_X1 U11704 ( .A1(n9775), .A2(n9774), .ZN(n11713) );
  OR2_X1 U11705 ( .A1(n9722), .A2(n11713), .ZN(n9777) );
  INV_X1 U11706 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11714) );
  OR2_X1 U11707 ( .A1(n9882), .A2(n11714), .ZN(n9776) );
  NAND4_X1 U11708 ( .A1(n9779), .A2(n9778), .A3(n9777), .A4(n9776), .ZN(n14739) );
  XNOR2_X1 U11709 ( .A(n11858), .B(n14739), .ZN(n11708) );
  NAND4_X1 U11710 ( .A1(n12003), .A2(n9780), .A3(n11854), .A4(n11708), .ZN(
        n9781) );
  NOR4_X1 U11711 ( .A1(n12624), .A2(n12355), .A3(n12096), .A4(n9781), .ZN(
        n9807) );
  NAND2_X1 U11712 ( .A1(n9782), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9783) );
  NOR2_X1 U11713 ( .A1(n7210), .A2(n11419), .ZN(n9784) );
  AOI21_X1 U11714 ( .B1(n14823), .B2(n7207), .A(n9784), .ZN(n9785) );
  NAND2_X1 U11715 ( .A1(n9894), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9794) );
  INV_X1 U11716 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9787) );
  OR2_X1 U11717 ( .A1(n9898), .A2(n9787), .ZN(n9793) );
  NAND2_X1 U11718 ( .A1(n9789), .A2(n9788), .ZN(n9790) );
  NAND2_X1 U11719 ( .A1(n9815), .A2(n9790), .ZN(n14609) );
  OR2_X1 U11720 ( .A1(n9722), .A2(n14609), .ZN(n9792) );
  INV_X1 U11721 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14836) );
  OR2_X1 U11722 ( .A1(n9882), .A2(n14836), .ZN(n9791) );
  NAND4_X1 U11723 ( .A1(n9794), .A2(n9793), .A3(n9792), .A4(n9791), .ZN(n15979) );
  XNOR2_X1 U11724 ( .A(n15950), .B(n15979), .ZN(n12631) );
  XNOR2_X1 U11725 ( .A(n9795), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U11726 ( .A1(n11463), .A2(n7207), .B1(n9832), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9796) );
  NAND2_X1 U11727 ( .A1(n9894), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9806) );
  INV_X1 U11728 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11885) );
  OR2_X1 U11729 ( .A1(n9898), .A2(n11885), .ZN(n9805) );
  INV_X1 U11730 ( .A(n9798), .ZN(n9802) );
  NAND2_X1 U11731 ( .A1(n9800), .A2(n9799), .ZN(n9801) );
  NAND2_X1 U11732 ( .A1(n9802), .A2(n9801), .ZN(n14647) );
  OR2_X1 U11733 ( .A1(n9722), .A2(n14647), .ZN(n9804) );
  INV_X1 U11734 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11892) );
  OR2_X1 U11735 ( .A1(n9882), .A2(n11892), .ZN(n9803) );
  NAND4_X1 U11736 ( .A1(n9806), .A2(n9805), .A3(n9804), .A4(n9803), .ZN(n14735) );
  XNOR2_X1 U11737 ( .A(n12915), .B(n14735), .ZN(n12419) );
  NAND4_X1 U11738 ( .A1(n15055), .A2(n9807), .A3(n12631), .A4(n12419), .ZN(
        n9822) );
  INV_X1 U11739 ( .A(n9621), .ZN(n9808) );
  OAI21_X1 U11740 ( .B1(n9809), .B2(n9808), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9811) );
  XNOR2_X1 U11741 ( .A(n9811), .B(n9810), .ZN(n14824) );
  AOI22_X1 U11742 ( .A1(n9832), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7207), 
        .B2(n15424), .ZN(n9812) );
  AND2_X1 U11743 ( .A1(n9815), .A2(n9814), .ZN(n9817) );
  OR2_X1 U11744 ( .A1(n9817), .A2(n9816), .ZN(n15987) );
  NAND2_X1 U11745 ( .A1(n9894), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U11746 ( .A1(n9721), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9818) );
  AND2_X1 U11747 ( .A1(n9819), .A2(n9818), .ZN(n9821) );
  NAND2_X1 U11748 ( .A1(n9893), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9820) );
  OAI211_X1 U11749 ( .C1(n15987), .C2(n9722), .A(n9821), .B(n9820), .ZN(n15058) );
  INV_X1 U11750 ( .A(n15058), .ZN(n14606) );
  XNOR2_X1 U11751 ( .A(n15077), .B(n14606), .ZN(n15081) );
  NOR2_X1 U11752 ( .A1(n9822), .A2(n15081), .ZN(n9845) );
  NAND2_X1 U11753 ( .A1(n9625), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9823) );
  XNOR2_X1 U11754 ( .A(n9823), .B(P1_IR_REG_17__SCAN_IN), .ZN(n15394) );
  AOI22_X1 U11755 ( .A1(n9832), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7207), 
        .B2(n15394), .ZN(n9824) );
  OR2_X1 U11756 ( .A1(n9826), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9827) );
  NAND2_X1 U11757 ( .A1(n9836), .A2(n9827), .ZN(n16030) );
  AOI22_X1 U11758 ( .A1(n9893), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9894), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n9829) );
  NAND2_X1 U11759 ( .A1(n9721), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9828) );
  OAI211_X1 U11760 ( .C1(n16030), .C2(n9722), .A(n9829), .B(n9828), .ZN(n15057) );
  XNOR2_X1 U11761 ( .A(n16026), .B(n15057), .ZN(n15039) );
  NAND2_X1 U11762 ( .A1(n9907), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9830) );
  MUX2_X1 U11763 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9830), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n9831) );
  NAND2_X1 U11764 ( .A1(n9831), .A2(n9909), .ZN(n14840) );
  INV_X1 U11765 ( .A(n14840), .ZN(n15404) );
  AOI22_X1 U11766 ( .A1(n9832), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7207), 
        .B2(n15404), .ZN(n9833) );
  NAND2_X1 U11767 ( .A1(n9836), .A2(n9835), .ZN(n9837) );
  NAND2_X1 U11768 ( .A1(n9838), .A2(n9837), .ZN(n15019) );
  OR2_X1 U11769 ( .A1(n15019), .A2(n9722), .ZN(n9843) );
  INV_X1 U11770 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15020) );
  NAND2_X1 U11771 ( .A1(n9894), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U11772 ( .A1(n9721), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9839) );
  OAI211_X1 U11773 ( .C1(n15020), .C2(n9882), .A(n9840), .B(n9839), .ZN(n9841)
         );
  INV_X1 U11774 ( .A(n9841), .ZN(n9842) );
  NAND2_X1 U11775 ( .A1(n15018), .A2(n16018), .ZN(n12868) );
  NAND2_X1 U11776 ( .A1(n15175), .A2(n15001), .ZN(n9844) );
  NAND2_X1 U11777 ( .A1(n12868), .A2(n9844), .ZN(n15026) );
  NAND4_X1 U11778 ( .A1(n7937), .A2(n9845), .A3(n15039), .A4(n15026), .ZN(
        n9846) );
  NOR4_X1 U11779 ( .A1(n14965), .A2(n9599), .A3(n14990), .A4(n9846), .ZN(n9877) );
  OR2_X1 U11780 ( .A1(n7210), .A2(n12907), .ZN(n9847) );
  NAND2_X1 U11781 ( .A1(n9894), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9855) );
  INV_X1 U11782 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9849) );
  OR2_X1 U11783 ( .A1(n9898), .A2(n9849), .ZN(n9854) );
  OAI21_X1 U11784 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n9851), .A(n9850), .ZN(
        n14916) );
  OR2_X1 U11785 ( .A1(n9722), .A2(n14916), .ZN(n9853) );
  INV_X1 U11786 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14917) );
  OR2_X1 U11787 ( .A1(n9882), .A2(n14917), .ZN(n9852) );
  NAND4_X1 U11788 ( .A1(n9855), .A2(n9854), .A3(n9853), .A4(n9852), .ZN(n14730) );
  XNOR2_X1 U11789 ( .A(n14919), .B(n14730), .ZN(n14914) );
  OR2_X1 U11790 ( .A1(n7210), .A2(n15234), .ZN(n9856) );
  OR2_X1 U11791 ( .A1(n9870), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9859) );
  AND2_X1 U11792 ( .A1(n9859), .A2(n9858), .ZN(n14933) );
  NAND2_X1 U11793 ( .A1(n14933), .A2(n9860), .ZN(n9866) );
  INV_X1 U11794 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U11795 ( .A1(n9894), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9862) );
  NAND2_X1 U11796 ( .A1(n9893), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9861) );
  OAI211_X1 U11797 ( .C1(n9898), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9864)
         );
  INV_X1 U11798 ( .A(n9864), .ZN(n9865) );
  XNOR2_X1 U11799 ( .A(n15135), .B(n14731), .ZN(n12871) );
  INV_X1 U11800 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12761) );
  OR2_X1 U11801 ( .A1(n7210), .A2(n12761), .ZN(n9867) );
  AND2_X1 U11802 ( .A1(n9869), .A2(n14616), .ZN(n9871) );
  OR2_X1 U11803 ( .A1(n9871), .A2(n9870), .ZN(n14945) );
  INV_X1 U11804 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U11805 ( .A1(n9893), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U11806 ( .A1(n9894), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9872) );
  OAI211_X1 U11807 ( .C1(n9898), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9875)
         );
  INV_X1 U11808 ( .A(n9875), .ZN(n9876) );
  XNOR2_X1 U11809 ( .A(n15141), .B(n14958), .ZN(n14942) );
  INV_X1 U11810 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15218) );
  OR2_X1 U11811 ( .A1(n7210), .A2(n15218), .ZN(n9880) );
  NAND2_X1 U11812 ( .A1(n9894), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9886) );
  NAND2_X1 U11813 ( .A1(n9721), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9885) );
  OR2_X1 U11814 ( .A1(n9722), .A2(n12889), .ZN(n9884) );
  INV_X1 U11815 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n12893) );
  OR2_X1 U11816 ( .A1(n9882), .A2(n12893), .ZN(n9883) );
  NAND4_X1 U11817 ( .A1(n9886), .A2(n9885), .A3(n9884), .A4(n9883), .ZN(n14726) );
  XNOR2_X1 U11818 ( .A(n9939), .B(n14726), .ZN(n12887) );
  INV_X1 U11819 ( .A(n9887), .ZN(n9888) );
  INV_X1 U11820 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15217) );
  OR2_X1 U11821 ( .A1(n7210), .A2(n15217), .ZN(n9891) );
  NAND2_X1 U11822 ( .A1(n9892), .A2(n9891), .ZN(n9923) );
  INV_X1 U11823 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U11824 ( .A1(n9893), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U11825 ( .A1(n9894), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9895) );
  OAI211_X1 U11826 ( .C1(n9898), .C2(n9897), .A(n9896), .B(n9895), .ZN(n14725)
         );
  XNOR2_X1 U11827 ( .A(n9923), .B(n14725), .ZN(n9899) );
  NAND2_X1 U11828 ( .A1(n10067), .A2(n8221), .ZN(n9900) );
  NAND2_X1 U11829 ( .A1(n9901), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U11830 ( .A1(n12729), .A2(n10719), .ZN(n10058) );
  NAND3_X1 U11831 ( .A1(n9905), .A2(n9911), .A3(n9904), .ZN(n9906) );
  OAI21_X1 U11832 ( .B1(n9907), .B2(n9906), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9908) );
  NAND2_X1 U11833 ( .A1(n9911), .A2(n9910), .ZN(n9914) );
  INV_X1 U11834 ( .A(n9912), .ZN(n9913) );
  NOR2_X1 U11835 ( .A1(n14855), .A2(n9949), .ZN(n9931) );
  NAND2_X2 U11836 ( .A1(n7968), .A2(n12485), .ZN(n10940) );
  OR2_X1 U11837 ( .A1(n10940), .A2(n12404), .ZN(n11530) );
  NAND2_X1 U11838 ( .A1(n9945), .A2(n15236), .ZN(n10725) );
  NAND2_X1 U11839 ( .A1(n12485), .A2(n10939), .ZN(n9916) );
  NAND2_X1 U11840 ( .A1(n10725), .A2(n9916), .ZN(n9917) );
  NAND2_X1 U11841 ( .A1(n11530), .A2(n9917), .ZN(n10065) );
  XOR2_X1 U11842 ( .A(n9931), .B(n10065), .Z(n9920) );
  NAND2_X1 U11843 ( .A1(n14855), .A2(n10053), .ZN(n9930) );
  XOR2_X1 U11844 ( .A(n10065), .B(n9930), .Z(n9918) );
  NAND2_X1 U11845 ( .A1(n15091), .A2(n9918), .ZN(n9919) );
  OAI211_X1 U11846 ( .C1(n15091), .C2(n9920), .A(n9919), .B(n10058), .ZN(n9921) );
  NAND2_X1 U11847 ( .A1(n9945), .A2(n10719), .ZN(n10943) );
  OAI21_X1 U11848 ( .B1(n14855), .B2(n10943), .A(n14725), .ZN(n9924) );
  INV_X1 U11849 ( .A(n9923), .ZN(n15094) );
  MUX2_X1 U11850 ( .A(n9924), .B(n15094), .S(n10053), .Z(n10081) );
  NAND2_X1 U11851 ( .A1(n9926), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9925) );
  MUX2_X1 U11852 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9925), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9928) );
  NAND2_X1 U11853 ( .A1(n9928), .A2(n10090), .ZN(n10873) );
  INV_X1 U11854 ( .A(n10873), .ZN(n9929) );
  NAND2_X1 U11855 ( .A1(n9929), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12759) );
  INV_X1 U11856 ( .A(n12759), .ZN(n10083) );
  NAND2_X1 U11857 ( .A1(n10081), .A2(n10083), .ZN(n9938) );
  INV_X1 U11858 ( .A(n9930), .ZN(n9934) );
  INV_X1 U11859 ( .A(n9931), .ZN(n9932) );
  NOR2_X1 U11860 ( .A1(n15091), .A2(n9932), .ZN(n9933) );
  AOI211_X1 U11861 ( .C1(n15091), .C2(n9934), .A(n10065), .B(n9933), .ZN(
        n10080) );
  INV_X1 U11862 ( .A(n10080), .ZN(n9937) );
  OAI21_X1 U11863 ( .B1(n14855), .B2(n12729), .A(n14725), .ZN(n9935) );
  MUX2_X1 U11864 ( .A(n9935), .B(n15094), .S(n10054), .Z(n10084) );
  NOR2_X1 U11865 ( .A1(n10084), .A2(n12759), .ZN(n10079) );
  INV_X1 U11866 ( .A(n10079), .ZN(n9936) );
  OAI22_X1 U11867 ( .A1(n10066), .A2(n9938), .B1(n9937), .B2(n9936), .ZN(
        n10072) );
  INV_X1 U11868 ( .A(n14726), .ZN(n13030) );
  MUX2_X1 U11869 ( .A(n13030), .B(n15099), .S(n10053), .Z(n10063) );
  MUX2_X1 U11870 ( .A(n14726), .B(n9939), .S(n10054), .Z(n10062) );
  NOR2_X1 U11871 ( .A1(n10063), .A2(n10062), .ZN(n10102) );
  MUX2_X1 U11872 ( .A(n14887), .B(n14868), .S(n10053), .Z(n9941) );
  INV_X1 U11873 ( .A(n14887), .ZN(n14727) );
  MUX2_X1 U11874 ( .A(n14727), .B(n15105), .S(n10054), .Z(n9940) );
  NAND2_X1 U11875 ( .A1(n9941), .A2(n9940), .ZN(n10105) );
  INV_X1 U11876 ( .A(n9940), .ZN(n9943) );
  INV_X1 U11877 ( .A(n9941), .ZN(n9942) );
  NAND2_X1 U11878 ( .A1(n9943), .A2(n9942), .ZN(n10077) );
  INV_X1 U11879 ( .A(n15000), .ZN(n14733) );
  MUX2_X1 U11880 ( .A(n14733), .B(n14988), .S(n10054), .Z(n10029) );
  INV_X1 U11881 ( .A(n11617), .ZN(n11499) );
  MUX2_X1 U11882 ( .A(n10943), .B(n9945), .S(n9944), .Z(n9947) );
  OAI21_X1 U11883 ( .B1(n11499), .B2(n10940), .A(n9947), .ZN(n9946) );
  AND2_X1 U11884 ( .A1(n14746), .A2(n9946), .ZN(n9953) );
  NAND2_X1 U11885 ( .A1(n11499), .A2(n9949), .ZN(n9948) );
  OAI22_X1 U11886 ( .A1(n14746), .A2(n9948), .B1(n11499), .B2(n9947), .ZN(
        n9952) );
  NAND2_X1 U11887 ( .A1(n14744), .A2(n9710), .ZN(n9950) );
  NAND2_X1 U11888 ( .A1(n9954), .A2(n9950), .ZN(n9951) );
  NOR2_X1 U11889 ( .A1(n10660), .A2(n9710), .ZN(n11500) );
  OAI21_X1 U11890 ( .B1(n9954), .B2(n11500), .A(n11837), .ZN(n9957) );
  MUX2_X1 U11891 ( .A(n14743), .B(n7476), .S(n10054), .Z(n9955) );
  OAI21_X1 U11892 ( .B1(n15686), .B2(n7516), .A(n9955), .ZN(n9956) );
  MUX2_X1 U11893 ( .A(n14742), .B(n14624), .S(n9949), .Z(n9959) );
  INV_X1 U11894 ( .A(n9959), .ZN(n9961) );
  MUX2_X1 U11895 ( .A(n14624), .B(n14742), .S(n9949), .Z(n9960) );
  NAND2_X1 U11896 ( .A1(n9962), .A2(n9961), .ZN(n9963) );
  MUX2_X1 U11897 ( .A(n14741), .B(n11531), .S(n10054), .Z(n9966) );
  MUX2_X1 U11898 ( .A(n14741), .B(n11531), .S(n9949), .Z(n9965) );
  INV_X1 U11899 ( .A(n9970), .ZN(n9968) );
  INV_X1 U11900 ( .A(n11686), .ZN(n14740) );
  MUX2_X1 U11901 ( .A(n11543), .B(n14740), .S(n10054), .Z(n9969) );
  INV_X1 U11902 ( .A(n9969), .ZN(n9967) );
  NAND2_X1 U11903 ( .A1(n9970), .A2(n9969), .ZN(n9972) );
  MUX2_X1 U11904 ( .A(n11543), .B(n14740), .S(n9949), .Z(n9971) );
  INV_X1 U11905 ( .A(n11709), .ZN(n11704) );
  MUX2_X1 U11906 ( .A(n11694), .B(n11704), .S(n9949), .Z(n9974) );
  MUX2_X1 U11907 ( .A(n11694), .B(n11704), .S(n10054), .Z(n9973) );
  MUX2_X1 U11908 ( .A(n11858), .B(n14739), .S(n10054), .Z(n9976) );
  MUX2_X1 U11909 ( .A(n11858), .B(n14739), .S(n9949), .Z(n9975) );
  MUX2_X1 U11910 ( .A(n14738), .B(n12198), .S(n10054), .Z(n9978) );
  MUX2_X1 U11911 ( .A(n12198), .B(n14738), .S(n10054), .Z(n9977) );
  MUX2_X1 U11912 ( .A(n12273), .B(n14737), .S(n10054), .Z(n9982) );
  NAND2_X1 U11913 ( .A1(n9981), .A2(n9982), .ZN(n9980) );
  MUX2_X1 U11914 ( .A(n12273), .B(n14737), .S(n10053), .Z(n9979) );
  NAND2_X1 U11915 ( .A1(n9980), .A2(n9979), .ZN(n9986) );
  NAND2_X1 U11916 ( .A1(n9984), .A2(n9983), .ZN(n9985) );
  MUX2_X1 U11917 ( .A(n12364), .B(n12565), .S(n10053), .Z(n9989) );
  MUX2_X1 U11918 ( .A(n12565), .B(n12364), .S(n10053), .Z(n9987) );
  MUX2_X1 U11919 ( .A(n14736), .B(n15900), .S(n9949), .Z(n9991) );
  MUX2_X1 U11920 ( .A(n14736), .B(n15900), .S(n10054), .Z(n9990) );
  INV_X1 U11921 ( .A(n9991), .ZN(n9992) );
  MUX2_X1 U11922 ( .A(n14735), .B(n12915), .S(n10054), .Z(n9996) );
  NAND2_X1 U11923 ( .A1(n9995), .A2(n9996), .ZN(n9994) );
  MUX2_X1 U11924 ( .A(n14735), .B(n12915), .S(n10053), .Z(n9993) );
  INV_X1 U11925 ( .A(n9995), .ZN(n9998) );
  INV_X1 U11926 ( .A(n9996), .ZN(n9997) );
  INV_X1 U11927 ( .A(n14649), .ZN(n14734) );
  MUX2_X1 U11928 ( .A(n12921), .B(n14734), .S(n10054), .Z(n10002) );
  NAND2_X1 U11929 ( .A1(n10001), .A2(n10002), .ZN(n10000) );
  MUX2_X1 U11930 ( .A(n14734), .B(n12921), .S(n10054), .Z(n9999) );
  MUX2_X1 U11931 ( .A(n15950), .B(n15979), .S(n10053), .Z(n10005) );
  MUX2_X1 U11932 ( .A(n15979), .B(n15950), .S(n10053), .Z(n10004) );
  MUX2_X1 U11933 ( .A(n15058), .B(n15077), .S(n10053), .Z(n10008) );
  MUX2_X1 U11934 ( .A(n15058), .B(n15077), .S(n10054), .Z(n10006) );
  MUX2_X1 U11935 ( .A(n16008), .B(n15977), .S(n10053), .Z(n10010) );
  MUX2_X1 U11936 ( .A(n16008), .B(n15977), .S(n10054), .Z(n10009) );
  INV_X1 U11937 ( .A(n10010), .ZN(n10011) );
  MUX2_X1 U11938 ( .A(n15057), .B(n16026), .S(n10053), .Z(n10015) );
  NAND2_X1 U11939 ( .A1(n10014), .A2(n10015), .ZN(n10013) );
  MUX2_X1 U11940 ( .A(n15057), .B(n16026), .S(n10054), .Z(n10012) );
  MUX2_X1 U11941 ( .A(n15175), .B(n15001), .S(n10053), .Z(n10019) );
  MUX2_X1 U11942 ( .A(n15001), .B(n15175), .S(n10053), .Z(n10018) );
  INV_X1 U11943 ( .A(n10019), .ZN(n10020) );
  MUX2_X1 U11944 ( .A(n15031), .B(n15170), .S(n10053), .Z(n10024) );
  NAND2_X1 U11945 ( .A1(n10023), .A2(n10024), .ZN(n10022) );
  MUX2_X1 U11946 ( .A(n15170), .B(n15031), .S(n10053), .Z(n10021) );
  INV_X1 U11947 ( .A(n10023), .ZN(n10026) );
  INV_X1 U11948 ( .A(n10024), .ZN(n10025) );
  MUX2_X1 U11949 ( .A(n14733), .B(n14988), .S(n10053), .Z(n10027) );
  INV_X1 U11950 ( .A(n14965), .ZN(n14953) );
  AND2_X1 U11951 ( .A1(n14984), .A2(n10053), .ZN(n10031) );
  OAI21_X1 U11952 ( .B1(n10053), .B2(n14984), .A(n15154), .ZN(n10030) );
  OAI21_X1 U11953 ( .B1(n10031), .B2(n15154), .A(n10030), .ZN(n10032) );
  MUX2_X1 U11954 ( .A(n10034), .B(n12884), .S(n10053), .Z(n10035) );
  MUX2_X1 U11955 ( .A(n14958), .B(n15141), .S(n10053), .Z(n10039) );
  MUX2_X1 U11956 ( .A(n14958), .B(n15141), .S(n10054), .Z(n10037) );
  MUX2_X1 U11957 ( .A(n14731), .B(n15135), .S(n10054), .Z(n10042) );
  MUX2_X1 U11958 ( .A(n14731), .B(n15135), .S(n10053), .Z(n10041) );
  MUX2_X1 U11959 ( .A(n14730), .B(n14919), .S(n10053), .Z(n10045) );
  MUX2_X1 U11960 ( .A(n14730), .B(n14919), .S(n10054), .Z(n10044) );
  INV_X1 U11961 ( .A(n14888), .ZN(n14729) );
  MUX2_X1 U11962 ( .A(n14729), .B(n15121), .S(n10054), .Z(n10049) );
  NAND2_X1 U11963 ( .A1(n10048), .A2(n10049), .ZN(n10047) );
  MUX2_X1 U11964 ( .A(n14729), .B(n15121), .S(n10053), .Z(n10046) );
  INV_X1 U11965 ( .A(n10048), .ZN(n10051) );
  INV_X1 U11966 ( .A(n10049), .ZN(n10050) );
  NAND2_X1 U11967 ( .A1(n10051), .A2(n10050), .ZN(n10052) );
  INV_X1 U11968 ( .A(n14904), .ZN(n14728) );
  MUX2_X1 U11969 ( .A(n15114), .B(n14728), .S(n10053), .Z(n10056) );
  MUX2_X1 U11970 ( .A(n15114), .B(n14728), .S(n10054), .Z(n10055) );
  NAND3_X1 U11971 ( .A1(n10067), .A2(n10065), .A3(n10058), .ZN(n10095) );
  INV_X1 U11972 ( .A(n10084), .ZN(n10059) );
  NAND2_X1 U11973 ( .A1(n10063), .A2(n10062), .ZN(n10070) );
  INV_X1 U11974 ( .A(n10078), .ZN(n10064) );
  NAND2_X1 U11975 ( .A1(n10064), .A2(n10105), .ZN(n10075) );
  INV_X1 U11976 ( .A(n10065), .ZN(n10068) );
  AOI211_X1 U11977 ( .C1(n10068), .C2(n10067), .A(n12759), .B(n10066), .ZN(
        n10069) );
  INV_X1 U11978 ( .A(n10069), .ZN(n10074) );
  INV_X1 U11979 ( .A(n10070), .ZN(n10071) );
  NAND2_X1 U11980 ( .A1(n10072), .A2(n10071), .ZN(n10073) );
  INV_X1 U11981 ( .A(n10081), .ZN(n10082) );
  NAND3_X1 U11982 ( .A1(n10084), .A2(n10083), .A3(n10082), .ZN(n10096) );
  NAND2_X1 U11983 ( .A1(n10087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10089) );
  OR2_X1 U11984 ( .A1(n10725), .A2(n10715), .ZN(n10928) );
  INV_X1 U11985 ( .A(n15227), .ZN(n15379) );
  INV_X1 U11986 ( .A(n10725), .ZN(n10874) );
  INV_X1 U11987 ( .A(n15223), .ZN(n10985) );
  NAND3_X1 U11988 ( .A1(n11494), .A2(n15379), .A3(n15075), .ZN(n10093) );
  OAI211_X1 U11989 ( .C1(n15236), .C2(n12759), .A(n10093), .B(P1_B_REG_SCAN_IN), .ZN(n10094) );
  OAI21_X1 U11990 ( .B1(n10096), .B2(n10095), .A(n10094), .ZN(n10097) );
  INV_X1 U11991 ( .A(n10097), .ZN(n10098) );
  NAND2_X1 U11992 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  AOI21_X1 U11993 ( .B1(n10102), .B2(n10101), .A(n10100), .ZN(n10103) );
  INV_X1 U11994 ( .A(n10107), .ZN(n10108) );
  NAND2_X1 U11995 ( .A1(n10109), .A2(n10108), .ZN(n10111) );
  NAND2_X1 U11996 ( .A1(n15221), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10110) );
  XNOR2_X1 U11997 ( .A(n15218), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n10115) );
  XNOR2_X1 U11998 ( .A(n10117), .B(n10115), .ZN(n13782) );
  NAND2_X1 U11999 ( .A1(n13782), .A2(n10142), .ZN(n10114) );
  NAND2_X1 U12000 ( .A1(n10112), .A2(SI_29_), .ZN(n10113) );
  NAND2_X1 U12001 ( .A1(n10114), .A2(n10113), .ZN(n10637) );
  OR2_X1 U12002 ( .A1(n10637), .A2(n13108), .ZN(n10287) );
  INV_X1 U12003 ( .A(n10115), .ZN(n10116) );
  NAND2_X1 U12004 ( .A1(n10117), .A2(n10116), .ZN(n10119) );
  NAND2_X1 U12005 ( .A1(n15218), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n10118) );
  NAND2_X1 U12006 ( .A1(n10119), .A2(n10118), .ZN(n10134) );
  XNOR2_X1 U12007 ( .A(n15217), .B(P1_DATAO_REG_30__SCAN_IN), .ZN(n10132) );
  XNOR2_X1 U12008 ( .A(n10134), .B(n10132), .ZN(n13034) );
  NAND2_X1 U12009 ( .A1(n13034), .A2(n10142), .ZN(n10121) );
  INV_X1 U12010 ( .A(SI_30_), .ZN(n13882) );
  OR2_X1 U12011 ( .A1(n7486), .A2(n13882), .ZN(n10120) );
  NAND2_X1 U12012 ( .A1(n10121), .A2(n10120), .ZN(n10131) );
  NAND2_X1 U12013 ( .A1(n10125), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U12014 ( .A1(n8558), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U12015 ( .A1(n10126), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10122) );
  NAND4_X1 U12016 ( .A1(n10130), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n13429) );
  NAND2_X1 U12017 ( .A1(n8558), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U12018 ( .A1(n10125), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n10128) );
  NAND2_X1 U12019 ( .A1(n10126), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n10127) );
  NAND2_X1 U12020 ( .A1(n10131), .A2(n10630), .ZN(n10298) );
  NAND2_X1 U12021 ( .A1(n10637), .A2(n13108), .ZN(n10284) );
  AND2_X1 U12022 ( .A1(n10298), .A2(n10284), .ZN(n10290) );
  OAI21_X1 U12023 ( .B1(n13708), .B2(n13429), .A(n10290), .ZN(n10143) );
  INV_X1 U12024 ( .A(n10132), .ZN(n10133) );
  NAND2_X1 U12025 ( .A1(n10134), .A2(n10133), .ZN(n10136) );
  NAND2_X1 U12026 ( .A1(n15217), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10135) );
  NAND2_X1 U12027 ( .A1(n10136), .A2(n10135), .ZN(n10139) );
  INV_X1 U12028 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10137) );
  XNOR2_X1 U12029 ( .A(n10137), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n10138) );
  XNOR2_X1 U12030 ( .A(n10139), .B(n10138), .ZN(n13780) );
  INV_X1 U12031 ( .A(SI_31_), .ZN(n13775) );
  NOR2_X1 U12032 ( .A1(n7486), .A2(n13775), .ZN(n10141) );
  AND2_X1 U12033 ( .A1(n13705), .A2(n13429), .ZN(n10296) );
  INV_X1 U12034 ( .A(n13705), .ZN(n10145) );
  INV_X1 U12035 ( .A(n13429), .ZN(n10144) );
  INV_X1 U12036 ( .A(n10630), .ZN(n13202) );
  AND2_X1 U12037 ( .A1(n13708), .A2(n13202), .ZN(n10317) );
  NAND2_X1 U12038 ( .A1(n10154), .A2(n10259), .ZN(n13468) );
  INV_X1 U12039 ( .A(n13503), .ZN(n13498) );
  NAND2_X1 U12040 ( .A1(n13482), .A2(n13498), .ZN(n10155) );
  NOR2_X1 U12041 ( .A1(n13468), .A2(n10155), .ZN(n10156) );
  NAND2_X1 U12042 ( .A1(n13224), .A2(n8118), .ZN(n10305) );
  NAND2_X1 U12043 ( .A1(n10157), .A2(n10305), .ZN(n10158) );
  NAND2_X1 U12044 ( .A1(n10162), .A2(n10158), .ZN(n10164) );
  OAI211_X1 U12045 ( .C1(n11818), .C2(n10164), .A(n10160), .B(n10159), .ZN(
        n10161) );
  NAND2_X1 U12046 ( .A1(n10161), .A2(n10166), .ZN(n10169) );
  NAND3_X1 U12047 ( .A1(n11739), .A2(n10162), .A3(n11900), .ZN(n10163) );
  NAND3_X1 U12048 ( .A1(n8773), .A2(n10164), .A3(n10163), .ZN(n10167) );
  AND3_X1 U12049 ( .A1(n10167), .A2(n10166), .A3(n10165), .ZN(n10168) );
  MUX2_X1 U12050 ( .A(n10169), .B(n10168), .S(n10276), .Z(n10172) );
  OR2_X1 U12051 ( .A1(n11443), .A2(n11040), .ZN(n10170) );
  NOR2_X1 U12052 ( .A1(n8398), .A2(n10170), .ZN(n10171) );
  OAI21_X1 U12053 ( .B1(n10172), .B2(n10171), .A(n12069), .ZN(n10176) );
  NAND2_X1 U12054 ( .A1(n13220), .A2(n15737), .ZN(n10173) );
  MUX2_X1 U12055 ( .A(n10174), .B(n10173), .S(n10276), .Z(n10175) );
  NAND3_X1 U12056 ( .A1(n10176), .A2(n12233), .A3(n10175), .ZN(n10180) );
  MUX2_X1 U12057 ( .A(n10178), .B(n10177), .S(n10276), .Z(n10179) );
  NAND3_X1 U12058 ( .A1(n10180), .A2(n12215), .A3(n10179), .ZN(n10184) );
  MUX2_X1 U12059 ( .A(n10182), .B(n10181), .S(n11040), .Z(n10183) );
  AOI21_X1 U12060 ( .B1(n10184), .B2(n10183), .A(n12123), .ZN(n10192) );
  MUX2_X1 U12061 ( .A(n10186), .B(n10185), .S(n11040), .Z(n10187) );
  NAND2_X1 U12062 ( .A1(n10187), .A2(n12299), .ZN(n10191) );
  INV_X1 U12063 ( .A(n12394), .ZN(n10307) );
  MUX2_X1 U12064 ( .A(n10189), .B(n10188), .S(n10276), .Z(n10190) );
  OAI211_X1 U12065 ( .C1(n10192), .C2(n10191), .A(n10307), .B(n10190), .ZN(
        n10196) );
  MUX2_X1 U12066 ( .A(n10194), .B(n10193), .S(n11040), .Z(n10195) );
  NAND2_X1 U12067 ( .A1(n10196), .A2(n10195), .ZN(n10201) );
  MUX2_X1 U12068 ( .A(n10198), .B(n10197), .S(n11040), .Z(n10199) );
  NAND2_X1 U12069 ( .A1(n10199), .A2(n12717), .ZN(n10200) );
  AOI21_X1 U12070 ( .B1(n10201), .B2(n8149), .A(n10200), .ZN(n10208) );
  NAND2_X1 U12071 ( .A1(n12734), .A2(n10202), .ZN(n10204) );
  NAND2_X1 U12072 ( .A1(n10205), .A2(n12778), .ZN(n10203) );
  MUX2_X1 U12073 ( .A(n10204), .B(n10203), .S(n11040), .Z(n10207) );
  INV_X1 U12074 ( .A(n12806), .ZN(n12737) );
  MUX2_X1 U12075 ( .A(n10205), .B(n12734), .S(n11040), .Z(n10206) );
  OAI211_X1 U12076 ( .C1(n10208), .C2(n10207), .A(n12737), .B(n10206), .ZN(
        n10209) );
  NAND2_X1 U12077 ( .A1(n10209), .A2(n12768), .ZN(n10218) );
  INV_X1 U12078 ( .A(n10210), .ZN(n10212) );
  OAI21_X1 U12079 ( .B1(n10218), .B2(n10212), .A(n10211), .ZN(n10215) );
  INV_X1 U12080 ( .A(n10213), .ZN(n10214) );
  AOI21_X1 U12081 ( .B1(n10215), .B2(n12822), .A(n10214), .ZN(n10223) );
  OAI21_X1 U12082 ( .B1(n10218), .B2(n8777), .A(n10217), .ZN(n10221) );
  INV_X1 U12083 ( .A(n10219), .ZN(n10220) );
  AOI21_X1 U12084 ( .B1(n10221), .B2(n12822), .A(n10220), .ZN(n10222) );
  MUX2_X1 U12085 ( .A(n10223), .B(n10222), .S(n11040), .Z(n10228) );
  MUX2_X1 U12086 ( .A(n10225), .B(n10224), .S(n10276), .Z(n10226) );
  INV_X1 U12087 ( .A(n10226), .ZN(n10227) );
  AOI21_X1 U12088 ( .B1(n10228), .B2(n13631), .A(n10227), .ZN(n10241) );
  NAND2_X1 U12089 ( .A1(n13593), .A2(n13612), .ZN(n10302) );
  INV_X1 U12090 ( .A(n10229), .ZN(n10230) );
  NAND2_X1 U12091 ( .A1(n10235), .A2(n10230), .ZN(n10231) );
  AND3_X1 U12092 ( .A1(n10300), .A2(n10234), .A3(n10231), .ZN(n10239) );
  INV_X1 U12093 ( .A(n10232), .ZN(n10233) );
  NAND2_X1 U12094 ( .A1(n10234), .A2(n10233), .ZN(n10236) );
  NAND2_X1 U12095 ( .A1(n10236), .A2(n10235), .ZN(n10237) );
  NOR2_X1 U12096 ( .A1(n10301), .A2(n10237), .ZN(n10238) );
  MUX2_X1 U12097 ( .A(n10239), .B(n10238), .S(n10276), .Z(n10240) );
  OAI21_X1 U12098 ( .B1(n10241), .B2(n10302), .A(n10240), .ZN(n10244) );
  INV_X1 U12099 ( .A(n10301), .ZN(n10242) );
  MUX2_X1 U12100 ( .A(n10300), .B(n10242), .S(n11040), .Z(n10243) );
  NAND3_X1 U12101 ( .A1(n10244), .A2(n8779), .A3(n10243), .ZN(n10248) );
  MUX2_X1 U12102 ( .A(n10246), .B(n10245), .S(n10276), .Z(n10247) );
  NAND3_X1 U12103 ( .A1(n10248), .A2(n13542), .A3(n10247), .ZN(n10252) );
  NAND2_X1 U12104 ( .A1(n13120), .A2(n13206), .ZN(n10250) );
  MUX2_X1 U12105 ( .A(n10250), .B(n10249), .S(n11040), .Z(n10251) );
  NAND3_X1 U12106 ( .A1(n10252), .A2(n7745), .A3(n10251), .ZN(n10256) );
  MUX2_X1 U12107 ( .A(n10254), .B(n10253), .S(n11040), .Z(n10255) );
  NAND3_X1 U12108 ( .A1(n10256), .A2(n13513), .A3(n10255), .ZN(n10257) );
  OAI21_X1 U12109 ( .B1(n11040), .B2(n13499), .A(n10257), .ZN(n10258) );
  NAND2_X1 U12110 ( .A1(n10299), .A2(n10258), .ZN(n10283) );
  INV_X1 U12111 ( .A(n13468), .ZN(n13470) );
  NAND2_X1 U12112 ( .A1(n10260), .A2(n10259), .ZN(n10262) );
  OR2_X1 U12113 ( .A1(n13463), .A2(n13100), .ZN(n10261) );
  NAND2_X1 U12114 ( .A1(n10262), .A2(n10261), .ZN(n10278) );
  NAND2_X1 U12115 ( .A1(n13104), .A2(n10263), .ZN(n10269) );
  NAND2_X1 U12116 ( .A1(n10265), .A2(n10264), .ZN(n10270) );
  AND4_X1 U12117 ( .A1(n13454), .A2(n13470), .A3(n10273), .A4(n10270), .ZN(
        n10268) );
  XNOR2_X1 U12118 ( .A(n10266), .B(n10276), .ZN(n10267) );
  OAI21_X1 U12119 ( .B1(n10269), .B2(n10268), .A(n10267), .ZN(n10282) );
  INV_X1 U12120 ( .A(n10269), .ZN(n10280) );
  INV_X1 U12121 ( .A(n10270), .ZN(n10275) );
  NAND2_X1 U12122 ( .A1(n10272), .A2(n10271), .ZN(n10274) );
  AOI21_X1 U12123 ( .B1(n10275), .B2(n10274), .A(n8127), .ZN(n10277) );
  AOI21_X1 U12124 ( .B1(n10278), .B2(n10277), .A(n10276), .ZN(n10279) );
  NAND2_X1 U12125 ( .A1(n10280), .A2(n10279), .ZN(n10281) );
  NAND3_X1 U12126 ( .A1(n10283), .A2(n10282), .A3(n10281), .ZN(n10286) );
  INV_X1 U12127 ( .A(n10635), .ZN(n10285) );
  NAND2_X1 U12128 ( .A1(n10286), .A2(n10285), .ZN(n10291) );
  INV_X1 U12129 ( .A(n10317), .ZN(n10292) );
  AND2_X1 U12130 ( .A1(n10292), .A2(n10287), .ZN(n10289) );
  INV_X1 U12131 ( .A(n10298), .ZN(n10288) );
  AOI21_X1 U12132 ( .B1(n10291), .B2(n10289), .A(n10288), .ZN(n10295) );
  NAND2_X1 U12133 ( .A1(n10291), .A2(n10290), .ZN(n10293) );
  NAND2_X1 U12134 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  INV_X1 U12135 ( .A(n10296), .ZN(n10319) );
  INV_X1 U12136 ( .A(n11821), .ZN(n10323) );
  NOR2_X1 U12137 ( .A1(n10301), .A2(n8151), .ZN(n13578) );
  INV_X1 U12138 ( .A(n10302), .ZN(n10314) );
  AND2_X1 U12139 ( .A1(n8773), .A2(n12233), .ZN(n10304) );
  NOR2_X1 U12140 ( .A1(n12218), .A2(n12123), .ZN(n10303) );
  NAND4_X1 U12141 ( .A1(n10304), .A2(n12069), .A3(n8149), .A4(n10303), .ZN(
        n10310) );
  NAND2_X1 U12142 ( .A1(n11739), .A2(n10305), .ZN(n11247) );
  NOR2_X1 U12143 ( .A1(n12140), .A2(n11247), .ZN(n10308) );
  INV_X1 U12144 ( .A(n10306), .ZN(n11740) );
  NAND4_X1 U12145 ( .A1(n10308), .A2(n12299), .A3(n10307), .A4(n11740), .ZN(
        n10309) );
  NOR2_X1 U12146 ( .A1(n10310), .A2(n10309), .ZN(n10311) );
  NAND4_X1 U12147 ( .A1(n10311), .A2(n12717), .A3(n12737), .A4(n12773), .ZN(
        n10312) );
  NOR3_X1 U12148 ( .A1(n12817), .A2(n12763), .A3(n10312), .ZN(n10313) );
  NAND4_X1 U12149 ( .A1(n13578), .A2(n13631), .A3(n10314), .A4(n10313), .ZN(
        n10315) );
  NOR2_X1 U12150 ( .A1(n13552), .A2(n10315), .ZN(n10316) );
  NAND3_X1 U12151 ( .A1(n10320), .A2(n10147), .A3(n10319), .ZN(n10321) );
  XNOR2_X1 U12152 ( .A(n10321), .B(n13412), .ZN(n10322) );
  OAI22_X1 U12153 ( .A1(n10326), .A2(n10323), .B1(n10322), .B2(n11295), .ZN(
        n10324) );
  OR2_X1 U12154 ( .A1(n11200), .A2(P3_U3151), .ZN(n12113) );
  NOR3_X1 U12155 ( .A1(n11215), .A2(n10329), .A3(n12903), .ZN(n10332) );
  OAI21_X1 U12156 ( .B1(n12113), .B2(n10330), .A(P3_B_REG_SCAN_IN), .ZN(n10331) );
  OR2_X1 U12157 ( .A1(n10332), .A2(n10331), .ZN(n10333) );
  NAND2_X1 U12158 ( .A1(n10345), .A2(n11383), .ZN(n10337) );
  NAND2_X1 U12159 ( .A1(n14193), .A2(n10375), .ZN(n10336) );
  NAND2_X1 U12160 ( .A1(n10345), .A2(n14193), .ZN(n10339) );
  NAND2_X1 U12161 ( .A1(n11383), .A2(n10375), .ZN(n10338) );
  NAND2_X1 U12162 ( .A1(n10345), .A2(n11397), .ZN(n10341) );
  NAND2_X1 U12163 ( .A1(n10335), .A2(n10348), .ZN(n10340) );
  NAND2_X1 U12164 ( .A1(n10344), .A2(n11292), .ZN(n10343) );
  INV_X1 U12165 ( .A(n11094), .ZN(n10583) );
  NAND2_X1 U12166 ( .A1(n10347), .A2(n10346), .ZN(n10351) );
  NAND2_X1 U12167 ( .A1(n10345), .A2(n10348), .ZN(n10350) );
  NAND2_X1 U12168 ( .A1(n10375), .A2(n11397), .ZN(n10349) );
  INV_X1 U12169 ( .A(n10353), .ZN(n10356) );
  INV_X1 U12170 ( .A(n10354), .ZN(n10355) );
  NAND2_X1 U12171 ( .A1(n10356), .A2(n10355), .ZN(n10357) );
  NAND2_X1 U12172 ( .A1(n11336), .A2(n10550), .ZN(n10359) );
  NAND2_X1 U12173 ( .A1(n14192), .A2(n10372), .ZN(n10358) );
  NAND2_X1 U12174 ( .A1(n10359), .A2(n10358), .ZN(n10364) );
  NAND2_X1 U12175 ( .A1(n10363), .A2(n10364), .ZN(n10362) );
  AOI22_X1 U12176 ( .A1(n11336), .A2(n10372), .B1(n14192), .B2(n10550), .ZN(
        n10360) );
  INV_X1 U12177 ( .A(n10360), .ZN(n10361) );
  NAND2_X1 U12178 ( .A1(n10362), .A2(n10361), .ZN(n10368) );
  NAND2_X1 U12179 ( .A1(n10366), .A2(n10365), .ZN(n10367) );
  NAND2_X1 U12180 ( .A1(n11473), .A2(n10372), .ZN(n10370) );
  NAND2_X1 U12181 ( .A1(n10396), .A2(n14191), .ZN(n10369) );
  NAND2_X1 U12182 ( .A1(n10370), .A2(n10369), .ZN(n10377) );
  NOR2_X1 U12183 ( .A1(n11429), .A2(n10550), .ZN(n10371) );
  AOI21_X1 U12184 ( .B1(n11405), .B2(n10396), .A(n10371), .ZN(n10380) );
  NAND2_X1 U12185 ( .A1(n11405), .A2(n10372), .ZN(n10374) );
  NAND2_X1 U12186 ( .A1(n10396), .A2(n14190), .ZN(n10373) );
  NAND2_X1 U12187 ( .A1(n10374), .A2(n10373), .ZN(n10379) );
  AOI22_X1 U12188 ( .A1(n11473), .A2(n10396), .B1(n10545), .B2(n14191), .ZN(
        n10376) );
  AOI21_X1 U12189 ( .B1(n10378), .B2(n10377), .A(n10376), .ZN(n10382) );
  NAND2_X1 U12190 ( .A1(n10380), .A2(n10379), .ZN(n10381) );
  NAND2_X1 U12191 ( .A1(n15801), .A2(n10554), .ZN(n10385) );
  NAND2_X1 U12192 ( .A1(n10396), .A2(n14189), .ZN(n10384) );
  NAND2_X1 U12193 ( .A1(n10385), .A2(n10384), .ZN(n10391) );
  NAND2_X1 U12194 ( .A1(n10390), .A2(n10391), .ZN(n10389) );
  NAND2_X1 U12195 ( .A1(n15801), .A2(n7394), .ZN(n10387) );
  NAND2_X1 U12196 ( .A1(n10554), .A2(n14189), .ZN(n10386) );
  NAND2_X1 U12197 ( .A1(n10387), .A2(n10386), .ZN(n10388) );
  NAND2_X1 U12198 ( .A1(n10389), .A2(n10388), .ZN(n10395) );
  INV_X1 U12199 ( .A(n10390), .ZN(n10393) );
  INV_X1 U12200 ( .A(n10391), .ZN(n10392) );
  NAND2_X1 U12201 ( .A1(n10393), .A2(n10392), .ZN(n10394) );
  NAND2_X1 U12202 ( .A1(n15831), .A2(n10396), .ZN(n10398) );
  NAND2_X1 U12203 ( .A1(n10554), .A2(n14188), .ZN(n10397) );
  AOI22_X1 U12204 ( .A1(n15831), .A2(n10554), .B1(n14188), .B2(n10550), .ZN(
        n10399) );
  NAND2_X1 U12205 ( .A1(n11654), .A2(n10554), .ZN(n10401) );
  NAND2_X1 U12206 ( .A1(n10396), .A2(n14187), .ZN(n10400) );
  NAND2_X1 U12207 ( .A1(n10401), .A2(n10400), .ZN(n10407) );
  NAND2_X1 U12208 ( .A1(n11654), .A2(n7394), .ZN(n10403) );
  NAND2_X1 U12209 ( .A1(n10554), .A2(n14187), .ZN(n10402) );
  NAND2_X1 U12210 ( .A1(n10403), .A2(n10402), .ZN(n10404) );
  NAND2_X1 U12211 ( .A1(n10405), .A2(n10404), .ZN(n10409) );
  INV_X1 U12212 ( .A(n10407), .ZN(n10408) );
  NAND2_X1 U12213 ( .A1(n11998), .A2(n7394), .ZN(n10411) );
  NAND2_X1 U12214 ( .A1(n10554), .A2(n14185), .ZN(n10410) );
  NAND2_X1 U12215 ( .A1(n10411), .A2(n10410), .ZN(n10413) );
  AOI22_X1 U12216 ( .A1(n11998), .A2(n10554), .B1(n14185), .B2(n10550), .ZN(
        n10412) );
  NAND2_X1 U12217 ( .A1(n12043), .A2(n10554), .ZN(n10415) );
  NAND2_X1 U12218 ( .A1(n10396), .A2(n14184), .ZN(n10414) );
  NAND2_X1 U12219 ( .A1(n10415), .A2(n10414), .ZN(n10421) );
  NAND2_X1 U12220 ( .A1(n12043), .A2(n7394), .ZN(n10417) );
  NAND2_X1 U12221 ( .A1(n10554), .A2(n14184), .ZN(n10416) );
  NAND2_X1 U12222 ( .A1(n10417), .A2(n10416), .ZN(n10418) );
  NAND2_X1 U12223 ( .A1(n10419), .A2(n10418), .ZN(n10425) );
  INV_X1 U12224 ( .A(n10420), .ZN(n10423) );
  INV_X1 U12225 ( .A(n10421), .ZN(n10422) );
  NAND2_X1 U12226 ( .A1(n10423), .A2(n10422), .ZN(n10424) );
  NAND2_X1 U12227 ( .A1(n12279), .A2(n7394), .ZN(n10427) );
  NAND2_X1 U12228 ( .A1(n10554), .A2(n14183), .ZN(n10426) );
  NAND2_X1 U12229 ( .A1(n10427), .A2(n10426), .ZN(n10429) );
  AOI22_X1 U12230 ( .A1(n12279), .A2(n10554), .B1(n14183), .B2(n10550), .ZN(
        n10428) );
  NAND2_X1 U12231 ( .A1(n15918), .A2(n10554), .ZN(n10431) );
  NAND2_X1 U12232 ( .A1(n10396), .A2(n14182), .ZN(n10430) );
  NAND2_X1 U12233 ( .A1(n10431), .A2(n10430), .ZN(n10437) );
  NAND2_X1 U12234 ( .A1(n15918), .A2(n7394), .ZN(n10433) );
  NAND2_X1 U12235 ( .A1(n10545), .A2(n14182), .ZN(n10432) );
  NAND2_X1 U12236 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  NAND2_X1 U12237 ( .A1(n10435), .A2(n10434), .ZN(n10441) );
  INV_X1 U12238 ( .A(n10436), .ZN(n10439) );
  INV_X1 U12239 ( .A(n10437), .ZN(n10438) );
  NAND2_X1 U12240 ( .A1(n10439), .A2(n10438), .ZN(n10440) );
  NAND2_X1 U12241 ( .A1(n12537), .A2(n7394), .ZN(n10443) );
  NAND2_X1 U12242 ( .A1(n10545), .A2(n14181), .ZN(n10442) );
  NAND2_X1 U12243 ( .A1(n10443), .A2(n10442), .ZN(n10445) );
  AOI22_X1 U12244 ( .A1(n12537), .A2(n10554), .B1(n14181), .B2(n10550), .ZN(
        n10444) );
  NAND2_X1 U12245 ( .A1(n12655), .A2(n10545), .ZN(n10449) );
  NAND2_X1 U12246 ( .A1(n10550), .A2(n14180), .ZN(n10448) );
  NAND2_X1 U12247 ( .A1(n10449), .A2(n10448), .ZN(n10451) );
  AOI22_X1 U12248 ( .A1(n12655), .A2(n7394), .B1(n10554), .B2(n14180), .ZN(
        n10450) );
  NAND2_X1 U12249 ( .A1(n15960), .A2(n7394), .ZN(n10454) );
  NAND2_X1 U12250 ( .A1(n14179), .A2(n10554), .ZN(n10453) );
  NAND2_X1 U12251 ( .A1(n10454), .A2(n10453), .ZN(n10458) );
  NAND2_X1 U12252 ( .A1(n15960), .A2(n10554), .ZN(n10456) );
  NAND2_X1 U12253 ( .A1(n14179), .A2(n10550), .ZN(n10455) );
  NAND2_X1 U12254 ( .A1(n14512), .A2(n10554), .ZN(n10460) );
  NAND2_X1 U12255 ( .A1(n14178), .A2(n7394), .ZN(n10459) );
  NAND2_X1 U12256 ( .A1(n10460), .A2(n10459), .ZN(n10465) );
  NAND2_X1 U12257 ( .A1(n10464), .A2(n10465), .ZN(n10463) );
  AOI22_X1 U12258 ( .A1(n14512), .A2(n7394), .B1(n10545), .B2(n14178), .ZN(
        n10461) );
  NAND2_X1 U12259 ( .A1(n10463), .A2(n10462), .ZN(n10469) );
  INV_X1 U12260 ( .A(n10464), .ZN(n10467) );
  INV_X1 U12261 ( .A(n10465), .ZN(n10466) );
  NAND2_X1 U12262 ( .A1(n10467), .A2(n10466), .ZN(n10468) );
  AND2_X1 U12263 ( .A1(n14177), .A2(n10545), .ZN(n10470) );
  AOI21_X1 U12264 ( .B1(n14557), .B2(n7394), .A(n10470), .ZN(n10471) );
  INV_X1 U12265 ( .A(n10471), .ZN(n10472) );
  NAND2_X1 U12266 ( .A1(n14557), .A2(n10554), .ZN(n10474) );
  NAND2_X1 U12267 ( .A1(n14500), .A2(n10545), .ZN(n10478) );
  NAND2_X1 U12268 ( .A1(n14176), .A2(n7394), .ZN(n10477) );
  NAND2_X1 U12269 ( .A1(n10478), .A2(n10477), .ZN(n10480) );
  AOI22_X1 U12270 ( .A1(n14500), .A2(n7394), .B1(n10554), .B2(n14176), .ZN(
        n10479) );
  NAND2_X1 U12271 ( .A1(n14405), .A2(n7394), .ZN(n10482) );
  NAND2_X1 U12272 ( .A1(n14175), .A2(n10554), .ZN(n10481) );
  NAND2_X1 U12273 ( .A1(n10482), .A2(n10481), .ZN(n10488) );
  NAND2_X1 U12274 ( .A1(n10487), .A2(n10488), .ZN(n10486) );
  NAND2_X1 U12275 ( .A1(n14405), .A2(n10554), .ZN(n10484) );
  NAND2_X1 U12276 ( .A1(n14175), .A2(n7394), .ZN(n10483) );
  NAND2_X1 U12277 ( .A1(n10484), .A2(n10483), .ZN(n10485) );
  NAND2_X1 U12278 ( .A1(n10486), .A2(n10485), .ZN(n10492) );
  INV_X1 U12279 ( .A(n10487), .ZN(n10490) );
  INV_X1 U12280 ( .A(n10488), .ZN(n10489) );
  NAND2_X1 U12281 ( .A1(n10490), .A2(n10489), .ZN(n10491) );
  NAND2_X1 U12282 ( .A1(n14392), .A2(n10554), .ZN(n10494) );
  NAND2_X1 U12283 ( .A1(n14174), .A2(n7394), .ZN(n10493) );
  NAND2_X1 U12284 ( .A1(n10494), .A2(n10493), .ZN(n10496) );
  AOI22_X1 U12285 ( .A1(n14392), .A2(n7394), .B1(n10545), .B2(n14174), .ZN(
        n10495) );
  NAND2_X1 U12286 ( .A1(n14376), .A2(n7394), .ZN(n10499) );
  NAND2_X1 U12287 ( .A1(n14173), .A2(n10545), .ZN(n10498) );
  NAND2_X1 U12288 ( .A1(n10499), .A2(n10498), .ZN(n10502) );
  NAND2_X1 U12289 ( .A1(n14376), .A2(n10554), .ZN(n10501) );
  NAND2_X1 U12290 ( .A1(n14173), .A2(n7394), .ZN(n10500) );
  NAND2_X1 U12291 ( .A1(n14540), .A2(n10554), .ZN(n10505) );
  NAND2_X1 U12292 ( .A1(n14172), .A2(n7394), .ZN(n10504) );
  AOI22_X1 U12293 ( .A1(n14540), .A2(n7394), .B1(n10545), .B2(n14172), .ZN(
        n10506) );
  NAND2_X1 U12294 ( .A1(n14469), .A2(n10550), .ZN(n10508) );
  NAND2_X1 U12295 ( .A1(n14171), .A2(n10554), .ZN(n10507) );
  NAND2_X1 U12296 ( .A1(n10508), .A2(n10507), .ZN(n10511) );
  AOI22_X1 U12297 ( .A1(n14469), .A2(n10554), .B1(n14171), .B2(n10550), .ZN(
        n10509) );
  AOI21_X1 U12298 ( .B1(n10512), .B2(n10511), .A(n10509), .ZN(n10510) );
  INV_X1 U12299 ( .A(n10510), .ZN(n10513) );
  NAND2_X1 U12300 ( .A1(n14466), .A2(n10545), .ZN(n10515) );
  NAND2_X1 U12301 ( .A1(n14170), .A2(n7394), .ZN(n10514) );
  NAND2_X1 U12302 ( .A1(n14466), .A2(n7394), .ZN(n10516) );
  OAI21_X1 U12303 ( .B1(n10517), .B2(n10396), .A(n10516), .ZN(n10518) );
  NAND2_X1 U12304 ( .A1(n14323), .A2(n10550), .ZN(n10520) );
  NAND2_X1 U12305 ( .A1(n14169), .A2(n10554), .ZN(n10519) );
  NAND2_X1 U12306 ( .A1(n10520), .A2(n10519), .ZN(n10521) );
  AOI22_X1 U12307 ( .A1(n14323), .A2(n10554), .B1(n14169), .B2(n10550), .ZN(
        n10523) );
  OAI22_X1 U12308 ( .A1(n14531), .A2(n10550), .B1(n14000), .B2(n10554), .ZN(
        n10525) );
  AOI22_X1 U12309 ( .A1(n7634), .A2(n7394), .B1(n10554), .B2(n14168), .ZN(
        n10524) );
  INV_X1 U12310 ( .A(n10525), .ZN(n10526) );
  NAND2_X1 U12311 ( .A1(n14561), .A2(n7478), .ZN(n10528) );
  NAND2_X1 U12312 ( .A1(n10534), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n10527) );
  INV_X1 U12313 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14436) );
  NAND2_X1 U12314 ( .A1(n7168), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n10531) );
  NAND2_X1 U12315 ( .A1(n10529), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n10530) );
  OAI211_X1 U12316 ( .C1(n10532), .C2(n14436), .A(n10531), .B(n10530), .ZN(
        n14247) );
  XNOR2_X1 U12317 ( .A(n10578), .B(n14247), .ZN(n10592) );
  NAND2_X1 U12318 ( .A1(n14567), .A2(n7478), .ZN(n10536) );
  NAND2_X1 U12319 ( .A1(n10534), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10535) );
  NAND2_X1 U12320 ( .A1(n10396), .A2(n14247), .ZN(n10577) );
  NAND2_X1 U12321 ( .A1(n10621), .A2(n11967), .ZN(n10587) );
  AND2_X1 U12322 ( .A1(n10537), .A2(n11390), .ZN(n10538) );
  AND2_X1 U12323 ( .A1(n10587), .A2(n10538), .ZN(n10540) );
  AOI21_X1 U12324 ( .B1(n10577), .B2(n10540), .A(n10539), .ZN(n10541) );
  AOI21_X1 U12325 ( .B1(n14524), .B2(n10545), .A(n10541), .ZN(n10571) );
  NAND2_X1 U12326 ( .A1(n14524), .A2(n7394), .ZN(n10543) );
  NAND2_X1 U12327 ( .A1(n10554), .A2(n14164), .ZN(n10542) );
  NAND2_X1 U12328 ( .A1(n10543), .A2(n10542), .ZN(n10570) );
  AND2_X1 U12329 ( .A1(n14165), .A2(n10550), .ZN(n10544) );
  AOI21_X1 U12330 ( .B1(n14262), .B2(n10554), .A(n10544), .ZN(n10568) );
  NAND2_X1 U12331 ( .A1(n14262), .A2(n7394), .ZN(n10547) );
  NAND2_X1 U12332 ( .A1(n14165), .A2(n10545), .ZN(n10546) );
  NAND2_X1 U12333 ( .A1(n10547), .A2(n10546), .ZN(n10567) );
  OAI22_X1 U12334 ( .A1(n10571), .A2(n10570), .B1(n10568), .B2(n10567), .ZN(
        n10548) );
  NAND2_X1 U12335 ( .A1(n10592), .A2(n10548), .ZN(n10573) );
  AND2_X1 U12336 ( .A1(n14166), .A2(n10554), .ZN(n10549) );
  AOI21_X1 U12337 ( .B1(n14444), .B2(n10550), .A(n10549), .ZN(n10564) );
  NAND2_X1 U12338 ( .A1(n14444), .A2(n10554), .ZN(n10552) );
  NAND2_X1 U12339 ( .A1(n14166), .A2(n7394), .ZN(n10551) );
  NAND2_X1 U12340 ( .A1(n10552), .A2(n10551), .ZN(n10563) );
  NAND2_X1 U12341 ( .A1(n10564), .A2(n10563), .ZN(n10553) );
  NAND2_X1 U12342 ( .A1(n14448), .A2(n10554), .ZN(n10556) );
  NAND2_X1 U12343 ( .A1(n14167), .A2(n7394), .ZN(n10555) );
  NAND2_X1 U12344 ( .A1(n10556), .A2(n10555), .ZN(n10560) );
  AND2_X1 U12345 ( .A1(n14167), .A2(n10554), .ZN(n10557) );
  AOI21_X1 U12346 ( .B1(n14448), .B2(n7394), .A(n10557), .ZN(n10559) );
  INV_X1 U12347 ( .A(n10559), .ZN(n10562) );
  INV_X1 U12348 ( .A(n10560), .ZN(n10561) );
  NAND2_X1 U12349 ( .A1(n10562), .A2(n10561), .ZN(n10575) );
  INV_X1 U12350 ( .A(n10563), .ZN(n10566) );
  INV_X1 U12351 ( .A(n10564), .ZN(n10565) );
  AOI22_X1 U12352 ( .A1(n10568), .A2(n10567), .B1(n10566), .B2(n10565), .ZN(
        n10569) );
  NAND2_X1 U12353 ( .A1(n10592), .A2(n10569), .ZN(n10572) );
  AOI22_X1 U12354 ( .A1(n10573), .A2(n10572), .B1(n10571), .B2(n10570), .ZN(
        n10574) );
  OAI21_X1 U12355 ( .B1(n10576), .B2(n10575), .A(n10574), .ZN(n10582) );
  NAND2_X1 U12356 ( .A1(n10554), .A2(n14247), .ZN(n10580) );
  NAND2_X1 U12357 ( .A1(n10577), .A2(n10396), .ZN(n10579) );
  MUX2_X1 U12358 ( .A(n10580), .B(n10579), .S(n10578), .Z(n10581) );
  AOI21_X1 U12359 ( .B1(n10583), .B2(n12792), .A(n9420), .ZN(n10584) );
  AOI21_X1 U12360 ( .B1(n7198), .B2(n12669), .A(n10584), .ZN(n10585) );
  INV_X1 U12361 ( .A(n10585), .ZN(n10590) );
  NAND3_X1 U12362 ( .A1(n11390), .A2(n15339), .A3(n7198), .ZN(n10586) );
  NAND2_X1 U12363 ( .A1(n10587), .A2(n10586), .ZN(n10588) );
  OAI21_X1 U12364 ( .B1(n10591), .B2(n10590), .A(n10589), .ZN(n10619) );
  INV_X1 U12365 ( .A(n10592), .ZN(n10613) );
  XNOR2_X1 U12366 ( .A(n14524), .B(n14164), .ZN(n10611) );
  XNOR2_X1 U12367 ( .A(n14323), .B(n14147), .ZN(n14320) );
  XOR2_X1 U12368 ( .A(n14174), .B(n14392), .Z(n14389) );
  OAI21_X1 U12369 ( .B1(n14194), .B2(n7629), .A(n11241), .ZN(n11971) );
  NAND4_X1 U12370 ( .A1(n11285), .A2(n7198), .A3(n10593), .A4(n11971), .ZN(
        n10594) );
  NOR2_X1 U12371 ( .A1(n11324), .A2(n10594), .ZN(n10595) );
  XNOR2_X1 U12372 ( .A(n11405), .B(n14190), .ZN(n11028) );
  NAND4_X1 U12373 ( .A1(n15795), .A2(n10595), .A3(n11479), .A4(n11028), .ZN(
        n10596) );
  NOR2_X1 U12374 ( .A1(n11633), .A2(n10596), .ZN(n10598) );
  NAND4_X1 U12375 ( .A1(n11793), .A2(n10598), .A3(n10597), .A4(n11656), .ZN(
        n10599) );
  NOR2_X1 U12376 ( .A1(n11974), .A2(n10599), .ZN(n10600) );
  NAND4_X1 U12377 ( .A1(n12380), .A2(n10600), .A3(n12521), .A4(n12511), .ZN(
        n10601) );
  NOR2_X1 U12378 ( .A1(n12592), .A2(n10601), .ZN(n10602) );
  NAND4_X1 U12379 ( .A1(n14420), .A2(n10602), .A3(n12671), .A4(n12434), .ZN(
        n10603) );
  NOR4_X1 U12380 ( .A1(n14389), .A2(n14370), .A3(n14411), .A4(n10603), .ZN(
        n10606) );
  NAND2_X1 U12381 ( .A1(n10605), .A2(n10604), .ZN(n14346) );
  NAND4_X1 U12382 ( .A1(n10607), .A2(n10606), .A3(n14346), .A4(n14357), .ZN(
        n10608) );
  NOR4_X1 U12383 ( .A1(n14274), .A2(n14320), .A3(n14303), .A4(n10608), .ZN(
        n10610) );
  NAND4_X1 U12384 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n14289), .ZN(
        n10612) );
  NOR2_X1 U12385 ( .A1(n10613), .A2(n10612), .ZN(n10614) );
  XNOR2_X1 U12386 ( .A(n10614), .B(n15339), .ZN(n10615) );
  OR2_X1 U12387 ( .A1(n10756), .A2(P2_U3088), .ZN(n12754) );
  NOR4_X1 U12388 ( .A1(n15247), .A2(n14580), .A3(n7526), .A4(n10620), .ZN(
        n10623) );
  OAI21_X1 U12389 ( .B1(n12754), .B2(n10621), .A(P2_B_REG_SCAN_IN), .ZN(n10622) );
  OR2_X1 U12390 ( .A1(n10623), .A2(n10622), .ZN(n10624) );
  NAND2_X1 U12391 ( .A1(n10625), .A2(n10624), .ZN(P2_U3328) );
  INV_X1 U12392 ( .A(n13072), .ZN(n13459) );
  AND2_X1 U12393 ( .A1(n11044), .A2(P3_B_REG_SCAN_IN), .ZN(n10629) );
  OR2_X1 U12394 ( .A1(n13629), .A2(n10629), .ZN(n13427) );
  OR2_X1 U12395 ( .A1(n10643), .A2(n15892), .ZN(n10642) );
  INV_X1 U12396 ( .A(n10637), .ZN(n13437) );
  INV_X1 U12397 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10638) );
  OR2_X1 U12398 ( .A1(n15894), .A2(n10638), .ZN(n10639) );
  OAI21_X1 U12399 ( .B1(n13437), .B2(n13694), .A(n10639), .ZN(n10640) );
  INV_X1 U12400 ( .A(n10640), .ZN(n10641) );
  NAND2_X1 U12401 ( .A1(n10642), .A2(n10641), .ZN(P3_U3488) );
  OR2_X1 U12402 ( .A1(n10643), .A2(n15895), .ZN(n10647) );
  INV_X1 U12403 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10644) );
  INV_X1 U12404 ( .A(n10645), .ZN(n10646) );
  NAND2_X1 U12405 ( .A1(n10647), .A2(n10646), .ZN(P3_U3456) );
  INV_X1 U12406 ( .A(n10756), .ZN(n10648) );
  INV_X1 U12407 ( .A(n11201), .ZN(n10650) );
  INV_X1 U12408 ( .A(n10940), .ZN(n10651) );
  NAND2_X1 U12409 ( .A1(n14746), .A2(n12999), .ZN(n10655) );
  OAI22_X1 U12410 ( .A1(n7171), .A2(n11617), .B1(n10652), .B2(n10714), .ZN(
        n10653) );
  INV_X1 U12411 ( .A(n10653), .ZN(n10654) );
  NAND2_X1 U12412 ( .A1(n10655), .A2(n10654), .ZN(n10927) );
  NAND2_X1 U12413 ( .A1(n12404), .A2(n15236), .ZN(n10656) );
  AND2_X2 U12414 ( .A1(n10940), .A2(n10656), .ZN(n13009) );
  INV_X1 U12415 ( .A(n14746), .ZN(n10963) );
  OAI22_X1 U12416 ( .A1(n13024), .A2(n11617), .B1(n7345), .B2(n10714), .ZN(
        n10658) );
  INV_X1 U12417 ( .A(n10658), .ZN(n10659) );
  NAND2_X1 U12418 ( .A1(n10660), .A2(n12999), .ZN(n10662) );
  NAND2_X1 U12419 ( .A1(n9710), .A2(n10680), .ZN(n10661) );
  NAND2_X1 U12420 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  XNOR2_X1 U12421 ( .A(n10663), .B(n13009), .ZN(n10668) );
  INV_X1 U12422 ( .A(n10668), .ZN(n10667) );
  NAND2_X1 U12423 ( .A1(n9710), .A2(n12999), .ZN(n10664) );
  AND2_X1 U12424 ( .A1(n10665), .A2(n10664), .ZN(n10669) );
  INV_X1 U12425 ( .A(n10669), .ZN(n10666) );
  NAND2_X1 U12426 ( .A1(n10667), .A2(n10666), .ZN(n10670) );
  NAND2_X1 U12427 ( .A1(n10669), .A2(n10668), .ZN(n10671) );
  NAND2_X1 U12428 ( .A1(n10670), .A2(n10671), .ZN(n10962) );
  INV_X1 U12429 ( .A(n10671), .ZN(n10672) );
  INV_X2 U12430 ( .A(n13009), .ZN(n13025) );
  INV_X2 U12431 ( .A(n13023), .ZN(n13018) );
  NAND2_X1 U12432 ( .A1(n13018), .A2(n14743), .ZN(n10675) );
  NAND2_X1 U12433 ( .A1(n7476), .A2(n12999), .ZN(n10674) );
  NAND2_X1 U12434 ( .A1(n10675), .A2(n10674), .ZN(n10677) );
  XNOR2_X1 U12435 ( .A(n10676), .B(n10677), .ZN(n11000) );
  INV_X1 U12436 ( .A(n10676), .ZN(n10679) );
  INV_X1 U12437 ( .A(n10677), .ZN(n10678) );
  AOI22_X1 U12438 ( .A1(n14624), .A2(n13019), .B1(n13018), .B2(n14742), .ZN(
        n10682) );
  INV_X2 U12439 ( .A(n7171), .ZN(n13014) );
  AOI22_X1 U12440 ( .A1(n14624), .A2(n13014), .B1(n13019), .B2(n14742), .ZN(
        n10681) );
  XNOR2_X1 U12441 ( .A(n10681), .B(n13025), .ZN(n10683) );
  XOR2_X1 U12442 ( .A(n10682), .B(n10683), .Z(n14622) );
  INV_X1 U12443 ( .A(n11531), .ZN(n15746) );
  INV_X1 U12444 ( .A(n14741), .ZN(n11532) );
  OAI22_X1 U12445 ( .A1(n15746), .A2(n13024), .B1(n11532), .B2(n13023), .ZN(
        n10685) );
  AOI22_X1 U12446 ( .A1(n11531), .A2(n13014), .B1(n13019), .B2(n14741), .ZN(
        n10686) );
  XNOR2_X1 U12447 ( .A(n10686), .B(n13025), .ZN(n11576) );
  NOR2_X1 U12448 ( .A1(n11686), .A2(n13024), .ZN(n10687) );
  AOI21_X1 U12449 ( .B1(n11543), .B2(n13014), .A(n10687), .ZN(n10688) );
  XNOR2_X1 U12450 ( .A(n10688), .B(n13025), .ZN(n10690) );
  NOR2_X1 U12451 ( .A1(n11686), .A2(n13023), .ZN(n10689) );
  AOI21_X1 U12452 ( .B1(n11543), .B2(n13019), .A(n10689), .ZN(n10691) );
  INV_X1 U12453 ( .A(n10690), .ZN(n10693) );
  INV_X1 U12454 ( .A(n10691), .ZN(n10692) );
  NAND2_X1 U12455 ( .A1(n10693), .A2(n10692), .ZN(n10736) );
  NAND2_X1 U12456 ( .A1(n7334), .A2(n10736), .ZN(n10694) );
  XNOR2_X1 U12457 ( .A(n10737), .B(n10694), .ZN(n10718) );
  INV_X1 U12458 ( .A(n15228), .ZN(n10695) );
  AND2_X1 U12459 ( .A1(n10696), .A2(n10695), .ZN(n10698) );
  NAND3_X1 U12460 ( .A1(n12906), .A2(P1_B_REG_SCAN_IN), .A3(n15231), .ZN(
        n10697) );
  INV_X1 U12461 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10699) );
  AND2_X1 U12462 ( .A1(n12906), .A2(n15228), .ZN(n10854) );
  AOI21_X1 U12463 ( .B1(n10700), .B2(n10699), .A(n10854), .ZN(n10948) );
  NOR2_X1 U12464 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n10704) );
  NOR4_X1 U12465 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10703) );
  NOR4_X1 U12466 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10702) );
  NOR4_X1 U12467 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10701) );
  NAND4_X1 U12468 ( .A1(n10704), .A2(n10703), .A3(n10702), .A4(n10701), .ZN(
        n10710) );
  NOR4_X1 U12469 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10708) );
  NOR4_X1 U12470 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10707) );
  NOR4_X1 U12471 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10706) );
  NOR4_X1 U12472 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10705) );
  NAND4_X1 U12473 ( .A1(n10708), .A2(n10707), .A3(n10706), .A4(n10705), .ZN(
        n10709) );
  NOR2_X1 U12474 ( .A1(n10710), .A2(n10709), .ZN(n10711) );
  OR2_X1 U12475 ( .A1(n10843), .A2(n10711), .ZN(n10946) );
  AND2_X1 U12476 ( .A1(n10948), .A2(n10946), .ZN(n11495) );
  OR2_X1 U12477 ( .A1(n10843), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10712) );
  NAND2_X1 U12478 ( .A1(n15231), .A2(n15228), .ZN(n10844) );
  NAND2_X1 U12479 ( .A1(n11495), .A2(n11493), .ZN(n10724) );
  INV_X1 U12480 ( .A(n10715), .ZN(n10716) );
  NAND3_X1 U12481 ( .A1(n11497), .A2(n10725), .A3(n15990), .ZN(n10717) );
  NOR2_X1 U12482 ( .A1(n10718), .A2(n16022), .ZN(n10730) );
  NAND2_X1 U12483 ( .A1(n15912), .A2(n12729), .ZN(n11496) );
  NAND2_X1 U12484 ( .A1(n10724), .A2(n11496), .ZN(n10721) );
  AND2_X1 U12485 ( .A1(n10721), .A2(n11497), .ZN(n10929) );
  AND2_X1 U12486 ( .A1(n11543), .A2(n15949), .ZN(n15776) );
  AND2_X1 U12487 ( .A1(n10929), .A2(n15776), .ZN(n10729) );
  NAND2_X1 U12488 ( .A1(n10721), .A2(n10720), .ZN(n10722) );
  NOR2_X1 U12489 ( .A1(n16031), .A2(n11544), .ZN(n10728) );
  INV_X1 U12490 ( .A(n11494), .ZN(n10723) );
  NAND2_X1 U12491 ( .A1(n16011), .A2(n15075), .ZN(n16016) );
  INV_X1 U12492 ( .A(n15042), .ZN(n15076) );
  AND2_X1 U12493 ( .A1(n16011), .A2(n15076), .ZN(n15978) );
  NAND2_X1 U12494 ( .A1(n15978), .A2(n11704), .ZN(n10726) );
  NAND2_X1 U12495 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10912) );
  OAI211_X1 U12496 ( .C1(n11532), .C2(n16016), .A(n10726), .B(n10912), .ZN(
        n10727) );
  OR4_X1 U12497 ( .A1(n10730), .A2(n10729), .A3(n10728), .A4(n10727), .ZN(
        P1_U3227) );
  NAND2_X1 U12498 ( .A1(n11694), .A2(n13014), .ZN(n10732) );
  OR2_X1 U12499 ( .A1(n11709), .A2(n13024), .ZN(n10731) );
  NAND2_X1 U12500 ( .A1(n10732), .A2(n10731), .ZN(n10733) );
  XNOR2_X1 U12501 ( .A(n10733), .B(n13025), .ZN(n10791) );
  NAND2_X1 U12502 ( .A1(n11694), .A2(n13019), .ZN(n10735) );
  OR2_X1 U12503 ( .A1(n11709), .A2(n13023), .ZN(n10734) );
  NAND2_X1 U12504 ( .A1(n10735), .A2(n10734), .ZN(n10738) );
  INV_X1 U12505 ( .A(n10738), .ZN(n10790) );
  AND2_X1 U12506 ( .A1(n13018), .A2(n14739), .ZN(n10740) );
  AOI21_X1 U12507 ( .B1(n11858), .B2(n13019), .A(n10740), .ZN(n12189) );
  AOI22_X1 U12508 ( .A1(n11858), .A2(n13014), .B1(n13019), .B2(n14739), .ZN(
        n10741) );
  XNOR2_X1 U12509 ( .A(n10741), .B(n13025), .ZN(n12190) );
  XOR2_X1 U12510 ( .A(n12189), .B(n12190), .Z(n12193) );
  XNOR2_X1 U12511 ( .A(n12194), .B(n12193), .ZN(n10742) );
  NOR2_X1 U12512 ( .A1(n10742), .A2(n16022), .ZN(n10747) );
  AND2_X1 U12513 ( .A1(n16027), .A2(n11858), .ZN(n10746) );
  NOR2_X1 U12514 ( .A1(n16031), .A2(n11713), .ZN(n10745) );
  NAND2_X1 U12515 ( .A1(n15978), .A2(n14738), .ZN(n10743) );
  NAND2_X1 U12516 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14782) );
  OAI211_X1 U12517 ( .C1(n11709), .C2(n16016), .A(n10743), .B(n14782), .ZN(
        n10744) );
  OR4_X1 U12518 ( .A1(n10747), .A2(n10746), .A3(n10745), .A4(n10744), .ZN(
        P1_U3213) );
  NAND2_X1 U12519 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n11352) );
  INV_X1 U12520 ( .A(n11352), .ZN(n10776) );
  INV_X1 U12521 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10748) );
  MUX2_X1 U12522 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10748), .S(n10780), .Z(
        n10761) );
  INV_X1 U12523 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n15720) );
  MUX2_X1 U12524 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n15720), .S(n14199), .Z(
        n14202) );
  INV_X1 U12525 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10749) );
  MUX2_X1 U12526 ( .A(n10749), .B(P2_REG2_REG_1__SCAN_IN), .S(n10802), .Z(
        n15261) );
  NAND2_X1 U12527 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15265) );
  INV_X1 U12528 ( .A(n15265), .ZN(n10750) );
  NAND2_X1 U12529 ( .A1(n15261), .A2(n10750), .ZN(n15262) );
  NAND2_X1 U12530 ( .A1(n15257), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10751) );
  NAND2_X1 U12531 ( .A1(n15262), .A2(n10751), .ZN(n14201) );
  NAND2_X1 U12532 ( .A1(n14202), .A2(n14201), .ZN(n14200) );
  NAND2_X1 U12533 ( .A1(n14199), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10752) );
  NAND2_X1 U12534 ( .A1(n14200), .A2(n10752), .ZN(n14216) );
  INV_X1 U12535 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10753) );
  MUX2_X1 U12536 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10753), .S(n14210), .Z(
        n14217) );
  NAND2_X1 U12537 ( .A1(n14216), .A2(n14217), .ZN(n14215) );
  NAND2_X1 U12538 ( .A1(n14210), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10754) );
  NAND2_X1 U12539 ( .A1(n14215), .A2(n10754), .ZN(n10760) );
  AOI21_X1 U12540 ( .B1(n11106), .B2(n10756), .A(n10755), .ZN(n10757) );
  OR2_X1 U12541 ( .A1(n10758), .A2(n10757), .ZN(n10772) );
  NOR2_X1 U12542 ( .A1(n7526), .A2(P2_U3088), .ZN(n14575) );
  INV_X1 U12543 ( .A(n14580), .ZN(n10759) );
  NAND2_X1 U12544 ( .A1(n10760), .A2(n10761), .ZN(n10782) );
  OAI211_X1 U12545 ( .C1(n10761), .C2(n10760), .A(n15333), .B(n10782), .ZN(
        n10762) );
  INV_X1 U12546 ( .A(n10762), .ZN(n10775) );
  INV_X1 U12547 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10763) );
  MUX2_X1 U12548 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10763), .S(n10802), .Z(
        n15259) );
  NAND2_X1 U12549 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15260) );
  NOR2_X1 U12550 ( .A1(n15259), .A2(n15260), .ZN(n15258) );
  AOI21_X1 U12551 ( .B1(n15257), .B2(P2_REG1_REG_1__SCAN_IN), .A(n15258), .ZN(
        n14197) );
  INV_X1 U12552 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10764) );
  MUX2_X1 U12553 ( .A(n10764), .B(P2_REG1_REG_2__SCAN_IN), .S(n14199), .Z(
        n14196) );
  INV_X1 U12554 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10765) );
  MUX2_X1 U12555 ( .A(n10765), .B(P2_REG1_REG_3__SCAN_IN), .S(n14210), .Z(
        n14212) );
  INV_X1 U12556 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10766) );
  MUX2_X1 U12557 ( .A(n10766), .B(P2_REG1_REG_4__SCAN_IN), .S(n10780), .Z(
        n10768) );
  AOI211_X1 U12558 ( .C1(n10769), .C2(n10768), .A(n10777), .B(n15368), .ZN(
        n10774) );
  INV_X1 U12559 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15465) );
  AND2_X1 U12560 ( .A1(n7526), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10771) );
  INV_X1 U12561 ( .A(n15374), .ZN(n15322) );
  INV_X1 U12562 ( .A(n10780), .ZN(n10824) );
  OAI22_X1 U12563 ( .A1(n15377), .A2(n15465), .B1(n15322), .B2(n10824), .ZN(
        n10773) );
  OR4_X1 U12564 ( .A1(n10776), .A2(n10775), .A3(n10774), .A4(n10773), .ZN(
        P2_U3218) );
  AND2_X1 U12565 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10789) );
  AOI21_X1 U12566 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n10780), .A(n10777), .ZN(
        n10779) );
  XNOR2_X1 U12567 ( .A(n11263), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n10778) );
  NOR2_X1 U12568 ( .A1(n10779), .A2(n10778), .ZN(n11262) );
  AOI211_X1 U12569 ( .C1(n10779), .C2(n10778), .A(n15368), .B(n11262), .ZN(
        n10788) );
  INV_X1 U12570 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11601) );
  XNOR2_X1 U12571 ( .A(n11263), .B(n11601), .ZN(n10784) );
  NAND2_X1 U12572 ( .A1(n10780), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U12573 ( .A1(n10782), .A2(n10781), .ZN(n10783) );
  NAND2_X1 U12574 ( .A1(n10783), .A2(n10784), .ZN(n11253) );
  OAI211_X1 U12575 ( .C1(n10784), .C2(n10783), .A(n15333), .B(n11253), .ZN(
        n10785) );
  INV_X1 U12576 ( .A(n10785), .ZN(n10787) );
  INV_X1 U12577 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15469) );
  INV_X1 U12578 ( .A(n11263), .ZN(n10822) );
  OAI22_X1 U12579 ( .A1(n15377), .A2(n15469), .B1(n15322), .B2(n10822), .ZN(
        n10786) );
  OR4_X1 U12580 ( .A1(n10789), .A2(n10788), .A3(n10787), .A4(n10786), .ZN(
        P2_U3219) );
  XNOR2_X1 U12581 ( .A(n10791), .B(n10790), .ZN(n10792) );
  XNOR2_X1 U12582 ( .A(n10793), .B(n10792), .ZN(n10794) );
  NOR2_X1 U12583 ( .A1(n10794), .A2(n16022), .ZN(n10800) );
  INV_X1 U12584 ( .A(n10929), .ZN(n10795) );
  NAND2_X1 U12585 ( .A1(n11694), .A2(n15949), .ZN(n15788) );
  NOR2_X1 U12586 ( .A1(n10795), .A2(n15788), .ZN(n10799) );
  NOR2_X1 U12587 ( .A1(n16031), .A2(n11690), .ZN(n10798) );
  NAND2_X1 U12588 ( .A1(n15978), .A2(n14739), .ZN(n10796) );
  NAND2_X1 U12589 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14770) );
  OAI211_X1 U12590 ( .C1(n11686), .C2(n16016), .A(n10796), .B(n14770), .ZN(
        n10797) );
  OR4_X1 U12591 ( .A1(n10800), .A2(n10799), .A3(n10798), .A4(n10797), .ZN(
        P1_U3239) );
  NOR2_X1 U12592 ( .A1(n10801), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14576) );
  INV_X2 U12593 ( .A(n14576), .ZN(n14592) );
  OAI222_X1 U12594 ( .A1(n14578), .A2(n10807), .B1(n14592), .B2(n10803), .C1(
        P2_U3088), .C2(n10802), .ZN(P2_U3326) );
  INV_X1 U12595 ( .A(n10804), .ZN(n10834) );
  OAI222_X1 U12596 ( .A1(n14592), .A2(n10805), .B1(n14578), .B2(n10834), .C1(
        n7464), .C2(P2_U3088), .ZN(P2_U3325) );
  NAND2_X1 U12597 ( .A1(n8863), .A2(P1_U3086), .ZN(n15235) );
  AND2_X1 U12598 ( .A1(n10806), .A2(P1_U3086), .ZN(n12757) );
  INV_X2 U12599 ( .A(n12757), .ZN(n15233) );
  OAI222_X1 U12600 ( .A1(n15235), .A2(n8846), .B1(n15233), .B2(n10807), .C1(
        P1_U3086), .C2(n10879), .ZN(P1_U3354) );
  INV_X1 U12601 ( .A(n10808), .ZN(n10830) );
  INV_X1 U12602 ( .A(n14210), .ZN(n10809) );
  OAI222_X1 U12603 ( .A1(n14592), .A2(n10810), .B1(n14578), .B2(n10830), .C1(
        n10809), .C2(P2_U3088), .ZN(P2_U3324) );
  NAND2_X1 U12604 ( .A1(n8863), .A2(P3_U3151), .ZN(n13787) );
  INV_X1 U12605 ( .A(SI_8_), .ZN(n10812) );
  NOR2_X1 U12606 ( .A1(n10801), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13779) );
  INV_X2 U12607 ( .A(n13779), .ZN(n13993) );
  OAI222_X1 U12608 ( .A1(P3_U3151), .A2(n12174), .B1(n13787), .B2(n10812), 
        .C1(n13993), .C2(n10811), .ZN(P3_U3287) );
  OAI222_X1 U12609 ( .A1(P3_U3151), .A2(n7498), .B1(n13787), .B2(n7509), .C1(
        n13993), .C2(n10813), .ZN(P3_U3293) );
  INV_X1 U12610 ( .A(SI_3_), .ZN(n13925) );
  OAI222_X1 U12611 ( .A1(P3_U3151), .A2(n11173), .B1(n13993), .B2(n10814), 
        .C1(n13787), .C2(n13925), .ZN(P3_U3292) );
  INV_X1 U12612 ( .A(SI_5_), .ZN(n13836) );
  OAI222_X1 U12613 ( .A1(P3_U3151), .A2(n11759), .B1(n13993), .B2(n10815), 
        .C1(n13787), .C2(n13836), .ZN(P3_U3290) );
  INV_X1 U12614 ( .A(n13236), .ZN(n11769) );
  INV_X1 U12615 ( .A(n10816), .ZN(n10817) );
  OAI222_X1 U12616 ( .A1(P3_U3151), .A2(n11769), .B1(n13993), .B2(n10817), 
        .C1(n13923), .C2(n13787), .ZN(P3_U3289) );
  INV_X1 U12617 ( .A(n10818), .ZN(n10820) );
  OAI222_X1 U12618 ( .A1(P3_U3151), .A2(n7493), .B1(n13993), .B2(n10820), .C1(
        n10819), .C2(n13787), .ZN(P3_U3294) );
  OAI222_X1 U12619 ( .A1(P2_U3088), .A2(n10822), .B1(n14578), .B2(n10832), 
        .C1(n10821), .C2(n14592), .ZN(P2_U3322) );
  INV_X1 U12620 ( .A(n10823), .ZN(n10826) );
  OAI222_X1 U12621 ( .A1(n14592), .A2(n10825), .B1(n14578), .B2(n10826), .C1(
        P2_U3088), .C2(n10824), .ZN(P2_U3323) );
  INV_X1 U12622 ( .A(n10885), .ZN(n11016) );
  OAI222_X1 U12623 ( .A1(n15235), .A2(n10827), .B1(n15233), .B2(n10826), .C1(
        n11016), .C2(P1_U3086), .ZN(P1_U3351) );
  OAI222_X1 U12624 ( .A1(n12687), .A2(P3_U3151), .B1(n13993), .B2(n10828), 
        .C1(n13787), .C2(n13912), .ZN(P3_U3284) );
  INV_X1 U12625 ( .A(n14760), .ZN(n10883) );
  INV_X1 U12626 ( .A(n15235), .ZN(n15212) );
  OAI222_X1 U12627 ( .A1(P1_U3086), .A2(n10883), .B1(n15233), .B2(n10830), 
        .C1(n10829), .C2(n15224), .ZN(P1_U3352) );
  INV_X1 U12628 ( .A(n10914), .ZN(n10886) );
  OAI222_X1 U12629 ( .A1(P1_U3086), .A2(n10886), .B1(n15233), .B2(n10832), 
        .C1(n10831), .C2(n15224), .ZN(P1_U3350) );
  INV_X1 U12630 ( .A(n10993), .ZN(n10881) );
  OAI222_X1 U12631 ( .A1(P1_U3086), .A2(n10881), .B1(n15233), .B2(n10834), 
        .C1(n10833), .C2(n15224), .ZN(P1_U3353) );
  INV_X1 U12632 ( .A(n14772), .ZN(n10888) );
  INV_X1 U12633 ( .A(n10835), .ZN(n10837) );
  OAI222_X1 U12634 ( .A1(P1_U3086), .A2(n10888), .B1(n15233), .B2(n10837), 
        .C1(n7462), .C2(n15224), .ZN(P1_U3349) );
  INV_X1 U12635 ( .A(n15270), .ZN(n10836) );
  OAI222_X1 U12636 ( .A1(n14592), .A2(n10953), .B1(n14578), .B2(n10837), .C1(
        n10836), .C2(P2_U3088), .ZN(P2_U3321) );
  INV_X1 U12637 ( .A(n13787), .ZN(n12117) );
  OAI222_X1 U12638 ( .A1(P3_U3151), .A2(n12335), .B1(n13995), .B2(n13915), 
        .C1(n13993), .C2(n10838), .ZN(P3_U3285) );
  OAI222_X1 U12639 ( .A1(P3_U3151), .A2(n11185), .B1(n13995), .B2(n10840), 
        .C1(n13993), .C2(n10839), .ZN(P3_U3291) );
  OAI222_X1 U12640 ( .A1(P3_U3151), .A2(n15642), .B1(n13995), .B2(n13827), 
        .C1(n13993), .C2(n10841), .ZN(P3_U3286) );
  OAI222_X1 U12641 ( .A1(n13993), .A2(n10842), .B1(n13995), .B2(n8324), .C1(
        n11757), .C2(P3_U3151), .ZN(P3_U3288) );
  NAND2_X2 U12642 ( .A1(n10843), .A2(n11497), .ZN(n15240) );
  INV_X1 U12643 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10847) );
  INV_X1 U12644 ( .A(n10844), .ZN(n10845) );
  AOI22_X1 U12645 ( .A1(n15240), .A2(n10847), .B1(n10846), .B2(n10845), .ZN(
        P1_U3445) );
  INV_X1 U12646 ( .A(n10848), .ZN(n10852) );
  INV_X1 U12647 ( .A(n14226), .ZN(n10849) );
  OAI222_X1 U12648 ( .A1(n14592), .A2(n10850), .B1(n14578), .B2(n10852), .C1(
        n10849), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U12649 ( .A(n14784), .ZN(n10889) );
  OAI222_X1 U12650 ( .A1(P1_U3086), .A2(n10889), .B1(n15233), .B2(n10852), 
        .C1(n10851), .C2(n15224), .ZN(P1_U3348) );
  NAND2_X1 U12651 ( .A1(n15240), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10853) );
  OAI21_X1 U12652 ( .B1(n15240), .B2(n10854), .A(n10853), .ZN(P1_U3446) );
  OAI222_X1 U12653 ( .A1(n14592), .A2(n10855), .B1(n14578), .B2(n10857), .C1(
        n14238), .C2(P2_U3088), .ZN(P2_U3319) );
  INV_X1 U12654 ( .A(n10890), .ZN(n10903) );
  INV_X1 U12655 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10856) );
  OAI222_X1 U12656 ( .A1(P1_U3086), .A2(n10903), .B1(n15233), .B2(n10857), 
        .C1(n10856), .C2(n15224), .ZN(P1_U3347) );
  INV_X1 U12657 ( .A(n10858), .ZN(n10859) );
  OAI222_X1 U12658 ( .A1(n13787), .A2(n13914), .B1(n13993), .B2(n10859), .C1(
        n13252), .C2(P3_U3151), .ZN(P3_U3283) );
  AND2_X1 U12659 ( .A1(n10861), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12660 ( .A1(n10861), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12661 ( .A1(n10861), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12662 ( .A1(n10861), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12663 ( .A1(n10861), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12664 ( .A1(n10861), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12665 ( .A1(n10861), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12666 ( .A1(n10861), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12667 ( .A1(n10861), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12668 ( .A1(n10861), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12669 ( .A1(n10861), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12670 ( .A1(n10861), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12671 ( .A1(n10861), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12672 ( .A1(n10861), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12673 ( .A1(n10861), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12674 ( .A1(n10861), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12675 ( .A1(n10861), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12676 ( .A1(n10861), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12677 ( .A1(n10861), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12678 ( .A1(n10861), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12679 ( .A1(n10861), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12680 ( .A1(n10861), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12681 ( .A1(n10861), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12682 ( .A1(n10861), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12683 ( .A1(n10861), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12684 ( .A1(n10861), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12685 ( .A1(n10861), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12686 ( .A1(n10861), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12687 ( .A1(n10861), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12688 ( .A1(n10861), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  MUX2_X1 U12689 ( .A(n10898), .B(P1_REG1_REG_8__SCAN_IN), .S(n10890), .Z(
        n10870) );
  INV_X1 U12690 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10867) );
  INV_X1 U12691 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10865) );
  INV_X1 U12692 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10864) );
  INV_X1 U12693 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10863) );
  INV_X1 U12694 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15676) );
  MUX2_X1 U12695 ( .A(n15676), .B(P1_REG1_REG_1__SCAN_IN), .S(n10879), .Z(
        n14752) );
  AND2_X1 U12696 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n14751) );
  NAND2_X1 U12697 ( .A1(n14752), .A2(n14751), .ZN(n14750) );
  INV_X1 U12698 ( .A(n10879), .ZN(n14753) );
  NAND2_X1 U12699 ( .A1(n14753), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U12700 ( .A1(n14750), .A2(n10862), .ZN(n10988) );
  XNOR2_X1 U12701 ( .A(n10883), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n14763) );
  NAND2_X1 U12702 ( .A1(n14762), .A2(n14763), .ZN(n14761) );
  OAI21_X1 U12703 ( .B1(n10864), .B2(n10883), .A(n14761), .ZN(n11008) );
  XNOR2_X1 U12704 ( .A(n11016), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U12705 ( .A1(n11008), .A2(n11009), .ZN(n11007) );
  OAI21_X1 U12706 ( .B1(n10865), .B2(n11016), .A(n11007), .ZN(n10910) );
  MUX2_X1 U12707 ( .A(n10866), .B(P1_REG1_REG_5__SCAN_IN), .S(n10914), .Z(
        n10911) );
  NOR2_X1 U12708 ( .A1(n10910), .A2(n10911), .ZN(n10909) );
  AOI21_X1 U12709 ( .B1(n10886), .B2(n10866), .A(n10909), .ZN(n14777) );
  XNOR2_X1 U12710 ( .A(n10888), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n14778) );
  NAND2_X1 U12711 ( .A1(n14777), .A2(n14778), .ZN(n14776) );
  OAI21_X1 U12712 ( .B1(n10867), .B2(n10888), .A(n14776), .ZN(n14790) );
  XNOR2_X1 U12713 ( .A(n10889), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n14789) );
  AOI21_X1 U12714 ( .B1(n10870), .B2(n10869), .A(n10897), .ZN(n10896) );
  INV_X1 U12715 ( .A(n11497), .ZN(n10871) );
  NAND2_X1 U12716 ( .A1(n10871), .A2(n12759), .ZN(n10877) );
  AOI21_X1 U12717 ( .B1(n10874), .B2(n10873), .A(n7207), .ZN(n10875) );
  NAND2_X1 U12718 ( .A1(n10877), .A2(n10875), .ZN(n15383) );
  INV_X1 U12719 ( .A(n10875), .ZN(n10876) );
  AND2_X1 U12720 ( .A1(n10877), .A2(n10876), .ZN(n15381) );
  INV_X1 U12721 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15498) );
  NAND2_X1 U12722 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n12207) );
  OAI21_X1 U12723 ( .B1(n15430), .B2(n15498), .A(n12207), .ZN(n10878) );
  AOI21_X1 U12724 ( .B1(n10890), .B2(n15423), .A(n10878), .ZN(n10895) );
  MUX2_X1 U12725 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10882), .S(n10993), .Z(
        n10992) );
  MUX2_X1 U12726 ( .A(n10880), .B(P1_REG2_REG_1__SCAN_IN), .S(n10879), .Z(
        n14749) );
  AND2_X1 U12727 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14748) );
  NAND2_X1 U12728 ( .A1(n14749), .A2(n14748), .ZN(n14747) );
  OAI21_X1 U12729 ( .B1(n10880), .B2(n10879), .A(n14747), .ZN(n10991) );
  NAND2_X1 U12730 ( .A1(n10992), .A2(n10991), .ZN(n10990) );
  OAI21_X1 U12731 ( .B1(n10882), .B2(n10881), .A(n10990), .ZN(n14765) );
  XOR2_X1 U12732 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14760), .Z(n14766) );
  NAND2_X1 U12733 ( .A1(n14765), .A2(n14766), .ZN(n14764) );
  OAI21_X1 U12734 ( .B1(n10884), .B2(n10883), .A(n14764), .ZN(n11013) );
  XOR2_X1 U12735 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10885), .Z(n11014) );
  NAND2_X1 U12736 ( .A1(n11013), .A2(n11014), .ZN(n11012) );
  OAI21_X1 U12737 ( .B1(n11517), .B2(n11016), .A(n11012), .ZN(n10916) );
  MUX2_X1 U12738 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10887), .S(n10914), .Z(
        n10917) );
  NAND2_X1 U12739 ( .A1(n10916), .A2(n10917), .ZN(n10915) );
  OAI21_X1 U12740 ( .B1(n10887), .B2(n10886), .A(n10915), .ZN(n14774) );
  XOR2_X1 U12741 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n14772), .Z(n14775) );
  NAND2_X1 U12742 ( .A1(n14774), .A2(n14775), .ZN(n14773) );
  OAI21_X1 U12743 ( .B1(n11691), .B2(n10888), .A(n14773), .ZN(n14786) );
  XOR2_X1 U12744 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n14784), .Z(n14787) );
  NAND2_X1 U12745 ( .A1(n14786), .A2(n14787), .ZN(n14785) );
  OAI21_X1 U12746 ( .B1(n11714), .B2(n10889), .A(n14785), .ZN(n10893) );
  MUX2_X1 U12747 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11869), .S(n10890), .Z(
        n10892) );
  NAND2_X1 U12748 ( .A1(n10893), .A2(n10892), .ZN(n10902) );
  OR2_X1 U12749 ( .A1(n15223), .A2(n15227), .ZN(n10891) );
  INV_X1 U12750 ( .A(n15413), .ZN(n15426) );
  OAI211_X1 U12751 ( .C1(n10893), .C2(n10892), .A(n10902), .B(n15426), .ZN(
        n10894) );
  OAI211_X1 U12752 ( .C1(n10896), .C2(n15397), .A(n10895), .B(n10894), .ZN(
        P1_U3251) );
  MUX2_X1 U12753 ( .A(n10969), .B(P1_REG1_REG_9__SCAN_IN), .S(n10922), .Z(
        n10900) );
  NOR2_X1 U12754 ( .A1(n10899), .A2(n10900), .ZN(n10968) );
  AOI21_X1 U12755 ( .B1(n10900), .B2(n10899), .A(n10968), .ZN(n10908) );
  NAND2_X1 U12756 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n12268) );
  OAI21_X1 U12757 ( .B1(n15430), .B2(n15510), .A(n12268), .ZN(n10901) );
  AOI21_X1 U12758 ( .B1(n10922), .B2(n15423), .A(n10901), .ZN(n10907) );
  OAI21_X1 U12759 ( .B1(n11869), .B2(n10903), .A(n10902), .ZN(n10905) );
  XOR2_X1 U12760 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10922), .Z(n10904) );
  NAND2_X1 U12761 ( .A1(n10905), .A2(n10904), .ZN(n10974) );
  OAI211_X1 U12762 ( .C1(n10905), .C2(n10904), .A(n10974), .B(n15426), .ZN(
        n10906) );
  OAI211_X1 U12763 ( .C1(n10908), .C2(n15397), .A(n10907), .B(n10906), .ZN(
        P1_U3252) );
  AOI21_X1 U12764 ( .B1(n10911), .B2(n10910), .A(n10909), .ZN(n10920) );
  INV_X1 U12765 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15475) );
  OAI21_X1 U12766 ( .B1(n15430), .B2(n15475), .A(n10912), .ZN(n10913) );
  AOI21_X1 U12767 ( .B1(n10914), .B2(n15423), .A(n10913), .ZN(n10919) );
  OAI211_X1 U12768 ( .C1(n10917), .C2(n10916), .A(n15426), .B(n10915), .ZN(
        n10918) );
  OAI211_X1 U12769 ( .C1(n10920), .C2(n15397), .A(n10919), .B(n10918), .ZN(
        P1_U3248) );
  OAI222_X1 U12770 ( .A1(P3_U3151), .A2(n13294), .B1(n13995), .B2(n13880), 
        .C1(n13993), .C2(n10921), .ZN(P3_U3282) );
  INV_X1 U12771 ( .A(n10922), .ZN(n10975) );
  OAI222_X1 U12772 ( .A1(n15235), .A2(n10923), .B1(n15233), .B2(n10925), .C1(
        P1_U3086), .C2(n10975), .ZN(P1_U3346) );
  INV_X1 U12773 ( .A(n11924), .ZN(n11913) );
  OAI222_X1 U12774 ( .A1(P2_U3088), .A2(n11913), .B1(n14578), .B2(n10925), 
        .C1(n10924), .C2(n14592), .ZN(P2_U3318) );
  XNOR2_X1 U12775 ( .A(n10926), .B(n10927), .ZN(n10983) );
  NAND2_X1 U12776 ( .A1(n10929), .A2(n10928), .ZN(n11004) );
  AOI22_X1 U12777 ( .A1(n15978), .A2(n14744), .B1(n11004), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10931) );
  NAND2_X1 U12778 ( .A1(n16027), .A2(n11499), .ZN(n10930) );
  OAI211_X1 U12779 ( .C1(n10983), .C2(n16022), .A(n10931), .B(n10930), .ZN(
        P1_U3232) );
  CLKBUF_X2 U12780 ( .A(P1_U4016), .Z(n14745) );
  NOR2_X1 U12781 ( .A1(n15381), .A2(n14745), .ZN(P1_U3085) );
  OAI222_X1 U12782 ( .A1(n13305), .A2(P3_U3151), .B1(n13993), .B2(n10932), 
        .C1(n13787), .C2(n8092), .ZN(P3_U3281) );
  INV_X1 U12783 ( .A(n10933), .ZN(n10936) );
  INV_X1 U12784 ( .A(n15373), .ZN(n10934) );
  OAI222_X1 U12785 ( .A1(n14592), .A2(n10951), .B1(n14578), .B2(n10936), .C1(
        n10934), .C2(P2_U3088), .ZN(P2_U3317) );
  INV_X1 U12786 ( .A(n14799), .ZN(n10976) );
  OAI222_X1 U12787 ( .A1(P1_U3086), .A2(n10976), .B1(n15233), .B2(n10936), 
        .C1(n10935), .C2(n15224), .ZN(P1_U3345) );
  INV_X1 U12788 ( .A(n10937), .ZN(n10958) );
  AOI22_X1 U12789 ( .A1(n12026), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n14576), .ZN(n10938) );
  OAI21_X1 U12790 ( .B1(n10958), .B2(n14578), .A(n10938), .ZN(P2_U3316) );
  INV_X1 U12791 ( .A(n10945), .ZN(n15663) );
  NOR2_X1 U12792 ( .A1(n11617), .A2(n11511), .ZN(n15657) );
  NOR2_X1 U12793 ( .A1(n10940), .A2(n10939), .ZN(n10941) );
  INV_X1 U12794 ( .A(n15671), .ZN(n15025) );
  NOR2_X1 U12795 ( .A1(n15025), .A2(n15993), .ZN(n10944) );
  OAI22_X1 U12796 ( .A1(n10945), .A2(n10944), .B1(n9711), .B2(n15042), .ZN(
        n15661) );
  AOI211_X1 U12797 ( .C1(n15912), .C2(n15663), .A(n15657), .B(n15661), .ZN(
        n15655) );
  NAND2_X1 U12798 ( .A1(n10946), .A2(n11496), .ZN(n10947) );
  NOR2_X1 U12799 ( .A1(n10948), .A2(n10947), .ZN(n10949) );
  AND2_X1 U12800 ( .A1(n10949), .A2(n11494), .ZN(n11880) );
  INV_X1 U12801 ( .A(n16001), .ZN(n15999) );
  NAND2_X1 U12802 ( .A1(n15999), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10950) );
  OAI21_X1 U12803 ( .B1(n15655), .B2(n15999), .A(n10950), .ZN(P1_U3528) );
  MUX2_X1 U12804 ( .A(n10951), .B(n12362), .S(n14745), .Z(n10952) );
  INV_X1 U12805 ( .A(n10952), .ZN(P1_U3570) );
  MUX2_X1 U12806 ( .A(n10953), .B(n11709), .S(n14745), .Z(n10954) );
  INV_X1 U12807 ( .A(n10954), .ZN(P1_U3566) );
  INV_X1 U12808 ( .A(n10955), .ZN(n10957) );
  OAI22_X1 U12809 ( .A1(n13346), .A2(P3_U3151), .B1(SI_15_), .B2(n13995), .ZN(
        n10956) );
  AOI21_X1 U12810 ( .B1(n10957), .B2(n13779), .A(n10956), .ZN(P3_U3280) );
  INV_X1 U12811 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10959) );
  INV_X1 U12812 ( .A(n10977), .ZN(n11457) );
  OAI222_X1 U12813 ( .A1(n15235), .A2(n10959), .B1(n15233), .B2(n10958), .C1(
        P1_U3086), .C2(n11457), .ZN(P1_U3344) );
  AOI21_X1 U12814 ( .B1(n10962), .B2(n10961), .A(n10960), .ZN(n10967) );
  INV_X1 U12815 ( .A(n15978), .ZN(n16019) );
  OAI22_X1 U12816 ( .A1(n16019), .A2(n7516), .B1(n10963), .B2(n16016), .ZN(
        n10965) );
  INV_X1 U12817 ( .A(n16027), .ZN(n15982) );
  NOR2_X1 U12818 ( .A1(n15982), .A2(n15670), .ZN(n10964) );
  AOI211_X1 U12819 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n11004), .A(n10965), .B(
        n10964), .ZN(n10966) );
  OAI21_X1 U12820 ( .B1(n10967), .B2(n16022), .A(n10966), .ZN(P1_U3222) );
  MUX2_X1 U12821 ( .A(n11456), .B(P1_REG1_REG_11__SCAN_IN), .S(n10977), .Z(
        n10972) );
  AOI21_X1 U12822 ( .B1(n10969), .B2(n10975), .A(n10968), .ZN(n14796) );
  MUX2_X1 U12823 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10970), .S(n14799), .Z(
        n14795) );
  NAND2_X1 U12824 ( .A1(n14796), .A2(n14795), .ZN(n14794) );
  OAI21_X1 U12825 ( .B1(n10976), .B2(n10970), .A(n14794), .ZN(n10971) );
  AOI21_X1 U12826 ( .B1(n10972), .B2(n10971), .A(n11455), .ZN(n10982) );
  INV_X1 U12827 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15528) );
  NAND2_X1 U12828 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n12562)
         );
  OAI21_X1 U12829 ( .B1(n15430), .B2(n15528), .A(n12562), .ZN(n10973) );
  AOI21_X1 U12830 ( .B1(n15423), .B2(n10977), .A(n10973), .ZN(n10981) );
  OAI21_X1 U12831 ( .B1(n10975), .B2(n12012), .A(n10974), .ZN(n14802) );
  MUX2_X1 U12832 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n12091), .S(n14799), .Z(
        n14801) );
  NAND2_X1 U12833 ( .A1(n14802), .A2(n14801), .ZN(n14800) );
  OAI21_X1 U12834 ( .B1(n10976), .B2(n12091), .A(n14800), .ZN(n10979) );
  XOR2_X1 U12835 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10977), .Z(n10978) );
  NAND2_X1 U12836 ( .A1(n10979), .A2(n10978), .ZN(n11450) );
  OAI211_X1 U12837 ( .C1(n10979), .C2(n10978), .A(n11450), .B(n15426), .ZN(
        n10980) );
  OAI211_X1 U12838 ( .C1(n10982), .C2(n15397), .A(n10981), .B(n10980), .ZN(
        P1_U3254) );
  MUX2_X1 U12839 ( .A(n14748), .B(n10983), .S(n15227), .Z(n10986) );
  INV_X1 U12840 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n15666) );
  AOI21_X1 U12841 ( .B1(n15379), .B2(n15666), .A(n15223), .ZN(n15378) );
  OAI21_X1 U12842 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n15378), .A(n14745), .ZN(
        n10984) );
  AOI21_X1 U12843 ( .B1(n10986), .B2(n10985), .A(n10984), .ZN(n11019) );
  INV_X1 U12844 ( .A(n15397), .ZN(n15427) );
  OAI211_X1 U12845 ( .C1(n10989), .C2(n10988), .A(n15427), .B(n10987), .ZN(
        n10997) );
  OAI211_X1 U12846 ( .C1(n10992), .C2(n10991), .A(n15426), .B(n10990), .ZN(
        n10996) );
  AOI22_X1 U12847 ( .A1(n15381), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10995) );
  NAND2_X1 U12848 ( .A1(n15423), .A2(n10993), .ZN(n10994) );
  NAND4_X1 U12849 ( .A1(n10997), .A2(n10996), .A3(n10995), .A4(n10994), .ZN(
        n10998) );
  OR2_X1 U12850 ( .A1(n11019), .A2(n10998), .ZN(P1_U3245) );
  AOI21_X1 U12851 ( .B1(n10999), .B2(n11000), .A(n11001), .ZN(n11006) );
  INV_X1 U12852 ( .A(n14742), .ZN(n11505) );
  OAI22_X1 U12853 ( .A1(n16019), .A2(n11505), .B1(n9711), .B2(n16016), .ZN(
        n11003) );
  NOR2_X1 U12854 ( .A1(n15982), .A2(n15686), .ZN(n11002) );
  AOI211_X1 U12855 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n11004), .A(n11003), .B(
        n11002), .ZN(n11005) );
  OAI21_X1 U12856 ( .B1(n11006), .B2(n16022), .A(n11005), .ZN(P1_U3237) );
  INV_X1 U12857 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n11011) );
  OAI211_X1 U12858 ( .C1(n11009), .C2(n11008), .A(n15427), .B(n11007), .ZN(
        n11010) );
  NAND2_X1 U12859 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n11578) );
  OAI211_X1 U12860 ( .C1(n15430), .C2(n11011), .A(n11010), .B(n11578), .ZN(
        n11018) );
  OAI211_X1 U12861 ( .C1(n11014), .C2(n11013), .A(n15426), .B(n11012), .ZN(
        n11015) );
  OAI21_X1 U12862 ( .B1(n14812), .B2(n11016), .A(n11015), .ZN(n11017) );
  OR3_X1 U12863 ( .A1(n11019), .A2(n11018), .A3(n11017), .ZN(P1_U3247) );
  INV_X1 U12864 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n11023) );
  INV_X1 U12865 ( .A(n11088), .ZN(n11021) );
  INV_X1 U12866 ( .A(n14423), .ZN(n12532) );
  NOR2_X1 U12867 ( .A1(n12532), .A2(n15797), .ZN(n11020) );
  INV_X1 U12868 ( .A(n10348), .ZN(n11097) );
  OR2_X1 U12869 ( .A1(n11097), .A2(n11977), .ZN(n11238) );
  OAI21_X1 U12870 ( .B1(n11020), .B2(n11971), .A(n11238), .ZN(n11964) );
  AOI21_X1 U12871 ( .B1(n7629), .B2(n11021), .A(n11964), .ZN(n11965) );
  OAI21_X1 U12872 ( .B1(n9421), .B2(n11971), .A(n11965), .ZN(n11338) );
  NAND2_X1 U12873 ( .A1(n15970), .A2(n11338), .ZN(n11022) );
  OAI21_X1 U12874 ( .B1(n15970), .B2(n11023), .A(n11022), .ZN(P2_U3499) );
  INV_X1 U12875 ( .A(SI_16_), .ZN(n13901) );
  OAI222_X1 U12876 ( .A1(P3_U3151), .A2(n13365), .B1(n13995), .B2(n13901), 
        .C1(n13993), .C2(n11024), .ZN(P3_U3279) );
  INV_X1 U12877 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11034) );
  XNOR2_X1 U12878 ( .A(n11025), .B(n11028), .ZN(n11607) );
  INV_X1 U12879 ( .A(n11026), .ZN(n11472) );
  INV_X1 U12880 ( .A(n11027), .ZN(n15805) );
  AOI211_X1 U12881 ( .C1(n11405), .C2(n11472), .A(n14360), .B(n15805), .ZN(
        n11605) );
  AOI21_X1 U12882 ( .B1(n15959), .B2(n11405), .A(n11605), .ZN(n11032) );
  XNOR2_X1 U12883 ( .A(n11029), .B(n11028), .ZN(n11031) );
  NAND2_X1 U12884 ( .A1(n14152), .A2(n14191), .ZN(n11030) );
  OAI21_X1 U12885 ( .B1(n11803), .B2(n11977), .A(n11030), .ZN(n11412) );
  AOI21_X1 U12886 ( .B1(n11031), .B2(n15797), .A(n11412), .ZN(n11610) );
  OAI211_X1 U12887 ( .C1(n15834), .C2(n11607), .A(n11032), .B(n11610), .ZN(
        n11361) );
  NAND2_X1 U12888 ( .A1(n11361), .A2(n15970), .ZN(n11033) );
  OAI21_X1 U12889 ( .B1(n15970), .B2(n11034), .A(n11033), .ZN(P2_U3504) );
  MUX2_X1 U12890 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n7206), .Z(n11179) );
  XOR2_X1 U12891 ( .A(n11185), .B(n11179), .Z(n11181) );
  INV_X1 U12892 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11046) );
  INV_X1 U12893 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11035) );
  MUX2_X1 U12894 ( .A(n11046), .B(n11035), .S(n7206), .Z(n11153) );
  NAND2_X1 U12895 ( .A1(n11153), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11114) );
  OAI22_X1 U12896 ( .A1(n11115), .A2(n11114), .B1(n11036), .B2(n7493), .ZN(
        n11132) );
  MUX2_X1 U12897 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n7166), .Z(n11037) );
  INV_X1 U12898 ( .A(n11037), .ZN(n11038) );
  MUX2_X1 U12899 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n7206), .Z(n11039) );
  XNOR2_X1 U12900 ( .A(n11039), .B(n11173), .ZN(n11164) );
  XOR2_X1 U12901 ( .A(n11181), .B(n11182), .Z(n11079) );
  INV_X1 U12902 ( .A(n11185), .ZN(n11191) );
  NAND2_X1 U12903 ( .A1(n11040), .A2(n11200), .ZN(n11041) );
  NAND2_X1 U12904 ( .A1(n11042), .A2(n11041), .ZN(n11073) );
  INV_X1 U12905 ( .A(n11073), .ZN(n11043) );
  NAND2_X1 U12906 ( .A1(n11220), .A2(n12113), .ZN(n11072) );
  INV_X1 U12907 ( .A(n11058), .ZN(n11057) );
  INV_X1 U12908 ( .A(P3_U3897), .ZN(n13223) );
  INV_X1 U12909 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11045) );
  MUX2_X1 U12910 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n11045), .S(n11062), .Z(
        n11136) );
  INV_X1 U12911 ( .A(n11156), .ZN(n11047) );
  NAND2_X1 U12912 ( .A1(n11129), .A2(n11047), .ZN(n11048) );
  NAND2_X1 U12913 ( .A1(n8375), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11049) );
  NAND2_X1 U12914 ( .A1(n11048), .A2(n11049), .ZN(n11117) );
  INV_X1 U12915 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11116) );
  NAND2_X1 U12916 ( .A1(n11119), .A2(n11049), .ZN(n11135) );
  NAND2_X1 U12917 ( .A1(n7498), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n11050) );
  NAND2_X1 U12918 ( .A1(n11134), .A2(n11050), .ZN(n11051) );
  NAND2_X1 U12919 ( .A1(n11051), .A2(n11173), .ZN(n11053) );
  INV_X1 U12920 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11168) );
  INV_X1 U12921 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11052) );
  MUX2_X1 U12922 ( .A(n11052), .B(P3_REG2_REG_4__SCAN_IN), .S(n11185), .Z(
        n11054) );
  AND3_X1 U12923 ( .A1(n11170), .A2(n11054), .A3(n11053), .ZN(n11055) );
  NOR2_X1 U12924 ( .A1(n11184), .A2(n11055), .ZN(n11076) );
  INV_X1 U12925 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15682) );
  NAND2_X1 U12926 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n11162), .ZN(n11059) );
  NAND2_X1 U12927 ( .A1(n11129), .A2(n11059), .ZN(n11060) );
  NAND2_X1 U12928 ( .A1(n8375), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11061) );
  NAND2_X1 U12929 ( .A1(n11060), .A2(n11061), .ZN(n11121) );
  INV_X1 U12930 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11748) );
  NAND2_X1 U12931 ( .A1(n7498), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n11063) );
  NAND2_X1 U12932 ( .A1(n11064), .A2(n11173), .ZN(n11066) );
  OAI21_X1 U12933 ( .B1(n11064), .B2(n11173), .A(n11066), .ZN(n11165) );
  INV_X1 U12934 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15727) );
  NAND2_X1 U12935 ( .A1(n11167), .A2(n11066), .ZN(n11065) );
  INV_X1 U12936 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15741) );
  MUX2_X1 U12937 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n15741), .S(n11185), .Z(
        n11067) );
  NAND2_X1 U12938 ( .A1(n11065), .A2(n11067), .ZN(n11190) );
  INV_X1 U12939 ( .A(n11066), .ZN(n11068) );
  NOR2_X1 U12940 ( .A1(n11068), .A2(n11067), .ZN(n11069) );
  NAND2_X1 U12941 ( .A1(n11167), .A2(n11069), .ZN(n11070) );
  NAND2_X1 U12942 ( .A1(n11190), .A2(n11070), .ZN(n11071) );
  NAND2_X1 U12943 ( .A1(n13422), .A2(n11071), .ZN(n11075) );
  INV_X1 U12944 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n13963) );
  NOR2_X1 U12945 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13963), .ZN(n11732) );
  AOI21_X1 U12946 ( .B1(n15246), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11732), .ZN(
        n11074) );
  OAI211_X1 U12947 ( .C1(n11076), .C2(n15636), .A(n11075), .B(n11074), .ZN(
        n11077) );
  AOI21_X1 U12948 ( .B1(n11191), .B2(n15618), .A(n11077), .ZN(n11078) );
  OAI21_X1 U12949 ( .B1(n11079), .B2(n13390), .A(n11078), .ZN(P3_U3186) );
  INV_X1 U12950 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n14207) );
  NAND2_X1 U12951 ( .A1(n11081), .A2(n11080), .ZN(n11386) );
  NOR2_X1 U12952 ( .A1(n15249), .A2(n11386), .ZN(n11086) );
  INV_X1 U12953 ( .A(n11086), .ZN(n11083) );
  INV_X1 U12954 ( .A(n11388), .ZN(n11082) );
  AOI21_X1 U12955 ( .B1(n11083), .B2(n11089), .A(n11082), .ZN(n11232) );
  NAND2_X1 U12956 ( .A1(n11232), .A2(n11084), .ZN(n11085) );
  AND2_X1 U12957 ( .A1(n11086), .A2(n15250), .ZN(n11108) );
  INV_X1 U12958 ( .A(n11087), .ZN(n12503) );
  NOR2_X1 U12959 ( .A1(n11088), .A2(n12503), .ZN(n15707) );
  NAND2_X1 U12960 ( .A1(n11108), .A2(n15707), .ZN(n11091) );
  INV_X1 U12961 ( .A(n11089), .ZN(n11090) );
  INV_X1 U12962 ( .A(n14152), .ZN(n11790) );
  OAI22_X1 U12963 ( .A1(n11790), .A2(n11228), .B1(n11341), .B2(n11977), .ZN(
        n11332) );
  AOI22_X1 U12964 ( .A1(n14095), .A2(n11332), .B1(P2_U3088), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n11093) );
  OAI21_X1 U12965 ( .B1(n11782), .B2(n14135), .A(n11093), .ZN(n11112) );
  NOR2_X1 U12966 ( .A1(n7209), .A2(n11228), .ZN(n11103) );
  NAND2_X1 U12967 ( .A1(n11094), .A2(n15339), .ZN(n11095) );
  XNOR2_X1 U12968 ( .A(n11383), .B(n14072), .ZN(n11101) );
  OR2_X1 U12969 ( .A1(n14308), .A2(n11097), .ZN(n11098) );
  INV_X1 U12970 ( .A(n11098), .ZN(n11100) );
  OR2_X1 U12971 ( .A1(n14308), .A2(n11241), .ZN(n11237) );
  NAND2_X1 U12972 ( .A1(n14072), .A2(n11292), .ZN(n11225) );
  AND2_X1 U12973 ( .A1(n11237), .A2(n11225), .ZN(n11099) );
  OAI21_X1 U12974 ( .B1(n11100), .B2(n11377), .A(n11227), .ZN(n11102) );
  XNOR2_X1 U12975 ( .A(n11101), .B(n11103), .ZN(n11378) );
  XNOR2_X1 U12976 ( .A(n11336), .B(n14038), .ZN(n11346) );
  NOR2_X1 U12977 ( .A1(n7209), .A2(n11104), .ZN(n11105) );
  NAND2_X1 U12978 ( .A1(n11346), .A2(n11105), .ZN(n11342) );
  OAI21_X1 U12979 ( .B1(n11346), .B2(n11105), .A(n11342), .ZN(n11109) );
  NOR2_X1 U12980 ( .A1(n15959), .A2(n11106), .ZN(n11107) );
  NAND2_X2 U12981 ( .A1(n11108), .A2(n11107), .ZN(n14163) );
  AOI211_X1 U12982 ( .C1(n11110), .C2(n11109), .A(n14163), .B(n11345), .ZN(
        n11111) );
  AOI211_X1 U12983 ( .C1(n14207), .C2(n14155), .A(n11112), .B(n11111), .ZN(
        n11113) );
  INV_X1 U12984 ( .A(n11113), .ZN(P2_U3190) );
  INV_X1 U12985 ( .A(n11114), .ZN(n11158) );
  XNOR2_X1 U12986 ( .A(n11115), .B(n11158), .ZN(n11131) );
  INV_X1 U12987 ( .A(n15636), .ZN(n13242) );
  NAND2_X1 U12988 ( .A1(n11117), .A2(n11116), .ZN(n11118) );
  NAND2_X1 U12989 ( .A1(n11119), .A2(n11118), .ZN(n11120) );
  NAND2_X1 U12990 ( .A1(n13242), .A2(n11120), .ZN(n11127) );
  NAND2_X1 U12991 ( .A1(n11121), .A2(n11748), .ZN(n11122) );
  NAND2_X1 U12992 ( .A1(n11123), .A2(n11122), .ZN(n11124) );
  NAND2_X1 U12993 ( .A1(n13422), .A2(n11124), .ZN(n11126) );
  AOI22_X1 U12994 ( .A1(n15246), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11125) );
  NAND3_X1 U12995 ( .A1(n11127), .A2(n11126), .A3(n11125), .ZN(n11128) );
  AOI21_X1 U12996 ( .B1(n11129), .B2(n15618), .A(n11128), .ZN(n11130) );
  OAI21_X1 U12997 ( .B1(n13390), .B2(n11131), .A(n11130), .ZN(P3_U3183) );
  XOR2_X1 U12998 ( .A(n11132), .B(n11133), .Z(n11147) );
  OAI21_X1 U12999 ( .B1(n11136), .B2(n11135), .A(n11134), .ZN(n11137) );
  NAND2_X1 U13000 ( .A1(n13242), .A2(n11137), .ZN(n11144) );
  OAI21_X1 U13001 ( .B1(n11140), .B2(n11139), .A(n11138), .ZN(n11141) );
  NAND2_X1 U13002 ( .A1(n13422), .A2(n11141), .ZN(n11143) );
  AOI22_X1 U13003 ( .A1(n15246), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11142) );
  NAND3_X1 U13004 ( .A1(n11144), .A2(n11143), .A3(n11142), .ZN(n11145) );
  AOI21_X1 U13005 ( .B1(n7409), .B2(n15618), .A(n11145), .ZN(n11146) );
  OAI21_X1 U13006 ( .B1(n11147), .B2(n13390), .A(n11146), .ZN(P3_U3184) );
  INV_X1 U13007 ( .A(SI_17_), .ZN(n13799) );
  OAI222_X1 U13008 ( .A1(n13787), .A2(n13799), .B1(n13993), .B2(n11148), .C1(
        n13386), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U13009 ( .A(n11463), .ZN(n11891) );
  INV_X1 U13010 ( .A(n11149), .ZN(n11151) );
  OAI222_X1 U13011 ( .A1(P1_U3086), .A2(n11891), .B1(n15233), .B2(n11151), 
        .C1(n11150), .C2(n15224), .ZN(P1_U3343) );
  INV_X1 U13012 ( .A(n12615), .ZN(n12604) );
  OAI222_X1 U13013 ( .A1(n14592), .A2(n11152), .B1(n14578), .B2(n11151), .C1(
        n12604), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U13014 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11224) );
  OAI22_X1 U13015 ( .A1(n15651), .A2(n15432), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11224), .ZN(n11155) );
  NOR2_X1 U13016 ( .A1(n13422), .A2(n15638), .ZN(n11157) );
  NOR3_X1 U13017 ( .A1(n11157), .A2(P3_IR_REG_0__SCAN_IN), .A3(n11153), .ZN(
        n11154) );
  AOI211_X1 U13018 ( .C1(n11156), .C2(n13242), .A(n11155), .B(n11154), .ZN(
        n11161) );
  INV_X1 U13019 ( .A(n11157), .ZN(n11159) );
  OAI21_X1 U13020 ( .B1(n11159), .B2(n13242), .A(n11158), .ZN(n11160) );
  OAI211_X1 U13021 ( .C1(n11162), .C2(n15641), .A(n11161), .B(n11160), .ZN(
        P3_U3182) );
  XOR2_X1 U13022 ( .A(n11164), .B(n11163), .Z(n11178) );
  NAND2_X1 U13023 ( .A1(n11165), .A2(n15727), .ZN(n11166) );
  NAND2_X1 U13024 ( .A1(n11167), .A2(n11166), .ZN(n11176) );
  AND2_X1 U13025 ( .A1(n11170), .A2(n11169), .ZN(n11172) );
  NOR2_X1 U13026 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13944), .ZN(n11442) );
  AOI21_X1 U13027 ( .B1(n15246), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n11442), .ZN(
        n11171) );
  OAI21_X1 U13028 ( .B1(n15636), .B2(n11172), .A(n11171), .ZN(n11175) );
  NOR2_X1 U13029 ( .A1(n15641), .A2(n11173), .ZN(n11174) );
  AOI211_X1 U13030 ( .C1(n13422), .C2(n11176), .A(n11175), .B(n11174), .ZN(
        n11177) );
  OAI21_X1 U13031 ( .B1(n11178), .B2(n13390), .A(n11177), .ZN(P3_U3185) );
  INV_X1 U13032 ( .A(n11179), .ZN(n11180) );
  MUX2_X1 U13033 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n7206), .Z(n11760) );
  XNOR2_X1 U13034 ( .A(n11760), .B(n11759), .ZN(n11761) );
  XNOR2_X1 U13035 ( .A(n11762), .B(n11761), .ZN(n11183) );
  NAND2_X1 U13036 ( .A1(n11183), .A2(n15638), .ZN(n11199) );
  INV_X1 U13037 ( .A(n11759), .ZN(n11186) );
  AOI21_X1 U13038 ( .B1(n11187), .B2(n11186), .A(n13240), .ZN(n11188) );
  OAI21_X1 U13039 ( .B1(n11188), .B2(P3_REG2_REG_5__SCAN_IN), .A(n13237), .ZN(
        n11197) );
  NOR2_X1 U13040 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8418), .ZN(n11908) );
  INV_X1 U13041 ( .A(n11908), .ZN(n11189) );
  OAI21_X1 U13042 ( .B1(n15651), .B2(n15476), .A(n11189), .ZN(n11196) );
  INV_X1 U13043 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15768) );
  OAI21_X1 U13044 ( .B1(n11191), .B2(n15741), .A(n11190), .ZN(n11192) );
  NAND2_X1 U13045 ( .A1(n11192), .A2(n11759), .ZN(n11768) );
  OAI21_X1 U13046 ( .B1(n11192), .B2(n11759), .A(n11768), .ZN(n11193) );
  AOI21_X1 U13047 ( .B1(n15768), .B2(n11193), .A(n13231), .ZN(n11194) );
  NOR2_X1 U13048 ( .A1(n15631), .A2(n11194), .ZN(n11195) );
  AOI211_X1 U13049 ( .C1(n13242), .C2(n11197), .A(n11196), .B(n11195), .ZN(
        n11198) );
  OAI211_X1 U13050 ( .C1(n15641), .C2(n11759), .A(n11199), .B(n11198), .ZN(
        P3_U3187) );
  INV_X1 U13051 ( .A(n11208), .ZN(n11204) );
  AND3_X1 U13052 ( .A1(n11317), .A2(n11201), .A3(n11200), .ZN(n11203) );
  OR2_X1 U13053 ( .A1(n11217), .A2(n11209), .ZN(n11202) );
  OAI211_X1 U13054 ( .C1(n11219), .C2(n11204), .A(n11203), .B(n11202), .ZN(
        n11205) );
  NAND2_X1 U13055 ( .A1(n11205), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11207) );
  OR2_X1 U13056 ( .A1(n11217), .A2(n11215), .ZN(n11206) );
  NOR2_X1 U13057 ( .A1(n13190), .A2(P3_U3151), .ZN(n11375) );
  NAND3_X1 U13058 ( .A1(n11219), .A2(n11208), .A3(n15886), .ZN(n11212) );
  INV_X1 U13059 ( .A(n11209), .ZN(n11210) );
  NAND2_X1 U13060 ( .A1(n11217), .A2(n11210), .ZN(n11211) );
  NAND2_X1 U13061 ( .A1(n11212), .A2(n11211), .ZN(n11214) );
  INV_X1 U13062 ( .A(n11215), .ZN(n11216) );
  AND2_X1 U13063 ( .A1(n11217), .A2(n11216), .ZN(n11308) );
  INV_X1 U13064 ( .A(n11308), .ZN(n11218) );
  OR2_X1 U13065 ( .A1(n11219), .A2(n11821), .ZN(n11221) );
  OAI22_X1 U13066 ( .A1(n11303), .A2(n13174), .B1(n13178), .B2(n8118), .ZN(
        n11222) );
  AOI21_X1 U13067 ( .B1(n13168), .B2(n11247), .A(n11222), .ZN(n11223) );
  OAI21_X1 U13068 ( .B1(n11375), .B2(n11224), .A(n11223), .ZN(P3_U3172) );
  OR2_X1 U13069 ( .A1(n14163), .A2(n14308), .ZN(n14146) );
  INV_X1 U13070 ( .A(n14146), .ZN(n14126) );
  INV_X1 U13071 ( .A(n11241), .ZN(n11281) );
  INV_X1 U13072 ( .A(n11225), .ZN(n11226) );
  AOI22_X1 U13073 ( .A1(n14126), .A2(n11281), .B1(n11226), .B2(n14102), .ZN(
        n11236) );
  INV_X1 U13074 ( .A(n11227), .ZN(n11379) );
  NAND2_X1 U13075 ( .A1(n14152), .A2(n14194), .ZN(n11230) );
  OR2_X1 U13076 ( .A1(n11228), .A2(n11977), .ZN(n11229) );
  AND2_X1 U13077 ( .A1(n11230), .A2(n11229), .ZN(n11288) );
  INV_X1 U13078 ( .A(n11288), .ZN(n11231) );
  AOI22_X1 U13079 ( .A1(n14102), .A2(n11379), .B1(n14095), .B2(n11231), .ZN(
        n11234) );
  AND2_X1 U13080 ( .A1(n11232), .A2(n15250), .ZN(n11376) );
  INV_X1 U13081 ( .A(n11376), .ZN(n11240) );
  AOI22_X1 U13082 ( .A1(n14159), .A2(n7436), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n11240), .ZN(n11233) );
  OAI211_X1 U13083 ( .C1(n11236), .C2(n11235), .A(n11234), .B(n11233), .ZN(
        P2_U3194) );
  AOI21_X1 U13084 ( .B1(n14102), .B2(n11237), .A(n14159), .ZN(n11244) );
  INV_X1 U13085 ( .A(n11238), .ZN(n11239) );
  AOI22_X1 U13086 ( .A1(n11240), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n14095), 
        .B2(n11239), .ZN(n11243) );
  NAND3_X1 U13087 ( .A1(n14126), .A2(n14194), .A3(n11241), .ZN(n11242) );
  OAI211_X1 U13088 ( .C1(n11244), .C2(n11292), .A(n11243), .B(n11242), .ZN(
        P2_U3204) );
  INV_X1 U13089 ( .A(n11245), .ZN(n11246) );
  NAND3_X1 U13090 ( .A1(n11247), .A2(n15886), .A3(n11246), .ZN(n11248) );
  OAI21_X1 U13091 ( .B1(n11303), .B2(n13629), .A(n11248), .ZN(n11446) );
  INV_X1 U13092 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11249) );
  OAI22_X1 U13093 ( .A1(n8118), .A2(n13767), .B1(n15898), .B2(n11249), .ZN(
        n11250) );
  AOI21_X1 U13094 ( .B1(n11446), .B2(n15898), .A(n11250), .ZN(n11251) );
  INV_X1 U13095 ( .A(n11251), .ZN(P3_U3390) );
  XNOR2_X1 U13096 ( .A(n11924), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n11261) );
  NAND2_X1 U13097 ( .A1(n11263), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n11252) );
  NAND2_X1 U13098 ( .A1(n11253), .A2(n11252), .ZN(n15276) );
  INV_X1 U13099 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11254) );
  XNOR2_X1 U13100 ( .A(n15270), .B(n11254), .ZN(n15277) );
  NAND2_X1 U13101 ( .A1(n15276), .A2(n15277), .ZN(n15275) );
  NAND2_X1 U13102 ( .A1(n15270), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n11255) );
  NAND2_X1 U13103 ( .A1(n15275), .A2(n11255), .ZN(n14228) );
  INV_X1 U13104 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11256) );
  MUX2_X1 U13105 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11256), .S(n14226), .Z(
        n14229) );
  NAND2_X1 U13106 ( .A1(n14228), .A2(n14229), .ZN(n14227) );
  NAND2_X1 U13107 ( .A1(n14226), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n11257) );
  NAND2_X1 U13108 ( .A1(n14227), .A2(n11257), .ZN(n14241) );
  INV_X1 U13109 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11650) );
  MUX2_X1 U13110 ( .A(n11650), .B(P2_REG2_REG_8__SCAN_IN), .S(n14238), .Z(
        n14242) );
  NAND2_X1 U13111 ( .A1(n14241), .A2(n14242), .ZN(n14240) );
  NAND2_X1 U13112 ( .A1(n11267), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11258) );
  NAND2_X1 U13113 ( .A1(n14240), .A2(n11258), .ZN(n11260) );
  OR2_X1 U13114 ( .A1(n11260), .A2(n11261), .ZN(n11915) );
  INV_X1 U13115 ( .A(n11915), .ZN(n11259) );
  AOI21_X1 U13116 ( .B1(n11261), .B2(n11260), .A(n11259), .ZN(n11276) );
  INV_X1 U13117 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n11264) );
  MUX2_X1 U13118 ( .A(n11264), .B(P2_REG1_REG_6__SCAN_IN), .S(n15270), .Z(
        n15273) );
  INV_X1 U13119 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11265) );
  MUX2_X1 U13120 ( .A(n11265), .B(P2_REG1_REG_7__SCAN_IN), .S(n14226), .Z(
        n14221) );
  AOI21_X1 U13121 ( .B1(n14226), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7239), .ZN(
        n14235) );
  INV_X1 U13122 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11266) );
  MUX2_X1 U13123 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n11266), .S(n14238), .Z(
        n14234) );
  INV_X1 U13124 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11268) );
  MUX2_X1 U13125 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n11268), .S(n11924), .Z(
        n11269) );
  OAI21_X1 U13126 ( .B1(n11270), .B2(n11269), .A(n11923), .ZN(n11271) );
  INV_X1 U13127 ( .A(n15368), .ZN(n15251) );
  NAND2_X1 U13128 ( .A1(n11271), .A2(n15251), .ZN(n11275) );
  NAND2_X1 U13129 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n11989) );
  INV_X1 U13130 ( .A(n11989), .ZN(n11273) );
  NOR2_X1 U13131 ( .A1(n15322), .A2(n11913), .ZN(n11272) );
  AOI211_X1 U13132 ( .C1(n15271), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n11273), .B(
        n11272), .ZN(n11274) );
  OAI211_X1 U13133 ( .C1(n11276), .C2(n15364), .A(n11275), .B(n11274), .ZN(
        P2_U3223) );
  INV_X1 U13134 ( .A(n11277), .ZN(n11280) );
  OAI222_X1 U13135 ( .A1(n14592), .A2(n11278), .B1(n14578), .B2(n11280), .C1(
        n12616), .C2(P2_U3088), .ZN(P2_U3314) );
  OAI222_X1 U13136 ( .A1(P1_U3086), .A2(n14811), .B1(n15233), .B2(n11280), 
        .C1(n11279), .C2(n15224), .ZN(P1_U3342) );
  NAND2_X1 U13137 ( .A1(n11285), .A2(n11281), .ZN(n11282) );
  NAND2_X1 U13138 ( .A1(n11283), .A2(n11282), .ZN(n11284) );
  INV_X1 U13139 ( .A(n11284), .ZN(n11401) );
  NAND2_X1 U13140 ( .A1(n11284), .A2(n12532), .ZN(n11290) );
  OAI21_X1 U13141 ( .B1(n11286), .B2(n11285), .A(n15697), .ZN(n11287) );
  NAND2_X1 U13142 ( .A1(n11287), .A2(n15797), .ZN(n11289) );
  AND3_X1 U13143 ( .A1(n11290), .A2(n11289), .A3(n11288), .ZN(n11398) );
  INV_X1 U13144 ( .A(n15695), .ZN(n11291) );
  OAI211_X1 U13145 ( .C1(n11569), .C2(n11292), .A(n11291), .B(n14308), .ZN(
        n11395) );
  OAI211_X1 U13146 ( .C1(n11401), .C2(n9421), .A(n11398), .B(n11395), .ZN(
        n11567) );
  NOR2_X1 U13147 ( .A1(n15970), .A2(n10763), .ZN(n11293) );
  AOI21_X1 U13148 ( .B1(n15970), .B2(n11567), .A(n11293), .ZN(n11294) );
  OAI21_X1 U13149 ( .B1(n11569), .B2(n14498), .A(n11294), .ZN(P2_U3500) );
  INV_X1 U13150 ( .A(n11295), .ZN(n11296) );
  NAND2_X1 U13151 ( .A1(n13773), .A2(n11296), .ZN(n11299) );
  NAND2_X1 U13152 ( .A1(n11820), .A2(n11787), .ZN(n11297) );
  NAND2_X1 U13153 ( .A1(n8118), .A2(n13103), .ZN(n11300) );
  NAND2_X1 U13154 ( .A1(n11737), .A2(n11300), .ZN(n11306) );
  XNOR2_X1 U13155 ( .A(n11301), .B(n7167), .ZN(n11302) );
  NAND2_X1 U13156 ( .A1(n11303), .A2(n11302), .ZN(n11366) );
  OAI21_X1 U13157 ( .B1(n11303), .B2(n11302), .A(n11366), .ZN(n11305) );
  INV_X1 U13158 ( .A(n11367), .ZN(n11304) );
  AOI21_X1 U13159 ( .B1(n11306), .B2(n11305), .A(n11304), .ZN(n11313) );
  OAI22_X1 U13160 ( .A1(n7398), .A2(n13174), .B1(n7432), .B2(n13178), .ZN(
        n11311) );
  INV_X1 U13161 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11309) );
  NOR2_X1 U13162 ( .A1(n11375), .A2(n11309), .ZN(n11310) );
  AOI211_X1 U13163 ( .C1(n13172), .C2(n13224), .A(n11311), .B(n11310), .ZN(
        n11312) );
  OAI21_X1 U13164 ( .B1(n11313), .B2(n13200), .A(n11312), .ZN(P3_U3162) );
  AOI21_X1 U13165 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n13634), .A(n11446), .ZN(
        n11323) );
  XNOR2_X1 U13166 ( .A(n11316), .B(n11315), .ZN(n11319) );
  NAND3_X1 U13167 ( .A1(n11319), .A2(n11318), .A3(n11317), .ZN(n11320) );
  OR2_X1 U13168 ( .A1(n11821), .A2(n15886), .ZN(n11940) );
  OAI22_X1 U13169 ( .A1(n8118), .A2(n13637), .B1(n13565), .B2(n11046), .ZN(
        n11321) );
  INV_X1 U13170 ( .A(n11321), .ZN(n11322) );
  OAI21_X1 U13171 ( .B1(n11323), .B2(n13635), .A(n11322), .ZN(P3_U3233) );
  OR2_X1 U13172 ( .A1(n11325), .A2(n11324), .ZN(n11326) );
  AND2_X1 U13173 ( .A1(n11327), .A2(n11326), .ZN(n11335) );
  INV_X1 U13174 ( .A(n11335), .ZN(n11630) );
  AOI21_X1 U13175 ( .B1(n11336), .B2(n15694), .A(n14360), .ZN(n11328) );
  AND2_X1 U13176 ( .A1(n11470), .A2(n11328), .ZN(n11626) );
  OAI21_X1 U13177 ( .B1(n11331), .B2(n11330), .A(n11329), .ZN(n11333) );
  AOI21_X1 U13178 ( .B1(n11333), .B2(n15797), .A(n11332), .ZN(n11334) );
  OAI21_X1 U13179 ( .B1(n11335), .B2(n14423), .A(n11334), .ZN(n11625) );
  AOI211_X1 U13180 ( .C1(n15758), .C2(n11630), .A(n11626), .B(n11625), .ZN(
        n11785) );
  AOI22_X1 U13181 ( .A1(n14510), .A2(n11336), .B1(n15968), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n11337) );
  OAI21_X1 U13182 ( .B1(n11785), .B2(n15968), .A(n11337), .ZN(P2_U3502) );
  INV_X1 U13183 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n11340) );
  NAND2_X1 U13184 ( .A1(n15973), .A2(n11338), .ZN(n11339) );
  OAI21_X1 U13185 ( .B1(n15973), .B2(n11340), .A(n11339), .ZN(P2_U3430) );
  XNOR2_X1 U13186 ( .A(n11473), .B(n14038), .ZN(n11408) );
  NOR2_X1 U13187 ( .A1(n7209), .A2(n11341), .ZN(n11402) );
  XNOR2_X1 U13188 ( .A(n11408), .B(n11402), .ZN(n11355) );
  INV_X1 U13189 ( .A(n11342), .ZN(n11343) );
  INV_X1 U13190 ( .A(n11411), .ZN(n11358) );
  NAND3_X1 U13191 ( .A1(n14126), .A2(n11346), .A3(n14192), .ZN(n11347) );
  OAI21_X1 U13192 ( .B1(n7885), .B2(n14163), .A(n11347), .ZN(n11356) );
  NOR2_X1 U13193 ( .A1(n14092), .A2(n11474), .ZN(n11354) );
  INV_X1 U13194 ( .A(n11473), .ZN(n15754) );
  NAND2_X1 U13195 ( .A1(n14153), .A2(n14190), .ZN(n11349) );
  NAND2_X1 U13196 ( .A1(n14152), .A2(n14192), .ZN(n11348) );
  AND2_X1 U13197 ( .A1(n11349), .A2(n11348), .ZN(n11482) );
  INV_X1 U13198 ( .A(n11482), .ZN(n11350) );
  NAND2_X1 U13199 ( .A1(n14095), .A2(n11350), .ZN(n11351) );
  OAI211_X1 U13200 ( .C1(n14135), .C2(n15754), .A(n11352), .B(n11351), .ZN(
        n11353) );
  AOI211_X1 U13201 ( .C1(n11356), .C2(n11355), .A(n11354), .B(n11353), .ZN(
        n11357) );
  OAI21_X1 U13202 ( .B1(n11358), .B2(n14163), .A(n11357), .ZN(P2_U3202) );
  OAI222_X1 U13203 ( .A1(n13993), .A2(n11360), .B1(n13995), .B2(n11359), .C1(
        P3_U3151), .C2(n13412), .ZN(P3_U3276) );
  NAND2_X1 U13204 ( .A1(n11361), .A2(n15973), .ZN(n11362) );
  OAI21_X1 U13205 ( .B1(n15973), .B2(n9053), .A(n11362), .ZN(P2_U3445) );
  INV_X1 U13206 ( .A(n13407), .ZN(n13398) );
  INV_X1 U13207 ( .A(n11363), .ZN(n11364) );
  OAI222_X1 U13208 ( .A1(P3_U3151), .A2(n13398), .B1(n13995), .B2(n13898), 
        .C1(n13993), .C2(n11364), .ZN(P3_U3277) );
  INV_X1 U13209 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n13878) );
  XNOR2_X1 U13210 ( .A(n11434), .B(n7398), .ZN(n11369) );
  NAND2_X1 U13211 ( .A1(n11367), .A2(n11366), .ZN(n11368) );
  NAND2_X1 U13212 ( .A1(n11368), .A2(n11369), .ZN(n11438) );
  OAI21_X1 U13213 ( .B1(n11369), .B2(n11368), .A(n11438), .ZN(n11370) );
  NAND2_X1 U13214 ( .A1(n11370), .A2(n13168), .ZN(n11374) );
  OAI22_X1 U13215 ( .A1(n8398), .A2(n13174), .B1(n13178), .B2(n15678), .ZN(
        n11372) );
  AOI21_X1 U13216 ( .B1(n13172), .B2(n11371), .A(n11372), .ZN(n11373) );
  OAI211_X1 U13217 ( .C1(n11375), .C2(n13878), .A(n11374), .B(n11373), .ZN(
        P3_U3177) );
  AOI22_X1 U13218 ( .A1(n14153), .A2(n14192), .B1(n14152), .B2(n10348), .ZN(
        n15701) );
  INV_X1 U13219 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n15715) );
  OAI22_X1 U13220 ( .A1(n14157), .A2(n15701), .B1(n11376), .B2(n15715), .ZN(
        n11382) );
  AOI22_X1 U13221 ( .A1(n14126), .A2(n10348), .B1(n14102), .B2(n11377), .ZN(
        n11380) );
  NOR3_X1 U13222 ( .A1(n11380), .A2(n11379), .A3(n11378), .ZN(n11381) );
  AOI211_X1 U13223 ( .C1(n11383), .C2(n14159), .A(n11382), .B(n11381), .ZN(
        n11384) );
  OAI21_X1 U13224 ( .B1(n11385), .B2(n14163), .A(n11384), .ZN(P2_U3209) );
  INV_X1 U13225 ( .A(n11386), .ZN(n11387) );
  AND2_X1 U13226 ( .A1(n11388), .A2(n11387), .ZN(n11389) );
  NAND3_X1 U13227 ( .A1(n15250), .A2(n11389), .A3(n15249), .ZN(n11392) );
  NAND2_X1 U13228 ( .A1(n11967), .A2(n11390), .ZN(n11606) );
  INV_X1 U13229 ( .A(n11606), .ZN(n11391) );
  NAND2_X1 U13230 ( .A1(n15721), .A2(n11391), .ZN(n14431) );
  INV_X1 U13231 ( .A(n11392), .ZN(n11393) );
  INV_X1 U13232 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11394) );
  OAI22_X1 U13233 ( .A1(n15717), .A2(n11395), .B1(n11394), .B2(n15714), .ZN(
        n11396) );
  AOI21_X1 U13234 ( .B1(n15917), .B2(n7436), .A(n11396), .ZN(n11400) );
  MUX2_X1 U13235 ( .A(n10749), .B(n11398), .S(n15721), .Z(n11399) );
  OAI211_X1 U13236 ( .C1(n11401), .C2(n14431), .A(n11400), .B(n11399), .ZN(
        P2_U3264) );
  INV_X1 U13237 ( .A(n11408), .ZN(n11404) );
  INV_X1 U13238 ( .A(n11402), .ZN(n11403) );
  XNOR2_X1 U13239 ( .A(n11405), .B(n14038), .ZN(n11422) );
  NOR2_X1 U13240 ( .A1(n7209), .A2(n11429), .ZN(n11421) );
  XNOR2_X1 U13241 ( .A(n11422), .B(n11421), .ZN(n11407) );
  INV_X1 U13242 ( .A(n11407), .ZN(n11410) );
  AOI22_X1 U13243 ( .A1(n14126), .A2(n14191), .B1(n14102), .B2(n11408), .ZN(
        n11409) );
  NOR3_X1 U13244 ( .A1(n11411), .A2(n11410), .A3(n11409), .ZN(n11416) );
  AOI22_X1 U13245 ( .A1(n14095), .A2(n11412), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11414) );
  OR2_X1 U13246 ( .A1(n14092), .A2(n11600), .ZN(n11413) );
  OAI211_X1 U13247 ( .C1(n11602), .C2(n14135), .A(n11414), .B(n11413), .ZN(
        n11415) );
  INV_X1 U13248 ( .A(n11417), .ZN(P2_U3199) );
  INV_X1 U13249 ( .A(n11418), .ZN(n11420) );
  INV_X1 U13250 ( .A(n12838), .ZN(n12613) );
  OAI222_X1 U13251 ( .A1(n14592), .A2(n8046), .B1(n14578), .B2(n11420), .C1(
        P2_U3088), .C2(n12613), .ZN(P2_U3313) );
  INV_X1 U13252 ( .A(n14823), .ZN(n14837) );
  OAI222_X1 U13253 ( .A1(n14837), .A2(P1_U3086), .B1(n15233), .B2(n11420), 
        .C1(n11419), .C2(n15224), .ZN(P1_U3341) );
  INV_X1 U13254 ( .A(n11421), .ZN(n11425) );
  INV_X1 U13255 ( .A(n11422), .ZN(n11424) );
  XNOR2_X1 U13256 ( .A(n15801), .B(n14072), .ZN(n11802) );
  OR2_X1 U13257 ( .A1(n11803), .A2(n14308), .ZN(n11426) );
  NOR2_X1 U13258 ( .A1(n11802), .A2(n11426), .ZN(n11583) );
  AOI21_X1 U13259 ( .B1(n11802), .B2(n11426), .A(n11583), .ZN(n11427) );
  NAND2_X1 U13260 ( .A1(n11428), .A2(n11427), .ZN(n11585) );
  OAI211_X1 U13261 ( .C1(n11428), .C2(n11427), .A(n11585), .B(n14102), .ZN(
        n11433) );
  OAI22_X1 U13262 ( .A1(n11790), .A2(n11429), .B1(n11595), .B2(n11977), .ZN(
        n15796) );
  AOI22_X1 U13263 ( .A1(n14095), .A2(n15796), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11430) );
  OAI21_X1 U13264 ( .B1(n15811), .B2(n14135), .A(n11430), .ZN(n11431) );
  INV_X1 U13265 ( .A(n11431), .ZN(n11432) );
  OAI211_X1 U13266 ( .C1(n14092), .C2(n15799), .A(n11433), .B(n11432), .ZN(
        P2_U3211) );
  INV_X1 U13267 ( .A(n13190), .ZN(n12585) );
  INV_X1 U13268 ( .A(n11434), .ZN(n11435) );
  NAND2_X1 U13269 ( .A1(n11435), .A2(n7398), .ZN(n11436) );
  AND2_X1 U13270 ( .A1(n11438), .A2(n11436), .ZN(n11440) );
  XNOR2_X1 U13271 ( .A(n11722), .B(n8398), .ZN(n11439) );
  AND2_X1 U13272 ( .A1(n11439), .A2(n11436), .ZN(n11437) );
  NAND2_X1 U13273 ( .A1(n11438), .A2(n11437), .ZN(n11724) );
  OAI211_X1 U13274 ( .C1(n11440), .C2(n11439), .A(n13168), .B(n11724), .ZN(
        n11445) );
  OAI22_X1 U13275 ( .A1(n13195), .A2(n7398), .B1(n12235), .B2(n13174), .ZN(
        n11441) );
  AOI211_X1 U13276 ( .C1(n13197), .C2(n11443), .A(n11442), .B(n11441), .ZN(
        n11444) );
  OAI211_X1 U13277 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12585), .A(n11445), .B(
        n11444), .ZN(P3_U3158) );
  INV_X1 U13278 ( .A(n11446), .ZN(n11449) );
  INV_X1 U13279 ( .A(n13694), .ZN(n13688) );
  AOI22_X1 U13280 ( .A1(n13688), .A2(n11447), .B1(n15892), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n11448) );
  OAI21_X1 U13281 ( .B1(n11449), .B2(n15892), .A(n11448), .ZN(P3_U3459) );
  MUX2_X1 U13282 ( .A(n11892), .B(P1_REG2_REG_12__SCAN_IN), .S(n11463), .Z(
        n11453) );
  OAI21_X1 U13283 ( .B1(n11457), .B2(n11451), .A(n11450), .ZN(n11452) );
  NOR2_X1 U13284 ( .A1(n11452), .A2(n11453), .ZN(n11890) );
  AOI21_X1 U13285 ( .B1(n11453), .B2(n11452), .A(n11890), .ZN(n11465) );
  INV_X1 U13286 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n11454) );
  NAND2_X1 U13287 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14648)
         );
  OAI21_X1 U13288 ( .B1(n15430), .B2(n11454), .A(n14648), .ZN(n11462) );
  MUX2_X1 U13289 ( .A(n11885), .B(P1_REG1_REG_12__SCAN_IN), .S(n11463), .Z(
        n11459) );
  AOI21_X1 U13290 ( .B1(n11459), .B2(n11458), .A(n11884), .ZN(n11460) );
  NOR2_X1 U13291 ( .A1(n11460), .A2(n15397), .ZN(n11461) );
  AOI211_X1 U13292 ( .C1(n15423), .C2(n11463), .A(n11462), .B(n11461), .ZN(
        n11464) );
  OAI21_X1 U13293 ( .B1(n11465), .B2(n15413), .A(n11464), .ZN(P1_U3255) );
  INV_X1 U13294 ( .A(n14431), .ZN(n15944) );
  OR2_X1 U13295 ( .A1(n11467), .A2(n11466), .ZN(n11468) );
  NAND2_X1 U13296 ( .A1(n11469), .A2(n11468), .ZN(n15757) );
  AOI21_X1 U13297 ( .B1(n11473), .B2(n11470), .A(n14360), .ZN(n11471) );
  NAND2_X1 U13298 ( .A1(n11472), .A2(n11471), .ZN(n15753) );
  NAND2_X1 U13299 ( .A1(n15917), .A2(n11473), .ZN(n11477) );
  INV_X1 U13300 ( .A(n15714), .ZN(n15936) );
  INV_X1 U13301 ( .A(n11474), .ZN(n11475) );
  NAND2_X1 U13302 ( .A1(n15936), .A2(n11475), .ZN(n11476) );
  OAI211_X1 U13303 ( .C1(n15753), .C2(n15717), .A(n11477), .B(n11476), .ZN(
        n11486) );
  NAND2_X1 U13304 ( .A1(n15757), .A2(n12532), .ZN(n11484) );
  OAI21_X1 U13305 ( .B1(n11480), .B2(n11479), .A(n11478), .ZN(n11481) );
  NAND2_X1 U13306 ( .A1(n11481), .A2(n15797), .ZN(n11483) );
  NAND3_X1 U13307 ( .A1(n11484), .A2(n11483), .A3(n11482), .ZN(n15755) );
  MUX2_X1 U13308 ( .A(n15755), .B(P2_REG2_REG_4__SCAN_IN), .S(n15947), .Z(
        n11485) );
  AOI211_X1 U13309 ( .C1(n15944), .C2(n15757), .A(n11486), .B(n11485), .ZN(
        n11487) );
  INV_X1 U13310 ( .A(n11487), .ZN(P2_U3261) );
  NAND2_X1 U13311 ( .A1(n7516), .A2(n7476), .ZN(n11489) );
  INV_X1 U13312 ( .A(n14624), .ZN(n15730) );
  NAND2_X1 U13313 ( .A1(n15730), .A2(n14742), .ZN(n11490) );
  NAND2_X1 U13314 ( .A1(n11555), .A2(n11490), .ZN(n11492) );
  NAND2_X1 U13315 ( .A1(n14624), .A2(n11505), .ZN(n11491) );
  NAND3_X1 U13316 ( .A1(n11495), .A2(n11494), .A3(n11879), .ZN(n12892) );
  INV_X1 U13317 ( .A(n11496), .ZN(n11498) );
  INV_X1 U13318 ( .A(n15083), .ZN(n15052) );
  AND2_X1 U13319 ( .A1(n14746), .A2(n11499), .ZN(n11621) );
  INV_X1 U13320 ( .A(n11500), .ZN(n11501) );
  NAND2_X1 U13321 ( .A1(n11835), .A2(n11834), .ZN(n11504) );
  OR2_X1 U13322 ( .A1(n7476), .A2(n14743), .ZN(n11503) );
  INV_X1 U13323 ( .A(n11554), .ZN(n11553) );
  NAND2_X1 U13324 ( .A1(n15730), .A2(n11505), .ZN(n11506) );
  XNOR2_X1 U13325 ( .A(n11524), .B(n11507), .ZN(n15751) );
  INV_X1 U13326 ( .A(n11508), .ZN(n12090) );
  INV_X1 U13327 ( .A(n15069), .ZN(n15088) );
  NAND2_X1 U13328 ( .A1(n15751), .A2(n15088), .ZN(n11523) );
  AND2_X1 U13329 ( .A1(n15670), .A2(n11617), .ZN(n11846) );
  INV_X1 U13330 ( .A(n11541), .ZN(n11542) );
  AOI21_X1 U13331 ( .B1(n11531), .B2(n11559), .A(n15731), .ZN(n11510) );
  NAND2_X1 U13332 ( .A1(n11542), .A2(n11510), .ZN(n15745) );
  INV_X1 U13333 ( .A(n15745), .ZN(n11521) );
  NOR2_X1 U13334 ( .A1(n11511), .A2(n12485), .ZN(n11512) );
  OR2_X1 U13335 ( .A1(n11686), .A2(n15042), .ZN(n11514) );
  NAND2_X1 U13336 ( .A1(n14742), .A2(n15075), .ZN(n11513) );
  AND2_X1 U13337 ( .A1(n11514), .A2(n11513), .ZN(n15744) );
  INV_X1 U13338 ( .A(n15744), .ZN(n11516) );
  INV_X1 U13339 ( .A(n11515), .ZN(n11580) );
  INV_X1 U13340 ( .A(n15660), .ZN(n15043) );
  AOI22_X1 U13341 ( .A1(n15021), .A2(n11516), .B1(n11580), .B2(n15043), .ZN(
        n11519) );
  OR2_X1 U13342 ( .A1(n15021), .A2(n11517), .ZN(n11518) );
  OAI211_X1 U13343 ( .C1(n15078), .C2(n15746), .A(n11519), .B(n11518), .ZN(
        n11520) );
  AOI21_X1 U13344 ( .B1(n15049), .B2(n11521), .A(n11520), .ZN(n11522) );
  OAI211_X1 U13345 ( .C1(n15748), .C2(n15052), .A(n11523), .B(n11522), .ZN(
        P1_U3289) );
  NAND2_X1 U13346 ( .A1(n11527), .A2(n11526), .ZN(n11528) );
  INV_X1 U13347 ( .A(n11534), .ZN(n11680) );
  NAND2_X1 U13348 ( .A1(n11528), .A2(n11680), .ZN(n11529) );
  NAND2_X1 U13349 ( .A1(n11678), .A2(n11529), .ZN(n11536) );
  INV_X1 U13350 ( .A(n11536), .ZN(n15774) );
  INV_X1 U13351 ( .A(n11530), .ZN(n15664) );
  AND2_X1 U13352 ( .A1(n15021), .A2(n15664), .ZN(n15034) );
  AND2_X1 U13353 ( .A1(n11531), .A2(n11532), .ZN(n11533) );
  XNOR2_X1 U13354 ( .A(n11681), .B(n11534), .ZN(n11535) );
  NAND2_X1 U13355 ( .A1(n11535), .A2(n15993), .ZN(n11539) );
  NAND2_X1 U13356 ( .A1(n11536), .A2(n15025), .ZN(n11538) );
  AOI22_X1 U13357 ( .A1(n11704), .A2(n15076), .B1(n15075), .B2(n14741), .ZN(
        n11537) );
  NAND3_X1 U13358 ( .A1(n11539), .A2(n11538), .A3(n11537), .ZN(n15777) );
  MUX2_X1 U13359 ( .A(n15777), .B(P1_REG2_REG_5__SCAN_IN), .S(n15667), .Z(
        n11540) );
  INV_X1 U13360 ( .A(n11540), .ZN(n11547) );
  INV_X1 U13361 ( .A(n11543), .ZN(n11682) );
  AOI211_X1 U13362 ( .C1(n11543), .C2(n11542), .A(n15731), .B(n7333), .ZN(
        n15775) );
  OAI22_X1 U13363 ( .A1(n15078), .A2(n11682), .B1(n15660), .B2(n11544), .ZN(
        n11545) );
  AOI21_X1 U13364 ( .B1(n15775), .B2(n15049), .A(n11545), .ZN(n11546) );
  OAI211_X1 U13365 ( .C1(n15774), .C2(n12432), .A(n11547), .B(n11546), .ZN(
        P1_U3288) );
  INV_X1 U13366 ( .A(n11548), .ZN(n11551) );
  OAI222_X1 U13367 ( .A1(n14592), .A2(n11549), .B1(n14578), .B2(n11551), .C1(
        n15289), .C2(P2_U3088), .ZN(P2_U3312) );
  OAI222_X1 U13368 ( .A1(P1_U3086), .A2(n14824), .B1(n15233), .B2(n11551), 
        .C1(n11550), .C2(n15224), .ZN(P1_U3340) );
  XNOR2_X1 U13369 ( .A(n11553), .B(n11552), .ZN(n15735) );
  INV_X1 U13370 ( .A(n15735), .ZN(n11564) );
  XNOR2_X1 U13371 ( .A(n11555), .B(n11554), .ZN(n11556) );
  NAND2_X1 U13372 ( .A1(n11556), .A2(n15993), .ZN(n11558) );
  AOI22_X1 U13373 ( .A1(n15075), .A2(n14743), .B1(n14741), .B2(n15076), .ZN(
        n11557) );
  NAND2_X1 U13374 ( .A1(n11558), .A2(n11557), .ZN(n15733) );
  INV_X1 U13375 ( .A(n11845), .ZN(n11560) );
  OAI21_X1 U13376 ( .B1(n15730), .B2(n11560), .A(n11559), .ZN(n15732) );
  OAI22_X1 U13377 ( .A1(n15732), .A2(n15063), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15660), .ZN(n11561) );
  OAI21_X1 U13378 ( .B1(n15733), .B2(n11561), .A(n15021), .ZN(n11563) );
  AOI22_X1 U13379 ( .A1(n15066), .A2(n14624), .B1(n15667), .B2(
        P1_REG2_REG_3__SCAN_IN), .ZN(n11562) );
  OAI211_X1 U13380 ( .C1(n15069), .C2(n11564), .A(n11563), .B(n11562), .ZN(
        P1_U3290) );
  INV_X1 U13381 ( .A(n14558), .ZN(n14553) );
  INV_X1 U13382 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11565) );
  NOR2_X1 U13383 ( .A1(n15973), .A2(n11565), .ZN(n11566) );
  AOI21_X1 U13384 ( .B1(n15973), .B2(n11567), .A(n11566), .ZN(n11568) );
  OAI21_X1 U13385 ( .B1(n11569), .B2(n14553), .A(n11568), .ZN(P2_U3433) );
  OAI222_X1 U13386 ( .A1(P1_U3086), .A2(n14827), .B1(n15233), .B2(n11572), 
        .C1(n11570), .C2(n15224), .ZN(P1_U3339) );
  INV_X1 U13387 ( .A(n15308), .ZN(n11571) );
  OAI222_X1 U13388 ( .A1(n14592), .A2(n11573), .B1(n14578), .B2(n11572), .C1(
        n11571), .C2(P2_U3088), .ZN(P2_U3311) );
  OAI21_X1 U13389 ( .B1(n11576), .B2(n11575), .A(n11574), .ZN(n11577) );
  NAND2_X1 U13390 ( .A1(n11577), .A2(n16010), .ZN(n11582) );
  INV_X1 U13391 ( .A(n16011), .ZN(n14689) );
  OAI21_X1 U13392 ( .B1(n14689), .B2(n15744), .A(n11578), .ZN(n11579) );
  AOI21_X1 U13393 ( .B1(n11580), .B2(n14721), .A(n11579), .ZN(n11581) );
  OAI211_X1 U13394 ( .C1(n15746), .C2(n15982), .A(n11582), .B(n11581), .ZN(
        P1_U3230) );
  NOR2_X1 U13395 ( .A1(n7209), .A2(n11595), .ZN(n11587) );
  XNOR2_X1 U13396 ( .A(n15831), .B(n14072), .ZN(n11594) );
  INV_X1 U13397 ( .A(n11594), .ZN(n11586) );
  XNOR2_X1 U13398 ( .A(n11594), .B(n11587), .ZN(n11815) );
  INV_X1 U13399 ( .A(n11583), .ZN(n11584) );
  NAND3_X1 U13400 ( .A1(n11585), .A2(n11815), .A3(n11584), .ZN(n11810) );
  OAI21_X1 U13401 ( .B1(n11587), .B2(n11586), .A(n11810), .ZN(n11588) );
  XNOR2_X1 U13402 ( .A(n11654), .B(n14072), .ZN(n11984) );
  NOR2_X1 U13403 ( .A1(n7209), .A2(n11637), .ZN(n11986) );
  XNOR2_X1 U13404 ( .A(n11984), .B(n11986), .ZN(n11593) );
  NAND2_X1 U13405 ( .A1(n11588), .A2(n11593), .ZN(n11985) );
  NOR2_X1 U13406 ( .A1(n14092), .A2(n11649), .ZN(n11592) );
  NAND2_X1 U13407 ( .A1(n14153), .A2(n14185), .ZN(n11590) );
  NAND2_X1 U13408 ( .A1(n14152), .A2(n14188), .ZN(n11589) );
  AND2_X1 U13409 ( .A1(n11590), .A2(n11589), .ZN(n11647) );
  NAND2_X1 U13410 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14237) );
  OAI21_X1 U13411 ( .B1(n14157), .B2(n11647), .A(n14237), .ZN(n11591) );
  AOI211_X1 U13412 ( .C1(n11654), .C2(n14159), .A(n11592), .B(n11591), .ZN(
        n11599) );
  INV_X1 U13413 ( .A(n11593), .ZN(n11597) );
  OAI22_X1 U13414 ( .A1(n11595), .A2(n14146), .B1(n11594), .B2(n14163), .ZN(
        n11596) );
  NAND3_X1 U13415 ( .A1(n11810), .A2(n11597), .A3(n11596), .ZN(n11598) );
  OAI211_X1 U13416 ( .C1(n11985), .C2(n14163), .A(n11599), .B(n11598), .ZN(
        P2_U3193) );
  OAI22_X1 U13417 ( .A1(n15721), .A2(n11601), .B1(n11600), .B2(n15714), .ZN(
        n11604) );
  NOR2_X1 U13418 ( .A1(n15940), .A2(n11602), .ZN(n11603) );
  AOI211_X1 U13419 ( .C1(n11605), .C2(n15934), .A(n11604), .B(n11603), .ZN(
        n11609) );
  NAND2_X1 U13420 ( .A1(n14423), .A2(n11606), .ZN(n15713) );
  OR2_X1 U13421 ( .A1(n11607), .A2(n14369), .ZN(n11608) );
  OAI211_X1 U13422 ( .C1(n15947), .C2(n11610), .A(n11609), .B(n11608), .ZN(
        P2_U3260) );
  OAI21_X1 U13423 ( .B1(n11612), .B2(n11502), .A(n11611), .ZN(n11613) );
  NAND2_X1 U13424 ( .A1(n11613), .A2(n15993), .ZN(n11615) );
  AOI22_X1 U13425 ( .A1(n15075), .A2(n14746), .B1(n14743), .B2(n15076), .ZN(
        n11614) );
  AND2_X1 U13426 ( .A1(n11615), .A2(n11614), .ZN(n15669) );
  OAI22_X1 U13427 ( .A1(n15021), .A2(n10880), .B1(n11616), .B2(n15660), .ZN(
        n11620) );
  OAI21_X1 U13428 ( .B1(n15670), .B2(n11617), .A(n15071), .ZN(n11618) );
  OR2_X1 U13429 ( .A1(n11846), .A2(n11618), .ZN(n15668) );
  NOR2_X1 U13430 ( .A1(n15086), .A2(n15668), .ZN(n11619) );
  AOI211_X1 U13431 ( .C1(n15066), .C2(n9710), .A(n11620), .B(n11619), .ZN(
        n11624) );
  AOI21_X1 U13432 ( .B1(n15025), .B2(n15021), .A(n15034), .ZN(n14897) );
  INV_X1 U13433 ( .A(n14897), .ZN(n11622) );
  XOR2_X1 U13434 ( .A(n11621), .B(n11502), .Z(n15672) );
  INV_X1 U13435 ( .A(n15672), .ZN(n15675) );
  NAND2_X1 U13436 ( .A1(n11622), .A2(n15675), .ZN(n11623) );
  OAI211_X1 U13437 ( .C1(n15667), .C2(n15669), .A(n11624), .B(n11623), .ZN(
        P1_U3292) );
  MUX2_X1 U13438 ( .A(n11625), .B(P2_REG2_REG_3__SCAN_IN), .S(n15947), .Z(
        n11629) );
  AOI22_X1 U13439 ( .A1(n15934), .A2(n11626), .B1(n15936), .B2(n14207), .ZN(
        n11627) );
  OAI21_X1 U13440 ( .B1(n11782), .B2(n15940), .A(n11627), .ZN(n11628) );
  AOI211_X1 U13441 ( .C1(n15944), .C2(n11630), .A(n11629), .B(n11628), .ZN(
        n11631) );
  INV_X1 U13442 ( .A(n11631), .ZN(P2_U3262) );
  INV_X1 U13443 ( .A(n11633), .ZN(n11634) );
  XNOR2_X1 U13444 ( .A(n11632), .B(n11634), .ZN(n15835) );
  XNOR2_X1 U13445 ( .A(n11635), .B(n11634), .ZN(n11638) );
  NAND2_X1 U13446 ( .A1(n14152), .A2(n14189), .ZN(n11636) );
  OAI21_X1 U13447 ( .B1(n11637), .B2(n11977), .A(n11636), .ZN(n11806) );
  AOI21_X1 U13448 ( .B1(n11638), .B2(n15797), .A(n11806), .ZN(n15838) );
  MUX2_X1 U13449 ( .A(n11256), .B(n15838), .S(n15721), .Z(n11644) );
  NAND2_X1 U13450 ( .A1(n15804), .A2(n15831), .ZN(n11639) );
  NAND2_X1 U13451 ( .A1(n11639), .A2(n7209), .ZN(n11640) );
  NOR2_X1 U13452 ( .A1(n11651), .A2(n11640), .ZN(n15833) );
  INV_X1 U13453 ( .A(n15831), .ZN(n11641) );
  OAI22_X1 U13454 ( .A1(n15940), .A2(n11641), .B1(n11809), .B2(n15714), .ZN(
        n11642) );
  AOI21_X1 U13455 ( .B1(n15833), .B2(n15934), .A(n11642), .ZN(n11643) );
  OAI211_X1 U13456 ( .C1(n14369), .C2(n15835), .A(n11644), .B(n11643), .ZN(
        P2_U3258) );
  INV_X1 U13457 ( .A(n11668), .ZN(n11645) );
  AOI21_X1 U13458 ( .B1(n9111), .B2(n11646), .A(n11645), .ZN(n11648) );
  OAI21_X1 U13459 ( .B1(n11648), .B2(n15702), .A(n11647), .ZN(n15854) );
  INV_X1 U13460 ( .A(n15854), .ZN(n11659) );
  OAI22_X1 U13461 ( .A1(n15721), .A2(n11650), .B1(n11649), .B2(n15714), .ZN(
        n11653) );
  OAI211_X1 U13462 ( .C1(n11651), .C2(n15852), .A(n14308), .B(n11663), .ZN(
        n15849) );
  NOR2_X1 U13463 ( .A1(n15849), .A2(n15717), .ZN(n11652) );
  AOI211_X1 U13464 ( .C1(n15917), .C2(n11654), .A(n11653), .B(n11652), .ZN(
        n11658) );
  NAND2_X1 U13465 ( .A1(n11655), .A2(n11656), .ZN(n15847) );
  NAND3_X1 U13466 ( .A1(n15848), .A2(n15847), .A3(n15807), .ZN(n11657) );
  OAI211_X1 U13467 ( .C1(n11659), .C2(n15947), .A(n11658), .B(n11657), .ZN(
        P2_U3257) );
  OR2_X1 U13468 ( .A1(n11669), .A2(n11660), .ZN(n11661) );
  NAND2_X1 U13469 ( .A1(n11662), .A2(n11661), .ZN(n11955) );
  AOI211_X1 U13470 ( .C1(n11998), .C2(n11663), .A(n14360), .B(n11794), .ZN(
        n11957) );
  INV_X1 U13471 ( .A(n11998), .ZN(n11664) );
  NOR2_X1 U13472 ( .A1(n11664), .A2(n15940), .ZN(n11666) );
  INV_X1 U13473 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11912) );
  OAI22_X1 U13474 ( .A1(n15721), .A2(n11912), .B1(n11991), .B2(n15714), .ZN(
        n11665) );
  AOI211_X1 U13475 ( .C1(n11957), .C2(n15934), .A(n11666), .B(n11665), .ZN(
        n11676) );
  NAND3_X1 U13476 ( .A1(n11669), .A2(n11668), .A3(n11667), .ZN(n11671) );
  AOI21_X1 U13477 ( .B1(n11671), .B2(n11670), .A(n15702), .ZN(n11673) );
  NAND2_X1 U13478 ( .A1(n14152), .A2(n14187), .ZN(n11672) );
  OAI21_X1 U13479 ( .B1(n12038), .B2(n11977), .A(n11672), .ZN(n11988) );
  NOR2_X1 U13480 ( .A1(n11673), .A2(n11988), .ZN(n11674) );
  OAI21_X1 U13481 ( .B1(n14423), .B2(n11955), .A(n11674), .ZN(n11956) );
  NAND2_X1 U13482 ( .A1(n11956), .A2(n15721), .ZN(n11675) );
  OAI211_X1 U13483 ( .C1(n11955), .C2(n14431), .A(n11676), .B(n11675), .ZN(
        P2_U3256) );
  NAND2_X1 U13484 ( .A1(n11682), .A2(n11686), .ZN(n11677) );
  OAI21_X1 U13485 ( .B1(n11679), .B2(n11685), .A(n11699), .ZN(n15792) );
  INV_X1 U13486 ( .A(n15792), .ZN(n11697) );
  NAND2_X1 U13487 ( .A1(n11681), .A2(n11680), .ZN(n11684) );
  NAND2_X1 U13488 ( .A1(n11682), .A2(n14740), .ZN(n11683) );
  INV_X1 U13489 ( .A(n11685), .ZN(n11702) );
  XNOR2_X1 U13490 ( .A(n11703), .B(n11702), .ZN(n11689) );
  INV_X1 U13491 ( .A(n14739), .ZN(n11857) );
  OAI22_X1 U13492 ( .A1(n11857), .A2(n15042), .B1(n11686), .B2(n15041), .ZN(
        n11687) );
  AOI21_X1 U13493 ( .B1(n15792), .B2(n15025), .A(n11687), .ZN(n11688) );
  OAI21_X1 U13494 ( .B1(n15747), .B2(n11689), .A(n11688), .ZN(n15790) );
  NAND2_X1 U13495 ( .A1(n15790), .A2(n15021), .ZN(n11696) );
  OAI22_X1 U13496 ( .A1(n15021), .A2(n11691), .B1(n11690), .B2(n15660), .ZN(
        n11693) );
  INV_X1 U13497 ( .A(n11694), .ZN(n11705) );
  OAI211_X1 U13498 ( .C1(n7333), .C2(n11705), .A(n15071), .B(n11715), .ZN(
        n15789) );
  NOR2_X1 U13499 ( .A1(n15789), .A2(n15086), .ZN(n11692) );
  AOI211_X1 U13500 ( .C1(n15066), .C2(n11694), .A(n11693), .B(n11692), .ZN(
        n11695) );
  OAI211_X1 U13501 ( .C1(n11697), .C2(n12432), .A(n11696), .B(n11695), .ZN(
        P1_U3287) );
  NAND2_X1 U13502 ( .A1(n11705), .A2(n11709), .ZN(n11698) );
  NAND2_X1 U13503 ( .A1(n11699), .A2(n11698), .ZN(n11701) );
  INV_X1 U13504 ( .A(n11708), .ZN(n11700) );
  NAND2_X1 U13505 ( .A1(n11701), .A2(n11700), .ZN(n11853) );
  OAI21_X1 U13506 ( .B1(n11701), .B2(n11700), .A(n11853), .ZN(n15828) );
  INV_X1 U13507 ( .A(n15828), .ZN(n11721) );
  NAND2_X1 U13508 ( .A1(n11703), .A2(n11702), .ZN(n11707) );
  NAND2_X1 U13509 ( .A1(n11705), .A2(n11704), .ZN(n11706) );
  XNOR2_X1 U13510 ( .A(n11861), .B(n11708), .ZN(n11712) );
  INV_X1 U13511 ( .A(n14738), .ZN(n12000) );
  OAI22_X1 U13512 ( .A1(n12000), .A2(n15042), .B1(n11709), .B2(n15041), .ZN(
        n11710) );
  AOI21_X1 U13513 ( .B1(n15828), .B2(n15025), .A(n11710), .ZN(n11711) );
  OAI21_X1 U13514 ( .B1(n15747), .B2(n11712), .A(n11711), .ZN(n15826) );
  NAND2_X1 U13515 ( .A1(n15826), .A2(n15021), .ZN(n11720) );
  OAI22_X1 U13516 ( .A1(n15021), .A2(n11714), .B1(n11713), .B2(n15660), .ZN(
        n11718) );
  INV_X1 U13517 ( .A(n11715), .ZN(n11716) );
  INV_X1 U13518 ( .A(n11867), .ZN(n11868) );
  OAI211_X1 U13519 ( .C1(n7583), .C2(n11716), .A(n11868), .B(n15071), .ZN(
        n15825) );
  NOR2_X1 U13520 ( .A1(n15825), .A2(n15086), .ZN(n11717) );
  AOI211_X1 U13521 ( .C1(n15066), .C2(n11858), .A(n11718), .B(n11717), .ZN(
        n11719) );
  OAI211_X1 U13522 ( .C1(n11721), .C2(n12432), .A(n11720), .B(n11719), .ZN(
        P1_U3286) );
  NAND2_X1 U13523 ( .A1(n13221), .A2(n11722), .ZN(n11723) );
  XNOR2_X1 U13524 ( .A(n15737), .B(n13041), .ZN(n11725) );
  NAND2_X1 U13525 ( .A1(n12235), .A2(n11725), .ZN(n11902) );
  INV_X1 U13526 ( .A(n11725), .ZN(n11726) );
  NAND2_X1 U13527 ( .A1(n11726), .A2(n13220), .ZN(n11727) );
  NAND2_X1 U13528 ( .A1(n11902), .A2(n11727), .ZN(n11729) );
  INV_X1 U13529 ( .A(n11903), .ZN(n11728) );
  AOI21_X1 U13530 ( .B1(n11730), .B2(n11729), .A(n11728), .ZN(n11735) );
  OAI22_X1 U13531 ( .A1(n13195), .A2(n8398), .B1(n12217), .B2(n13174), .ZN(
        n11731) );
  AOI211_X1 U13532 ( .C1(n13197), .C2(n12082), .A(n11732), .B(n11731), .ZN(
        n11734) );
  NAND2_X1 U13533 ( .A1(n13190), .A2(n12081), .ZN(n11733) );
  OAI211_X1 U13534 ( .C1(n11735), .C2(n13200), .A(n11734), .B(n11733), .ZN(
        P3_U3170) );
  OAI21_X1 U13535 ( .B1(n11737), .B2(n10306), .A(n11826), .ZN(n11743) );
  OAI22_X1 U13536 ( .A1(n11738), .A2(n13627), .B1(n7398), .B2(n13629), .ZN(
        n11742) );
  XNOR2_X1 U13537 ( .A(n11740), .B(n11739), .ZN(n11945) );
  NOR2_X1 U13538 ( .A1(n11945), .A2(n15764), .ZN(n11741) );
  AOI211_X1 U13539 ( .C1(n13604), .C2(n11743), .A(n11742), .B(n11741), .ZN(
        n11939) );
  INV_X1 U13540 ( .A(n11945), .ZN(n11750) );
  INV_X1 U13541 ( .A(n15873), .ZN(n15858) );
  INV_X1 U13542 ( .A(n13749), .ZN(n11746) );
  INV_X1 U13543 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n11744) );
  OAI22_X1 U13544 ( .A1(n7432), .A2(n13767), .B1(n15898), .B2(n11744), .ZN(
        n11745) );
  AOI21_X1 U13545 ( .B1(n11750), .B2(n11746), .A(n11745), .ZN(n11747) );
  OAI21_X1 U13546 ( .B1(n11939), .B2(n15895), .A(n11747), .ZN(P3_U3393) );
  NAND2_X1 U13547 ( .A1(n15894), .A2(n15873), .ZN(n13673) );
  INV_X1 U13548 ( .A(n13673), .ZN(n15766) );
  OAI22_X1 U13549 ( .A1(n13694), .A2(n7432), .B1(n15894), .B2(n11748), .ZN(
        n11749) );
  AOI21_X1 U13550 ( .B1(n11750), .B2(n15766), .A(n11749), .ZN(n11751) );
  OAI21_X1 U13551 ( .B1(n11939), .B2(n15892), .A(n11751), .ZN(P3_U3460) );
  INV_X1 U13552 ( .A(n13240), .ZN(n11752) );
  INV_X1 U13553 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n12224) );
  MUX2_X1 U13554 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n12224), .S(n13236), .Z(
        n13238) );
  INV_X1 U13555 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15612) );
  XNOR2_X1 U13556 ( .A(n15617), .B(n11753), .ZN(n15611) );
  INV_X1 U13557 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12309) );
  MUX2_X1 U13558 ( .A(n12309), .B(P3_REG2_REG_8__SCAN_IN), .S(n12174), .Z(
        n11755) );
  INV_X1 U13559 ( .A(n12155), .ZN(n11754) );
  AOI21_X1 U13560 ( .B1(n11756), .B2(n11755), .A(n11754), .ZN(n11780) );
  INV_X1 U13561 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11772) );
  MUX2_X1 U13562 ( .A(n12309), .B(n11772), .S(n7165), .Z(n12169) );
  XNOR2_X1 U13563 ( .A(n12169), .B(n12174), .ZN(n11766) );
  MUX2_X1 U13564 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n7206), .Z(n11758) );
  OR2_X1 U13565 ( .A1(n11758), .A2(n11757), .ZN(n11764) );
  XNOR2_X1 U13566 ( .A(n11758), .B(n15617), .ZN(n15614) );
  MUX2_X1 U13567 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n7166), .Z(n11763) );
  XNOR2_X1 U13568 ( .A(n11763), .B(n13236), .ZN(n13226) );
  OAI22_X1 U13569 ( .A1(n11762), .A2(n11761), .B1(n11760), .B2(n11759), .ZN(
        n13227) );
  NAND2_X1 U13570 ( .A1(n13226), .A2(n13227), .ZN(n13225) );
  OAI21_X1 U13571 ( .B1(n11763), .B2(n11769), .A(n13225), .ZN(n15615) );
  NAND2_X1 U13572 ( .A1(n15614), .A2(n15615), .ZN(n15613) );
  OAI21_X1 U13573 ( .B1(n11766), .B2(n11765), .A(n12166), .ZN(n11778) );
  NOR2_X1 U13574 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13857), .ZN(n12248) );
  AOI21_X1 U13575 ( .B1(n15246), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12248), .ZN(
        n11767) );
  OAI21_X1 U13576 ( .B1(n15641), .B2(n12174), .A(n11767), .ZN(n11777) );
  INV_X1 U13577 ( .A(n11768), .ZN(n13230) );
  INV_X1 U13578 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15785) );
  MUX2_X1 U13579 ( .A(n15785), .B(P3_REG1_REG_6__SCAN_IN), .S(n13236), .Z(
        n13229) );
  NOR2_X1 U13580 ( .A1(n15617), .A2(n11770), .ZN(n11771) );
  INV_X1 U13581 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15822) );
  NOR2_X1 U13582 ( .A1(n11771), .A2(n15621), .ZN(n11774) );
  MUX2_X1 U13583 ( .A(n11772), .B(P3_REG1_REG_8__SCAN_IN), .S(n12174), .Z(
        n11773) );
  OR2_X2 U13584 ( .A1(n11774), .A2(n11773), .ZN(n12176) );
  NAND2_X1 U13585 ( .A1(n11774), .A2(n11773), .ZN(n11775) );
  AOI21_X1 U13586 ( .B1(n12176), .B2(n11775), .A(n15631), .ZN(n11776) );
  AOI211_X1 U13587 ( .C1(n15638), .C2(n11778), .A(n11777), .B(n11776), .ZN(
        n11779) );
  OAI21_X1 U13588 ( .B1(n11780), .B2(n15636), .A(n11779), .ZN(P3_U3190) );
  INV_X1 U13589 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11781) );
  OAI22_X1 U13590 ( .A1(n14553), .A2(n11782), .B1(n15973), .B2(n11781), .ZN(
        n11783) );
  INV_X1 U13591 ( .A(n11783), .ZN(n11784) );
  OAI21_X1 U13592 ( .B1(n11785), .B2(n15971), .A(n11784), .ZN(P2_U3439) );
  INV_X1 U13593 ( .A(n11786), .ZN(n11788) );
  INV_X1 U13594 ( .A(SI_20_), .ZN(n13896) );
  OAI222_X1 U13595 ( .A1(n13993), .A2(n11788), .B1(n13995), .B2(n13896), .C1(
        P3_U3151), .C2(n11787), .ZN(P3_U3275) );
  XNOR2_X1 U13596 ( .A(n11789), .B(n11793), .ZN(n11791) );
  OAI22_X1 U13597 ( .A1(n11790), .A2(n12044), .B1(n12280), .B2(n11977), .ZN(
        n12039) );
  AOI21_X1 U13598 ( .B1(n11791), .B2(n15797), .A(n12039), .ZN(n11947) );
  XOR2_X1 U13599 ( .A(n11793), .B(n11792), .Z(n11948) );
  INV_X1 U13600 ( .A(n11948), .ZN(n11800) );
  INV_X1 U13601 ( .A(n11794), .ZN(n11795) );
  AOI21_X1 U13602 ( .B1(n11795), .B2(n12043), .A(n14360), .ZN(n11796) );
  NAND2_X1 U13603 ( .A1(n11796), .A2(n11979), .ZN(n11946) );
  INV_X1 U13604 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11916) );
  OAI22_X1 U13605 ( .A1(n15721), .A2(n11916), .B1(n12041), .B2(n15714), .ZN(
        n11797) );
  AOI21_X1 U13606 ( .B1(n12043), .B2(n15917), .A(n11797), .ZN(n11798) );
  OAI21_X1 U13607 ( .B1(n11946), .B2(n15717), .A(n11798), .ZN(n11799) );
  AOI21_X1 U13608 ( .B1(n11800), .B2(n15807), .A(n11799), .ZN(n11801) );
  OAI21_X1 U13609 ( .B1(n15947), .B2(n11947), .A(n11801), .ZN(P2_U3255) );
  INV_X1 U13610 ( .A(n11585), .ZN(n11805) );
  NOR3_X1 U13611 ( .A1(n14146), .A2(n11803), .A3(n11802), .ZN(n11804) );
  AOI21_X1 U13612 ( .B1(n11805), .B2(n14102), .A(n11804), .ZN(n11814) );
  NAND2_X1 U13613 ( .A1(n14095), .A2(n11806), .ZN(n11808) );
  NAND2_X1 U13614 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n11807) );
  OAI211_X1 U13615 ( .C1(n14092), .C2(n11809), .A(n11808), .B(n11807), .ZN(
        n11812) );
  NOR2_X1 U13616 ( .A1(n11810), .A2(n14163), .ZN(n11811) );
  AOI211_X1 U13617 ( .C1(n15831), .C2(n14159), .A(n11812), .B(n11811), .ZN(
        n11813) );
  OAI21_X1 U13618 ( .B1(n11815), .B2(n11814), .A(n11813), .ZN(P2_U3185) );
  INV_X1 U13619 ( .A(n11816), .ZN(n11817) );
  AOI21_X1 U13620 ( .B1(n11819), .B2(n11818), .A(n11817), .ZN(n15679) );
  AND2_X1 U13621 ( .A1(n11821), .A2(n11820), .ZN(n11822) );
  AND2_X1 U13622 ( .A1(n13565), .A2(n11822), .ZN(n12467) );
  AOI22_X1 U13623 ( .A1(n13609), .A2(n11371), .B1(n13221), .B2(n13606), .ZN(
        n11830) );
  INV_X1 U13624 ( .A(n11824), .ZN(n11828) );
  AND3_X1 U13625 ( .A1(n11826), .A2(n8773), .A3(n11825), .ZN(n11827) );
  OAI21_X1 U13626 ( .B1(n11828), .B2(n11827), .A(n13604), .ZN(n11829) );
  OAI211_X1 U13627 ( .C1(n15679), .C2(n15764), .A(n11830), .B(n11829), .ZN(
        n15681) );
  OAI22_X1 U13628 ( .A1(n15678), .A2(n11940), .B1(n13878), .B2(n13520), .ZN(
        n11831) );
  NOR2_X1 U13629 ( .A1(n15681), .A2(n11831), .ZN(n11832) );
  MUX2_X1 U13630 ( .A(n11045), .B(n11832), .S(n13565), .Z(n11833) );
  OAI21_X1 U13631 ( .B1(n15679), .B2(n13571), .A(n11833), .ZN(P3_U3231) );
  XNOR2_X1 U13632 ( .A(n11835), .B(n11834), .ZN(n15688) );
  NAND2_X1 U13633 ( .A1(n15688), .A2(n15025), .ZN(n11844) );
  OAI21_X1 U13634 ( .B1(n11838), .B2(n11837), .A(n11836), .ZN(n11842) );
  NAND2_X1 U13635 ( .A1(n14744), .A2(n15075), .ZN(n11840) );
  NAND2_X1 U13636 ( .A1(n14742), .A2(n15076), .ZN(n11839) );
  NAND2_X1 U13637 ( .A1(n11840), .A2(n11839), .ZN(n11841) );
  AOI21_X1 U13638 ( .B1(n11842), .B2(n15993), .A(n11841), .ZN(n11843) );
  AND2_X1 U13639 ( .A1(n11844), .A2(n11843), .ZN(n15690) );
  OAI211_X1 U13640 ( .C1(n15686), .C2(n11846), .A(n15071), .B(n11845), .ZN(
        n15685) );
  OAI22_X1 U13641 ( .A1(n15021), .A2(n10882), .B1(n11847), .B2(n15660), .ZN(
        n11848) );
  AOI21_X1 U13642 ( .B1(n15066), .B2(n7476), .A(n11848), .ZN(n11849) );
  OAI21_X1 U13643 ( .B1(n15086), .B2(n15685), .A(n11849), .ZN(n11850) );
  AOI21_X1 U13644 ( .B1(n15034), .B2(n15688), .A(n11850), .ZN(n11851) );
  OAI21_X1 U13645 ( .B1(n15667), .B2(n15690), .A(n11851), .ZN(P1_U3291) );
  OR2_X1 U13646 ( .A1(n11858), .A2(n14739), .ZN(n11852) );
  NAND2_X1 U13647 ( .A1(n11853), .A2(n11852), .ZN(n11855) );
  NAND2_X1 U13648 ( .A1(n11855), .A2(n11863), .ZN(n12002) );
  OAI21_X1 U13649 ( .B1(n11855), .B2(n11863), .A(n12002), .ZN(n11856) );
  INV_X1 U13650 ( .A(n11856), .ZN(n11877) );
  NOR2_X1 U13651 ( .A1(n11858), .A2(n11857), .ZN(n11860) );
  NAND2_X1 U13652 ( .A1(n11858), .A2(n11857), .ZN(n11859) );
  AOI21_X1 U13653 ( .B1(n11862), .B2(n11863), .A(n15747), .ZN(n11864) );
  AOI22_X1 U13654 ( .A1(n11864), .A2(n12005), .B1(n15075), .B2(n14739), .ZN(
        n11875) );
  AND2_X1 U13655 ( .A1(n14737), .A2(n15076), .ZN(n11874) );
  INV_X1 U13656 ( .A(n11874), .ZN(n11865) );
  OAI211_X1 U13657 ( .C1(n15660), .C2(n12206), .A(n11875), .B(n11865), .ZN(
        n11866) );
  NAND2_X1 U13658 ( .A1(n11866), .A2(n15021), .ZN(n11872) );
  INV_X1 U13659 ( .A(n12013), .ZN(n12015) );
  AOI211_X1 U13660 ( .C1(n12198), .C2(n11868), .A(n15731), .B(n12015), .ZN(
        n11873) );
  OAI22_X1 U13661 ( .A1(n12213), .A2(n15078), .B1(n15021), .B2(n11869), .ZN(
        n11870) );
  AOI21_X1 U13662 ( .B1(n11873), .B2(n15049), .A(n11870), .ZN(n11871) );
  OAI211_X1 U13663 ( .C1(n14897), .C2(n11877), .A(n11872), .B(n11871), .ZN(
        P1_U3285) );
  INV_X1 U13664 ( .A(n15912), .ZN(n15773) );
  AOI211_X1 U13665 ( .C1(n15949), .C2(n12198), .A(n11874), .B(n11873), .ZN(
        n11876) );
  OAI211_X1 U13666 ( .C1(n15953), .C2(n11877), .A(n11876), .B(n11875), .ZN(
        n11881) );
  NAND2_X1 U13667 ( .A1(n11881), .A2(n16001), .ZN(n11878) );
  OAI21_X1 U13668 ( .B1(n16001), .B2(n10898), .A(n11878), .ZN(P1_U3536) );
  INV_X1 U13669 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11883) );
  NAND2_X1 U13670 ( .A1(n11881), .A2(n16005), .ZN(n11882) );
  OAI21_X1 U13671 ( .B1(n16005), .B2(n11883), .A(n11882), .ZN(P1_U3483) );
  INV_X1 U13672 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n15931) );
  MUX2_X1 U13673 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15931), .S(n11893), .Z(
        n14807) );
  NAND2_X1 U13674 ( .A1(n14808), .A2(n14807), .ZN(n14806) );
  OAI21_X1 U13675 ( .B1(n14811), .B2(n15931), .A(n14806), .ZN(n14822) );
  XNOR2_X1 U13676 ( .A(n14822), .B(n14823), .ZN(n11887) );
  INV_X1 U13677 ( .A(n11887), .ZN(n11886) );
  OAI21_X1 U13678 ( .B1(n11886), .B2(P1_REG1_REG_14__SCAN_IN), .A(n15427), 
        .ZN(n11899) );
  NOR2_X1 U13679 ( .A1(n11887), .A2(n9787), .ZN(n14821) );
  INV_X1 U13680 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n11888) );
  NAND2_X1 U13681 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14605)
         );
  OAI21_X1 U13682 ( .B1(n15430), .B2(n11888), .A(n14605), .ZN(n11889) );
  AOI21_X1 U13683 ( .B1(n14823), .B2(n15423), .A(n11889), .ZN(n11898) );
  AOI21_X1 U13684 ( .B1(n11892), .B2(n11891), .A(n11890), .ZN(n14816) );
  MUX2_X1 U13685 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11894), .S(n11893), .Z(
        n14815) );
  NAND2_X1 U13686 ( .A1(n14816), .A2(n14815), .ZN(n14814) );
  OAI21_X1 U13687 ( .B1(n14811), .B2(n11894), .A(n14814), .ZN(n11896) );
  MUX2_X1 U13688 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n14836), .S(n14823), .Z(
        n11895) );
  NAND2_X1 U13689 ( .A1(n11896), .A2(n11895), .ZN(n14835) );
  OAI211_X1 U13690 ( .C1(n11896), .C2(n11895), .A(n14835), .B(n15426), .ZN(
        n11897) );
  OAI211_X1 U13691 ( .C1(n11899), .C2(n14821), .A(n11898), .B(n11897), .ZN(
        P1_U3257) );
  INV_X1 U13692 ( .A(SI_21_), .ZN(n13895) );
  OAI222_X1 U13693 ( .A1(n13993), .A2(n11901), .B1(n13995), .B2(n13895), .C1(
        P3_U3151), .C2(n11900), .ZN(P3_U3274) );
  INV_X1 U13694 ( .A(n12239), .ZN(n11911) );
  XNOR2_X1 U13695 ( .A(n15762), .B(n13041), .ZN(n12059) );
  XNOR2_X1 U13696 ( .A(n12059), .B(n12217), .ZN(n11905) );
  OAI21_X1 U13697 ( .B1(n11905), .B2(n11904), .A(n12062), .ZN(n11906) );
  NAND2_X1 U13698 ( .A1(n11906), .A2(n13168), .ZN(n11910) );
  OAI22_X1 U13699 ( .A1(n13195), .A2(n12235), .B1(n12236), .B2(n13174), .ZN(
        n11907) );
  AOI211_X1 U13700 ( .C1(n13197), .C2(n15762), .A(n11908), .B(n11907), .ZN(
        n11909) );
  OAI211_X1 U13701 ( .C1(n11911), .C2(n12585), .A(n11910), .B(n11909), .ZN(
        P3_U3167) );
  XNOR2_X1 U13702 ( .A(n12026), .B(P2_REG2_REG_11__SCAN_IN), .ZN(n11920) );
  NAND2_X1 U13703 ( .A1(n11913), .A2(n11912), .ZN(n11914) );
  NAND2_X1 U13704 ( .A1(n11915), .A2(n11914), .ZN(n15365) );
  MUX2_X1 U13705 ( .A(n11916), .B(P2_REG2_REG_10__SCAN_IN), .S(n15373), .Z(
        n15366) );
  NAND2_X1 U13706 ( .A1(n15373), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11917) );
  NAND2_X1 U13707 ( .A1(n15362), .A2(n11917), .ZN(n11919) );
  INV_X1 U13708 ( .A(n12028), .ZN(n11918) );
  AOI21_X1 U13709 ( .B1(n11920), .B2(n11919), .A(n11918), .ZN(n11932) );
  INV_X1 U13710 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n11922) );
  AND2_X1 U13711 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12286) );
  INV_X1 U13712 ( .A(n12286), .ZN(n11921) );
  OAI21_X1 U13713 ( .B1(n15377), .B2(n11922), .A(n11921), .ZN(n11930) );
  INV_X1 U13714 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11925) );
  MUX2_X1 U13715 ( .A(n11925), .B(P2_REG1_REG_10__SCAN_IN), .S(n15373), .Z(
        n15370) );
  INV_X1 U13716 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11926) );
  MUX2_X1 U13717 ( .A(n11926), .B(P2_REG1_REG_11__SCAN_IN), .S(n12026), .Z(
        n11927) );
  AOI211_X1 U13718 ( .C1(n11928), .C2(n11927), .A(n15368), .B(n12021), .ZN(
        n11929) );
  AOI211_X1 U13719 ( .C1(n15374), .C2(n12026), .A(n11930), .B(n11929), .ZN(
        n11931) );
  OAI21_X1 U13720 ( .B1(n11932), .B2(n15364), .A(n11931), .ZN(P2_U3225) );
  INV_X1 U13721 ( .A(n11933), .ZN(n11937) );
  INV_X1 U13722 ( .A(n15323), .ZN(n11934) );
  OAI222_X1 U13723 ( .A1(n14592), .A2(n11935), .B1(n14578), .B2(n11937), .C1(
        P2_U3088), .C2(n11934), .ZN(P2_U3310) );
  INV_X1 U13724 ( .A(n15394), .ZN(n11938) );
  OAI222_X1 U13725 ( .A1(n11938), .A2(P1_U3086), .B1(n15233), .B2(n11937), 
        .C1(n11936), .C2(n15224), .ZN(P1_U3338) );
  OAI21_X1 U13726 ( .B1(n7432), .B2(n11940), .A(n11939), .ZN(n11942) );
  NAND2_X1 U13727 ( .A1(n11942), .A2(n13565), .ZN(n11944) );
  AOI22_X1 U13728 ( .A1(n13635), .A2(P3_REG2_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(n13634), .ZN(n11943) );
  OAI211_X1 U13729 ( .C1(n11945), .C2(n13571), .A(n11944), .B(n11943), .ZN(
        P3_U3232) );
  OAI211_X1 U13730 ( .C1(n11948), .C2(n15834), .A(n11947), .B(n11946), .ZN(
        n11951) );
  NAND2_X1 U13731 ( .A1(n11951), .A2(n15970), .ZN(n11950) );
  NAND2_X1 U13732 ( .A1(n12043), .A2(n14510), .ZN(n11949) );
  OAI211_X1 U13733 ( .C1(n15970), .C2(n11925), .A(n11950), .B(n11949), .ZN(
        P2_U3509) );
  INV_X1 U13734 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11954) );
  NAND2_X1 U13735 ( .A1(n11951), .A2(n15973), .ZN(n11953) );
  NAND2_X1 U13736 ( .A1(n12043), .A2(n14558), .ZN(n11952) );
  OAI211_X1 U13737 ( .C1(n15973), .C2(n11954), .A(n11953), .B(n11952), .ZN(
        P2_U3460) );
  INV_X1 U13738 ( .A(n11955), .ZN(n11958) );
  AOI211_X1 U13739 ( .C1(n11958), .C2(n15758), .A(n11957), .B(n11956), .ZN(
        n11963) );
  AOI22_X1 U13740 ( .A1(n11998), .A2(n14510), .B1(n15968), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11959) );
  OAI21_X1 U13741 ( .B1(n11963), .B2(n15968), .A(n11959), .ZN(P2_U3508) );
  INV_X1 U13742 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11960) );
  NOR2_X1 U13743 ( .A1(n15973), .A2(n11960), .ZN(n11961) );
  AOI21_X1 U13744 ( .B1(n11998), .B2(n14558), .A(n11961), .ZN(n11962) );
  OAI21_X1 U13745 ( .B1(n11963), .B2(n15971), .A(n11962), .ZN(P2_U3457) );
  INV_X1 U13746 ( .A(n11964), .ZN(n11966) );
  AOI21_X1 U13747 ( .B1(n15936), .B2(P2_REG3_REG_0__SCAN_IN), .A(n11968), .ZN(
        n11970) );
  NAND2_X1 U13748 ( .A1(n15947), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n11969) );
  OAI211_X1 U13749 ( .C1(n14431), .C2(n11971), .A(n11970), .B(n11969), .ZN(
        P2_U3265) );
  INV_X1 U13750 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11983) );
  OAI21_X1 U13751 ( .B1(n8015), .B2(n11974), .A(n11973), .ZN(n12053) );
  XNOR2_X1 U13752 ( .A(n11975), .B(n11974), .ZN(n11978) );
  NAND2_X1 U13753 ( .A1(n14152), .A2(n14184), .ZN(n11976) );
  OAI21_X1 U13754 ( .B1(n12312), .B2(n11977), .A(n11976), .ZN(n12287) );
  AOI21_X1 U13755 ( .B1(n11978), .B2(n15797), .A(n12287), .ZN(n12058) );
  AOI21_X1 U13756 ( .B1(n11979), .B2(n12279), .A(n14360), .ZN(n11980) );
  AND2_X1 U13757 ( .A1(n11980), .A2(n12509), .ZN(n12056) );
  AOI21_X1 U13758 ( .B1(n15959), .B2(n12279), .A(n12056), .ZN(n11981) );
  OAI211_X1 U13759 ( .C1(n12053), .C2(n15834), .A(n12058), .B(n11981), .ZN(
        n14518) );
  NAND2_X1 U13760 ( .A1(n14518), .A2(n15973), .ZN(n11982) );
  OAI21_X1 U13761 ( .B1(n15973), .B2(n11983), .A(n11982), .ZN(P2_U3463) );
  INV_X1 U13762 ( .A(n11984), .ZN(n11992) );
  OAI21_X1 U13763 ( .B1(n11986), .B2(n11992), .A(n11985), .ZN(n11987) );
  XNOR2_X1 U13764 ( .A(n11998), .B(n14072), .ZN(n12045) );
  NOR2_X1 U13765 ( .A1(n7209), .A2(n12044), .ZN(n12036) );
  XNOR2_X1 U13766 ( .A(n12045), .B(n12036), .ZN(n11994) );
  NAND2_X1 U13767 ( .A1(n14095), .A2(n11988), .ZN(n11990) );
  OAI211_X1 U13768 ( .C1(n14092), .C2(n11991), .A(n11990), .B(n11989), .ZN(
        n11997) );
  INV_X1 U13769 ( .A(n11985), .ZN(n11995) );
  AOI22_X1 U13770 ( .A1(n11992), .A2(n14102), .B1(n14126), .B2(n14187), .ZN(
        n11993) );
  NOR3_X1 U13771 ( .A1(n11995), .A2(n11994), .A3(n11993), .ZN(n11996) );
  AOI211_X1 U13772 ( .C1(n11998), .C2(n14159), .A(n11997), .B(n11996), .ZN(
        n11999) );
  OAI21_X1 U13773 ( .B1(n12048), .B2(n14163), .A(n11999), .ZN(P2_U3203) );
  NAND2_X1 U13774 ( .A1(n12213), .A2(n12000), .ZN(n12001) );
  NAND2_X1 U13775 ( .A1(n12002), .A2(n12001), .ZN(n12004) );
  NAND2_X1 U13776 ( .A1(n12004), .A2(n12008), .ZN(n12086) );
  OAI21_X1 U13777 ( .B1(n12004), .B2(n12008), .A(n12086), .ZN(n15868) );
  INV_X1 U13778 ( .A(n15868), .ZN(n12020) );
  INV_X1 U13779 ( .A(n12095), .ZN(n12006) );
  AOI21_X1 U13780 ( .B1(n12008), .B2(n12007), .A(n12006), .ZN(n12011) );
  AOI22_X1 U13781 ( .A1(n12565), .A2(n15076), .B1(n15075), .B2(n14738), .ZN(
        n12010) );
  NAND2_X1 U13782 ( .A1(n15868), .A2(n15025), .ZN(n12009) );
  OAI211_X1 U13783 ( .C1(n12011), .C2(n15747), .A(n12010), .B(n12009), .ZN(
        n15866) );
  NAND2_X1 U13784 ( .A1(n15866), .A2(n15021), .ZN(n12019) );
  OAI22_X1 U13785 ( .A1(n15021), .A2(n12012), .B1(n12271), .B2(n15660), .ZN(
        n12017) );
  INV_X1 U13786 ( .A(n12273), .ZN(n15865) );
  INV_X1 U13787 ( .A(n12349), .ZN(n12014) );
  OAI211_X1 U13788 ( .C1(n15865), .C2(n12015), .A(n12014), .B(n15071), .ZN(
        n15864) );
  NOR2_X1 U13789 ( .A1(n15864), .A2(n15086), .ZN(n12016) );
  AOI211_X1 U13790 ( .C1(n15066), .C2(n12273), .A(n12017), .B(n12016), .ZN(
        n12018) );
  OAI211_X1 U13791 ( .C1(n12020), .C2(n12432), .A(n12019), .B(n12018), .ZN(
        P1_U3284) );
  INV_X1 U13792 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n12022) );
  MUX2_X1 U13793 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n12022), .S(n12615), .Z(
        n12023) );
  OAI21_X1 U13794 ( .B1(n12024), .B2(n12023), .A(n12614), .ZN(n12025) );
  INV_X1 U13795 ( .A(n12025), .ZN(n12035) );
  INV_X1 U13796 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12603) );
  XNOR2_X1 U13797 ( .A(n12615), .B(n12603), .ZN(n12030) );
  OR2_X1 U13798 ( .A1(n12026), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n12027) );
  NAND2_X1 U13799 ( .A1(n12028), .A2(n12027), .ZN(n12029) );
  NAND2_X1 U13800 ( .A1(n12029), .A2(n12030), .ZN(n12606) );
  OAI21_X1 U13801 ( .B1(n12030), .B2(n12029), .A(n12606), .ZN(n12033) );
  NAND2_X1 U13802 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n12321)
         );
  NAND2_X1 U13803 ( .A1(n15271), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n12031) );
  OAI211_X1 U13804 ( .C1(n15322), .C2(n12604), .A(n12321), .B(n12031), .ZN(
        n12032) );
  AOI21_X1 U13805 ( .B1(n12033), .B2(n15333), .A(n12032), .ZN(n12034) );
  OAI21_X1 U13806 ( .B1(n12035), .B2(n15368), .A(n12034), .ZN(P2_U3226) );
  INV_X1 U13807 ( .A(n12036), .ZN(n12037) );
  NOR2_X1 U13808 ( .A1(n7209), .A2(n12038), .ZN(n12276) );
  XNOR2_X1 U13809 ( .A(n12043), .B(n14072), .ZN(n12278) );
  XOR2_X1 U13810 ( .A(n12276), .B(n12278), .Z(n12047) );
  AOI22_X1 U13811 ( .A1(n14095), .A2(n12039), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12040) );
  OAI21_X1 U13812 ( .B1(n12041), .B2(n14092), .A(n12040), .ZN(n12042) );
  AOI21_X1 U13813 ( .B1(n12043), .B2(n14159), .A(n12042), .ZN(n12050) );
  OAI22_X1 U13814 ( .A1(n12045), .A2(n14163), .B1(n12044), .B2(n14146), .ZN(
        n12046) );
  NAND3_X1 U13815 ( .A1(n12048), .A2(n12047), .A3(n12046), .ZN(n12049) );
  OAI211_X1 U13816 ( .C1(n7335), .C2(n14163), .A(n12050), .B(n12049), .ZN(
        P2_U3189) );
  NAND2_X1 U13817 ( .A1(n12279), .A2(n15917), .ZN(n12052) );
  NAND2_X1 U13818 ( .A1(n15947), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n12051) );
  OAI211_X1 U13819 ( .C1(n15714), .C2(n12284), .A(n12052), .B(n12051), .ZN(
        n12055) );
  NOR2_X1 U13820 ( .A1(n12053), .A2(n14369), .ZN(n12054) );
  AOI211_X1 U13821 ( .C1(n12056), .C2(n15934), .A(n12055), .B(n12054), .ZN(
        n12057) );
  OAI21_X1 U13822 ( .B1(n15947), .B2(n12058), .A(n12057), .ZN(P2_U3254) );
  INV_X1 U13823 ( .A(n12225), .ZN(n12068) );
  INV_X1 U13824 ( .A(n12059), .ZN(n12060) );
  NAND2_X1 U13825 ( .A1(n12060), .A2(n12217), .ZN(n12061) );
  XNOR2_X1 U13826 ( .A(n15781), .B(n13041), .ZN(n12103) );
  XNOR2_X1 U13827 ( .A(n12236), .B(n12103), .ZN(n12063) );
  OAI211_X1 U13828 ( .C1(n12064), .C2(n12063), .A(n12105), .B(n13168), .ZN(
        n12067) );
  INV_X1 U13829 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n13978) );
  NOR2_X1 U13830 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13978), .ZN(n13235) );
  OAI22_X1 U13831 ( .A1(n13195), .A2(n12217), .B1(n12302), .B2(n13174), .ZN(
        n12065) );
  AOI211_X1 U13832 ( .C1(n13197), .C2(n15781), .A(n13235), .B(n12065), .ZN(
        n12066) );
  OAI211_X1 U13833 ( .C1(n12068), .C2(n12585), .A(n12067), .B(n12066), .ZN(
        P3_U3179) );
  OR2_X1 U13834 ( .A1(n12070), .A2(n12069), .ZN(n12071) );
  NAND2_X1 U13835 ( .A1(n12072), .A2(n12071), .ZN(n12075) );
  INV_X1 U13836 ( .A(n12075), .ZN(n15738) );
  XNOR2_X1 U13837 ( .A(n12073), .B(n12074), .ZN(n12079) );
  NAND2_X1 U13838 ( .A1(n12075), .A2(n13556), .ZN(n12078) );
  OAI22_X1 U13839 ( .A1(n8398), .A2(n13627), .B1(n12217), .B2(n13629), .ZN(
        n12076) );
  INV_X1 U13840 ( .A(n12076), .ZN(n12077) );
  OAI211_X1 U13841 ( .C1(n12079), .C2(n13625), .A(n12078), .B(n12077), .ZN(
        n15739) );
  MUX2_X1 U13842 ( .A(n15739), .B(P3_REG2_REG_4__SCAN_IN), .S(n13635), .Z(
        n12080) );
  INV_X1 U13843 ( .A(n12080), .ZN(n12084) );
  AOI22_X1 U13844 ( .A1(n13568), .A2(n12082), .B1(n13634), .B2(n12081), .ZN(
        n12083) );
  OAI211_X1 U13845 ( .C1(n15738), .C2(n13571), .A(n12084), .B(n12083), .ZN(
        P3_U3229) );
  INV_X1 U13846 ( .A(n14737), .ZN(n12208) );
  NAND2_X1 U13847 ( .A1(n15865), .A2(n12208), .ZN(n12085) );
  OAI21_X1 U13848 ( .B1(n12087), .B2(n12096), .A(n12354), .ZN(n15883) );
  XNOR2_X1 U13849 ( .A(n12364), .B(n12349), .ZN(n12088) );
  AOI22_X1 U13850 ( .A1(n12088), .A2(n15071), .B1(n15076), .B2(n14736), .ZN(
        n15879) );
  INV_X1 U13851 ( .A(n15879), .ZN(n12089) );
  AOI21_X1 U13852 ( .B1(n15883), .B2(n12090), .A(n12089), .ZN(n12102) );
  NOR2_X1 U13853 ( .A1(n15880), .A2(n15078), .ZN(n12093) );
  OAI22_X1 U13854 ( .A1(n15021), .A2(n12091), .B1(n12368), .B2(n15660), .ZN(
        n12092) );
  AOI211_X1 U13855 ( .C1(n15883), .C2(n15034), .A(n12093), .B(n12092), .ZN(
        n12101) );
  NAND2_X1 U13856 ( .A1(n12273), .A2(n12208), .ZN(n12094) );
  INV_X1 U13857 ( .A(n12096), .ZN(n12097) );
  OAI211_X1 U13858 ( .C1(n12098), .C2(n12097), .A(n12347), .B(n15993), .ZN(
        n12099) );
  OAI21_X1 U13859 ( .B1(n12208), .B2(n15041), .A(n12099), .ZN(n15881) );
  NAND2_X1 U13860 ( .A1(n15881), .A2(n15021), .ZN(n12100) );
  OAI211_X1 U13861 ( .C1(n12102), .C2(n15086), .A(n12101), .B(n12100), .ZN(
        P1_U3283) );
  NAND2_X1 U13862 ( .A1(n13218), .A2(n12103), .ZN(n12104) );
  NAND2_X1 U13863 ( .A1(n12105), .A2(n12104), .ZN(n12243) );
  XNOR2_X1 U13864 ( .A(n12132), .B(n13041), .ZN(n12244) );
  XNOR2_X1 U13865 ( .A(n12244), .B(n12302), .ZN(n12242) );
  XNOR2_X1 U13866 ( .A(n12243), .B(n12242), .ZN(n12111) );
  NAND2_X1 U13867 ( .A1(n13216), .A2(n13191), .ZN(n12108) );
  NAND2_X1 U13868 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n15626) );
  INV_X1 U13869 ( .A(n15626), .ZN(n12106) );
  AOI21_X1 U13870 ( .B1(n13197), .B2(n12132), .A(n12106), .ZN(n12107) );
  OAI211_X1 U13871 ( .C1(n12236), .C2(n13195), .A(n12108), .B(n12107), .ZN(
        n12109) );
  AOI21_X1 U13872 ( .B1(n12131), .B2(n13190), .A(n12109), .ZN(n12110) );
  OAI21_X1 U13873 ( .B1(n12111), .B2(n13200), .A(n12110), .ZN(P3_U3153) );
  INV_X1 U13874 ( .A(SI_23_), .ZN(n12115) );
  NAND2_X1 U13875 ( .A1(n12112), .A2(n13779), .ZN(n12114) );
  OAI211_X1 U13876 ( .C1(n12115), .C2(n13995), .A(n12114), .B(n12113), .ZN(
        P3_U3272) );
  INV_X1 U13877 ( .A(n12116), .ZN(n12118) );
  AOI222_X1 U13878 ( .A1(n12119), .A2(P3_STATE_REG_SCAN_IN), .B1(n12118), .B2(
        n13779), .C1(n12117), .C2(n9283), .ZN(P3_U3273) );
  NAND2_X1 U13879 ( .A1(n12296), .A2(n12121), .ZN(n12122) );
  XNOR2_X1 U13880 ( .A(n12123), .B(n12122), .ZN(n12130) );
  OR2_X1 U13881 ( .A1(n12125), .A2(n12124), .ZN(n12126) );
  NAND2_X1 U13882 ( .A1(n12127), .A2(n12126), .ZN(n15821) );
  OAI22_X1 U13883 ( .A1(n12247), .A2(n13629), .B1(n12236), .B2(n13627), .ZN(
        n12128) );
  AOI21_X1 U13884 ( .B1(n15821), .B2(n13556), .A(n12128), .ZN(n12129) );
  OAI21_X1 U13885 ( .B1(n13625), .B2(n12130), .A(n12129), .ZN(n15819) );
  INV_X1 U13886 ( .A(n15819), .ZN(n12136) );
  AOI22_X1 U13887 ( .A1(n13568), .A2(n12132), .B1(n13634), .B2(n12131), .ZN(
        n12133) );
  OAI21_X1 U13888 ( .B1(n15612), .B2(n13565), .A(n12133), .ZN(n12134) );
  AOI21_X1 U13889 ( .B1(n15821), .B2(n12467), .A(n12134), .ZN(n12135) );
  OAI21_X1 U13890 ( .B1(n12136), .B2(n13635), .A(n12135), .ZN(P3_U3226) );
  OAI21_X1 U13891 ( .B1(n12139), .B2(n12138), .A(n12137), .ZN(n15726) );
  OAI22_X1 U13892 ( .A1(n13637), .A2(n15723), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n13520), .ZN(n12148) );
  AOI21_X1 U13893 ( .B1(n11824), .B2(n12141), .A(n12140), .ZN(n12146) );
  NAND2_X1 U13894 ( .A1(n12142), .A2(n13604), .ZN(n12145) );
  NAND2_X1 U13895 ( .A1(n15726), .A2(n13556), .ZN(n12144) );
  AOI22_X1 U13896 ( .A1(n13222), .A2(n13609), .B1(n13606), .B2(n13220), .ZN(
        n12143) );
  OAI211_X1 U13897 ( .C1(n12146), .C2(n12145), .A(n12144), .B(n12143), .ZN(
        n15724) );
  MUX2_X1 U13898 ( .A(n15724), .B(P3_REG2_REG_3__SCAN_IN), .S(n13635), .Z(
        n12147) );
  AOI211_X1 U13899 ( .C1(n12467), .C2(n15726), .A(n12148), .B(n12147), .ZN(
        n12149) );
  INV_X1 U13900 ( .A(n12149), .ZN(P3_U3230) );
  INV_X1 U13901 ( .A(n12150), .ZN(n12152) );
  OAI222_X1 U13902 ( .A1(P1_U3086), .A2(n14840), .B1(n15233), .B2(n12152), 
        .C1(n12151), .C2(n15224), .ZN(P1_U3337) );
  INV_X1 U13903 ( .A(n15326), .ZN(n15343) );
  OAI222_X1 U13904 ( .A1(n14592), .A2(n12153), .B1(n14578), .B2(n12152), .C1(
        n15343), .C2(P2_U3088), .ZN(P2_U3309) );
  NAND2_X1 U13905 ( .A1(n12174), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n12154) );
  NOR2_X1 U13906 ( .A1(n12178), .A2(n12156), .ZN(n12157) );
  INV_X1 U13907 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15635) );
  INV_X1 U13908 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12465) );
  MUX2_X1 U13909 ( .A(n12465), .B(P3_REG2_REG_10__SCAN_IN), .S(n12335), .Z(
        n12159) );
  INV_X1 U13910 ( .A(n12337), .ZN(n12158) );
  AOI21_X1 U13911 ( .B1(n12160), .B2(n12159), .A(n12158), .ZN(n12188) );
  MUX2_X1 U13912 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n7165), .Z(n12330) );
  INV_X1 U13913 ( .A(n12335), .ZN(n12161) );
  XNOR2_X1 U13914 ( .A(n12330), .B(n12161), .ZN(n12172) );
  INV_X1 U13915 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12162) );
  MUX2_X1 U13916 ( .A(n15635), .B(n12162), .S(n7165), .Z(n12163) );
  NOR2_X1 U13917 ( .A1(n12163), .A2(n12178), .ZN(n12170) );
  INV_X1 U13918 ( .A(n12163), .ZN(n12164) );
  NOR2_X1 U13919 ( .A1(n12164), .A2(n15642), .ZN(n12165) );
  NOR2_X1 U13920 ( .A1(n12170), .A2(n12165), .ZN(n15640) );
  INV_X1 U13921 ( .A(n12166), .ZN(n12167) );
  NOR2_X1 U13922 ( .A1(n12170), .A2(n15643), .ZN(n12171) );
  OAI21_X1 U13923 ( .B1(n12172), .B2(n12171), .A(n12331), .ZN(n12186) );
  INV_X1 U13924 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n13935) );
  NOR2_X1 U13925 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13935), .ZN(n12582) );
  AOI21_X1 U13926 ( .B1(n15246), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n12582), 
        .ZN(n12173) );
  OAI21_X1 U13927 ( .B1(n15641), .B2(n12335), .A(n12173), .ZN(n12185) );
  NAND2_X1 U13928 ( .A1(n12174), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n12175) );
  NOR2_X1 U13929 ( .A1(n12178), .A2(n12177), .ZN(n12179) );
  INV_X1 U13930 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12180) );
  MUX2_X1 U13931 ( .A(n12180), .B(P3_REG1_REG_10__SCAN_IN), .S(n12335), .Z(
        n12181) );
  OR2_X2 U13932 ( .A1(n12182), .A2(n12181), .ZN(n12327) );
  NAND2_X1 U13933 ( .A1(n12182), .A2(n12181), .ZN(n12183) );
  AOI21_X1 U13934 ( .B1(n12327), .B2(n12183), .A(n15631), .ZN(n12184) );
  AOI211_X1 U13935 ( .C1(n15638), .C2(n12186), .A(n12185), .B(n12184), .ZN(
        n12187) );
  OAI21_X1 U13936 ( .B1(n12188), .B2(n15636), .A(n12187), .ZN(P3_U3192) );
  INV_X1 U13937 ( .A(n12189), .ZN(n12192) );
  INV_X1 U13938 ( .A(n12190), .ZN(n12191) );
  NAND2_X1 U13939 ( .A1(n12198), .A2(n13014), .ZN(n12196) );
  NAND2_X1 U13940 ( .A1(n14738), .A2(n12999), .ZN(n12195) );
  NAND2_X1 U13941 ( .A1(n12196), .A2(n12195), .ZN(n12197) );
  XNOR2_X1 U13942 ( .A(n12197), .B(n13025), .ZN(n12202) );
  NAND2_X1 U13943 ( .A1(n12198), .A2(n13019), .ZN(n12200) );
  NAND2_X1 U13944 ( .A1(n13018), .A2(n14738), .ZN(n12199) );
  NAND2_X1 U13945 ( .A1(n12200), .A2(n12199), .ZN(n12201) );
  NOR2_X1 U13946 ( .A1(n12202), .A2(n12201), .ZN(n12255) );
  AOI21_X1 U13947 ( .B1(n12202), .B2(n12201), .A(n12255), .ZN(n12203) );
  OAI21_X1 U13948 ( .B1(n12204), .B2(n12203), .A(n12257), .ZN(n12205) );
  NAND2_X1 U13949 ( .A1(n12205), .A2(n16010), .ZN(n12212) );
  NOR2_X1 U13950 ( .A1(n16031), .A2(n12206), .ZN(n12210) );
  OAI21_X1 U13951 ( .B1(n16019), .B2(n12208), .A(n12207), .ZN(n12209) );
  AOI211_X1 U13952 ( .C1(n15980), .C2(n14739), .A(n12210), .B(n12209), .ZN(
        n12211) );
  OAI211_X1 U13953 ( .C1(n12213), .C2(n15982), .A(n12212), .B(n12211), .ZN(
        P1_U3221) );
  OAI21_X1 U13954 ( .B1(n12216), .B2(n12215), .A(n12214), .ZN(n15782) );
  INV_X1 U13955 ( .A(n15782), .ZN(n12228) );
  OAI22_X1 U13956 ( .A1(n12217), .A2(n13627), .B1(n12302), .B2(n13629), .ZN(
        n12223) );
  INV_X1 U13957 ( .A(n12296), .ZN(n12221) );
  AOI21_X1 U13958 ( .B1(n12230), .B2(n12219), .A(n12218), .ZN(n12220) );
  NOR3_X1 U13959 ( .A1(n12221), .A2(n12220), .A3(n13625), .ZN(n12222) );
  AOI211_X1 U13960 ( .C1(n13556), .C2(n15782), .A(n12223), .B(n12222), .ZN(
        n15784) );
  MUX2_X1 U13961 ( .A(n12224), .B(n15784), .S(n13565), .Z(n12227) );
  AOI22_X1 U13962 ( .A1(n13568), .A2(n15781), .B1(n13634), .B2(n12225), .ZN(
        n12226) );
  OAI211_X1 U13963 ( .C1(n12228), .C2(n13571), .A(n12227), .B(n12226), .ZN(
        P3_U3227) );
  AOI21_X1 U13964 ( .B1(n13556), .B2(n13565), .A(n12467), .ZN(n13512) );
  XOR2_X1 U13965 ( .A(n12229), .B(n12233), .Z(n15765) );
  INV_X1 U13966 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n12238) );
  INV_X1 U13967 ( .A(n12230), .ZN(n12231) );
  AOI21_X1 U13968 ( .B1(n12233), .B2(n12232), .A(n12231), .ZN(n12234) );
  OAI222_X1 U13969 ( .A1(n13629), .A2(n12236), .B1(n13627), .B2(n12235), .C1(
        n13625), .C2(n12234), .ZN(n15761) );
  INV_X1 U13970 ( .A(n15761), .ZN(n12237) );
  MUX2_X1 U13971 ( .A(n12238), .B(n12237), .S(n13565), .Z(n12241) );
  AOI22_X1 U13972 ( .A1(n13568), .A2(n15762), .B1(n13634), .B2(n12239), .ZN(
        n12240) );
  OAI211_X1 U13973 ( .C1(n13512), .C2(n15765), .A(n12241), .B(n12240), .ZN(
        P3_U3228) );
  NAND2_X1 U13974 ( .A1(n12243), .A2(n12242), .ZN(n12246) );
  NAND2_X1 U13975 ( .A1(n13217), .A2(n12244), .ZN(n12245) );
  NAND2_X1 U13976 ( .A1(n12246), .A2(n12245), .ZN(n12471) );
  XNOR2_X1 U13977 ( .A(n15841), .B(n13041), .ZN(n12472) );
  XNOR2_X1 U13978 ( .A(n12247), .B(n12472), .ZN(n12470) );
  XNOR2_X1 U13979 ( .A(n12471), .B(n12470), .ZN(n12254) );
  INV_X1 U13980 ( .A(n12248), .ZN(n12249) );
  OAI21_X1 U13981 ( .B1(n13178), .B2(n12250), .A(n12249), .ZN(n12252) );
  OAI22_X1 U13982 ( .A1(n13195), .A2(n12302), .B1(n12580), .B2(n13174), .ZN(
        n12251) );
  AOI211_X1 U13983 ( .C1(n12307), .C2(n13190), .A(n12252), .B(n12251), .ZN(
        n12253) );
  OAI21_X1 U13984 ( .B1(n12254), .B2(n13200), .A(n12253), .ZN(P3_U3161) );
  INV_X1 U13985 ( .A(n12255), .ZN(n12256) );
  NAND2_X1 U13986 ( .A1(n12273), .A2(n13014), .ZN(n12259) );
  NAND2_X1 U13987 ( .A1(n14737), .A2(n13019), .ZN(n12258) );
  NAND2_X1 U13988 ( .A1(n12259), .A2(n12258), .ZN(n12260) );
  XNOR2_X1 U13989 ( .A(n12260), .B(n13009), .ZN(n12262) );
  AND2_X1 U13990 ( .A1(n13018), .A2(n14737), .ZN(n12261) );
  AOI21_X1 U13991 ( .B1(n12273), .B2(n13019), .A(n12261), .ZN(n12263) );
  AND2_X1 U13992 ( .A1(n12262), .A2(n12263), .ZN(n12359) );
  INV_X1 U13993 ( .A(n12359), .ZN(n12266) );
  INV_X1 U13994 ( .A(n12262), .ZN(n12265) );
  INV_X1 U13995 ( .A(n12263), .ZN(n12264) );
  NAND2_X1 U13996 ( .A1(n12265), .A2(n12264), .ZN(n12360) );
  NAND2_X1 U13997 ( .A1(n12266), .A2(n12360), .ZN(n12267) );
  XNOR2_X1 U13998 ( .A(n12361), .B(n12267), .ZN(n12275) );
  OAI21_X1 U13999 ( .B1(n16019), .B2(n12362), .A(n12268), .ZN(n12269) );
  AOI21_X1 U14000 ( .B1(n15980), .B2(n14738), .A(n12269), .ZN(n12270) );
  OAI21_X1 U14001 ( .B1(n12271), .B2(n16031), .A(n12270), .ZN(n12272) );
  AOI21_X1 U14002 ( .B1(n16027), .B2(n12273), .A(n12272), .ZN(n12274) );
  OAI21_X1 U14003 ( .B1(n12275), .B2(n16022), .A(n12274), .ZN(P1_U3231) );
  INV_X1 U14004 ( .A(n12276), .ZN(n12277) );
  XNOR2_X1 U14005 ( .A(n12279), .B(n14072), .ZN(n12316) );
  OR2_X1 U14006 ( .A1(n12280), .A2(n14308), .ZN(n12281) );
  NOR2_X1 U14007 ( .A1(n12316), .A2(n12281), .ZN(n12313) );
  AOI21_X1 U14008 ( .B1(n12316), .B2(n12281), .A(n12313), .ZN(n12282) );
  OAI211_X1 U14009 ( .C1(n12283), .C2(n12282), .A(n12317), .B(n14102), .ZN(
        n12289) );
  NOR2_X1 U14010 ( .A1(n14092), .A2(n12284), .ZN(n12285) );
  AOI211_X1 U14011 ( .C1(n14095), .C2(n12287), .A(n12286), .B(n12285), .ZN(
        n12288) );
  OAI211_X1 U14012 ( .C1(n7632), .C2(n14135), .A(n12289), .B(n12288), .ZN(
        P2_U3208) );
  OR2_X1 U14013 ( .A1(n12291), .A2(n12299), .ZN(n12292) );
  NAND2_X1 U14014 ( .A1(n12290), .A2(n12292), .ZN(n15842) );
  NAND2_X1 U14015 ( .A1(n15842), .A2(n13556), .ZN(n12306) );
  NAND2_X1 U14016 ( .A1(n12296), .A2(n12293), .ZN(n12392) );
  AND2_X1 U14017 ( .A1(n12392), .A2(n12294), .ZN(n12390) );
  NAND2_X1 U14018 ( .A1(n12296), .A2(n12295), .ZN(n12298) );
  AND2_X1 U14019 ( .A1(n12297), .A2(n12298), .ZN(n12300) );
  NAND2_X1 U14020 ( .A1(n12300), .A2(n12299), .ZN(n12301) );
  NAND2_X1 U14021 ( .A1(n12390), .A2(n12301), .ZN(n12304) );
  OAI22_X1 U14022 ( .A1(n12302), .A2(n13627), .B1(n12580), .B2(n13629), .ZN(
        n12303) );
  AOI21_X1 U14023 ( .B1(n12304), .B2(n13604), .A(n12303), .ZN(n12305) );
  AND2_X1 U14024 ( .A1(n12306), .A2(n12305), .ZN(n15844) );
  AOI22_X1 U14025 ( .A1(n13568), .A2(n15841), .B1(n13634), .B2(n12307), .ZN(
        n12308) );
  OAI21_X1 U14026 ( .B1(n12309), .B2(n13565), .A(n12308), .ZN(n12310) );
  AOI21_X1 U14027 ( .B1(n15842), .B2(n12467), .A(n12310), .ZN(n12311) );
  OAI21_X1 U14028 ( .B1(n15844), .B2(n13635), .A(n12311), .ZN(P3_U3225) );
  XNOR2_X1 U14029 ( .A(n15918), .B(n14072), .ZN(n12486) );
  NOR2_X1 U14030 ( .A1(n7209), .A2(n12312), .ZN(n12487) );
  XNOR2_X1 U14031 ( .A(n12486), .B(n12487), .ZN(n12318) );
  INV_X1 U14032 ( .A(n12313), .ZN(n12314) );
  NAND3_X1 U14033 ( .A1(n12317), .A2(n12318), .A3(n12314), .ZN(n12490) );
  NAND2_X1 U14034 ( .A1(n14126), .A2(n14183), .ZN(n12315) );
  OAI22_X1 U14035 ( .A1(n12317), .A2(n14163), .B1(n12316), .B2(n12315), .ZN(
        n12320) );
  INV_X1 U14036 ( .A(n12318), .ZN(n12319) );
  NAND2_X1 U14037 ( .A1(n12320), .A2(n12319), .ZN(n12325) );
  NOR2_X1 U14038 ( .A1(n14092), .A2(n15915), .ZN(n12323) );
  AOI22_X1 U14039 ( .A1(n14153), .A2(n14181), .B1(n14152), .B2(n14183), .ZN(
        n12512) );
  OAI21_X1 U14040 ( .B1(n14157), .B2(n12512), .A(n12321), .ZN(n12322) );
  AOI211_X1 U14041 ( .C1(n15918), .C2(n14159), .A(n12323), .B(n12322), .ZN(
        n12324) );
  OAI211_X1 U14042 ( .C1(n12490), .C2(n14163), .A(n12325), .B(n12324), .ZN(
        P2_U3196) );
  INV_X1 U14043 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n15893) );
  NAND2_X1 U14044 ( .A1(n12335), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n12326) );
  NOR2_X1 U14045 ( .A1(n15893), .A2(n12328), .ZN(n12696) );
  AOI21_X1 U14046 ( .B1(n15893), .B2(n12328), .A(n12696), .ZN(n12345) );
  INV_X1 U14047 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12329) );
  MUX2_X1 U14048 ( .A(n12329), .B(n15893), .S(n7206), .Z(n12702) );
  XNOR2_X1 U14049 ( .A(n12702), .B(n12687), .ZN(n12334) );
  OR2_X1 U14050 ( .A1(n12330), .A2(n12335), .ZN(n12332) );
  NAND2_X1 U14051 ( .A1(n12334), .A2(n12333), .ZN(n12700) );
  OAI21_X1 U14052 ( .B1(n12334), .B2(n12333), .A(n12700), .ZN(n12343) );
  INV_X1 U14053 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n13793) );
  NOR2_X1 U14054 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13793), .ZN(n12718) );
  NAND2_X1 U14055 ( .A1(n12335), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n12336) );
  AOI21_X1 U14056 ( .B1(n12338), .B2(n12329), .A(n12689), .ZN(n12339) );
  NOR2_X1 U14057 ( .A1(n15636), .A2(n12339), .ZN(n12340) );
  AOI211_X1 U14058 ( .C1(n15246), .C2(P3_ADDR_REG_11__SCAN_IN), .A(n12718), 
        .B(n12340), .ZN(n12341) );
  OAI21_X1 U14059 ( .B1(n12687), .B2(n15641), .A(n12341), .ZN(n12342) );
  AOI21_X1 U14060 ( .B1(n15638), .B2(n12343), .A(n12342), .ZN(n12344) );
  OAI21_X1 U14061 ( .B1(n12345), .B2(n15631), .A(n12344), .ZN(P3_U3193) );
  NAND2_X1 U14062 ( .A1(n15880), .A2(n12565), .ZN(n12346) );
  XNOR2_X1 U14063 ( .A(n12409), .B(n12355), .ZN(n12348) );
  AOI222_X1 U14064 ( .A1(n15993), .A2(n12348), .B1(n14735), .B2(n15076), .C1(
        n12565), .C2(n15075), .ZN(n15902) );
  AOI211_X1 U14065 ( .C1(n15900), .C2(n12350), .A(n15731), .B(n7234), .ZN(
        n15899) );
  INV_X1 U14066 ( .A(n12567), .ZN(n12351) );
  AOI22_X1 U14067 ( .A1(n15667), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12351), 
        .B2(n15043), .ZN(n12352) );
  OAI21_X1 U14068 ( .B1(n7586), .B2(n15078), .A(n12352), .ZN(n12357) );
  NAND2_X1 U14069 ( .A1(n15880), .A2(n12362), .ZN(n12353) );
  XOR2_X1 U14070 ( .A(n12405), .B(n12355), .Z(n15903) );
  NOR2_X1 U14071 ( .A1(n15903), .A2(n14897), .ZN(n12356) );
  AOI211_X1 U14072 ( .C1(n15899), .C2(n15049), .A(n12357), .B(n12356), .ZN(
        n12358) );
  OAI21_X1 U14073 ( .B1(n15667), .B2(n15902), .A(n12358), .ZN(P1_U3282) );
  NOR2_X1 U14074 ( .A1(n12362), .A2(n13023), .ZN(n12363) );
  AOI21_X1 U14075 ( .B1(n12364), .B2(n13019), .A(n12363), .ZN(n12559) );
  AOI22_X1 U14076 ( .A1(n12364), .A2(n13014), .B1(n13019), .B2(n12565), .ZN(
        n12365) );
  XNOR2_X1 U14077 ( .A(n12365), .B(n13025), .ZN(n12558) );
  XOR2_X1 U14078 ( .A(n12559), .B(n12558), .Z(n12366) );
  OAI211_X1 U14079 ( .C1(n12367), .C2(n12366), .A(n12557), .B(n16010), .ZN(
        n12372) );
  NOR2_X1 U14080 ( .A1(n16031), .A2(n12368), .ZN(n12370) );
  NAND2_X1 U14081 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n14797)
         );
  OAI21_X1 U14082 ( .B1(n16019), .B2(n12423), .A(n14797), .ZN(n12369) );
  AOI211_X1 U14083 ( .C1(n15980), .C2(n14737), .A(n12370), .B(n12369), .ZN(
        n12371) );
  OAI211_X1 U14084 ( .C1(n15880), .C2(n15982), .A(n12372), .B(n12371), .ZN(
        P1_U3217) );
  XOR2_X1 U14085 ( .A(n12373), .B(n12380), .Z(n12374) );
  AOI22_X1 U14086 ( .A1(n14179), .A2(n14153), .B1(n14152), .B2(n14181), .ZN(
        n12652) );
  OAI21_X1 U14087 ( .B1(n12374), .B2(n15702), .A(n12652), .ZN(n12548) );
  INV_X1 U14088 ( .A(n12548), .ZN(n12384) );
  INV_X1 U14089 ( .A(n12444), .ZN(n12375) );
  AOI211_X1 U14090 ( .C1(n12655), .C2(n12524), .A(n14360), .B(n12375), .ZN(
        n12549) );
  INV_X1 U14091 ( .A(n12655), .ZN(n12376) );
  NOR2_X1 U14092 ( .A1(n12376), .A2(n15940), .ZN(n12379) );
  INV_X1 U14093 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12377) );
  OAI22_X1 U14094 ( .A1(n15721), .A2(n12377), .B1(n12650), .B2(n15714), .ZN(
        n12378) );
  AOI211_X1 U14095 ( .C1(n12549), .C2(n15934), .A(n12379), .B(n12378), .ZN(
        n12383) );
  XNOR2_X1 U14096 ( .A(n12381), .B(n12380), .ZN(n12550) );
  NAND2_X1 U14097 ( .A1(n12550), .A2(n15807), .ZN(n12382) );
  OAI211_X1 U14098 ( .C1(n15947), .C2(n12384), .A(n12383), .B(n12382), .ZN(
        P2_U3251) );
  INV_X1 U14099 ( .A(n12290), .ZN(n12386) );
  OAI21_X1 U14100 ( .B1(n12386), .B2(n12385), .A(n12394), .ZN(n12388) );
  NAND2_X1 U14101 ( .A1(n12388), .A2(n7411), .ZN(n15859) );
  AOI22_X1 U14102 ( .A1(n13609), .A2(n13216), .B1(n13214), .B2(n13606), .ZN(
        n12397) );
  AND2_X1 U14103 ( .A1(n12390), .A2(n12389), .ZN(n12395) );
  NAND2_X1 U14104 ( .A1(n12392), .A2(n12391), .ZN(n12393) );
  OAI211_X1 U14105 ( .C1(n12395), .C2(n12394), .A(n12393), .B(n13604), .ZN(
        n12396) );
  OAI211_X1 U14106 ( .C1(n15859), .C2(n15764), .A(n12397), .B(n12396), .ZN(
        n15861) );
  NAND2_X1 U14107 ( .A1(n15861), .A2(n13565), .ZN(n12401) );
  INV_X1 U14108 ( .A(n12479), .ZN(n12398) );
  OAI22_X1 U14109 ( .A1(n13637), .A2(n15857), .B1(n12398), .B2(n13520), .ZN(
        n12399) );
  AOI21_X1 U14110 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n13635), .A(n12399), .ZN(
        n12400) );
  OAI211_X1 U14111 ( .C1(n15859), .C2(n13571), .A(n12401), .B(n12400), .ZN(
        P3_U3224) );
  INV_X1 U14112 ( .A(n12402), .ZN(n12899) );
  OAI222_X1 U14113 ( .A1(P1_U3086), .A2(n12404), .B1(n15233), .B2(n12899), 
        .C1(n12403), .C2(n15224), .ZN(P1_U3336) );
  INV_X1 U14114 ( .A(n12419), .ZN(n12421) );
  OR2_X1 U14115 ( .A1(n12915), .A2(n14735), .ZN(n12406) );
  XNOR2_X1 U14116 ( .A(n12625), .B(n8112), .ZN(n15927) );
  NAND2_X1 U14117 ( .A1(n15900), .A2(n12423), .ZN(n12408) );
  OR2_X1 U14118 ( .A1(n15900), .A2(n12423), .ZN(n12410) );
  INV_X1 U14119 ( .A(n14735), .ZN(n12563) );
  OR2_X1 U14120 ( .A1(n12915), .A2(n12563), .ZN(n12411) );
  XNOR2_X1 U14121 ( .A(n12628), .B(n12624), .ZN(n15930) );
  NAND2_X1 U14122 ( .A1(n15930), .A2(n15083), .ZN(n12418) );
  OAI211_X1 U14123 ( .C1(n15926), .C2(n12427), .A(n15071), .B(n12636), .ZN(
        n15925) );
  INV_X1 U14124 ( .A(n15925), .ZN(n12416) );
  AOI22_X1 U14125 ( .A1(n15075), .A2(n14735), .B1(n15979), .B2(n15076), .ZN(
        n15924) );
  OAI22_X1 U14126 ( .A1(n15667), .A2(n15924), .B1(n14687), .B2(n15660), .ZN(
        n12413) );
  AOI21_X1 U14127 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n15667), .A(n12413), 
        .ZN(n12414) );
  OAI21_X1 U14128 ( .B1(n15926), .B2(n15078), .A(n12414), .ZN(n12415) );
  AOI21_X1 U14129 ( .B1(n12416), .B2(n15049), .A(n12415), .ZN(n12417) );
  OAI211_X1 U14130 ( .C1(n15927), .C2(n15069), .A(n12418), .B(n12417), .ZN(
        P1_U3280) );
  XNOR2_X1 U14131 ( .A(n12420), .B(n12419), .ZN(n15907) );
  XNOR2_X1 U14132 ( .A(n12422), .B(n12421), .ZN(n12425) );
  OAI22_X1 U14133 ( .A1(n12423), .A2(n15041), .B1(n14649), .B2(n15042), .ZN(
        n12424) );
  AOI21_X1 U14134 ( .B1(n12425), .B2(n15993), .A(n12424), .ZN(n12426) );
  OAI21_X1 U14135 ( .B1(n15671), .B2(n15907), .A(n12426), .ZN(n15909) );
  NAND2_X1 U14136 ( .A1(n15909), .A2(n15021), .ZN(n12431) );
  OAI22_X1 U14137 ( .A1(n15021), .A2(n11892), .B1(n14647), .B2(n15660), .ZN(
        n12429) );
  OAI211_X1 U14138 ( .C1(n7584), .C2(n7234), .A(n7587), .B(n15071), .ZN(n15908) );
  NOR2_X1 U14139 ( .A1(n15908), .A2(n15086), .ZN(n12428) );
  AOI211_X1 U14140 ( .C1(n15066), .C2(n12915), .A(n12429), .B(n12428), .ZN(
        n12430) );
  OAI211_X1 U14141 ( .C1(n15907), .C2(n12432), .A(n12431), .B(n12430), .ZN(
        P1_U3281) );
  XNOR2_X1 U14142 ( .A(n12434), .B(n12433), .ZN(n12435) );
  OR2_X1 U14143 ( .A1(n12435), .A2(n15702), .ZN(n12439) );
  NAND2_X1 U14144 ( .A1(n14178), .A2(n14153), .ZN(n12437) );
  NAND2_X1 U14145 ( .A1(n14152), .A2(n14180), .ZN(n12436) );
  NAND2_X1 U14146 ( .A1(n12437), .A2(n12436), .ZN(n12748) );
  INV_X1 U14147 ( .A(n12748), .ZN(n12438) );
  OR2_X1 U14148 ( .A1(n12441), .A2(n12440), .ZN(n12442) );
  NAND2_X1 U14149 ( .A1(n12443), .A2(n12442), .ZN(n15965) );
  NAND2_X1 U14150 ( .A1(n15960), .A2(n12444), .ZN(n12445) );
  NAND2_X1 U14151 ( .A1(n12445), .A2(n7209), .ZN(n12446) );
  OR2_X1 U14152 ( .A1(n12597), .A2(n12446), .ZN(n15962) );
  INV_X1 U14153 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12447) );
  OAI22_X1 U14154 ( .A1(n15721), .A2(n12447), .B1(n12750), .B2(n15714), .ZN(
        n12448) );
  AOI21_X1 U14155 ( .B1(n15960), .B2(n15917), .A(n12448), .ZN(n12449) );
  OAI21_X1 U14156 ( .B1(n15962), .B2(n15717), .A(n12449), .ZN(n12450) );
  AOI21_X1 U14157 ( .B1(n15965), .B2(n15807), .A(n12450), .ZN(n12451) );
  OAI21_X1 U14158 ( .B1(n15967), .B2(n15947), .A(n12451), .ZN(P2_U3250) );
  NAND2_X1 U14159 ( .A1(n12453), .A2(n12452), .ZN(n12454) );
  NAND2_X1 U14160 ( .A1(n12455), .A2(n12454), .ZN(n15874) );
  NAND2_X1 U14161 ( .A1(n15874), .A2(n13556), .ZN(n12463) );
  AND2_X1 U14162 ( .A1(n12457), .A2(n12456), .ZN(n12458) );
  XNOR2_X1 U14163 ( .A(n12458), .B(n8149), .ZN(n12461) );
  NAND2_X1 U14164 ( .A1(n13213), .A2(n13606), .ZN(n12459) );
  OAI21_X1 U14165 ( .B1(n12580), .B2(n13627), .A(n12459), .ZN(n12460) );
  AOI21_X1 U14166 ( .B1(n12461), .B2(n13604), .A(n12460), .ZN(n12462) );
  AND2_X1 U14167 ( .A1(n12463), .A2(n12462), .ZN(n15876) );
  AOI22_X1 U14168 ( .A1(n13568), .A2(n15871), .B1(n13634), .B2(n12571), .ZN(
        n12464) );
  OAI21_X1 U14169 ( .B1(n12465), .B2(n13565), .A(n12464), .ZN(n12466) );
  AOI21_X1 U14170 ( .B1(n15874), .B2(n12467), .A(n12466), .ZN(n12468) );
  OAI21_X1 U14171 ( .B1(n15876), .B2(n13635), .A(n12468), .ZN(P3_U3223) );
  XNOR2_X1 U14172 ( .A(n12469), .B(n13103), .ZN(n12572) );
  XNOR2_X1 U14173 ( .A(n12572), .B(n12580), .ZN(n12477) );
  NAND2_X1 U14174 ( .A1(n13216), .A2(n12472), .ZN(n12473) );
  INV_X1 U14175 ( .A(n12477), .ZN(n12474) );
  INV_X1 U14176 ( .A(n12576), .ZN(n12475) );
  AOI21_X1 U14177 ( .B1(n12477), .B2(n12476), .A(n12475), .ZN(n12482) );
  NOR2_X1 U14178 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8262), .ZN(n15648) );
  OAI22_X1 U14179 ( .A1(n12573), .A2(n13174), .B1(n13178), .B2(n15857), .ZN(
        n12478) );
  AOI211_X1 U14180 ( .C1(n13172), .C2(n13216), .A(n15648), .B(n12478), .ZN(
        n12481) );
  NAND2_X1 U14181 ( .A1(n13190), .A2(n12479), .ZN(n12480) );
  OAI211_X1 U14182 ( .C1(n12482), .C2(n13200), .A(n12481), .B(n12480), .ZN(
        P3_U3171) );
  INV_X1 U14183 ( .A(n12483), .ZN(n12502) );
  OAI222_X1 U14184 ( .A1(n12485), .A2(P1_U3086), .B1(n15233), .B2(n12502), 
        .C1(n12484), .C2(n15224), .ZN(P1_U3335) );
  NAND2_X1 U14185 ( .A1(n12486), .A2(n12488), .ZN(n12489) );
  XNOR2_X1 U14186 ( .A(n12537), .B(n14038), .ZN(n12494) );
  NOR2_X1 U14187 ( .A1(n7209), .A2(n12491), .ZN(n12493) );
  NOR2_X1 U14188 ( .A1(n12494), .A2(n12493), .ZN(n12646) );
  INV_X1 U14189 ( .A(n12646), .ZN(n12495) );
  NAND2_X1 U14190 ( .A1(n12494), .A2(n12493), .ZN(n12645) );
  NAND2_X1 U14191 ( .A1(n12495), .A2(n12645), .ZN(n12496) );
  XNOR2_X1 U14192 ( .A(n12647), .B(n12496), .ZN(n12501) );
  AOI22_X1 U14193 ( .A1(n14153), .A2(n14180), .B1(n14152), .B2(n14182), .ZN(
        n12529) );
  OAI22_X1 U14194 ( .A1(n14157), .A2(n12529), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12497), .ZN(n12499) );
  NOR2_X1 U14195 ( .A1(n15941), .A2(n14135), .ZN(n12498) );
  AOI211_X1 U14196 ( .C1(n14155), .C2(n15937), .A(n12499), .B(n12498), .ZN(
        n12500) );
  OAI21_X1 U14197 ( .B1(n12501), .B2(n14163), .A(n12500), .ZN(P2_U3206) );
  OAI222_X1 U14198 ( .A1(n14592), .A2(n12504), .B1(P2_U3088), .B2(n12503), 
        .C1(n14578), .C2(n12502), .ZN(P2_U3307) );
  INV_X1 U14199 ( .A(SI_24_), .ZN(n13887) );
  INV_X1 U14200 ( .A(n12505), .ZN(n12506) );
  OAI222_X1 U14201 ( .A1(P3_U3151), .A2(n12507), .B1(n13995), .B2(n13887), 
        .C1(n13993), .C2(n12506), .ZN(P3_U3271) );
  XNOR2_X1 U14202 ( .A(n12508), .B(n12511), .ZN(n15919) );
  AOI211_X1 U14203 ( .C1(n15918), .C2(n12509), .A(n14360), .B(n12523), .ZN(
        n15920) );
  XOR2_X1 U14204 ( .A(n12511), .B(n12510), .Z(n12513) );
  OAI21_X1 U14205 ( .B1(n12513), .B2(n15702), .A(n12512), .ZN(n12514) );
  AOI21_X1 U14206 ( .B1(n12532), .B2(n15919), .A(n12514), .ZN(n15923) );
  INV_X1 U14207 ( .A(n15923), .ZN(n12515) );
  AOI211_X1 U14208 ( .C1(n15758), .C2(n15919), .A(n15920), .B(n12515), .ZN(
        n12520) );
  AOI22_X1 U14209 ( .A1(n15918), .A2(n14510), .B1(n15968), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n12516) );
  OAI21_X1 U14210 ( .B1(n12520), .B2(n15968), .A(n12516), .ZN(P2_U3511) );
  INV_X1 U14211 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n12517) );
  NOR2_X1 U14212 ( .A1(n15973), .A2(n12517), .ZN(n12518) );
  AOI21_X1 U14213 ( .B1(n15918), .B2(n14558), .A(n12518), .ZN(n12519) );
  OAI21_X1 U14214 ( .B1(n12520), .B2(n15971), .A(n12519), .ZN(P2_U3466) );
  XNOR2_X1 U14215 ( .A(n12522), .B(n12521), .ZN(n15943) );
  INV_X1 U14216 ( .A(n12523), .ZN(n12526) );
  INV_X1 U14217 ( .A(n12524), .ZN(n12525) );
  AOI211_X1 U14218 ( .C1(n12537), .C2(n12526), .A(n14360), .B(n12525), .ZN(
        n15935) );
  XNOR2_X1 U14219 ( .A(n12528), .B(n12527), .ZN(n12530) );
  OAI21_X1 U14220 ( .B1(n12530), .B2(n15702), .A(n12529), .ZN(n12531) );
  AOI21_X1 U14221 ( .B1(n12532), .B2(n15943), .A(n12531), .ZN(n15946) );
  INV_X1 U14222 ( .A(n15946), .ZN(n12533) );
  AOI211_X1 U14223 ( .C1(n15758), .C2(n15943), .A(n15935), .B(n12533), .ZN(
        n12539) );
  INV_X1 U14224 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n12534) );
  OAI22_X1 U14225 ( .A1(n15941), .A2(n14553), .B1(n15973), .B2(n12534), .ZN(
        n12535) );
  INV_X1 U14226 ( .A(n12535), .ZN(n12536) );
  OAI21_X1 U14227 ( .B1(n12539), .B2(n15971), .A(n12536), .ZN(P2_U3469) );
  INV_X1 U14228 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U14229 ( .A1(n12537), .A2(n14510), .B1(n15968), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n12538) );
  OAI21_X1 U14230 ( .B1(n12539), .B2(n15968), .A(n12538), .ZN(P2_U3512) );
  XOR2_X1 U14231 ( .A(n12540), .B(n12717), .Z(n12541) );
  OAI222_X1 U14232 ( .A1(n13629), .A2(n12804), .B1(n13627), .B2(n12573), .C1(
        n12541), .C2(n13625), .ZN(n15888) );
  INV_X1 U14233 ( .A(n15888), .ZN(n12547) );
  OAI21_X1 U14234 ( .B1(n12543), .B2(n12717), .A(n12542), .ZN(n15890) );
  AOI22_X1 U14235 ( .A1(n13635), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n13634), 
        .B2(n12719), .ZN(n12544) );
  OAI21_X1 U14236 ( .B1(n15887), .B2(n13637), .A(n12544), .ZN(n12545) );
  AOI21_X1 U14237 ( .B1(n15890), .B2(n13639), .A(n12545), .ZN(n12546) );
  OAI21_X1 U14238 ( .B1(n12547), .B2(n13635), .A(n12546), .ZN(P3_U3222) );
  AOI211_X1 U14239 ( .C1(n15964), .C2(n12550), .A(n12549), .B(n12548), .ZN(
        n12555) );
  INV_X1 U14240 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n12551) );
  NOR2_X1 U14241 ( .A1(n15973), .A2(n12551), .ZN(n12552) );
  AOI21_X1 U14242 ( .B1(n12655), .B2(n14558), .A(n12552), .ZN(n12553) );
  OAI21_X1 U14243 ( .B1(n12555), .B2(n15971), .A(n12553), .ZN(P2_U3472) );
  AOI22_X1 U14244 ( .A1(n12655), .A2(n14510), .B1(n15968), .B2(
        P2_REG1_REG_14__SCAN_IN), .ZN(n12554) );
  OAI21_X1 U14245 ( .B1(n12555), .B2(n15968), .A(n12554), .ZN(P2_U3513) );
  AOI22_X1 U14246 ( .A1(n15900), .A2(n13014), .B1(n13019), .B2(n14736), .ZN(
        n12556) );
  XNOR2_X1 U14247 ( .A(n12556), .B(n13025), .ZN(n12909) );
  AOI22_X1 U14248 ( .A1(n15900), .A2(n13019), .B1(n13018), .B2(n14736), .ZN(
        n12910) );
  XNOR2_X1 U14249 ( .A(n12909), .B(n12910), .ZN(n12561) );
  AOI21_X1 U14250 ( .B1(n12561), .B2(n12560), .A(n12908), .ZN(n12570) );
  OAI21_X1 U14251 ( .B1(n16019), .B2(n12563), .A(n12562), .ZN(n12564) );
  AOI21_X1 U14252 ( .B1(n15980), .B2(n12565), .A(n12564), .ZN(n12566) );
  OAI21_X1 U14253 ( .B1(n12567), .B2(n16031), .A(n12566), .ZN(n12568) );
  AOI21_X1 U14254 ( .B1(n15900), .B2(n16027), .A(n12568), .ZN(n12569) );
  OAI21_X1 U14255 ( .B1(n12570), .B2(n16022), .A(n12569), .ZN(P1_U3236) );
  INV_X1 U14256 ( .A(n12571), .ZN(n12586) );
  NAND2_X1 U14257 ( .A1(n12572), .A2(n12580), .ZN(n12574) );
  AND2_X1 U14258 ( .A1(n12576), .A2(n12574), .ZN(n12578) );
  XNOR2_X1 U14259 ( .A(n15871), .B(n13041), .ZN(n12714) );
  XNOR2_X1 U14260 ( .A(n12714), .B(n12573), .ZN(n12577) );
  AND2_X1 U14261 ( .A1(n12577), .A2(n12574), .ZN(n12575) );
  NAND2_X1 U14262 ( .A1(n12576), .A2(n12575), .ZN(n12716) );
  OAI211_X1 U14263 ( .C1(n12578), .C2(n12577), .A(n13168), .B(n12716), .ZN(
        n12584) );
  OAI22_X1 U14264 ( .A1(n13195), .A2(n12580), .B1(n12579), .B2(n13178), .ZN(
        n12581) );
  AOI211_X1 U14265 ( .C1(n13191), .C2(n13213), .A(n12582), .B(n12581), .ZN(
        n12583) );
  OAI211_X1 U14266 ( .C1(n12586), .C2(n12585), .A(n12584), .B(n12583), .ZN(
        P3_U3157) );
  NAND2_X1 U14267 ( .A1(n12588), .A2(n12587), .ZN(n12589) );
  NAND2_X1 U14268 ( .A1(n12590), .A2(n12589), .ZN(n14515) );
  AND2_X1 U14269 ( .A1(n14179), .A2(n14152), .ZN(n12591) );
  AOI21_X1 U14270 ( .B1(n14177), .B2(n14153), .A(n12591), .ZN(n12858) );
  XNOR2_X1 U14271 ( .A(n12593), .B(n12592), .ZN(n12594) );
  NAND2_X1 U14272 ( .A1(n12594), .A2(n15797), .ZN(n12595) );
  OAI211_X1 U14273 ( .C1(n14515), .C2(n14423), .A(n12858), .B(n12595), .ZN(
        n14517) );
  NAND2_X1 U14274 ( .A1(n14517), .A2(n15721), .ZN(n12601) );
  INV_X1 U14275 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12596) );
  OAI22_X1 U14276 ( .A1(n15721), .A2(n12596), .B1(n12857), .B2(n15714), .ZN(
        n12599) );
  OAI211_X1 U14277 ( .C1(n12863), .C2(n12597), .A(n7209), .B(n12678), .ZN(
        n14513) );
  NOR2_X1 U14278 ( .A1(n14513), .A2(n15717), .ZN(n12598) );
  AOI211_X1 U14279 ( .C1(n15917), .C2(n14512), .A(n12599), .B(n12598), .ZN(
        n12600) );
  OAI211_X1 U14280 ( .C1(n14515), .C2(n14431), .A(n12601), .B(n12600), .ZN(
        P2_U3249) );
  NAND2_X1 U14281 ( .A1(n12838), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n12602) );
  OAI21_X1 U14282 ( .B1(n12838), .B2(P2_REG2_REG_14__SCAN_IN), .A(n12602), 
        .ZN(n12610) );
  NAND2_X1 U14283 ( .A1(n12604), .A2(n12603), .ZN(n12605) );
  NAND2_X1 U14284 ( .A1(n12606), .A2(n12605), .ZN(n15351) );
  INV_X1 U14285 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12607) );
  MUX2_X1 U14286 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n12607), .S(n12616), .Z(
        n15352) );
  NAND2_X1 U14287 ( .A1(n15358), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12608) );
  NAND2_X1 U14288 ( .A1(n15349), .A2(n12608), .ZN(n12609) );
  NOR2_X1 U14289 ( .A1(n12609), .A2(n12610), .ZN(n12836) );
  AOI21_X1 U14290 ( .B1(n12610), .B2(n12609), .A(n12836), .ZN(n12623) );
  NAND2_X1 U14291 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n12611)
         );
  OAI21_X1 U14292 ( .B1(n15322), .B2(n12613), .A(n12611), .ZN(n12621) );
  NOR2_X1 U14293 ( .A1(n12613), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n12612) );
  AOI21_X1 U14294 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n12613), .A(n12612), 
        .ZN(n12619) );
  OAI21_X1 U14295 ( .B1(n12615), .B2(P2_REG1_REG_12__SCAN_IN), .A(n12614), 
        .ZN(n15354) );
  MUX2_X1 U14296 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n12617), .S(n12616), .Z(
        n15355) );
  AOI211_X1 U14297 ( .C1(n12619), .C2(n12618), .A(n15368), .B(n12834), .ZN(
        n12620) );
  AOI211_X1 U14298 ( .C1(n15271), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n12621), 
        .B(n12620), .ZN(n12622) );
  OAI21_X1 U14299 ( .B1(n12623), .B2(n15364), .A(n12622), .ZN(P2_U3228) );
  NAND2_X1 U14300 ( .A1(n15926), .A2(n14649), .ZN(n12626) );
  INV_X1 U14301 ( .A(n12631), .ZN(n12627) );
  OAI21_X1 U14302 ( .B1(n7323), .B2(n12627), .A(n12865), .ZN(n15954) );
  NAND2_X1 U14303 ( .A1(n12628), .A2(n8112), .ZN(n12630) );
  NAND2_X1 U14304 ( .A1(n15926), .A2(n14734), .ZN(n12629) );
  XOR2_X1 U14305 ( .A(n12877), .B(n12631), .Z(n15956) );
  NAND2_X1 U14306 ( .A1(n15956), .A2(n15083), .ZN(n12641) );
  OR2_X1 U14307 ( .A1(n14649), .A2(n15041), .ZN(n12633) );
  NAND2_X1 U14308 ( .A1(n15058), .A2(n15076), .ZN(n12632) );
  NAND2_X1 U14309 ( .A1(n12633), .A2(n12632), .ZN(n15948) );
  INV_X1 U14310 ( .A(n14609), .ZN(n12634) );
  AOI22_X1 U14311 ( .A1(n15021), .A2(n15948), .B1(n12634), .B2(n15043), .ZN(
        n12635) );
  OAI21_X1 U14312 ( .B1(n14836), .B2(n15021), .A(n12635), .ZN(n12639) );
  OR2_X1 U14313 ( .A1(n15950), .A2(n12636), .ZN(n15070) );
  NAND2_X1 U14314 ( .A1(n12636), .A2(n15950), .ZN(n12637) );
  NAND3_X1 U14315 ( .A1(n15070), .A2(n15071), .A3(n12637), .ZN(n15951) );
  NOR2_X1 U14316 ( .A1(n15951), .A2(n15086), .ZN(n12638) );
  AOI211_X1 U14317 ( .C1(n15066), .C2(n15950), .A(n12639), .B(n12638), .ZN(
        n12640) );
  OAI211_X1 U14318 ( .C1(n15954), .C2(n15069), .A(n12641), .B(n12640), .ZN(
        P1_U3279) );
  XNOR2_X1 U14319 ( .A(n12655), .B(n14072), .ZN(n12644) );
  OR2_X1 U14320 ( .A1(n12642), .A2(n14308), .ZN(n12643) );
  NAND2_X1 U14321 ( .A1(n12644), .A2(n12643), .ZN(n12745) );
  OAI21_X1 U14322 ( .B1(n12644), .B2(n12643), .A(n12745), .ZN(n12649) );
  OAI21_X2 U14323 ( .B1(n12647), .B2(n12646), .A(n12645), .ZN(n12648) );
  AOI21_X1 U14324 ( .B1(n12649), .B2(n12648), .A(n12747), .ZN(n12657) );
  NOR2_X1 U14325 ( .A1(n14092), .A2(n12650), .ZN(n12654) );
  OAI22_X1 U14326 ( .A1(n14157), .A2(n12652), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12651), .ZN(n12653) );
  AOI211_X1 U14327 ( .C1(n12655), .C2(n14159), .A(n12654), .B(n12653), .ZN(
        n12656) );
  OAI21_X1 U14328 ( .B1(n12657), .B2(n14163), .A(n12656), .ZN(P2_U3187) );
  NAND2_X1 U14329 ( .A1(n12658), .A2(n12773), .ZN(n12659) );
  NAND3_X1 U14330 ( .A1(n12660), .A2(n13604), .A3(n12659), .ZN(n12662) );
  AOI22_X1 U14331 ( .A1(n13211), .A2(n13606), .B1(n13609), .B2(n13213), .ZN(
        n12661) );
  OR2_X1 U14332 ( .A1(n12663), .A2(n12773), .ZN(n12664) );
  NAND2_X1 U14333 ( .A1(n12735), .A2(n12664), .ZN(n12795) );
  AOI22_X1 U14334 ( .A1(n13635), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n13634), 
        .B2(n12783), .ZN(n12665) );
  OAI21_X1 U14335 ( .B1(n12803), .B2(n13637), .A(n12665), .ZN(n12666) );
  AOI21_X1 U14336 ( .B1(n12795), .B2(n13639), .A(n12666), .ZN(n12667) );
  OAI21_X1 U14337 ( .B1(n13635), .B2(n12796), .A(n12667), .ZN(P3_U3221) );
  INV_X1 U14338 ( .A(n12668), .ZN(n12728) );
  OAI222_X1 U14339 ( .A1(n14592), .A2(n12670), .B1(n14578), .B2(n12728), .C1(
        n12669), .C2(P2_U3088), .ZN(P2_U3306) );
  XNOR2_X1 U14340 ( .A(n12672), .B(n12671), .ZN(n12673) );
  OR2_X1 U14341 ( .A1(n12673), .A2(n15702), .ZN(n12675) );
  AND2_X1 U14342 ( .A1(n14178), .A2(n14152), .ZN(n12674) );
  AOI21_X1 U14343 ( .B1(n14176), .B2(n14153), .A(n12674), .ZN(n14104) );
  NAND2_X1 U14344 ( .A1(n12675), .A2(n14104), .ZN(n14505) );
  INV_X1 U14345 ( .A(n14505), .ZN(n12686) );
  XNOR2_X1 U14346 ( .A(n12677), .B(n12676), .ZN(n14506) );
  INV_X1 U14347 ( .A(n14557), .ZN(n14109) );
  NAND2_X1 U14348 ( .A1(n14557), .A2(n12678), .ZN(n12679) );
  NAND2_X1 U14349 ( .A1(n12679), .A2(n7209), .ZN(n12680) );
  NOR2_X1 U14350 ( .A1(n14426), .A2(n12680), .ZN(n14504) );
  NAND2_X1 U14351 ( .A1(n14504), .A2(n15934), .ZN(n12683) );
  INV_X1 U14352 ( .A(n12681), .ZN(n14106) );
  AOI22_X1 U14353 ( .A1(n15947), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14106), 
        .B2(n15936), .ZN(n12682) );
  OAI211_X1 U14354 ( .C1(n14109), .C2(n15940), .A(n12683), .B(n12682), .ZN(
        n12684) );
  AOI21_X1 U14355 ( .B1(n14506), .B2(n15807), .A(n12684), .ZN(n12685) );
  OAI21_X1 U14356 ( .B1(n15947), .B2(n12686), .A(n12685), .ZN(P2_U3248) );
  NOR2_X1 U14357 ( .A1(n7941), .A2(n12688), .ZN(n12690) );
  INV_X1 U14358 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12691) );
  MUX2_X1 U14359 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n12691), .S(n13252), .Z(
        n12704) );
  INV_X1 U14360 ( .A(n12704), .ZN(n12693) );
  INV_X1 U14361 ( .A(n13261), .ZN(n12692) );
  AOI21_X1 U14362 ( .B1(n12694), .B2(n12693), .A(n12692), .ZN(n12713) );
  NOR2_X1 U14363 ( .A1(n7941), .A2(n12695), .ZN(n12697) );
  INV_X1 U14364 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12801) );
  NAND2_X1 U14365 ( .A1(n12698), .A2(n12801), .ZN(n12699) );
  NAND2_X1 U14366 ( .A1(n13252), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n13253) );
  AND2_X1 U14367 ( .A1(n12699), .A2(n13253), .ZN(n12703) );
  OAI21_X1 U14368 ( .B1(n7772), .B2(n12703), .A(n13249), .ZN(n12711) );
  INV_X1 U14369 ( .A(n12700), .ZN(n12701) );
  MUX2_X1 U14370 ( .A(n12704), .B(n12703), .S(n7166), .Z(n12706) );
  INV_X1 U14371 ( .A(n13257), .ZN(n12705) );
  OAI211_X1 U14372 ( .C1(n12707), .C2(n12706), .A(n12705), .B(n15638), .ZN(
        n12709) );
  INV_X1 U14373 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13858) );
  NOR2_X1 U14374 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13858), .ZN(n12782) );
  AOI21_X1 U14375 ( .B1(n15246), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12782), 
        .ZN(n12708) );
  OAI211_X1 U14376 ( .C1(n15641), .C2(n13252), .A(n12709), .B(n12708), .ZN(
        n12710) );
  AOI21_X1 U14377 ( .B1(n12711), .B2(n13422), .A(n12710), .ZN(n12712) );
  OAI21_X1 U14378 ( .B1(n12713), .B2(n15636), .A(n12712), .ZN(P3_U3194) );
  NAND2_X1 U14379 ( .A1(n13214), .A2(n12714), .ZN(n12715) );
  NAND2_X1 U14380 ( .A1(n12716), .A2(n12715), .ZN(n12775) );
  XNOR2_X1 U14381 ( .A(n12717), .B(n13103), .ZN(n12774) );
  XOR2_X1 U14382 ( .A(n12775), .B(n12774), .Z(n12725) );
  AOI21_X1 U14383 ( .B1(n13212), .B2(n13191), .A(n12718), .ZN(n12723) );
  NAND2_X1 U14384 ( .A1(n13197), .A2(n12776), .ZN(n12722) );
  NAND2_X1 U14385 ( .A1(n13190), .A2(n12719), .ZN(n12721) );
  NAND2_X1 U14386 ( .A1(n13214), .A2(n13172), .ZN(n12720) );
  NAND4_X1 U14387 ( .A1(n12723), .A2(n12722), .A3(n12721), .A4(n12720), .ZN(
        n12724) );
  AOI21_X1 U14388 ( .B1(n12725), .B2(n13168), .A(n12724), .ZN(n12726) );
  INV_X1 U14389 ( .A(n12726), .ZN(P3_U3176) );
  OAI211_X1 U14390 ( .C1(n12731), .C2(n12806), .A(n12730), .B(n13604), .ZN(
        n12733) );
  AOI22_X1 U14391 ( .A1(n13212), .A2(n13609), .B1(n13606), .B2(n13210), .ZN(
        n12732) );
  NAND2_X1 U14392 ( .A1(n12733), .A2(n12732), .ZN(n12827) );
  INV_X1 U14393 ( .A(n12827), .ZN(n12742) );
  NAND2_X1 U14394 ( .A1(n12735), .A2(n12734), .ZN(n12738) );
  NAND2_X1 U14395 ( .A1(n12738), .A2(n12737), .ZN(n12736) );
  OAI21_X1 U14396 ( .B1(n12738), .B2(n12737), .A(n12736), .ZN(n12828) );
  AOI22_X1 U14397 ( .A1(n13635), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n13634), 
        .B2(n12813), .ZN(n12739) );
  OAI21_X1 U14398 ( .B1(n12833), .B2(n13637), .A(n12739), .ZN(n12740) );
  AOI21_X1 U14399 ( .B1(n12828), .B2(n13639), .A(n12740), .ZN(n12741) );
  OAI21_X1 U14400 ( .B1(n12742), .B2(n13635), .A(n12741), .ZN(P3_U3220) );
  INV_X1 U14401 ( .A(n12743), .ZN(n12744) );
  OAI222_X1 U14402 ( .A1(n7456), .A2(P3_U3151), .B1(n13993), .B2(n12744), .C1(
        n13812), .C2(n13787), .ZN(P3_U3269) );
  INV_X1 U14403 ( .A(n12745), .ZN(n12746) );
  NAND2_X1 U14404 ( .A1(n14360), .A2(n14179), .ZN(n12849) );
  XNOR2_X1 U14405 ( .A(n15960), .B(n14072), .ZN(n12848) );
  XOR2_X1 U14406 ( .A(n12849), .B(n12848), .Z(n12852) );
  XNOR2_X1 U14407 ( .A(n12853), .B(n12852), .ZN(n12753) );
  AOI22_X1 U14408 ( .A1(n14095), .A2(n12748), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12749) );
  OAI21_X1 U14409 ( .B1(n12750), .B2(n14092), .A(n12749), .ZN(n12751) );
  AOI21_X1 U14410 ( .B1(n15960), .B2(n14159), .A(n12751), .ZN(n12752) );
  OAI21_X1 U14411 ( .B1(n12753), .B2(n14163), .A(n12752), .ZN(P2_U3213) );
  INV_X1 U14412 ( .A(n12758), .ZN(n12756) );
  NAND2_X1 U14413 ( .A1(n14576), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12755) );
  OAI211_X1 U14414 ( .C1(n12756), .C2(n14578), .A(n12755), .B(n12754), .ZN(
        P2_U3304) );
  NAND2_X1 U14415 ( .A1(n12758), .A2(n12757), .ZN(n12760) );
  OAI211_X1 U14416 ( .C1(n12761), .C2(n15235), .A(n12760), .B(n12759), .ZN(
        P1_U3332) );
  OAI211_X1 U14417 ( .C1(n12764), .C2(n12763), .A(n12762), .B(n13604), .ZN(
        n12766) );
  AOI22_X1 U14418 ( .A1(n13211), .A2(n13609), .B1(n13606), .B2(n13209), .ZN(
        n12765) );
  AND2_X1 U14419 ( .A1(n12766), .A2(n12765), .ZN(n13700) );
  OAI21_X1 U14420 ( .B1(n12769), .B2(n12768), .A(n12767), .ZN(n13699) );
  AOI22_X1 U14421 ( .A1(n13635), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n13634), 
        .B2(n13079), .ZN(n12770) );
  OAI21_X1 U14422 ( .B1(n13702), .B2(n13637), .A(n12770), .ZN(n12771) );
  AOI21_X1 U14423 ( .B1(n13699), .B2(n13639), .A(n12771), .ZN(n12772) );
  OAI21_X1 U14424 ( .B1(n13635), .B2(n13700), .A(n12772), .ZN(P3_U3219) );
  XNOR2_X1 U14425 ( .A(n12773), .B(n13041), .ZN(n12805) );
  NAND2_X1 U14426 ( .A1(n13213), .A2(n12776), .ZN(n12777) );
  MUX2_X1 U14427 ( .A(n12778), .B(n12777), .S(n13041), .Z(n12779) );
  INV_X1 U14428 ( .A(n12809), .ZN(n12780) );
  AOI21_X1 U14429 ( .B1(n12805), .B2(n12781), .A(n12780), .ZN(n12790) );
  AOI21_X1 U14430 ( .B1(n13211), .B2(n13191), .A(n12782), .ZN(n12785) );
  NAND2_X1 U14431 ( .A1(n13190), .A2(n12783), .ZN(n12784) );
  OAI211_X1 U14432 ( .C1(n12786), .C2(n13195), .A(n12785), .B(n12784), .ZN(
        n12787) );
  AOI21_X1 U14433 ( .B1(n13197), .B2(n12788), .A(n12787), .ZN(n12789) );
  OAI21_X1 U14434 ( .B1(n12790), .B2(n13200), .A(n12789), .ZN(P3_U3164) );
  INV_X1 U14435 ( .A(n12791), .ZN(n12793) );
  OAI222_X1 U14436 ( .A1(n14592), .A2(n12794), .B1(n14578), .B2(n12793), .C1(
        n12792), .C2(P2_U3088), .ZN(P2_U3305) );
  NAND2_X1 U14437 ( .A1(n12795), .A2(n15891), .ZN(n12797) );
  AND2_X1 U14438 ( .A1(n12797), .A2(n12796), .ZN(n12800) );
  INV_X1 U14439 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n12798) );
  MUX2_X1 U14440 ( .A(n12800), .B(n12798), .S(n15895), .Z(n12799) );
  OAI21_X1 U14441 ( .B1(n12803), .B2(n13767), .A(n12799), .ZN(P3_U3426) );
  MUX2_X1 U14442 ( .A(n12801), .B(n12800), .S(n15894), .Z(n12802) );
  OAI21_X1 U14443 ( .B1(n12803), .B2(n13694), .A(n12802), .ZN(P3_U3471) );
  NAND2_X1 U14444 ( .A1(n12805), .A2(n12804), .ZN(n12807) );
  AND2_X1 U14445 ( .A1(n12809), .A2(n12807), .ZN(n12810) );
  XNOR2_X1 U14446 ( .A(n12806), .B(n13041), .ZN(n13037) );
  AND2_X1 U14447 ( .A1(n13037), .A2(n12807), .ZN(n12808) );
  OAI211_X1 U14448 ( .C1(n12810), .C2(n13037), .A(n13168), .B(n13040), .ZN(
        n12815) );
  INV_X1 U14449 ( .A(n13210), .ZN(n13194) );
  NOR2_X1 U14450 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8502), .ZN(n13266) );
  AOI21_X1 U14451 ( .B1(n13212), .B2(n13172), .A(n13266), .ZN(n12811) );
  OAI21_X1 U14452 ( .B1(n13194), .B2(n13174), .A(n12811), .ZN(n12812) );
  AOI21_X1 U14453 ( .B1(n12813), .B2(n13190), .A(n12812), .ZN(n12814) );
  OAI211_X1 U14454 ( .C1(n13178), .C2(n12833), .A(n12815), .B(n12814), .ZN(
        P3_U3174) );
  OAI211_X1 U14455 ( .C1(n12818), .C2(n12817), .A(n12816), .B(n13604), .ZN(
        n12820) );
  AOI22_X1 U14456 ( .A1(n13609), .A2(n13210), .B1(n13608), .B2(n13606), .ZN(
        n12819) );
  AND2_X1 U14457 ( .A1(n12820), .A2(n12819), .ZN(n13696) );
  OAI21_X1 U14458 ( .B1(n12823), .B2(n12822), .A(n12821), .ZN(n13695) );
  AOI22_X1 U14459 ( .A1(n13635), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n13634), 
        .B2(n13189), .ZN(n12824) );
  OAI21_X1 U14460 ( .B1(n13698), .B2(n13637), .A(n12824), .ZN(n12825) );
  AOI21_X1 U14461 ( .B1(n13695), .B2(n13639), .A(n12825), .ZN(n12826) );
  OAI21_X1 U14462 ( .B1(n13635), .B2(n13696), .A(n12826), .ZN(P3_U3218) );
  INV_X1 U14463 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12829) );
  AOI21_X1 U14464 ( .B1(n15891), .B2(n12828), .A(n12827), .ZN(n12831) );
  MUX2_X1 U14465 ( .A(n12829), .B(n12831), .S(n15898), .Z(n12830) );
  OAI21_X1 U14466 ( .B1(n13767), .B2(n12833), .A(n12830), .ZN(P3_U3429) );
  INV_X1 U14467 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13251) );
  MUX2_X1 U14468 ( .A(n13251), .B(n12831), .S(n15894), .Z(n12832) );
  OAI21_X1 U14469 ( .B1(n13694), .B2(n12833), .A(n12832), .ZN(P3_U3472) );
  INV_X1 U14470 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15969) );
  AOI211_X1 U14471 ( .C1(n12835), .C2(n15969), .A(n15284), .B(n15368), .ZN(
        n12845) );
  INV_X1 U14472 ( .A(n12836), .ZN(n12837) );
  OAI21_X1 U14473 ( .B1(n12838), .B2(P2_REG2_REG_14__SCAN_IN), .A(n12837), 
        .ZN(n15288) );
  XOR2_X1 U14474 ( .A(n12839), .B(n15288), .Z(n12840) );
  NOR2_X1 U14475 ( .A1(n12447), .A2(n12840), .ZN(n15290) );
  AOI211_X1 U14476 ( .C1(n12447), .C2(n12840), .A(n15290), .B(n15364), .ZN(
        n12844) );
  NAND2_X1 U14477 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n12842)
         );
  NAND2_X1 U14478 ( .A1(n15271), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n12841) );
  OAI211_X1 U14479 ( .C1(n15322), .C2(n15289), .A(n12842), .B(n12841), .ZN(
        n12843) );
  OR3_X1 U14480 ( .A1(n12845), .A2(n12844), .A3(n12843), .ZN(P2_U3229) );
  XNOR2_X1 U14481 ( .A(n14512), .B(n14038), .ZN(n12847) );
  AND2_X1 U14482 ( .A1(n14178), .A2(n14360), .ZN(n12846) );
  NOR2_X1 U14483 ( .A1(n12847), .A2(n12846), .ZN(n14001) );
  AOI21_X1 U14484 ( .B1(n12847), .B2(n12846), .A(n14001), .ZN(n12855) );
  INV_X1 U14485 ( .A(n12848), .ZN(n12851) );
  INV_X1 U14486 ( .A(n12849), .ZN(n12850) );
  OAI21_X1 U14487 ( .B1(n12855), .B2(n12854), .A(n14003), .ZN(n12856) );
  NAND2_X1 U14488 ( .A1(n12856), .A2(n14102), .ZN(n12862) );
  INV_X1 U14489 ( .A(n12857), .ZN(n12860) );
  NAND2_X1 U14490 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n15297)
         );
  OAI21_X1 U14491 ( .B1(n14157), .B2(n12858), .A(n15297), .ZN(n12859) );
  AOI21_X1 U14492 ( .B1(n12860), .B2(n14155), .A(n12859), .ZN(n12861) );
  OAI211_X1 U14493 ( .C1(n12863), .C2(n14135), .A(n12862), .B(n12861), .ZN(
        P2_U3198) );
  NAND2_X1 U14494 ( .A1(n15950), .A2(n15979), .ZN(n12864) );
  INV_X1 U14495 ( .A(n15977), .ZN(n16017) );
  NAND2_X1 U14496 ( .A1(n15189), .A2(n16017), .ZN(n12866) );
  NAND2_X1 U14497 ( .A1(n16026), .A2(n15057), .ZN(n12867) );
  OR2_X1 U14498 ( .A1(n15154), .A2(n14984), .ZN(n12870) );
  INV_X1 U14499 ( .A(n14942), .ZN(n14939) );
  INV_X1 U14500 ( .A(n14730), .ZN(n14926) );
  NAND2_X1 U14501 ( .A1(n15106), .A2(n8230), .ZN(n12873) );
  XNOR2_X1 U14502 ( .A(n12873), .B(n12872), .ZN(n15103) );
  INV_X1 U14503 ( .A(n15979), .ZN(n12874) );
  NOR2_X1 U14504 ( .A1(n15950), .A2(n12874), .ZN(n12876) );
  NAND2_X1 U14505 ( .A1(n15950), .A2(n12874), .ZN(n12875) );
  OR2_X1 U14506 ( .A1(n15077), .A2(n14606), .ZN(n12878) );
  NAND2_X1 U14507 ( .A1(n16008), .A2(n16017), .ZN(n12879) );
  INV_X1 U14508 ( .A(n15057), .ZN(n12880) );
  NAND2_X1 U14509 ( .A1(n16026), .A2(n12880), .ZN(n12882) );
  NOR2_X1 U14510 ( .A1(n16026), .A2(n12880), .ZN(n12881) );
  INV_X1 U14511 ( .A(n15026), .ZN(n12883) );
  INV_X1 U14512 ( .A(n15170), .ZN(n15009) );
  INV_X1 U14513 ( .A(n14984), .ZN(n14699) );
  NAND2_X1 U14514 ( .A1(n14943), .A2(n14942), .ZN(n14941) );
  OAI21_X1 U14515 ( .B1(n14949), .B2(n14958), .A(n14941), .ZN(n14928) );
  NAND2_X1 U14516 ( .A1(n14866), .A2(n12886), .ZN(n12888) );
  XNOR2_X1 U14517 ( .A(n12888), .B(n12872), .ZN(n15095) );
  NAND2_X1 U14518 ( .A1(n15095), .A2(n15083), .ZN(n12898) );
  NAND2_X1 U14519 ( .A1(n15161), .A2(n14999), .ZN(n14981) );
  NAND2_X1 U14520 ( .A1(n14932), .A2(n15128), .ZN(n14915) );
  OAI21_X1 U14521 ( .B1(n15099), .B2(n14869), .A(n14852), .ZN(n15096) );
  NAND2_X1 U14522 ( .A1(n14727), .A2(n15075), .ZN(n15098) );
  INV_X1 U14523 ( .A(n12889), .ZN(n12890) );
  NAND2_X1 U14524 ( .A1(n15043), .A2(n12890), .ZN(n12891) );
  OAI211_X1 U14525 ( .C1(n15096), .C2(n15063), .A(n15098), .B(n12891), .ZN(
        n12896) );
  NOR2_X1 U14526 ( .A1(n15099), .A2(n15078), .ZN(n12895) );
  AOI21_X1 U14527 ( .B1(n15379), .B2(P1_B_REG_SCAN_IN), .A(n15042), .ZN(n14854) );
  NAND2_X1 U14528 ( .A1(n14725), .A2(n14854), .ZN(n15097) );
  OAI22_X1 U14529 ( .A1(n15021), .A2(n12893), .B1(n15097), .B2(n12892), .ZN(
        n12894) );
  AOI211_X1 U14530 ( .C1(n12896), .C2(n15021), .A(n12895), .B(n12894), .ZN(
        n12897) );
  OAI211_X1 U14531 ( .C1(n15103), .C2(n15069), .A(n12898), .B(n12897), .ZN(
        P1_U3356) );
  OAI222_X1 U14532 ( .A1(n14592), .A2(n12900), .B1(n14578), .B2(n12899), .C1(
        n9420), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U14533 ( .A(SI_28_), .ZN(n12904) );
  INV_X1 U14534 ( .A(n12901), .ZN(n12902) );
  OAI222_X1 U14535 ( .A1(n13787), .A2(n12904), .B1(P3_U3151), .B2(n12903), 
        .C1(n13993), .C2(n12902), .ZN(P3_U3267) );
  INV_X1 U14536 ( .A(n12905), .ZN(n14587) );
  OAI222_X1 U14537 ( .A1(n15235), .A2(n12907), .B1(n15233), .B2(n14587), .C1(
        n12906), .C2(P1_U3086), .ZN(P1_U3330) );
  NAND2_X1 U14538 ( .A1(n12915), .A2(n13014), .ZN(n12912) );
  NAND2_X1 U14539 ( .A1(n14735), .A2(n13019), .ZN(n12911) );
  NAND2_X1 U14540 ( .A1(n12912), .A2(n12911), .ZN(n12913) );
  XNOR2_X1 U14541 ( .A(n12913), .B(n13025), .ZN(n12916) );
  AND2_X1 U14542 ( .A1(n13018), .A2(n14735), .ZN(n12914) );
  AOI21_X1 U14543 ( .B1(n12915), .B2(n12999), .A(n12914), .ZN(n12917) );
  XNOR2_X1 U14544 ( .A(n12916), .B(n12917), .ZN(n14646) );
  NOR2_X1 U14545 ( .A1(n14649), .A2(n13023), .ZN(n12920) );
  AOI21_X1 U14546 ( .B1(n12921), .B2(n13019), .A(n12920), .ZN(n12923) );
  AOI22_X1 U14547 ( .A1(n12921), .A2(n13014), .B1(n12999), .B2(n14734), .ZN(
        n12922) );
  XNOR2_X1 U14548 ( .A(n12922), .B(n13025), .ZN(n12924) );
  XOR2_X1 U14549 ( .A(n12923), .B(n12924), .Z(n14685) );
  OR2_X1 U14550 ( .A1(n12924), .A2(n12923), .ZN(n12925) );
  AOI22_X1 U14551 ( .A1(n15950), .A2(n12999), .B1(n13018), .B2(n15979), .ZN(
        n12930) );
  NAND2_X1 U14552 ( .A1(n15950), .A2(n13014), .ZN(n12927) );
  NAND2_X1 U14553 ( .A1(n15979), .A2(n12999), .ZN(n12926) );
  NAND2_X1 U14554 ( .A1(n12927), .A2(n12926), .ZN(n12928) );
  XNOR2_X1 U14555 ( .A(n12928), .B(n13025), .ZN(n12932) );
  XOR2_X1 U14556 ( .A(n12930), .B(n12932), .Z(n14604) );
  INV_X1 U14557 ( .A(n12930), .ZN(n12931) );
  NAND2_X1 U14558 ( .A1(n15077), .A2(n13014), .ZN(n12935) );
  NAND2_X1 U14559 ( .A1(n15058), .A2(n12999), .ZN(n12934) );
  NAND2_X1 U14560 ( .A1(n12935), .A2(n12934), .ZN(n12936) );
  XNOR2_X1 U14561 ( .A(n12936), .B(n13025), .ZN(n12937) );
  AOI22_X1 U14562 ( .A1(n15077), .A2(n13019), .B1(n13018), .B2(n15058), .ZN(
        n15976) );
  NAND2_X1 U14563 ( .A1(n16008), .A2(n13014), .ZN(n12940) );
  NAND2_X1 U14564 ( .A1(n15977), .A2(n13019), .ZN(n12939) );
  NAND2_X1 U14565 ( .A1(n12940), .A2(n12939), .ZN(n12941) );
  XNOR2_X1 U14566 ( .A(n12941), .B(n13025), .ZN(n12942) );
  AOI22_X1 U14567 ( .A1(n16008), .A2(n13019), .B1(n13018), .B2(n15977), .ZN(
        n12943) );
  XNOR2_X1 U14568 ( .A(n12942), .B(n12943), .ZN(n16007) );
  INV_X1 U14569 ( .A(n12942), .ZN(n12944) );
  NAND2_X1 U14570 ( .A1(n12944), .A2(n12943), .ZN(n12945) );
  NAND2_X1 U14571 ( .A1(n16026), .A2(n13014), .ZN(n12947) );
  NAND2_X1 U14572 ( .A1(n15057), .A2(n13019), .ZN(n12946) );
  NAND2_X1 U14573 ( .A1(n12947), .A2(n12946), .ZN(n12948) );
  XNOR2_X1 U14574 ( .A(n12948), .B(n13025), .ZN(n12949) );
  AOI22_X1 U14575 ( .A1(n16026), .A2(n13019), .B1(n13018), .B2(n15057), .ZN(
        n12950) );
  XNOR2_X1 U14576 ( .A(n12949), .B(n12950), .ZN(n16020) );
  INV_X1 U14577 ( .A(n12949), .ZN(n12951) );
  NAND2_X1 U14578 ( .A1(n12951), .A2(n12950), .ZN(n12952) );
  OAI22_X1 U14579 ( .A1(n15018), .A2(n13024), .B1(n16018), .B2(n13023), .ZN(
        n12954) );
  OAI22_X1 U14580 ( .A1(n15018), .A2(n7171), .B1(n16018), .B2(n13024), .ZN(
        n12953) );
  XNOR2_X1 U14581 ( .A(n12953), .B(n13025), .ZN(n12955) );
  XOR2_X1 U14582 ( .A(n12954), .B(n12955), .Z(n14705) );
  OR2_X1 U14583 ( .A1(n12955), .A2(n12954), .ZN(n12956) );
  NAND2_X1 U14584 ( .A1(n15170), .A2(n13014), .ZN(n12958) );
  NAND2_X1 U14585 ( .A1(n15031), .A2(n12999), .ZN(n12957) );
  NAND2_X1 U14586 ( .A1(n12958), .A2(n12957), .ZN(n12959) );
  XNOR2_X1 U14587 ( .A(n12959), .B(n13025), .ZN(n12960) );
  AOI22_X1 U14588 ( .A1(n15170), .A2(n12999), .B1(n13018), .B2(n15031), .ZN(
        n12961) );
  XNOR2_X1 U14589 ( .A(n12960), .B(n12961), .ZN(n14629) );
  INV_X1 U14590 ( .A(n12960), .ZN(n12962) );
  NAND2_X1 U14591 ( .A1(n12962), .A2(n12961), .ZN(n12963) );
  NOR2_X1 U14592 ( .A1(n15000), .A2(n13023), .ZN(n12964) );
  AOI21_X1 U14593 ( .B1(n14988), .B2(n13019), .A(n12964), .ZN(n12969) );
  NAND2_X1 U14594 ( .A1(n14988), .A2(n13014), .ZN(n12966) );
  OR2_X1 U14595 ( .A1(n15000), .A2(n13024), .ZN(n12965) );
  NAND2_X1 U14596 ( .A1(n12966), .A2(n12965), .ZN(n12967) );
  XNOR2_X1 U14597 ( .A(n12967), .B(n13025), .ZN(n12968) );
  XOR2_X1 U14598 ( .A(n12969), .B(n12968), .Z(n14676) );
  INV_X1 U14599 ( .A(n12968), .ZN(n12970) );
  OR2_X1 U14600 ( .A1(n12970), .A2(n12969), .ZN(n12971) );
  AOI22_X1 U14601 ( .A1(n15154), .A2(n13014), .B1(n13019), .B2(n14984), .ZN(
        n12972) );
  XNOR2_X1 U14602 ( .A(n12972), .B(n13025), .ZN(n12975) );
  AOI22_X1 U14603 ( .A1(n15154), .A2(n12999), .B1(n13018), .B2(n14984), .ZN(
        n12974) );
  XNOR2_X1 U14604 ( .A(n12975), .B(n12974), .ZN(n14639) );
  INV_X1 U14605 ( .A(n14639), .ZN(n12973) );
  NAND2_X1 U14606 ( .A1(n12975), .A2(n12974), .ZN(n12976) );
  NAND2_X1 U14607 ( .A1(n14959), .A2(n13014), .ZN(n12978) );
  NAND2_X1 U14608 ( .A1(n14732), .A2(n12999), .ZN(n12977) );
  NAND2_X1 U14609 ( .A1(n12978), .A2(n12977), .ZN(n12979) );
  XNOR2_X1 U14610 ( .A(n12979), .B(n13009), .ZN(n12982) );
  NOR2_X1 U14611 ( .A1(n14972), .A2(n13023), .ZN(n12980) );
  AOI21_X1 U14612 ( .B1(n14959), .B2(n13019), .A(n12980), .ZN(n12981) );
  OR2_X1 U14613 ( .A1(n12982), .A2(n12981), .ZN(n14695) );
  NAND2_X1 U14614 ( .A1(n14697), .A2(n14695), .ZN(n12983) );
  NAND2_X1 U14615 ( .A1(n12982), .A2(n12981), .ZN(n14694) );
  AOI22_X1 U14616 ( .A1(n15141), .A2(n13014), .B1(n12999), .B2(n14958), .ZN(
        n12984) );
  XOR2_X1 U14617 ( .A(n13025), .B(n12984), .Z(n12986) );
  INV_X1 U14618 ( .A(n14958), .ZN(n14927) );
  OAI22_X1 U14619 ( .A1(n14949), .A2(n13024), .B1(n14927), .B2(n13023), .ZN(
        n12985) );
  NOR2_X1 U14620 ( .A1(n12986), .A2(n12985), .ZN(n14666) );
  AOI21_X1 U14621 ( .B1(n12986), .B2(n12985), .A(n14666), .ZN(n14614) );
  INV_X1 U14622 ( .A(n14666), .ZN(n12987) );
  NAND2_X1 U14623 ( .A1(n15135), .A2(n13014), .ZN(n12989) );
  NAND2_X1 U14624 ( .A1(n14731), .A2(n12999), .ZN(n12988) );
  NAND2_X1 U14625 ( .A1(n12989), .A2(n12988), .ZN(n12990) );
  XNOR2_X1 U14626 ( .A(n12990), .B(n13009), .ZN(n12992) );
  AND2_X1 U14627 ( .A1(n14731), .A2(n13018), .ZN(n12991) );
  AOI21_X1 U14628 ( .B1(n15135), .B2(n13019), .A(n12991), .ZN(n12993) );
  NAND2_X1 U14629 ( .A1(n12992), .A2(n12993), .ZN(n12998) );
  INV_X1 U14630 ( .A(n12992), .ZN(n12995) );
  INV_X1 U14631 ( .A(n12993), .ZN(n12994) );
  NAND2_X1 U14632 ( .A1(n12995), .A2(n12994), .ZN(n12996) );
  NAND2_X1 U14633 ( .A1(n14919), .A2(n13014), .ZN(n13001) );
  NAND2_X1 U14634 ( .A1(n14730), .A2(n12999), .ZN(n13000) );
  NAND2_X1 U14635 ( .A1(n13001), .A2(n13000), .ZN(n13002) );
  XNOR2_X1 U14636 ( .A(n13002), .B(n13025), .ZN(n13003) );
  AOI22_X1 U14637 ( .A1(n14919), .A2(n13019), .B1(n13018), .B2(n14730), .ZN(
        n13004) );
  XNOR2_X1 U14638 ( .A(n13003), .B(n13004), .ZN(n14656) );
  INV_X1 U14639 ( .A(n13003), .ZN(n13005) );
  NAND2_X1 U14640 ( .A1(n13005), .A2(n13004), .ZN(n13006) );
  NAND2_X1 U14641 ( .A1(n15121), .A2(n13014), .ZN(n13008) );
  OR2_X1 U14642 ( .A1(n14888), .A2(n13024), .ZN(n13007) );
  NAND2_X1 U14643 ( .A1(n13008), .A2(n13007), .ZN(n13010) );
  XNOR2_X1 U14644 ( .A(n13010), .B(n13009), .ZN(n13013) );
  NOR2_X1 U14645 ( .A1(n14888), .A2(n13023), .ZN(n13011) );
  AOI21_X1 U14646 ( .B1(n15121), .B2(n13019), .A(n13011), .ZN(n13012) );
  OR2_X1 U14647 ( .A1(n13013), .A2(n13012), .ZN(n14714) );
  NAND2_X1 U14648 ( .A1(n14713), .A2(n14714), .ZN(n14712) );
  NAND2_X1 U14649 ( .A1(n13013), .A2(n13012), .ZN(n14715) );
  NAND2_X1 U14650 ( .A1(n15114), .A2(n13014), .ZN(n13016) );
  OR2_X1 U14651 ( .A1(n14904), .A2(n13024), .ZN(n13015) );
  NAND2_X1 U14652 ( .A1(n13016), .A2(n13015), .ZN(n13017) );
  XNOR2_X1 U14653 ( .A(n13017), .B(n13025), .ZN(n13020) );
  AOI22_X1 U14654 ( .A1(n15114), .A2(n13019), .B1(n13018), .B2(n14728), .ZN(
        n13021) );
  XNOR2_X1 U14655 ( .A(n13020), .B(n13021), .ZN(n14595) );
  INV_X1 U14656 ( .A(n13020), .ZN(n13022) );
  OAI22_X1 U14657 ( .A1(n14868), .A2(n7171), .B1(n14887), .B2(n13024), .ZN(
        n13028) );
  OAI22_X1 U14658 ( .A1(n14868), .A2(n13024), .B1(n14887), .B2(n13023), .ZN(
        n13026) );
  XNOR2_X1 U14659 ( .A(n13026), .B(n13025), .ZN(n13027) );
  XOR2_X1 U14660 ( .A(n13028), .B(n13027), .Z(n13029) );
  OAI22_X1 U14661 ( .A1(n13030), .A2(n15042), .B1(n14904), .B2(n15041), .ZN(
        n14865) );
  AOI22_X1 U14662 ( .A1(n16011), .A2(n14865), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13031) );
  OAI21_X1 U14663 ( .B1(n14873), .B2(n16031), .A(n13031), .ZN(n13032) );
  AOI21_X1 U14664 ( .B1(n15105), .B2(n16027), .A(n13032), .ZN(n13033) );
  INV_X1 U14665 ( .A(n13034), .ZN(n13035) );
  OAI222_X1 U14666 ( .A1(n13036), .A2(P3_U3151), .B1(n13787), .B2(n13882), 
        .C1(n13993), .C2(n13035), .ZN(P3_U3265) );
  XNOR2_X1 U14667 ( .A(n13463), .B(n13103), .ZN(n13099) );
  XNOR2_X1 U14668 ( .A(n13099), .B(n13473), .ZN(n13101) );
  INV_X1 U14669 ( .A(n13037), .ZN(n13038) );
  NAND2_X1 U14670 ( .A1(n13038), .A2(n13211), .ZN(n13039) );
  NAND2_X1 U14671 ( .A1(n13040), .A2(n13039), .ZN(n13078) );
  XNOR2_X1 U14672 ( .A(n13702), .B(n13041), .ZN(n13042) );
  XNOR2_X1 U14673 ( .A(n13042), .B(n13210), .ZN(n13077) );
  NAND2_X1 U14674 ( .A1(n13078), .A2(n13077), .ZN(n13045) );
  INV_X1 U14675 ( .A(n13042), .ZN(n13043) );
  NAND2_X1 U14676 ( .A1(n13043), .A2(n13210), .ZN(n13044) );
  XNOR2_X1 U14677 ( .A(n13698), .B(n13103), .ZN(n13186) );
  INV_X1 U14678 ( .A(n13186), .ZN(n13046) );
  XNOR2_X1 U14679 ( .A(n13768), .B(n13103), .ZN(n13047) );
  XNOR2_X1 U14680 ( .A(n13047), .B(n13139), .ZN(n13129) );
  NAND2_X1 U14681 ( .A1(n13047), .A2(n13608), .ZN(n13048) );
  NAND2_X1 U14682 ( .A1(n13128), .A2(n13048), .ZN(n13137) );
  XNOR2_X1 U14683 ( .A(n13618), .B(n13103), .ZN(n13049) );
  XNOR2_X1 U14684 ( .A(n13049), .B(n13628), .ZN(n13136) );
  NAND2_X1 U14685 ( .A1(n13137), .A2(n13136), .ZN(n13135) );
  NAND2_X1 U14686 ( .A1(n13049), .A2(n13588), .ZN(n13050) );
  NAND2_X1 U14687 ( .A1(n13135), .A2(n13050), .ZN(n13171) );
  XNOR2_X1 U14688 ( .A(n13599), .B(n13103), .ZN(n13051) );
  XNOR2_X1 U14689 ( .A(n13051), .B(n13574), .ZN(n13170) );
  NAND2_X1 U14690 ( .A1(n13171), .A2(n13170), .ZN(n13169) );
  NAND2_X1 U14691 ( .A1(n13051), .A2(n13607), .ZN(n13052) );
  NAND2_X1 U14692 ( .A1(n13169), .A2(n13052), .ZN(n13094) );
  XNOR2_X1 U14693 ( .A(n13582), .B(n13103), .ZN(n13053) );
  XNOR2_X1 U14694 ( .A(n13053), .B(n13590), .ZN(n13093) );
  NAND2_X1 U14695 ( .A1(n13094), .A2(n13093), .ZN(n13092) );
  NAND2_X1 U14696 ( .A1(n13053), .A2(n13208), .ZN(n13054) );
  NAND2_X1 U14697 ( .A1(n13092), .A2(n13054), .ZN(n13156) );
  XNOR2_X1 U14698 ( .A(n13746), .B(n13103), .ZN(n13055) );
  XNOR2_X1 U14699 ( .A(n13055), .B(n13207), .ZN(n13155) );
  NAND2_X1 U14700 ( .A1(n13156), .A2(n13155), .ZN(n13154) );
  INV_X1 U14701 ( .A(n13055), .ZN(n13056) );
  NAND2_X1 U14702 ( .A1(n13056), .A2(n13207), .ZN(n13057) );
  NAND2_X1 U14703 ( .A1(n13154), .A2(n13057), .ZN(n13115) );
  XNOR2_X1 U14704 ( .A(n13120), .B(n13103), .ZN(n13058) );
  XNOR2_X1 U14705 ( .A(n13058), .B(n13560), .ZN(n13114) );
  NAND2_X1 U14706 ( .A1(n13115), .A2(n13114), .ZN(n13113) );
  NAND2_X1 U14707 ( .A1(n13058), .A2(n13206), .ZN(n13059) );
  XNOR2_X1 U14708 ( .A(n13734), .B(n13103), .ZN(n13060) );
  INV_X1 U14709 ( .A(n13060), .ZN(n13061) );
  NOR2_X1 U14710 ( .A1(n13062), .A2(n13061), .ZN(n13063) );
  XNOR2_X1 U14711 ( .A(n13654), .B(n13103), .ZN(n13146) );
  XNOR2_X1 U14712 ( .A(n13657), .B(n13103), .ZN(n13065) );
  OAI22_X1 U14713 ( .A1(n13146), .A2(n13515), .B1(n13528), .B2(n13065), .ZN(
        n13066) );
  INV_X1 U14714 ( .A(n13065), .ZN(n13143) );
  OAI21_X1 U14715 ( .B1(n13143), .B2(n13204), .A(n13487), .ZN(n13064) );
  XNOR2_X1 U14716 ( .A(n13493), .B(n13103), .ZN(n13067) );
  XNOR2_X1 U14717 ( .A(n13067), .B(n13472), .ZN(n13122) );
  XNOR2_X1 U14718 ( .A(n13647), .B(n13103), .ZN(n13069) );
  XNOR2_X1 U14719 ( .A(n13069), .B(n13068), .ZN(n13180) );
  INV_X1 U14720 ( .A(n13069), .ZN(n13070) );
  XOR2_X1 U14721 ( .A(n13101), .B(n13102), .Z(n13076) );
  AOI22_X1 U14722 ( .A1(n13172), .A2(n13486), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13071) );
  OAI21_X1 U14723 ( .B1(n13072), .B2(n13174), .A(n13071), .ZN(n13074) );
  INV_X1 U14724 ( .A(n13463), .ZN(n13710) );
  NOR2_X1 U14725 ( .A1(n13710), .A2(n13178), .ZN(n13073) );
  AOI211_X1 U14726 ( .C1(n13462), .C2(n13190), .A(n13074), .B(n13073), .ZN(
        n13075) );
  OAI21_X1 U14727 ( .B1(n13076), .B2(n13200), .A(n13075), .ZN(P3_U3154) );
  XNOR2_X1 U14728 ( .A(n13078), .B(n13077), .ZN(n13086) );
  NAND2_X1 U14729 ( .A1(n13190), .A2(n13079), .ZN(n13081) );
  INV_X1 U14730 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13936) );
  NOR2_X1 U14731 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13936), .ZN(n13302) );
  AOI21_X1 U14732 ( .B1(n13191), .B2(n13209), .A(n13302), .ZN(n13080) );
  OAI211_X1 U14733 ( .C1(n13195), .C2(n13082), .A(n13081), .B(n13080), .ZN(
        n13083) );
  AOI21_X1 U14734 ( .B1(n13084), .B2(n13197), .A(n13083), .ZN(n13085) );
  OAI21_X1 U14735 ( .B1(n13086), .B2(n13200), .A(n13085), .ZN(P3_U3155) );
  XNOR2_X1 U14736 ( .A(n13144), .B(n13143), .ZN(n13145) );
  XNOR2_X1 U14737 ( .A(n13145), .B(n13528), .ZN(n13091) );
  AOI22_X1 U14738 ( .A1(n13191), .A2(n13487), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13088) );
  NAND2_X1 U14739 ( .A1(n13190), .A2(n13519), .ZN(n13087) );
  OAI211_X1 U14740 ( .C1(n13541), .C2(n13195), .A(n13088), .B(n13087), .ZN(
        n13089) );
  AOI21_X1 U14741 ( .B1(n13657), .B2(n13197), .A(n13089), .ZN(n13090) );
  OAI21_X1 U14742 ( .B1(n13091), .B2(n13200), .A(n13090), .ZN(P3_U3156) );
  OAI211_X1 U14743 ( .C1(n13094), .C2(n13093), .A(n13092), .B(n13168), .ZN(
        n13098) );
  NAND2_X1 U14744 ( .A1(n13172), .A2(n13607), .ZN(n13095) );
  NAND2_X1 U14745 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13413)
         );
  OAI211_X1 U14746 ( .C1(n13575), .C2(n13174), .A(n13095), .B(n13413), .ZN(
        n13096) );
  AOI21_X1 U14747 ( .B1(n13580), .B2(n13190), .A(n13096), .ZN(n13097) );
  OAI211_X1 U14748 ( .C1(n13178), .C2(n13582), .A(n13098), .B(n13097), .ZN(
        P3_U3159) );
  AOI22_X1 U14749 ( .A1(n13102), .A2(n13101), .B1(n13100), .B2(n13099), .ZN(
        n13106) );
  XNOR2_X1 U14750 ( .A(n13104), .B(n13103), .ZN(n13105) );
  XNOR2_X1 U14751 ( .A(n13106), .B(n13105), .ZN(n13112) );
  AOI22_X1 U14752 ( .A1(n13172), .A2(n13473), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13107) );
  OAI21_X1 U14753 ( .B1(n13108), .B2(n13174), .A(n13107), .ZN(n13110) );
  NOR2_X1 U14754 ( .A1(n13446), .A2(n13178), .ZN(n13109) );
  AOI211_X1 U14755 ( .C1(n13444), .C2(n13190), .A(n13110), .B(n13109), .ZN(
        n13111) );
  OAI21_X1 U14756 ( .B1(n13112), .B2(n13200), .A(n13111), .ZN(P3_U3160) );
  OAI211_X1 U14757 ( .C1(n13115), .C2(n13114), .A(n13113), .B(n13168), .ZN(
        n13119) );
  AOI22_X1 U14758 ( .A1(n13207), .A2(n13172), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13116) );
  OAI21_X1 U14759 ( .B1(n13541), .B2(n13174), .A(n13116), .ZN(n13117) );
  AOI21_X1 U14760 ( .B1(n13549), .B2(n13190), .A(n13117), .ZN(n13118) );
  OAI211_X1 U14761 ( .C1(n13120), .C2(n13178), .A(n13119), .B(n13118), .ZN(
        P3_U3163) );
  XOR2_X1 U14762 ( .A(n13122), .B(n13121), .Z(n13127) );
  AOI22_X1 U14763 ( .A1(n13191), .A2(n13486), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13124) );
  NAND2_X1 U14764 ( .A1(n13190), .A2(n13492), .ZN(n13123) );
  OAI211_X1 U14765 ( .C1(n13515), .C2(n13195), .A(n13124), .B(n13123), .ZN(
        n13125) );
  AOI21_X1 U14766 ( .B1(n13493), .B2(n13197), .A(n13125), .ZN(n13126) );
  OAI21_X1 U14767 ( .B1(n13127), .B2(n13200), .A(n13126), .ZN(P3_U3165) );
  OAI211_X1 U14768 ( .C1(n13130), .C2(n13129), .A(n13128), .B(n13168), .ZN(
        n13134) );
  NAND2_X1 U14769 ( .A1(n13172), .A2(n13209), .ZN(n13131) );
  NAND2_X1 U14770 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13342)
         );
  OAI211_X1 U14771 ( .C1(n13628), .C2(n13174), .A(n13131), .B(n13342), .ZN(
        n13132) );
  AOI21_X1 U14772 ( .B1(n13633), .B2(n13190), .A(n13132), .ZN(n13133) );
  OAI211_X1 U14773 ( .C1(n13768), .C2(n13178), .A(n13134), .B(n13133), .ZN(
        P3_U3166) );
  OAI211_X1 U14774 ( .C1(n13137), .C2(n13136), .A(n13135), .B(n13168), .ZN(
        n13142) );
  AND2_X1 U14775 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13373) );
  AOI21_X1 U14776 ( .B1(n13191), .B2(n13607), .A(n13373), .ZN(n13138) );
  OAI21_X1 U14777 ( .B1(n13195), .B2(n13139), .A(n13138), .ZN(n13140) );
  AOI21_X1 U14778 ( .B1(n13616), .B2(n13190), .A(n13140), .ZN(n13141) );
  OAI211_X1 U14779 ( .C1(n13618), .C2(n13178), .A(n13142), .B(n13141), .ZN(
        P3_U3168) );
  OAI22_X1 U14780 ( .A1(n13145), .A2(n13204), .B1(n13144), .B2(n13143), .ZN(
        n13148) );
  XNOR2_X1 U14781 ( .A(n13146), .B(n13515), .ZN(n13147) );
  XNOR2_X1 U14782 ( .A(n13148), .B(n13147), .ZN(n13153) );
  AOI22_X1 U14783 ( .A1(n13191), .A2(n13472), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13150) );
  NAND2_X1 U14784 ( .A1(n13190), .A2(n13506), .ZN(n13149) );
  OAI211_X1 U14785 ( .C1(n13528), .C2(n13195), .A(n13150), .B(n13149), .ZN(
        n13151) );
  AOI21_X1 U14786 ( .B1(n13654), .B2(n13197), .A(n13151), .ZN(n13152) );
  OAI21_X1 U14787 ( .B1(n13153), .B2(n13200), .A(n13152), .ZN(P3_U3169) );
  INV_X1 U14788 ( .A(n13746), .ZN(n13161) );
  OAI211_X1 U14789 ( .C1(n13156), .C2(n13155), .A(n13154), .B(n13168), .ZN(
        n13160) );
  NOR2_X1 U14790 ( .A1(n13195), .A2(n13590), .ZN(n13158) );
  OAI22_X1 U14791 ( .A1(n13560), .A2(n13174), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13971), .ZN(n13157) );
  AOI211_X1 U14792 ( .C1(n13567), .C2(n13190), .A(n13158), .B(n13157), .ZN(
        n13159) );
  OAI211_X1 U14793 ( .C1(n13161), .C2(n13178), .A(n13160), .B(n13159), .ZN(
        P3_U3173) );
  XNOR2_X1 U14794 ( .A(n13162), .B(n13205), .ZN(n13167) );
  AOI22_X1 U14795 ( .A1(n13206), .A2(n13172), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13164) );
  NAND2_X1 U14796 ( .A1(n13190), .A2(n13537), .ZN(n13163) );
  OAI211_X1 U14797 ( .C1(n13528), .C2(n13174), .A(n13164), .B(n13163), .ZN(
        n13165) );
  AOI21_X1 U14798 ( .B1(n13734), .B2(n13197), .A(n13165), .ZN(n13166) );
  OAI21_X1 U14799 ( .B1(n13167), .B2(n13200), .A(n13166), .ZN(P3_U3175) );
  OAI211_X1 U14800 ( .C1(n13171), .C2(n13170), .A(n13169), .B(n13168), .ZN(
        n13177) );
  NAND2_X1 U14801 ( .A1(n13172), .A2(n13588), .ZN(n13173) );
  NAND2_X1 U14802 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13384)
         );
  OAI211_X1 U14803 ( .C1(n13590), .C2(n13174), .A(n13173), .B(n13384), .ZN(
        n13175) );
  AOI21_X1 U14804 ( .B1(n13597), .B2(n13190), .A(n13175), .ZN(n13176) );
  OAI211_X1 U14805 ( .C1(n13599), .C2(n13178), .A(n13177), .B(n13176), .ZN(
        P3_U3178) );
  XOR2_X1 U14806 ( .A(n13180), .B(n13179), .Z(n13185) );
  AOI22_X1 U14807 ( .A1(n13191), .A2(n13473), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13182) );
  NAND2_X1 U14808 ( .A1(n13190), .A2(n13477), .ZN(n13181) );
  OAI211_X1 U14809 ( .C1(n13505), .C2(n13195), .A(n13182), .B(n13181), .ZN(
        n13183) );
  AOI21_X1 U14810 ( .B1(n13647), .B2(n13197), .A(n13183), .ZN(n13184) );
  OAI21_X1 U14811 ( .B1(n13185), .B2(n13200), .A(n13184), .ZN(P3_U3180) );
  XNOR2_X1 U14812 ( .A(n13186), .B(n13626), .ZN(n13187) );
  XNOR2_X1 U14813 ( .A(n13188), .B(n13187), .ZN(n13201) );
  NAND2_X1 U14814 ( .A1(n13190), .A2(n13189), .ZN(n13193) );
  AND2_X1 U14815 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13317) );
  AOI21_X1 U14816 ( .B1(n13191), .B2(n13608), .A(n13317), .ZN(n13192) );
  OAI211_X1 U14817 ( .C1(n13195), .C2(n13194), .A(n13193), .B(n13192), .ZN(
        n13196) );
  AOI21_X1 U14818 ( .B1(n13198), .B2(n13197), .A(n13196), .ZN(n13199) );
  OAI21_X1 U14819 ( .B1(n13201), .B2(n13200), .A(n13199), .ZN(P3_U3181) );
  MUX2_X1 U14820 ( .A(n13429), .B(P3_DATAO_REG_31__SCAN_IN), .S(n13223), .Z(
        P3_U3522) );
  MUX2_X1 U14821 ( .A(n13202), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13223), .Z(
        P3_U3521) );
  MUX2_X1 U14822 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n13203), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14823 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13459), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14824 ( .A(n13473), .B(P3_DATAO_REG_27__SCAN_IN), .S(n13223), .Z(
        P3_U3518) );
  MUX2_X1 U14825 ( .A(n13486), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13223), .Z(
        P3_U3517) );
  MUX2_X1 U14826 ( .A(n13472), .B(P3_DATAO_REG_25__SCAN_IN), .S(n13223), .Z(
        P3_U3516) );
  MUX2_X1 U14827 ( .A(n13487), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13223), .Z(
        P3_U3515) );
  MUX2_X1 U14828 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13204), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14829 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13205), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14830 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13206), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14831 ( .A(n13207), .B(P3_DATAO_REG_20__SCAN_IN), .S(n13223), .Z(
        P3_U3511) );
  MUX2_X1 U14832 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13208), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14833 ( .A(n13607), .B(P3_DATAO_REG_18__SCAN_IN), .S(n13223), .Z(
        P3_U3509) );
  MUX2_X1 U14834 ( .A(n13588), .B(P3_DATAO_REG_17__SCAN_IN), .S(n13223), .Z(
        P3_U3508) );
  MUX2_X1 U14835 ( .A(n13608), .B(P3_DATAO_REG_16__SCAN_IN), .S(n13223), .Z(
        P3_U3507) );
  MUX2_X1 U14836 ( .A(n13209), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13223), .Z(
        P3_U3506) );
  MUX2_X1 U14837 ( .A(n13210), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13223), .Z(
        P3_U3505) );
  MUX2_X1 U14838 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13211), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14839 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13212), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14840 ( .A(n13213), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13223), .Z(
        P3_U3502) );
  MUX2_X1 U14841 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13214), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14842 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13215), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14843 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13216), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14844 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13217), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14845 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13218), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14846 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13219), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14847 ( .A(n13220), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13223), .Z(
        P3_U3495) );
  MUX2_X1 U14848 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13221), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14849 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13222), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14850 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n11371), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14851 ( .A(n13224), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13223), .Z(
        P3_U3491) );
  OAI21_X1 U14852 ( .B1(n13227), .B2(n13226), .A(n13225), .ZN(n13228) );
  NAND2_X1 U14853 ( .A1(n13228), .A2(n15638), .ZN(n13248) );
  OR3_X1 U14854 ( .A1(n13231), .A2(n13230), .A3(n13229), .ZN(n13232) );
  AOI21_X1 U14855 ( .B1(n13233), .B2(n13232), .A(n15631), .ZN(n13234) );
  AOI211_X1 U14856 ( .C1(n15246), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n13235), .B(
        n13234), .ZN(n13247) );
  NAND2_X1 U14857 ( .A1(n15618), .A2(n13236), .ZN(n13246) );
  INV_X1 U14858 ( .A(n13237), .ZN(n13241) );
  INV_X1 U14859 ( .A(n13238), .ZN(n13239) );
  NOR3_X1 U14860 ( .A1(n13241), .A2(n13240), .A3(n13239), .ZN(n13243) );
  OAI21_X1 U14861 ( .B1(n13244), .B2(n13243), .A(n13242), .ZN(n13245) );
  NAND4_X1 U14862 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        P3_U3188) );
  NOR2_X1 U14863 ( .A1(n13251), .A2(n13250), .ZN(n13281) );
  AOI21_X1 U14864 ( .B1(n13251), .B2(n13250), .A(n13281), .ZN(n13271) );
  NAND2_X1 U14865 ( .A1(n13252), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13260) );
  INV_X1 U14866 ( .A(n13260), .ZN(n13255) );
  INV_X1 U14867 ( .A(n13253), .ZN(n13254) );
  MUX2_X1 U14868 ( .A(n13255), .B(n13254), .S(n7165), .Z(n13256) );
  MUX2_X1 U14869 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n7206), .Z(n13295) );
  INV_X1 U14870 ( .A(n13294), .ZN(n13280) );
  XNOR2_X1 U14871 ( .A(n13295), .B(n13280), .ZN(n13258) );
  NAND2_X1 U14872 ( .A1(n13259), .A2(n13258), .ZN(n13296) );
  OAI21_X1 U14873 ( .B1(n13259), .B2(n13258), .A(n13296), .ZN(n13269) );
  INV_X1 U14874 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13262) );
  AOI21_X1 U14875 ( .B1(n13263), .B2(n13262), .A(n13273), .ZN(n13264) );
  NOR2_X1 U14876 ( .A1(n15636), .A2(n13264), .ZN(n13265) );
  AOI211_X1 U14877 ( .C1(n15246), .C2(P3_ADDR_REG_13__SCAN_IN), .A(n13266), 
        .B(n13265), .ZN(n13267) );
  OAI21_X1 U14878 ( .B1(n13294), .B2(n15641), .A(n13267), .ZN(n13268) );
  AOI21_X1 U14879 ( .B1(n15638), .B2(n13269), .A(n13268), .ZN(n13270) );
  OAI21_X1 U14880 ( .B1(n13271), .B2(n15631), .A(n13270), .ZN(P3_U3195) );
  NOR2_X1 U14881 ( .A1(n13280), .A2(n13272), .ZN(n13274) );
  NAND2_X1 U14882 ( .A1(n13305), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13313) );
  OR2_X1 U14883 ( .A1(n13305), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13275) );
  NAND2_X1 U14884 ( .A1(n13313), .A2(n13275), .ZN(n13277) );
  OR2_X2 U14885 ( .A1(n13278), .A2(n13277), .ZN(n13314) );
  INV_X1 U14886 ( .A(n13314), .ZN(n13276) );
  AOI21_X1 U14887 ( .B1(n13278), .B2(n13277), .A(n13276), .ZN(n13309) );
  NOR2_X1 U14888 ( .A1(n13280), .A2(n13279), .ZN(n13282) );
  NOR2_X1 U14889 ( .A1(n13282), .A2(n13281), .ZN(n13285) );
  INV_X1 U14890 ( .A(n13285), .ZN(n13287) );
  NAND2_X1 U14891 ( .A1(n13305), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13310) );
  OR2_X1 U14892 ( .A1(n13305), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13283) );
  NAND2_X1 U14893 ( .A1(n13310), .A2(n13283), .ZN(n13284) );
  INV_X1 U14894 ( .A(n13284), .ZN(n13286) );
  OR2_X2 U14895 ( .A1(n13285), .A2(n13284), .ZN(n13311) );
  OAI21_X1 U14896 ( .B1(n13287), .B2(n13286), .A(n13311), .ZN(n13307) );
  INV_X1 U14897 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13289) );
  INV_X1 U14898 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13288) );
  MUX2_X1 U14899 ( .A(n13289), .B(n13288), .S(n7206), .Z(n13291) );
  INV_X1 U14900 ( .A(n13291), .ZN(n13293) );
  INV_X1 U14901 ( .A(n13305), .ZN(n13290) );
  NOR2_X1 U14902 ( .A1(n13291), .A2(n13290), .ZN(n13319) );
  INV_X1 U14903 ( .A(n13319), .ZN(n13292) );
  OAI21_X1 U14904 ( .B1(n13293), .B2(n13305), .A(n13292), .ZN(n13299) );
  OR2_X1 U14905 ( .A1(n13295), .A2(n13294), .ZN(n13297) );
  NAND2_X1 U14906 ( .A1(n13299), .A2(n13298), .ZN(n13301) );
  INV_X1 U14907 ( .A(n13318), .ZN(n13300) );
  NAND3_X1 U14908 ( .A1(n13301), .A2(n15638), .A3(n13300), .ZN(n13304) );
  AOI21_X1 U14909 ( .B1(n15246), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13302), 
        .ZN(n13303) );
  OAI211_X1 U14910 ( .C1(n15641), .C2(n13305), .A(n13304), .B(n13303), .ZN(
        n13306) );
  AOI21_X1 U14911 ( .B1(n13307), .B2(n13422), .A(n13306), .ZN(n13308) );
  OAI21_X1 U14912 ( .B1(n13309), .B2(n15636), .A(n13308), .ZN(P3_U3196) );
  INV_X1 U14913 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13321) );
  INV_X1 U14914 ( .A(n13346), .ZN(n13320) );
  AOI21_X1 U14915 ( .B1(n13321), .B2(n13312), .A(n13331), .ZN(n13330) );
  INV_X1 U14916 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13315) );
  AOI21_X1 U14917 ( .B1(n13316), .B2(n13315), .A(n13347), .ZN(n13327) );
  AOI21_X1 U14918 ( .B1(n15246), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13317), 
        .ZN(n13326) );
  MUX2_X1 U14919 ( .A(n13315), .B(n13321), .S(n7166), .Z(n13322) );
  NAND2_X1 U14920 ( .A1(n13322), .A2(n13323), .ZN(n13337) );
  OAI21_X1 U14921 ( .B1(n13323), .B2(n13322), .A(n13337), .ZN(n13324) );
  NAND2_X1 U14922 ( .A1(n13324), .A2(n15638), .ZN(n13325) );
  OAI211_X1 U14923 ( .C1(n15636), .C2(n13327), .A(n13326), .B(n13325), .ZN(
        n13328) );
  AOI21_X1 U14924 ( .B1(n13346), .B2(n15618), .A(n13328), .ZN(n13329) );
  OAI21_X1 U14925 ( .B1(n13330), .B2(n15631), .A(n13329), .ZN(P3_U3197) );
  NOR2_X1 U14926 ( .A1(n13346), .A2(n7267), .ZN(n13332) );
  NAND2_X1 U14927 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13365), .ZN(n13333) );
  OAI21_X1 U14928 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n13365), .A(n13333), 
        .ZN(n13334) );
  AOI21_X1 U14929 ( .B1(n13335), .B2(n13334), .A(n13361), .ZN(n13357) );
  NAND2_X1 U14930 ( .A1(n13346), .A2(n13336), .ZN(n13338) );
  NAND2_X1 U14931 ( .A1(n13338), .A2(n13337), .ZN(n13340) );
  MUX2_X1 U14932 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n7206), .Z(n13366) );
  XNOR2_X1 U14933 ( .A(n13366), .B(n13341), .ZN(n13339) );
  NAND2_X1 U14934 ( .A1(n13339), .A2(n13340), .ZN(n13367) );
  OAI21_X1 U14935 ( .B1(n13340), .B2(n13339), .A(n13367), .ZN(n13355) );
  INV_X1 U14936 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n13344) );
  NAND2_X1 U14937 ( .A1(n15618), .A2(n13341), .ZN(n13343) );
  OAI211_X1 U14938 ( .C1(n13344), .C2(n15651), .A(n13343), .B(n13342), .ZN(
        n13354) );
  NOR2_X1 U14939 ( .A1(n13346), .A2(n13345), .ZN(n13348) );
  NAND2_X1 U14940 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13365), .ZN(n13349) );
  OAI21_X1 U14941 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13365), .A(n13349), 
        .ZN(n13350) );
  AOI21_X1 U14942 ( .B1(n13351), .B2(n13350), .A(n13358), .ZN(n13352) );
  NOR2_X1 U14943 ( .A1(n13352), .A2(n15636), .ZN(n13353) );
  AOI211_X1 U14944 ( .C1(n15638), .C2(n13355), .A(n13354), .B(n13353), .ZN(
        n13356) );
  OAI21_X1 U14945 ( .B1(n13357), .B2(n15631), .A(n13356), .ZN(P3_U3198) );
  INV_X1 U14946 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13359) );
  AOI21_X1 U14947 ( .B1(n13360), .B2(n13359), .A(n13381), .ZN(n13379) );
  INV_X1 U14948 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13363) );
  AOI21_X1 U14949 ( .B1(n13363), .B2(n13362), .A(n13396), .ZN(n13364) );
  INV_X1 U14950 ( .A(n13364), .ZN(n13377) );
  MUX2_X1 U14951 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n7165), .Z(n13387) );
  XNOR2_X1 U14952 ( .A(n13387), .B(n13386), .ZN(n13369) );
  OR2_X1 U14953 ( .A1(n13366), .A2(n13365), .ZN(n13368) );
  NAND2_X1 U14954 ( .A1(n13368), .A2(n13367), .ZN(n13370) );
  NAND2_X1 U14955 ( .A1(n13369), .A2(n13370), .ZN(n13372) );
  INV_X1 U14956 ( .A(n13385), .ZN(n13371) );
  NAND3_X1 U14957 ( .A1(n13372), .A2(n15638), .A3(n13371), .ZN(n13375) );
  AOI21_X1 U14958 ( .B1(n15246), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13373), 
        .ZN(n13374) );
  OAI211_X1 U14959 ( .C1(n15641), .C2(n13386), .A(n13375), .B(n13374), .ZN(
        n13376) );
  AOI21_X1 U14960 ( .B1(n13377), .B2(n13422), .A(n13376), .ZN(n13378) );
  OAI21_X1 U14961 ( .B1(n13379), .B2(n15636), .A(n13378), .ZN(P3_U3199) );
  NAND2_X1 U14962 ( .A1(n13398), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13404) );
  OAI21_X1 U14963 ( .B1(n13398), .B2(P3_REG2_REG_18__SCAN_IN), .A(n13404), 
        .ZN(n13382) );
  AOI21_X1 U14964 ( .B1(n13383), .B2(n13382), .A(n13405), .ZN(n13403) );
  INV_X1 U14965 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15600) );
  OAI21_X1 U14966 ( .B1(n15651), .B2(n15600), .A(n13384), .ZN(n13393) );
  MUX2_X1 U14967 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n7206), .Z(n13389) );
  XNOR2_X1 U14968 ( .A(n13408), .B(n13407), .ZN(n13388) );
  NOR2_X1 U14969 ( .A1(n13391), .A2(n13390), .ZN(n13392) );
  NOR2_X1 U14970 ( .A1(n13395), .A2(n13394), .ZN(n13397) );
  NAND2_X1 U14971 ( .A1(n13398), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13417) );
  OAI21_X1 U14972 ( .B1(n13398), .B2(P3_REG1_REG_18__SCAN_IN), .A(n13417), 
        .ZN(n13399) );
  AND2_X1 U14973 ( .A1(n7301), .A2(n13399), .ZN(n13400) );
  OAI21_X1 U14974 ( .B1(n13419), .B2(n13400), .A(n13422), .ZN(n13401) );
  XNOR2_X1 U14975 ( .A(n13412), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13409) );
  AOI21_X1 U14976 ( .B1(n13408), .B2(n13407), .A(n13406), .ZN(n13411) );
  XNOR2_X1 U14977 ( .A(n13412), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13420) );
  MUX2_X1 U14978 ( .A(n13409), .B(n13420), .S(n7166), .Z(n13410) );
  XNOR2_X1 U14979 ( .A(n13411), .B(n13410), .ZN(n13416) );
  NOR2_X1 U14980 ( .A1(n15641), .A2(n13412), .ZN(n13415) );
  OAI21_X1 U14981 ( .B1(n15651), .B2(n8276), .A(n13413), .ZN(n13414) );
  INV_X1 U14982 ( .A(n13417), .ZN(n13418) );
  XNOR2_X1 U14983 ( .A(n13421), .B(n13420), .ZN(n13423) );
  NAND2_X1 U14984 ( .A1(n13423), .A2(n13422), .ZN(n13424) );
  OAI211_X1 U14985 ( .C1(n13426), .C2(n15636), .A(n13425), .B(n13424), .ZN(
        P3_U3201) );
  INV_X1 U14986 ( .A(n13427), .ZN(n13428) );
  NAND2_X1 U14987 ( .A1(n13429), .A2(n13428), .ZN(n13703) );
  INV_X1 U14988 ( .A(n13703), .ZN(n13431) );
  AND2_X1 U14989 ( .A1(n13634), .A2(n13430), .ZN(n13439) );
  NOR3_X1 U14990 ( .A1(n13431), .A2(n13635), .A3(n13439), .ZN(n13434) );
  NOR2_X1 U14991 ( .A1(n13565), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13432) );
  OAI22_X1 U14992 ( .A1(n13705), .A2(n13637), .B1(n13434), .B2(n13432), .ZN(
        P3_U3202) );
  NOR2_X1 U14993 ( .A1(n13565), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13433) );
  OAI22_X1 U14994 ( .A1(n13708), .A2(n13637), .B1(n13434), .B2(n13433), .ZN(
        P3_U3203) );
  INV_X1 U14995 ( .A(n13435), .ZN(n13442) );
  NAND2_X1 U14996 ( .A1(n13436), .A2(n13565), .ZN(n13441) );
  NOR2_X1 U14997 ( .A1(n13437), .A2(n13637), .ZN(n13438) );
  AOI211_X1 U14998 ( .C1(n13635), .C2(P3_REG2_REG_29__SCAN_IN), .A(n13439), 
        .B(n13438), .ZN(n13440) );
  OAI211_X1 U14999 ( .C1(n13512), .C2(n13442), .A(n13441), .B(n13440), .ZN(
        P3_U3204) );
  INV_X1 U15000 ( .A(n13443), .ZN(n13450) );
  AOI22_X1 U15001 ( .A1(n13635), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n13634), 
        .B2(n13444), .ZN(n13445) );
  OAI21_X1 U15002 ( .B1(n13446), .B2(n13637), .A(n13445), .ZN(n13447) );
  AOI21_X1 U15003 ( .B1(n13448), .B2(n13639), .A(n13447), .ZN(n13449) );
  OAI21_X1 U15004 ( .B1(n13450), .B2(n13635), .A(n13449), .ZN(P3_U3205) );
  OR2_X1 U15005 ( .A1(n13451), .A2(n13454), .ZN(n13452) );
  NAND2_X1 U15006 ( .A1(n13455), .A2(n13454), .ZN(n13456) );
  NAND2_X1 U15007 ( .A1(n13457), .A2(n13456), .ZN(n13458) );
  NAND2_X1 U15008 ( .A1(n13458), .A2(n13604), .ZN(n13461) );
  AOI22_X1 U15009 ( .A1(n13459), .A2(n13606), .B1(n13609), .B2(n13486), .ZN(
        n13460) );
  OAI211_X1 U15010 ( .C1(n15764), .C2(n13711), .A(n13461), .B(n13460), .ZN(
        n13709) );
  MUX2_X1 U15011 ( .A(n13709), .B(P3_REG2_REG_27__SCAN_IN), .S(n13635), .Z(
        n13466) );
  AOI22_X1 U15012 ( .A1(n13463), .A2(n13568), .B1(n13634), .B2(n13462), .ZN(
        n13464) );
  OAI21_X1 U15013 ( .B1(n13711), .B2(n13571), .A(n13464), .ZN(n13465) );
  XNOR2_X1 U15014 ( .A(n13469), .B(n13470), .ZN(n13471) );
  NAND2_X1 U15015 ( .A1(n13471), .A2(n13604), .ZN(n13475) );
  AOI22_X1 U15016 ( .A1(n13606), .A2(n13473), .B1(n13472), .B2(n13609), .ZN(
        n13474) );
  OAI211_X1 U15017 ( .C1(n15764), .C2(n13716), .A(n13475), .B(n13474), .ZN(
        n13714) );
  MUX2_X1 U15018 ( .A(n13714), .B(P3_REG2_REG_26__SCAN_IN), .S(n13635), .Z(
        n13476) );
  INV_X1 U15019 ( .A(n13476), .ZN(n13479) );
  AOI22_X1 U15020 ( .A1(n13647), .A2(n13568), .B1(n13634), .B2(n13477), .ZN(
        n13478) );
  OAI211_X1 U15021 ( .C1(n13716), .C2(n13571), .A(n13479), .B(n13478), .ZN(
        P3_U3207) );
  XNOR2_X1 U15022 ( .A(n13480), .B(n13482), .ZN(n13485) );
  INV_X1 U15023 ( .A(n13485), .ZN(n13721) );
  NAND2_X1 U15024 ( .A1(n13481), .A2(n13482), .ZN(n13483) );
  NAND3_X1 U15025 ( .A1(n13484), .A2(n13604), .A3(n13483), .ZN(n13490) );
  NAND2_X1 U15026 ( .A1(n13485), .A2(n13556), .ZN(n13489) );
  AOI22_X1 U15027 ( .A1(n13609), .A2(n13487), .B1(n13486), .B2(n13606), .ZN(
        n13488) );
  NAND3_X1 U15028 ( .A1(n13490), .A2(n13489), .A3(n13488), .ZN(n13719) );
  MUX2_X1 U15029 ( .A(n13719), .B(P3_REG2_REG_25__SCAN_IN), .S(n13635), .Z(
        n13491) );
  INV_X1 U15030 ( .A(n13491), .ZN(n13495) );
  AOI22_X1 U15031 ( .A1(n13493), .A2(n13568), .B1(n13634), .B2(n13492), .ZN(
        n13494) );
  OAI211_X1 U15032 ( .C1(n13721), .C2(n13571), .A(n13495), .B(n13494), .ZN(
        P3_U3208) );
  INV_X1 U15033 ( .A(n13496), .ZN(n13501) );
  AOI21_X1 U15034 ( .B1(n13659), .B2(n13499), .A(n13498), .ZN(n13500) );
  XNOR2_X1 U15035 ( .A(n13502), .B(n13503), .ZN(n13504) );
  OAI222_X1 U15036 ( .A1(n13629), .A2(n13505), .B1(n13627), .B2(n13528), .C1(
        n13504), .C2(n13625), .ZN(n13652) );
  NAND2_X1 U15037 ( .A1(n13652), .A2(n13565), .ZN(n13511) );
  INV_X1 U15038 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13508) );
  INV_X1 U15039 ( .A(n13506), .ZN(n13507) );
  OAI22_X1 U15040 ( .A1(n13565), .A2(n13508), .B1(n13507), .B2(n13520), .ZN(
        n13509) );
  AOI21_X1 U15041 ( .B1(n13654), .B2(n13568), .A(n13509), .ZN(n13510) );
  OAI211_X1 U15042 ( .C1(n13512), .C2(n13727), .A(n13511), .B(n13510), .ZN(
        P3_U3209) );
  AOI21_X1 U15043 ( .B1(n13514), .B2(n8783), .A(n13625), .ZN(n13518) );
  OAI22_X1 U15044 ( .A1(n13541), .A2(n13627), .B1(n13515), .B2(n13629), .ZN(
        n13516) );
  AOI21_X1 U15045 ( .B1(n13518), .B2(n13517), .A(n13516), .ZN(n13661) );
  INV_X1 U15046 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13522) );
  INV_X1 U15047 ( .A(n13519), .ZN(n13521) );
  OAI22_X1 U15048 ( .A1(n13565), .A2(n13522), .B1(n13521), .B2(n13520), .ZN(
        n13523) );
  AOI21_X1 U15049 ( .B1(n13657), .B2(n13568), .A(n13523), .ZN(n13526) );
  NAND2_X1 U15050 ( .A1(n13524), .A2(n7747), .ZN(n13658) );
  NAND3_X1 U15051 ( .A1(n13659), .A2(n13639), .A3(n13658), .ZN(n13525) );
  OAI211_X1 U15052 ( .C1(n13661), .C2(n13635), .A(n13526), .B(n13525), .ZN(
        P3_U3210) );
  XNOR2_X1 U15053 ( .A(n13527), .B(n7745), .ZN(n13535) );
  INV_X1 U15054 ( .A(n13535), .ZN(n13737) );
  INV_X1 U15055 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13536) );
  OAI22_X1 U15056 ( .A1(n13560), .A2(n13627), .B1(n13528), .B2(n13629), .ZN(
        n13534) );
  NAND3_X1 U15057 ( .A1(n13529), .A2(n7745), .A3(n13530), .ZN(n13531) );
  AOI21_X1 U15058 ( .B1(n13532), .B2(n13531), .A(n13625), .ZN(n13533) );
  AOI211_X1 U15059 ( .C1(n13535), .C2(n13556), .A(n13534), .B(n13533), .ZN(
        n13732) );
  MUX2_X1 U15060 ( .A(n13536), .B(n13732), .S(n13565), .Z(n13539) );
  AOI22_X1 U15061 ( .A1(n13734), .A2(n13568), .B1(n13634), .B2(n13537), .ZN(
        n13538) );
  OAI211_X1 U15062 ( .C1(n13737), .C2(n13571), .A(n13539), .B(n13538), .ZN(
        P3_U3211) );
  XNOR2_X1 U15063 ( .A(n13540), .B(n13542), .ZN(n13547) );
  INV_X1 U15064 ( .A(n13547), .ZN(n13743) );
  INV_X1 U15065 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13548) );
  OAI22_X1 U15066 ( .A1(n13541), .A2(n13629), .B1(n13575), .B2(n13627), .ZN(
        n13546) );
  NAND2_X1 U15067 ( .A1(n13543), .A2(n13542), .ZN(n13544) );
  AOI21_X1 U15068 ( .B1(n13529), .B2(n13544), .A(n13625), .ZN(n13545) );
  AOI211_X1 U15069 ( .C1(n13556), .C2(n13547), .A(n13546), .B(n13545), .ZN(
        n13738) );
  MUX2_X1 U15070 ( .A(n13548), .B(n13738), .S(n13565), .Z(n13551) );
  AOI22_X1 U15071 ( .A1(n13740), .A2(n13568), .B1(n13634), .B2(n13549), .ZN(
        n13550) );
  OAI211_X1 U15072 ( .C1(n13743), .C2(n13571), .A(n13551), .B(n13550), .ZN(
        P3_U3212) );
  NAND2_X1 U15073 ( .A1(n13553), .A2(n13552), .ZN(n13554) );
  NAND2_X1 U15074 ( .A1(n13555), .A2(n13554), .ZN(n13557) );
  INV_X1 U15075 ( .A(n13557), .ZN(n13750) );
  INV_X1 U15076 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13566) );
  NAND2_X1 U15077 ( .A1(n13557), .A2(n13556), .ZN(n13564) );
  XNOR2_X1 U15078 ( .A(n13558), .B(n8779), .ZN(n13559) );
  NAND2_X1 U15079 ( .A1(n13559), .A2(n13604), .ZN(n13563) );
  OAI22_X1 U15080 ( .A1(n13560), .A2(n13629), .B1(n13590), .B2(n13627), .ZN(
        n13561) );
  INV_X1 U15081 ( .A(n13561), .ZN(n13562) );
  MUX2_X1 U15082 ( .A(n13566), .B(n13744), .S(n13565), .Z(n13570) );
  AOI22_X1 U15083 ( .A1(n13746), .A2(n13568), .B1(n13634), .B2(n13567), .ZN(
        n13569) );
  OAI211_X1 U15084 ( .C1(n13750), .C2(n13571), .A(n13570), .B(n13569), .ZN(
        P3_U3213) );
  INV_X1 U15085 ( .A(n13578), .ZN(n13572) );
  XNOR2_X1 U15086 ( .A(n13573), .B(n13572), .ZN(n13577) );
  OAI22_X1 U15087 ( .A1(n13575), .A2(n13629), .B1(n13574), .B2(n13627), .ZN(
        n13576) );
  AOI21_X1 U15088 ( .B1(n13577), .B2(n13604), .A(n13576), .ZN(n13676) );
  XNOR2_X1 U15089 ( .A(n13579), .B(n13578), .ZN(n13674) );
  AOI22_X1 U15090 ( .A1(n13635), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n13634), 
        .B2(n13580), .ZN(n13581) );
  OAI21_X1 U15091 ( .B1(n13582), .B2(n13637), .A(n13581), .ZN(n13583) );
  AOI21_X1 U15092 ( .B1(n13674), .B2(n13639), .A(n13583), .ZN(n13584) );
  OAI21_X1 U15093 ( .B1(n13676), .B2(n13635), .A(n13584), .ZN(P3_U3214) );
  NAND2_X1 U15094 ( .A1(n13585), .A2(n13593), .ZN(n13586) );
  NAND2_X1 U15095 ( .A1(n13587), .A2(n13586), .ZN(n13592) );
  NAND2_X1 U15096 ( .A1(n13588), .A2(n13609), .ZN(n13589) );
  OAI21_X1 U15097 ( .B1(n13590), .B2(n13629), .A(n13589), .ZN(n13591) );
  AOI21_X1 U15098 ( .B1(n13592), .B2(n13604), .A(n13591), .ZN(n13681) );
  OR2_X1 U15099 ( .A1(n13594), .A2(n13593), .ZN(n13595) );
  NAND2_X1 U15100 ( .A1(n13596), .A2(n13595), .ZN(n13679) );
  AOI22_X1 U15101 ( .A1(n13635), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n13634), 
        .B2(n13597), .ZN(n13598) );
  OAI21_X1 U15102 ( .B1(n13599), .B2(n13637), .A(n13598), .ZN(n13600) );
  AOI21_X1 U15103 ( .B1(n13679), .B2(n13639), .A(n13600), .ZN(n13601) );
  OAI21_X1 U15104 ( .B1(n13681), .B2(n13635), .A(n13601), .ZN(P3_U3215) );
  NAND2_X1 U15105 ( .A1(n13602), .A2(n13612), .ZN(n13603) );
  NAND3_X1 U15106 ( .A1(n13605), .A2(n13604), .A3(n13603), .ZN(n13611) );
  AOI22_X1 U15107 ( .A1(n13609), .A2(n13608), .B1(n13607), .B2(n13606), .ZN(
        n13610) );
  OR2_X1 U15108 ( .A1(n13613), .A2(n13612), .ZN(n13614) );
  NAND2_X1 U15109 ( .A1(n13615), .A2(n13614), .ZN(n13684) );
  AOI22_X1 U15110 ( .A1(n13635), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n13634), 
        .B2(n13616), .ZN(n13617) );
  OAI21_X1 U15111 ( .B1(n13618), .B2(n13637), .A(n13617), .ZN(n13619) );
  AOI21_X1 U15112 ( .B1(n13684), .B2(n13639), .A(n13619), .ZN(n13620) );
  OAI21_X1 U15113 ( .B1(n13686), .B2(n13635), .A(n13620), .ZN(P3_U3216) );
  INV_X1 U15114 ( .A(n13621), .ZN(n13622) );
  AOI21_X1 U15115 ( .B1(n13631), .B2(n13623), .A(n13622), .ZN(n13624) );
  OAI222_X1 U15116 ( .A1(n13629), .A2(n13628), .B1(n13627), .B2(n13626), .C1(
        n13625), .C2(n13624), .ZN(n13690) );
  INV_X1 U15117 ( .A(n13690), .ZN(n13641) );
  OAI21_X1 U15118 ( .B1(n13632), .B2(n13631), .A(n13630), .ZN(n13691) );
  AOI22_X1 U15119 ( .A1(n13635), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n13634), 
        .B2(n13633), .ZN(n13636) );
  OAI21_X1 U15120 ( .B1(n13768), .B2(n13637), .A(n13636), .ZN(n13638) );
  AOI21_X1 U15121 ( .B1(n13691), .B2(n13639), .A(n13638), .ZN(n13640) );
  OAI21_X1 U15122 ( .B1(n13641), .B2(n13635), .A(n13640), .ZN(P3_U3217) );
  NOR2_X1 U15123 ( .A1(n15892), .A2(n13703), .ZN(n13643) );
  AOI21_X1 U15124 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15892), .A(n13643), 
        .ZN(n13642) );
  OAI21_X1 U15125 ( .B1(n13705), .B2(n13694), .A(n13642), .ZN(P3_U3490) );
  AOI21_X1 U15126 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15892), .A(n13643), 
        .ZN(n13644) );
  OAI21_X1 U15127 ( .B1(n13708), .B2(n13694), .A(n13644), .ZN(P3_U3489) );
  MUX2_X1 U15128 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13709), .S(n15894), .Z(
        n13646) );
  OAI22_X1 U15129 ( .A1(n13711), .A2(n13673), .B1(n13710), .B2(n13694), .ZN(
        n13645) );
  OR2_X1 U15130 ( .A1(n13646), .A2(n13645), .ZN(P3_U3486) );
  MUX2_X1 U15131 ( .A(n13714), .B(P3_REG1_REG_26__SCAN_IN), .S(n15892), .Z(
        n13649) );
  INV_X1 U15132 ( .A(n13647), .ZN(n13715) );
  OAI22_X1 U15133 ( .A1(n13716), .A2(n13673), .B1(n13715), .B2(n13694), .ZN(
        n13648) );
  OR2_X1 U15134 ( .A1(n13649), .A2(n13648), .ZN(P3_U3485) );
  MUX2_X1 U15135 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13719), .S(n15894), .Z(
        n13651) );
  OAI22_X1 U15136 ( .A1(n13721), .A2(n13673), .B1(n13720), .B2(n13694), .ZN(
        n13650) );
  OR2_X1 U15137 ( .A1(n13651), .A2(n13650), .ZN(P3_U3484) );
  INV_X1 U15138 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13655) );
  NOR2_X1 U15139 ( .A1(n13727), .A2(n15764), .ZN(n13653) );
  AOI211_X1 U15140 ( .C1(n15872), .C2(n13654), .A(n13653), .B(n13652), .ZN(
        n13724) );
  MUX2_X1 U15141 ( .A(n13655), .B(n13724), .S(n15894), .Z(n13656) );
  OAI21_X1 U15142 ( .B1(n13727), .B2(n13673), .A(n13656), .ZN(P3_U3483) );
  INV_X1 U15143 ( .A(n13657), .ZN(n13731) );
  NAND3_X1 U15144 ( .A1(n13659), .A2(n15891), .A3(n13658), .ZN(n13660) );
  AND2_X1 U15145 ( .A1(n13661), .A2(n13660), .ZN(n13729) );
  INV_X1 U15146 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13662) );
  MUX2_X1 U15147 ( .A(n13729), .B(n13662), .S(n15892), .Z(n13663) );
  OAI21_X1 U15148 ( .B1(n13731), .B2(n13694), .A(n13663), .ZN(P3_U3482) );
  INV_X1 U15149 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13664) );
  MUX2_X1 U15150 ( .A(n13664), .B(n13732), .S(n15894), .Z(n13666) );
  NAND2_X1 U15151 ( .A1(n13734), .A2(n13688), .ZN(n13665) );
  OAI211_X1 U15152 ( .C1(n13737), .C2(n13673), .A(n13666), .B(n13665), .ZN(
        P3_U3481) );
  INV_X1 U15153 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13667) );
  MUX2_X1 U15154 ( .A(n13667), .B(n13738), .S(n15894), .Z(n13669) );
  NAND2_X1 U15155 ( .A1(n13740), .A2(n13688), .ZN(n13668) );
  OAI211_X1 U15156 ( .C1(n13743), .C2(n13673), .A(n13669), .B(n13668), .ZN(
        P3_U3480) );
  INV_X1 U15157 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13670) );
  MUX2_X1 U15158 ( .A(n13670), .B(n13744), .S(n15894), .Z(n13672) );
  NAND2_X1 U15159 ( .A1(n13746), .A2(n13688), .ZN(n13671) );
  OAI211_X1 U15160 ( .C1(n13750), .C2(n13673), .A(n13672), .B(n13671), .ZN(
        P3_U3479) );
  NAND2_X1 U15161 ( .A1(n13674), .A2(n15891), .ZN(n13675) );
  NAND2_X1 U15162 ( .A1(n13676), .A2(n13675), .ZN(n13751) );
  MUX2_X1 U15163 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13751), .S(n15894), .Z(
        n13677) );
  AOI21_X1 U15164 ( .B1(n13688), .B2(n13753), .A(n13677), .ZN(n13678) );
  INV_X1 U15165 ( .A(n13678), .ZN(P3_U3478) );
  NAND2_X1 U15166 ( .A1(n13679), .A2(n15891), .ZN(n13680) );
  NAND2_X1 U15167 ( .A1(n13681), .A2(n13680), .ZN(n13755) );
  MUX2_X1 U15168 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13755), .S(n15894), .Z(
        n13682) );
  AOI21_X1 U15169 ( .B1(n13688), .B2(n13757), .A(n13682), .ZN(n13683) );
  INV_X1 U15170 ( .A(n13683), .ZN(P3_U3477) );
  NAND2_X1 U15171 ( .A1(n13684), .A2(n15891), .ZN(n13685) );
  NAND2_X1 U15172 ( .A1(n13686), .A2(n13685), .ZN(n13759) );
  MUX2_X1 U15173 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13759), .S(n15894), .Z(
        n13687) );
  AOI21_X1 U15174 ( .B1(n13688), .B2(n13761), .A(n13687), .ZN(n13689) );
  INV_X1 U15175 ( .A(n13689), .ZN(P3_U3476) );
  INV_X1 U15176 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13692) );
  AOI21_X1 U15177 ( .B1(n15891), .B2(n13691), .A(n13690), .ZN(n13764) );
  MUX2_X1 U15178 ( .A(n13692), .B(n13764), .S(n15894), .Z(n13693) );
  OAI21_X1 U15179 ( .B1(n13768), .B2(n13694), .A(n13693), .ZN(P3_U3475) );
  NAND2_X1 U15180 ( .A1(n13695), .A2(n15891), .ZN(n13697) );
  OAI211_X1 U15181 ( .C1(n13698), .C2(n15886), .A(n13697), .B(n13696), .ZN(
        n13769) );
  MUX2_X1 U15182 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13769), .S(n15894), .Z(
        P3_U3474) );
  NAND2_X1 U15183 ( .A1(n13699), .A2(n15891), .ZN(n13701) );
  OAI211_X1 U15184 ( .C1(n13702), .C2(n15886), .A(n13701), .B(n13700), .ZN(
        n13770) );
  MUX2_X1 U15185 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n13770), .S(n15894), .Z(
        P3_U3473) );
  NOR2_X1 U15186 ( .A1(n13703), .A2(n15895), .ZN(n13706) );
  AOI21_X1 U15187 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15895), .A(n13706), 
        .ZN(n13704) );
  OAI21_X1 U15188 ( .B1(n13705), .B2(n13767), .A(n13704), .ZN(P3_U3458) );
  AOI21_X1 U15189 ( .B1(n15895), .B2(P3_REG0_REG_30__SCAN_IN), .A(n13706), 
        .ZN(n13707) );
  OAI21_X1 U15190 ( .B1(n13708), .B2(n13767), .A(n13707), .ZN(P3_U3457) );
  MUX2_X1 U15191 ( .A(n13709), .B(P3_REG0_REG_27__SCAN_IN), .S(n15895), .Z(
        n13713) );
  OAI22_X1 U15192 ( .A1(n13711), .A2(n13749), .B1(n13710), .B2(n13767), .ZN(
        n13712) );
  MUX2_X1 U15193 ( .A(n13714), .B(P3_REG0_REG_26__SCAN_IN), .S(n15895), .Z(
        n13718) );
  OAI22_X1 U15194 ( .A1(n13716), .A2(n13749), .B1(n13715), .B2(n13767), .ZN(
        n13717) );
  OR2_X1 U15195 ( .A1(n13718), .A2(n13717), .ZN(P3_U3453) );
  MUX2_X1 U15196 ( .A(n13719), .B(P3_REG0_REG_25__SCAN_IN), .S(n15895), .Z(
        n13723) );
  OAI22_X1 U15197 ( .A1(n13721), .A2(n13749), .B1(n13720), .B2(n13767), .ZN(
        n13722) );
  OR2_X1 U15198 ( .A1(n13723), .A2(n13722), .ZN(P3_U3452) );
  INV_X1 U15199 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13725) );
  MUX2_X1 U15200 ( .A(n13725), .B(n13724), .S(n15898), .Z(n13726) );
  OAI21_X1 U15201 ( .B1(n13727), .B2(n13749), .A(n13726), .ZN(P3_U3451) );
  INV_X1 U15202 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13728) );
  MUX2_X1 U15203 ( .A(n13729), .B(n13728), .S(n15895), .Z(n13730) );
  OAI21_X1 U15204 ( .B1(n13731), .B2(n13767), .A(n13730), .ZN(P3_U3450) );
  INV_X1 U15205 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13733) );
  MUX2_X1 U15206 ( .A(n13733), .B(n13732), .S(n15898), .Z(n13736) );
  INV_X1 U15207 ( .A(n13767), .ZN(n13762) );
  NAND2_X1 U15208 ( .A1(n13734), .A2(n13762), .ZN(n13735) );
  OAI211_X1 U15209 ( .C1(n13737), .C2(n13749), .A(n13736), .B(n13735), .ZN(
        P3_U3449) );
  INV_X1 U15210 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13739) );
  MUX2_X1 U15211 ( .A(n13739), .B(n13738), .S(n15898), .Z(n13742) );
  NAND2_X1 U15212 ( .A1(n13740), .A2(n13762), .ZN(n13741) );
  OAI211_X1 U15213 ( .C1(n13743), .C2(n13749), .A(n13742), .B(n13741), .ZN(
        P3_U3448) );
  INV_X1 U15214 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13745) );
  MUX2_X1 U15215 ( .A(n13745), .B(n13744), .S(n15898), .Z(n13748) );
  NAND2_X1 U15216 ( .A1(n13746), .A2(n13762), .ZN(n13747) );
  OAI211_X1 U15217 ( .C1(n13750), .C2(n13749), .A(n13748), .B(n13747), .ZN(
        P3_U3447) );
  MUX2_X1 U15218 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13751), .S(n15898), .Z(
        n13752) );
  AOI21_X1 U15219 ( .B1(n13762), .B2(n13753), .A(n13752), .ZN(n13754) );
  INV_X1 U15220 ( .A(n13754), .ZN(P3_U3446) );
  MUX2_X1 U15221 ( .A(n13755), .B(P3_REG0_REG_18__SCAN_IN), .S(n15895), .Z(
        n13756) );
  AOI21_X1 U15222 ( .B1(n13762), .B2(n13757), .A(n13756), .ZN(n13758) );
  INV_X1 U15223 ( .A(n13758), .ZN(P3_U3444) );
  MUX2_X1 U15224 ( .A(n13759), .B(P3_REG0_REG_17__SCAN_IN), .S(n15895), .Z(
        n13760) );
  AOI21_X1 U15225 ( .B1(n13762), .B2(n13761), .A(n13760), .ZN(n13763) );
  INV_X1 U15226 ( .A(n13763), .ZN(P3_U3441) );
  INV_X1 U15227 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13765) );
  MUX2_X1 U15228 ( .A(n13765), .B(n13764), .S(n15898), .Z(n13766) );
  OAI21_X1 U15229 ( .B1(n13768), .B2(n13767), .A(n13766), .ZN(P3_U3438) );
  MUX2_X1 U15230 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13769), .S(n15898), .Z(
        P3_U3435) );
  MUX2_X1 U15231 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n13770), .S(n15898), .Z(
        P3_U3432) );
  MUX2_X1 U15232 ( .A(P3_D_REG_1__SCAN_IN), .B(n13771), .S(n13772), .Z(
        P3_U3377) );
  MUX2_X1 U15233 ( .A(P3_D_REG_0__SCAN_IN), .B(n13773), .S(n13772), .Z(
        P3_U3376) );
  INV_X1 U15234 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13774) );
  NAND3_X1 U15235 ( .A1(n13774), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13776) );
  OAI22_X1 U15236 ( .A1(n13777), .A2(n13776), .B1(n13775), .B2(n13995), .ZN(
        n13778) );
  AOI21_X1 U15237 ( .B1(n13780), .B2(n13779), .A(n13778), .ZN(n13781) );
  INV_X1 U15238 ( .A(n13781), .ZN(P3_U3264) );
  INV_X1 U15239 ( .A(n13782), .ZN(n13783) );
  OAI222_X1 U15240 ( .A1(n13787), .A2(n13785), .B1(P3_U3151), .B2(n13784), 
        .C1(n13993), .C2(n13783), .ZN(P3_U3266) );
  INV_X1 U15241 ( .A(n13786), .ZN(n13788) );
  XNOR2_X1 U15242 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n13991)
         );
  OAI22_X1 U15243 ( .A1(n13878), .A2(keyinput_59), .B1(keyinput_60), .B2(
        P3_REG3_REG_18__SCAN_IN), .ZN(n13790) );
  AOI221_X1 U15244 ( .B1(n13878), .B2(keyinput_59), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_60), .A(n13790), .ZN(n13875) );
  OAI22_X1 U15245 ( .A1(n8502), .A2(keyinput_56), .B1(keyinput_54), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n13791) );
  AOI221_X1 U15246 ( .B1(n8502), .B2(keyinput_56), .C1(P3_REG3_REG_0__SCAN_IN), 
        .C2(keyinput_54), .A(n13791), .ZN(n13873) );
  OAI22_X1 U15247 ( .A1(n13793), .A2(keyinput_58), .B1(keyinput_55), .B2(
        P3_REG3_REG_20__SCAN_IN), .ZN(n13792) );
  AOI221_X1 U15248 ( .B1(n13793), .B2(keyinput_58), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_55), .A(n13792), .ZN(n13872) );
  OAI22_X1 U15249 ( .A1(n13972), .A2(keyinput_57), .B1(n8262), .B2(keyinput_53), .ZN(n13794) );
  AOI221_X1 U15250 ( .B1(n13972), .B2(keyinput_57), .C1(keyinput_53), .C2(
        n8262), .A(n13794), .ZN(n13871) );
  XNOR2_X1 U15251 ( .A(keyinput_49), .B(n8418), .ZN(n13869) );
  OAI22_X1 U15252 ( .A1(n13963), .A2(keyinput_52), .B1(keyinput_51), .B2(
        P3_REG3_REG_24__SCAN_IN), .ZN(n13795) );
  AOI221_X1 U15253 ( .B1(n13963), .B2(keyinput_52), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_51), .A(n13795), .ZN(n13868) );
  OAI22_X1 U15254 ( .A1(n13961), .A2(keyinput_48), .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_50), .ZN(n13796) );
  AOI221_X1 U15255 ( .B1(n13961), .B2(keyinput_48), .C1(keyinput_50), .C2(
        P3_REG3_REG_17__SCAN_IN), .A(n13796), .ZN(n13867) );
  INV_X1 U15256 ( .A(keyinput_47), .ZN(n13865) );
  INV_X1 U15257 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n13947) );
  INV_X1 U15258 ( .A(keyinput_41), .ZN(n13855) );
  OAI22_X1 U15259 ( .A1(SI_0_), .A2(keyinput_32), .B1(keyinput_33), .B2(
        P3_RD_REG_SCAN_IN), .ZN(n13797) );
  AOI221_X1 U15260 ( .B1(SI_0_), .B2(keyinput_32), .C1(P3_RD_REG_SCAN_IN), 
        .C2(keyinput_33), .A(n13797), .ZN(n13849) );
  INV_X1 U15261 ( .A(keyinput_25), .ZN(n13834) );
  AND2_X1 U15262 ( .A1(keyinput_25), .A2(n8324), .ZN(n13833) );
  AOI22_X1 U15263 ( .A1(n13799), .A2(keyinput_15), .B1(n13898), .B2(
        keyinput_14), .ZN(n13798) );
  OAI221_X1 U15264 ( .B1(n13799), .B2(keyinput_15), .C1(n13898), .C2(
        keyinput_14), .A(n13798), .ZN(n13806) );
  AOI22_X1 U15265 ( .A1(n9283), .A2(keyinput_10), .B1(keyinput_12), .B2(n13896), .ZN(n13800) );
  OAI221_X1 U15266 ( .B1(n9283), .B2(keyinput_10), .C1(n13896), .C2(
        keyinput_12), .A(n13800), .ZN(n13805) );
  AOI22_X1 U15267 ( .A1(SI_16_), .A2(keyinput_16), .B1(SI_19_), .B2(
        keyinput_13), .ZN(n13801) );
  OAI221_X1 U15268 ( .B1(SI_16_), .B2(keyinput_16), .C1(SI_19_), .C2(
        keyinput_13), .A(n13801), .ZN(n13804) );
  AOI22_X1 U15269 ( .A1(SI_21_), .A2(keyinput_11), .B1(SI_23_), .B2(keyinput_9), .ZN(n13802) );
  OAI221_X1 U15270 ( .B1(SI_21_), .B2(keyinput_11), .C1(SI_23_), .C2(
        keyinput_9), .A(n13802), .ZN(n13803) );
  NOR4_X1 U15271 ( .A1(n13806), .A2(n13805), .A3(n13804), .A4(n13803), .ZN(
        n13819) );
  INV_X1 U15272 ( .A(keyinput_1), .ZN(n13809) );
  AOI22_X1 U15273 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_30_), .B2(
        keyinput_2), .ZN(n13807) );
  OAI221_X1 U15274 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_30_), 
        .C2(keyinput_2), .A(n13807), .ZN(n13808) );
  AOI221_X1 U15275 ( .B1(SI_31_), .B2(keyinput_1), .C1(n13775), .C2(n13809), 
        .A(n13808), .ZN(n13817) );
  AOI22_X1 U15276 ( .A1(SI_28_), .A2(keyinput_4), .B1(SI_29_), .B2(keyinput_3), 
        .ZN(n13810) );
  OAI221_X1 U15277 ( .B1(SI_28_), .B2(keyinput_4), .C1(SI_29_), .C2(keyinput_3), .A(n13810), .ZN(n13816) );
  OAI22_X1 U15278 ( .A1(n13812), .A2(keyinput_6), .B1(keyinput_8), .B2(SI_24_), 
        .ZN(n13811) );
  AOI221_X1 U15279 ( .B1(n13812), .B2(keyinput_6), .C1(SI_24_), .C2(keyinput_8), .A(n13811), .ZN(n13815) );
  OAI22_X1 U15280 ( .A1(SI_27_), .A2(keyinput_5), .B1(keyinput_7), .B2(SI_25_), 
        .ZN(n13813) );
  AOI221_X1 U15281 ( .B1(SI_27_), .B2(keyinput_5), .C1(SI_25_), .C2(keyinput_7), .A(n13813), .ZN(n13814) );
  OAI211_X1 U15282 ( .C1(n13817), .C2(n13816), .A(n13815), .B(n13814), .ZN(
        n13818) );
  AOI22_X1 U15283 ( .A1(n13819), .A2(n13818), .B1(keyinput_17), .B2(n13821), 
        .ZN(n13820) );
  OAI21_X1 U15284 ( .B1(keyinput_17), .B2(n13821), .A(n13820), .ZN(n13824) );
  AOI22_X1 U15285 ( .A1(SI_13_), .A2(keyinput_19), .B1(SI_14_), .B2(
        keyinput_18), .ZN(n13822) );
  OAI221_X1 U15286 ( .B1(SI_13_), .B2(keyinput_19), .C1(SI_14_), .C2(
        keyinput_18), .A(n13822), .ZN(n13823) );
  OAI22_X1 U15287 ( .A1(n13824), .A2(n13823), .B1(SI_10_), .B2(keyinput_22), 
        .ZN(n13825) );
  AOI21_X1 U15288 ( .B1(SI_10_), .B2(keyinput_22), .A(n13825), .ZN(n13831) );
  OAI22_X1 U15289 ( .A1(SI_12_), .A2(keyinput_20), .B1(SI_11_), .B2(
        keyinput_21), .ZN(n13826) );
  AOI221_X1 U15290 ( .B1(SI_12_), .B2(keyinput_20), .C1(keyinput_21), .C2(
        SI_11_), .A(n13826), .ZN(n13830) );
  XNOR2_X1 U15291 ( .A(n13827), .B(keyinput_23), .ZN(n13829) );
  XNOR2_X1 U15292 ( .A(SI_8_), .B(keyinput_24), .ZN(n13828) );
  AOI211_X1 U15293 ( .C1(n13831), .C2(n13830), .A(n13829), .B(n13828), .ZN(
        n13832) );
  AOI211_X1 U15294 ( .C1(SI_7_), .C2(n13834), .A(n13833), .B(n13832), .ZN(
        n13843) );
  AOI22_X1 U15295 ( .A1(SI_6_), .A2(keyinput_26), .B1(n13836), .B2(keyinput_27), .ZN(n13835) );
  OAI221_X1 U15296 ( .B1(SI_6_), .B2(keyinput_26), .C1(n13836), .C2(
        keyinput_27), .A(n13835), .ZN(n13842) );
  OAI22_X1 U15297 ( .A1(n13925), .A2(keyinput_29), .B1(n10819), .B2(
        keyinput_31), .ZN(n13837) );
  AOI221_X1 U15298 ( .B1(n13925), .B2(keyinput_29), .C1(keyinput_31), .C2(
        n10819), .A(n13837), .ZN(n13841) );
  XNOR2_X1 U15299 ( .A(n7509), .B(keyinput_30), .ZN(n13839) );
  XNOR2_X1 U15300 ( .A(SI_4_), .B(keyinput_28), .ZN(n13838) );
  NOR2_X1 U15301 ( .A1(n13839), .A2(n13838), .ZN(n13840) );
  OAI211_X1 U15302 ( .C1(n13843), .C2(n13842), .A(n13841), .B(n13840), .ZN(
        n13848) );
  AOI22_X1 U15303 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_36), .B1(
        P3_U3151), .B2(keyinput_34), .ZN(n13844) );
  OAI221_X1 U15304 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .C1(
        P3_U3151), .C2(keyinput_34), .A(n13844), .ZN(n13847) );
  AOI22_X1 U15305 ( .A1(n13935), .A2(keyinput_39), .B1(n13936), .B2(
        keyinput_37), .ZN(n13845) );
  OAI221_X1 U15306 ( .B1(n13935), .B2(keyinput_39), .C1(n13936), .C2(
        keyinput_37), .A(n13845), .ZN(n13846) );
  AOI211_X1 U15307 ( .C1(n13849), .C2(n13848), .A(n13847), .B(n13846), .ZN(
        n13853) );
  OAI22_X1 U15308 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_38), .B1(
        keyinput_35), .B2(P3_REG3_REG_7__SCAN_IN), .ZN(n13850) );
  AOI221_X1 U15309 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput_35), .A(n13850), .ZN(n13852) );
  NOR2_X1 U15310 ( .A1(n13944), .A2(keyinput_40), .ZN(n13851) );
  AOI221_X1 U15311 ( .B1(n13853), .B2(n13852), .C1(keyinput_40), .C2(n13944), 
        .A(n13851), .ZN(n13854) );
  AOI221_X1 U15312 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_41), .C1(
        n13947), .C2(n13855), .A(n13854), .ZN(n13863) );
  XNOR2_X1 U15313 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n13862)
         );
  OAI22_X1 U15314 ( .A1(n13858), .A2(keyinput_46), .B1(n13857), .B2(
        keyinput_43), .ZN(n13856) );
  AOI221_X1 U15315 ( .B1(n13858), .B2(keyinput_46), .C1(keyinput_43), .C2(
        n13857), .A(n13856), .ZN(n13861) );
  OAI22_X1 U15316 ( .A1(n8641), .A2(keyinput_45), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(keyinput_44), .ZN(n13859) );
  AOI221_X1 U15317 ( .B1(n8641), .B2(keyinput_45), .C1(keyinput_44), .C2(
        P3_REG3_REG_1__SCAN_IN), .A(n13859), .ZN(n13860) );
  OAI211_X1 U15318 ( .C1(n13863), .C2(n13862), .A(n13861), .B(n13860), .ZN(
        n13864) );
  OAI221_X1 U15319 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n13865), .C1(n13957), 
        .C2(keyinput_47), .A(n13864), .ZN(n13866) );
  NAND4_X1 U15320 ( .A1(n13869), .A2(n13868), .A3(n13867), .A4(n13866), .ZN(
        n13870) );
  NAND4_X1 U15321 ( .A1(n13873), .A2(n13872), .A3(n13871), .A4(n13870), .ZN(
        n13874) );
  AOI22_X1 U15322 ( .A1(n13875), .A2(n13874), .B1(keyinput_61), .B2(
        P3_REG3_REG_6__SCAN_IN), .ZN(n13876) );
  OAI21_X1 U15323 ( .B1(keyinput_61), .B2(P3_REG3_REG_6__SCAN_IN), .A(n13876), 
        .ZN(n13990) );
  INV_X1 U15324 ( .A(keyinput_126), .ZN(n13983) );
  AOI22_X1 U15325 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_124), .B1(
        n13878), .B2(keyinput_123), .ZN(n13877) );
  OAI221_X1 U15326 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .C1(
        n13878), .C2(keyinput_123), .A(n13877), .ZN(n13980) );
  XOR2_X1 U15327 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_115), .Z(n13967)
         );
  INV_X1 U15328 ( .A(keyinput_111), .ZN(n13958) );
  INV_X1 U15329 ( .A(keyinput_105), .ZN(n13948) );
  INV_X1 U15330 ( .A(keyinput_104), .ZN(n13945) );
  INV_X1 U15331 ( .A(keyinput_89), .ZN(n13921) );
  OAI22_X1 U15332 ( .A1(n8092), .A2(keyinput_82), .B1(n13880), .B2(keyinput_83), .ZN(n13879) );
  AOI221_X1 U15333 ( .B1(n8092), .B2(keyinput_82), .C1(keyinput_83), .C2(
        n13880), .A(n13879), .ZN(n13910) );
  INV_X1 U15334 ( .A(keyinput_65), .ZN(n13884) );
  AOI22_X1 U15335 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(n13882), 
        .B2(keyinput_66), .ZN(n13881) );
  OAI221_X1 U15336 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(n13882), 
        .C2(keyinput_66), .A(n13881), .ZN(n13883) );
  AOI221_X1 U15337 ( .B1(SI_31_), .B2(keyinput_65), .C1(n13775), .C2(n13884), 
        .A(n13883), .ZN(n13893) );
  AOI22_X1 U15338 ( .A1(SI_29_), .A2(keyinput_67), .B1(n12904), .B2(
        keyinput_68), .ZN(n13885) );
  OAI221_X1 U15339 ( .B1(SI_29_), .B2(keyinput_67), .C1(n12904), .C2(
        keyinput_68), .A(n13885), .ZN(n13892) );
  OAI22_X1 U15340 ( .A1(n13888), .A2(keyinput_69), .B1(n13887), .B2(
        keyinput_72), .ZN(n13886) );
  AOI221_X1 U15341 ( .B1(n13888), .B2(keyinput_69), .C1(keyinput_72), .C2(
        n13887), .A(n13886), .ZN(n13891) );
  OAI22_X1 U15342 ( .A1(SI_26_), .A2(keyinput_70), .B1(keyinput_71), .B2(
        SI_25_), .ZN(n13889) );
  AOI221_X1 U15343 ( .B1(SI_26_), .B2(keyinput_70), .C1(SI_25_), .C2(
        keyinput_71), .A(n13889), .ZN(n13890) );
  OAI211_X1 U15344 ( .C1(n13893), .C2(n13892), .A(n13891), .B(n13890), .ZN(
        n13908) );
  AOI22_X1 U15345 ( .A1(n13896), .A2(keyinput_76), .B1(n13895), .B2(
        keyinput_75), .ZN(n13894) );
  OAI221_X1 U15346 ( .B1(n13896), .B2(keyinput_76), .C1(n13895), .C2(
        keyinput_75), .A(n13894), .ZN(n13905) );
  AOI22_X1 U15347 ( .A1(n9283), .A2(keyinput_74), .B1(keyinput_78), .B2(n13898), .ZN(n13897) );
  OAI221_X1 U15348 ( .B1(n9283), .B2(keyinput_74), .C1(n13898), .C2(
        keyinput_78), .A(n13897), .ZN(n13904) );
  AOI22_X1 U15349 ( .A1(SI_17_), .A2(keyinput_79), .B1(SI_19_), .B2(
        keyinput_77), .ZN(n13899) );
  OAI221_X1 U15350 ( .B1(SI_17_), .B2(keyinput_79), .C1(SI_19_), .C2(
        keyinput_77), .A(n13899), .ZN(n13903) );
  AOI22_X1 U15351 ( .A1(SI_23_), .A2(keyinput_73), .B1(n13901), .B2(
        keyinput_80), .ZN(n13900) );
  OAI221_X1 U15352 ( .B1(SI_23_), .B2(keyinput_73), .C1(n13901), .C2(
        keyinput_80), .A(n13900), .ZN(n13902) );
  NOR4_X1 U15353 ( .A1(n13905), .A2(n13904), .A3(n13903), .A4(n13902), .ZN(
        n13907) );
  NOR2_X1 U15354 ( .A1(keyinput_81), .A2(SI_15_), .ZN(n13906) );
  AOI221_X1 U15355 ( .B1(n13908), .B2(n13907), .C1(SI_15_), .C2(keyinput_81), 
        .A(n13906), .ZN(n13909) );
  AOI22_X1 U15356 ( .A1(n13910), .A2(n13909), .B1(keyinput_85), .B2(n13912), 
        .ZN(n13911) );
  OAI21_X1 U15357 ( .B1(keyinput_85), .B2(n13912), .A(n13911), .ZN(n13919) );
  AOI22_X1 U15358 ( .A1(n13915), .A2(keyinput_86), .B1(n13914), .B2(
        keyinput_84), .ZN(n13913) );
  OAI221_X1 U15359 ( .B1(n13915), .B2(keyinput_86), .C1(n13914), .C2(
        keyinput_84), .A(n13913), .ZN(n13918) );
  OAI22_X1 U15360 ( .A1(SI_9_), .A2(keyinput_87), .B1(keyinput_88), .B2(SI_8_), 
        .ZN(n13916) );
  AOI221_X1 U15361 ( .B1(SI_9_), .B2(keyinput_87), .C1(SI_8_), .C2(keyinput_88), .A(n13916), .ZN(n13917) );
  OAI21_X1 U15362 ( .B1(n13919), .B2(n13918), .A(n13917), .ZN(n13920) );
  OAI221_X1 U15363 ( .B1(SI_7_), .B2(keyinput_89), .C1(n8324), .C2(n13921), 
        .A(n13920), .ZN(n13931) );
  OAI22_X1 U15364 ( .A1(n13923), .A2(keyinput_90), .B1(SI_5_), .B2(keyinput_91), .ZN(n13922) );
  AOI221_X1 U15365 ( .B1(n13923), .B2(keyinput_90), .C1(keyinput_91), .C2(
        SI_5_), .A(n13922), .ZN(n13930) );
  AOI22_X1 U15366 ( .A1(SI_4_), .A2(keyinput_92), .B1(n13925), .B2(keyinput_93), .ZN(n13924) );
  OAI221_X1 U15367 ( .B1(SI_4_), .B2(keyinput_92), .C1(n13925), .C2(
        keyinput_93), .A(n13924), .ZN(n13929) );
  XOR2_X1 U15368 ( .A(n10819), .B(keyinput_95), .Z(n13927) );
  XNOR2_X1 U15369 ( .A(SI_2_), .B(keyinput_94), .ZN(n13926) );
  NAND2_X1 U15370 ( .A1(n13927), .A2(n13926), .ZN(n13928) );
  AOI211_X1 U15371 ( .C1(n13931), .C2(n13930), .A(n13929), .B(n13928), .ZN(
        n13940) );
  INV_X1 U15372 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15653) );
  AOI22_X1 U15373 ( .A1(n9713), .A2(keyinput_96), .B1(keyinput_97), .B2(n15653), .ZN(n13932) );
  OAI221_X1 U15374 ( .B1(n9713), .B2(keyinput_96), .C1(n15653), .C2(
        keyinput_97), .A(n13932), .ZN(n13939) );
  OAI22_X1 U15375 ( .A1(P3_U3151), .A2(keyinput_98), .B1(keyinput_102), .B2(
        P3_REG3_REG_23__SCAN_IN), .ZN(n13933) );
  AOI221_X1 U15376 ( .B1(P3_U3151), .B2(keyinput_98), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_102), .A(n13933), .ZN(n13938)
         );
  OAI22_X1 U15377 ( .A1(n13936), .A2(keyinput_101), .B1(n13935), .B2(
        keyinput_103), .ZN(n13934) );
  AOI221_X1 U15378 ( .B1(n13936), .B2(keyinput_101), .C1(keyinput_103), .C2(
        n13935), .A(n13934), .ZN(n13937) );
  OAI211_X1 U15379 ( .C1(n13940), .C2(n13939), .A(n13938), .B(n13937), .ZN(
        n13943) );
  AOI22_X1 U15380 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_99), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .ZN(n13941) );
  OAI221_X1 U15381 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_100), .A(n13941), .ZN(n13942)
         );
  OAI222_X1 U15382 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(n13945), .B1(n13944), 
        .B2(keyinput_104), .C1(n13943), .C2(n13942), .ZN(n13946) );
  OAI221_X1 U15383 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(n13948), .C1(n13947), 
        .C2(keyinput_105), .A(n13946), .ZN(n13955) );
  XOR2_X1 U15384 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_106), .Z(n13954)
         );
  AOI22_X1 U15385 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(n8641), 
        .B2(keyinput_109), .ZN(n13949) );
  OAI221_X1 U15386 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(n8641), .C2(keyinput_109), .A(n13949), .ZN(n13953) );
  XNOR2_X1 U15387 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_108), .ZN(n13951)
         );
  XNOR2_X1 U15388 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_110), .ZN(n13950)
         );
  NAND2_X1 U15389 ( .A1(n13951), .A2(n13950), .ZN(n13952) );
  AOI211_X1 U15390 ( .C1(n13955), .C2(n13954), .A(n13953), .B(n13952), .ZN(
        n13956) );
  AOI221_X1 U15391 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n13958), .C1(n13957), 
        .C2(keyinput_111), .A(n13956), .ZN(n13966) );
  AOI22_X1 U15392 ( .A1(n13961), .A2(keyinput_112), .B1(n13960), .B2(
        keyinput_114), .ZN(n13959) );
  OAI221_X1 U15393 ( .B1(n13961), .B2(keyinput_112), .C1(n13960), .C2(
        keyinput_114), .A(n13959), .ZN(n13965) );
  AOI22_X1 U15394 ( .A1(n8418), .A2(keyinput_113), .B1(keyinput_116), .B2(
        n13963), .ZN(n13962) );
  OAI221_X1 U15395 ( .B1(n8418), .B2(keyinput_113), .C1(n13963), .C2(
        keyinput_116), .A(n13962), .ZN(n13964) );
  NOR4_X1 U15396 ( .A1(n13967), .A2(n13966), .A3(n13965), .A4(n13964), .ZN(
        n13976) );
  AOI22_X1 U15397 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_122), .B1(
        P3_REG3_REG_13__SCAN_IN), .B2(keyinput_120), .ZN(n13968) );
  OAI221_X1 U15398 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_120), .A(n13968), .ZN(n13975)
         );
  AOI22_X1 U15399 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_118), .B1(n8262), 
        .B2(keyinput_117), .ZN(n13969) );
  OAI221_X1 U15400 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .C1(n8262), .C2(keyinput_117), .A(n13969), .ZN(n13974) );
  AOI22_X1 U15401 ( .A1(n13972), .A2(keyinput_121), .B1(keyinput_119), .B2(
        n13971), .ZN(n13970) );
  OAI221_X1 U15402 ( .B1(n13972), .B2(keyinput_121), .C1(n13971), .C2(
        keyinput_119), .A(n13970), .ZN(n13973) );
  NOR4_X1 U15403 ( .A1(n13976), .A2(n13975), .A3(n13974), .A4(n13973), .ZN(
        n13979) );
  NAND2_X1 U15404 ( .A1(n13978), .A2(keyinput_125), .ZN(n13977) );
  OAI221_X1 U15405 ( .B1(n13980), .B2(n13979), .C1(n13978), .C2(keyinput_125), 
        .A(n13977), .ZN(n13981) );
  OAI221_X1 U15406 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(n13983), .C1(n13982), 
        .C2(keyinput_126), .A(n13981), .ZN(n13985) );
  INV_X1 U15407 ( .A(keyinput_63), .ZN(n13987) );
  AOI21_X1 U15408 ( .B1(keyinput_127), .B2(n13985), .A(n13987), .ZN(n13988) );
  INV_X1 U15409 ( .A(keyinput_127), .ZN(n13984) );
  AOI21_X1 U15410 ( .B1(n13985), .B2(n13984), .A(P3_REG3_REG_15__SCAN_IN), 
        .ZN(n13986) );
  AOI22_X1 U15411 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(n13988), .B1(n13987), 
        .B2(n13986), .ZN(n13989) );
  AOI21_X1 U15412 ( .B1(n13991), .B2(n13990), .A(n13989), .ZN(n13998) );
  OAI222_X1 U15413 ( .A1(P3_U3151), .A2(n13996), .B1(n13995), .B2(n13994), 
        .C1(n13993), .C2(n13992), .ZN(n13997) );
  XOR2_X1 U15414 ( .A(n13998), .B(n13997), .Z(P3_U3270) );
  MUX2_X1 U15415 ( .A(n13999), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  INV_X1 U15416 ( .A(n14448), .ZN(n14051) );
  NOR2_X1 U15417 ( .A1(n14000), .A2(n7209), .ZN(n14037) );
  XNOR2_X1 U15418 ( .A(n14531), .B(n14072), .ZN(n14036) );
  INV_X1 U15419 ( .A(n14001), .ZN(n14002) );
  NAND2_X1 U15420 ( .A1(n14003), .A2(n14002), .ZN(n14100) );
  XNOR2_X1 U15421 ( .A(n14557), .B(n14038), .ZN(n14005) );
  AND2_X1 U15422 ( .A1(n14177), .A2(n14360), .ZN(n14004) );
  NOR2_X1 U15423 ( .A1(n14005), .A2(n14004), .ZN(n14006) );
  AOI21_X1 U15424 ( .B1(n14005), .B2(n14004), .A(n14006), .ZN(n14101) );
  NAND2_X1 U15425 ( .A1(n14100), .A2(n14101), .ZN(n14099) );
  INV_X1 U15426 ( .A(n14006), .ZN(n14007) );
  NAND2_X1 U15427 ( .A1(n14099), .A2(n14007), .ZN(n14138) );
  NOR2_X1 U15428 ( .A1(n14008), .A2(n7209), .ZN(n14009) );
  XNOR2_X1 U15429 ( .A(n14500), .B(n14072), .ZN(n14011) );
  XOR2_X1 U15430 ( .A(n14009), .B(n14011), .Z(n14137) );
  INV_X1 U15431 ( .A(n14009), .ZN(n14010) );
  XNOR2_X1 U15432 ( .A(n14405), .B(n14072), .ZN(n14013) );
  NAND2_X1 U15433 ( .A1(n14175), .A2(n14360), .ZN(n14012) );
  NAND2_X1 U15434 ( .A1(n14013), .A2(n14012), .ZN(n14014) );
  OAI21_X1 U15435 ( .B1(n14013), .B2(n14012), .A(n14014), .ZN(n14063) );
  XNOR2_X1 U15436 ( .A(n14392), .B(n14038), .ZN(n14016) );
  AND2_X1 U15437 ( .A1(n14174), .A2(n14360), .ZN(n14015) );
  NAND2_X1 U15438 ( .A1(n14016), .A2(n14015), .ZN(n14117) );
  XNOR2_X1 U15439 ( .A(n14376), .B(n14072), .ZN(n14020) );
  NOR2_X1 U15440 ( .A1(n14017), .A2(n7209), .ZN(n14018) );
  XNOR2_X1 U15441 ( .A(n14020), .B(n14018), .ZN(n14081) );
  NAND2_X1 U15442 ( .A1(n14082), .A2(n14081), .ZN(n14080) );
  INV_X1 U15443 ( .A(n14018), .ZN(n14019) );
  NOR2_X1 U15444 ( .A1(n14022), .A2(n7209), .ZN(n14125) );
  XNOR2_X1 U15445 ( .A(n14469), .B(n14072), .ZN(n14025) );
  NOR2_X1 U15446 ( .A1(n14056), .A2(n7209), .ZN(n14055) );
  INV_X1 U15447 ( .A(n14024), .ZN(n14027) );
  INV_X1 U15448 ( .A(n14025), .ZN(n14026) );
  NAND2_X1 U15449 ( .A1(n14170), .A2(n14360), .ZN(n14029) );
  XNOR2_X1 U15450 ( .A(n14466), .B(n14072), .ZN(n14028) );
  XOR2_X1 U15451 ( .A(n14029), .B(n14028), .Z(n14111) );
  INV_X1 U15452 ( .A(n14028), .ZN(n14031) );
  INV_X1 U15453 ( .A(n14029), .ZN(n14030) );
  NOR2_X1 U15454 ( .A1(n14031), .A2(n14030), .ZN(n14032) );
  AOI21_X2 U15455 ( .B1(n14110), .B2(n14111), .A(n14032), .ZN(n14090) );
  XNOR2_X1 U15456 ( .A(n14323), .B(n14072), .ZN(n14148) );
  NAND2_X1 U15457 ( .A1(n14169), .A2(n14360), .ZN(n14033) );
  NOR2_X1 U15458 ( .A1(n14148), .A2(n14033), .ZN(n14034) );
  AOI21_X1 U15459 ( .B1(n14148), .B2(n14033), .A(n14034), .ZN(n14089) );
  NAND2_X1 U15460 ( .A1(n14090), .A2(n14089), .ZN(n14145) );
  XNOR2_X1 U15461 ( .A(n14036), .B(n14037), .ZN(n14149) );
  NOR2_X1 U15462 ( .A1(n14149), .A2(n14034), .ZN(n14035) );
  XNOR2_X1 U15463 ( .A(n14448), .B(n14038), .ZN(n14040) );
  AND2_X1 U15464 ( .A1(n14167), .A2(n14360), .ZN(n14039) );
  NAND2_X1 U15465 ( .A1(n14040), .A2(n14039), .ZN(n14070) );
  OAI21_X1 U15466 ( .B1(n14040), .B2(n14039), .A(n14070), .ZN(n14041) );
  AOI21_X1 U15467 ( .B1(n14042), .B2(n14041), .A(n14163), .ZN(n14043) );
  NAND2_X1 U15468 ( .A1(n14043), .A2(n14071), .ZN(n14050) );
  NAND2_X1 U15469 ( .A1(n14166), .A2(n14153), .ZN(n14045) );
  NAND2_X1 U15470 ( .A1(n14168), .A2(n14152), .ZN(n14044) );
  NAND2_X1 U15471 ( .A1(n14045), .A2(n14044), .ZN(n14287) );
  INV_X1 U15472 ( .A(n14296), .ZN(n14047) );
  OAI22_X1 U15473 ( .A1(n14047), .A2(n14092), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14046), .ZN(n14048) );
  AOI21_X1 U15474 ( .B1(n14287), .B2(n14095), .A(n14048), .ZN(n14049) );
  OAI211_X1 U15475 ( .C1(n14051), .C2(n14135), .A(n14050), .B(n14049), .ZN(
        P2_U3186) );
  NAND2_X1 U15476 ( .A1(n14170), .A2(n14153), .ZN(n14053) );
  NAND2_X1 U15477 ( .A1(n14172), .A2(n14152), .ZN(n14052) );
  NAND2_X1 U15478 ( .A1(n14053), .A2(n14052), .ZN(n14344) );
  AOI22_X1 U15479 ( .A1(n14344), .A2(n14095), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14054) );
  OAI21_X1 U15480 ( .B1(n14349), .B2(n14092), .A(n14054), .ZN(n14061) );
  NOR2_X1 U15481 ( .A1(n14055), .A2(n14163), .ZN(n14059) );
  NOR2_X1 U15482 ( .A1(n14056), .A2(n14146), .ZN(n14058) );
  MUX2_X1 U15483 ( .A(n14059), .B(n14058), .S(n14057), .Z(n14060) );
  AOI211_X1 U15484 ( .C1(n14469), .C2(n14159), .A(n14061), .B(n14060), .ZN(
        n14062) );
  INV_X1 U15485 ( .A(n14062), .ZN(P2_U3188) );
  AOI21_X1 U15486 ( .B1(n14064), .B2(n14063), .A(n7321), .ZN(n14069) );
  NOR2_X1 U15487 ( .A1(n14092), .A2(n14406), .ZN(n14067) );
  AND2_X1 U15488 ( .A1(n14176), .A2(n14152), .ZN(n14065) );
  AOI21_X1 U15489 ( .B1(n14174), .B2(n14153), .A(n14065), .ZN(n14414) );
  NAND2_X1 U15490 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n15348)
         );
  OAI21_X1 U15491 ( .B1(n14157), .B2(n14414), .A(n15348), .ZN(n14066) );
  AOI211_X1 U15492 ( .C1(n14405), .C2(n14159), .A(n14067), .B(n14066), .ZN(
        n14068) );
  OAI21_X1 U15493 ( .B1(n14069), .B2(n14163), .A(n14068), .ZN(P2_U3191) );
  MUX2_X1 U15494 ( .A(n14274), .B(n14444), .S(n14308), .Z(n14073) );
  NAND2_X1 U15495 ( .A1(n14165), .A2(n14153), .ZN(n14075) );
  NAND2_X1 U15496 ( .A1(n14167), .A2(n14152), .ZN(n14074) );
  NAND2_X1 U15497 ( .A1(n14075), .A2(n14074), .ZN(n14270) );
  OAI22_X1 U15498 ( .A1(n14279), .A2(n14092), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14076), .ZN(n14078) );
  NOR2_X1 U15499 ( .A1(n14283), .A2(n14135), .ZN(n14077) );
  AOI211_X1 U15500 ( .C1(n14095), .C2(n14270), .A(n14078), .B(n14077), .ZN(
        n14079) );
  OAI211_X1 U15501 ( .C1(n14082), .C2(n14081), .A(n14080), .B(n14102), .ZN(
        n14088) );
  INV_X1 U15502 ( .A(n14373), .ZN(n14086) );
  AND2_X1 U15503 ( .A1(n14174), .A2(n14152), .ZN(n14083) );
  AOI21_X1 U15504 ( .B1(n14172), .B2(n14153), .A(n14083), .ZN(n14381) );
  OAI22_X1 U15505 ( .A1(n14381), .A2(n14157), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14084), .ZN(n14085) );
  AOI21_X1 U15506 ( .B1(n14086), .B2(n14155), .A(n14085), .ZN(n14087) );
  OAI211_X1 U15507 ( .C1(n14545), .C2(n14135), .A(n14088), .B(n14087), .ZN(
        P2_U3195) );
  OAI211_X1 U15508 ( .C1(n14090), .C2(n14089), .A(n14145), .B(n14102), .ZN(
        n14098) );
  AOI22_X1 U15509 ( .A1(n14168), .A2(n14153), .B1(n14152), .B2(n14170), .ZN(
        n14318) );
  INV_X1 U15510 ( .A(n14318), .ZN(n14096) );
  INV_X1 U15511 ( .A(n14324), .ZN(n14093) );
  OAI22_X1 U15512 ( .A1(n14093), .A2(n14092), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14091), .ZN(n14094) );
  AOI21_X1 U15513 ( .B1(n14096), .B2(n14095), .A(n14094), .ZN(n14097) );
  OAI211_X1 U15514 ( .C1(n14535), .C2(n14135), .A(n14098), .B(n14097), .ZN(
        P2_U3197) );
  OAI21_X1 U15515 ( .B1(n14101), .B2(n14100), .A(n14099), .ZN(n14103) );
  NAND2_X1 U15516 ( .A1(n14103), .A2(n14102), .ZN(n14108) );
  NAND2_X1 U15517 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n15316)
         );
  OAI21_X1 U15518 ( .B1(n14157), .B2(n14104), .A(n15316), .ZN(n14105) );
  AOI21_X1 U15519 ( .B1(n14106), .B2(n14155), .A(n14105), .ZN(n14107) );
  OAI211_X1 U15520 ( .C1(n14109), .C2(n14135), .A(n14108), .B(n14107), .ZN(
        P2_U3200) );
  XOR2_X1 U15521 ( .A(n14111), .B(n14110), .Z(n14116) );
  AND2_X1 U15522 ( .A1(n14171), .A2(n14152), .ZN(n14112) );
  AOI21_X1 U15523 ( .B1(n14169), .B2(n14153), .A(n14112), .ZN(n14333) );
  AOI22_X1 U15524 ( .A1(n14337), .A2(n14155), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14113) );
  OAI21_X1 U15525 ( .B1(n14333), .B2(n14157), .A(n14113), .ZN(n14114) );
  AOI21_X1 U15526 ( .B1(n14466), .B2(n14159), .A(n14114), .ZN(n14115) );
  OAI21_X1 U15527 ( .B1(n14116), .B2(n14163), .A(n14115), .ZN(P2_U3201) );
  NAND2_X1 U15528 ( .A1(n7316), .A2(n14117), .ZN(n14118) );
  XNOR2_X1 U15529 ( .A(n14119), .B(n14118), .ZN(n14124) );
  AOI22_X1 U15530 ( .A1(n14173), .A2(n14153), .B1(n14152), .B2(n14175), .ZN(
        n14387) );
  OAI22_X1 U15531 ( .A1(n14387), .A2(n14157), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14120), .ZN(n14122) );
  NOR2_X1 U15532 ( .A1(n14549), .A2(n14135), .ZN(n14121) );
  AOI211_X1 U15533 ( .C1(n14155), .C2(n14393), .A(n14122), .B(n14121), .ZN(
        n14123) );
  OAI21_X1 U15534 ( .B1(n14124), .B2(n14163), .A(n14123), .ZN(P2_U3205) );
  INV_X1 U15535 ( .A(n14540), .ZN(n14136) );
  OR2_X1 U15536 ( .A1(n14125), .A2(n14163), .ZN(n14129) );
  NAND2_X1 U15537 ( .A1(n14126), .A2(n14172), .ZN(n14128) );
  MUX2_X1 U15538 ( .A(n14129), .B(n14128), .S(n14127), .Z(n14134) );
  AND2_X1 U15539 ( .A1(n14173), .A2(n14152), .ZN(n14130) );
  AOI21_X1 U15540 ( .B1(n14171), .B2(n14153), .A(n14130), .ZN(n14358) );
  OAI22_X1 U15541 ( .A1(n14358), .A2(n14157), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14131), .ZN(n14132) );
  AOI21_X1 U15542 ( .B1(n14363), .B2(n14155), .A(n14132), .ZN(n14133) );
  OAI211_X1 U15543 ( .C1(n14136), .C2(n14135), .A(n14134), .B(n14133), .ZN(
        P2_U3207) );
  XNOR2_X1 U15544 ( .A(n14138), .B(n14137), .ZN(n14144) );
  AND2_X1 U15545 ( .A1(n14177), .A2(n14152), .ZN(n14139) );
  AOI21_X1 U15546 ( .B1(n14175), .B2(n14153), .A(n14139), .ZN(n14422) );
  NAND2_X1 U15547 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n15334)
         );
  INV_X1 U15548 ( .A(n14140), .ZN(n14429) );
  NAND2_X1 U15549 ( .A1(n14155), .A2(n14429), .ZN(n14141) );
  OAI211_X1 U15550 ( .C1(n14157), .C2(n14422), .A(n15334), .B(n14141), .ZN(
        n14142) );
  AOI21_X1 U15551 ( .B1(n14500), .B2(n14159), .A(n14142), .ZN(n14143) );
  OAI21_X1 U15552 ( .B1(n14144), .B2(n14163), .A(n14143), .ZN(P2_U3210) );
  NOR2_X1 U15553 ( .A1(n14145), .A2(n14163), .ZN(n14151) );
  NOR3_X1 U15554 ( .A1(n14148), .A2(n14147), .A3(n14146), .ZN(n14150) );
  OAI21_X1 U15555 ( .B1(n14151), .B2(n14150), .A(n14149), .ZN(n14161) );
  AOI22_X1 U15556 ( .A1(n14167), .A2(n14153), .B1(n14152), .B2(n14169), .ZN(
        n14304) );
  INV_X1 U15557 ( .A(n14154), .ZN(n14311) );
  AOI22_X1 U15558 ( .A1(n14311), .A2(n14155), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14156) );
  OAI21_X1 U15559 ( .B1(n14304), .B2(n14157), .A(n14156), .ZN(n14158) );
  AOI21_X1 U15560 ( .B1(n7634), .B2(n14159), .A(n14158), .ZN(n14160) );
  OAI211_X1 U15561 ( .C1(n14163), .C2(n14162), .A(n14161), .B(n14160), .ZN(
        P2_U3212) );
  INV_X2 U15562 ( .A(P2_U3947), .ZN(n14186) );
  MUX2_X1 U15563 ( .A(n14247), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14186), .Z(
        P2_U3562) );
  MUX2_X1 U15564 ( .A(n14164), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14186), .Z(
        P2_U3561) );
  MUX2_X1 U15565 ( .A(n14165), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14186), .Z(
        P2_U3560) );
  MUX2_X1 U15566 ( .A(n14166), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14186), .Z(
        P2_U3559) );
  MUX2_X1 U15567 ( .A(n14167), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14186), .Z(
        P2_U3558) );
  MUX2_X1 U15568 ( .A(n14168), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14186), .Z(
        P2_U3557) );
  MUX2_X1 U15569 ( .A(n14169), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14186), .Z(
        P2_U3556) );
  MUX2_X1 U15570 ( .A(n14170), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14186), .Z(
        P2_U3555) );
  MUX2_X1 U15571 ( .A(n14171), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14186), .Z(
        P2_U3554) );
  MUX2_X1 U15572 ( .A(n14172), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14186), .Z(
        P2_U3553) );
  MUX2_X1 U15573 ( .A(n14173), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14186), .Z(
        P2_U3552) );
  MUX2_X1 U15574 ( .A(n14174), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14186), .Z(
        P2_U3551) );
  MUX2_X1 U15575 ( .A(n14175), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14186), .Z(
        P2_U3550) );
  MUX2_X1 U15576 ( .A(n14176), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14186), .Z(
        P2_U3549) );
  MUX2_X1 U15577 ( .A(n14177), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14186), .Z(
        P2_U3548) );
  MUX2_X1 U15578 ( .A(n14178), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14186), .Z(
        P2_U3547) );
  MUX2_X1 U15579 ( .A(n14179), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14186), .Z(
        P2_U3546) );
  MUX2_X1 U15580 ( .A(n14180), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14186), .Z(
        P2_U3545) );
  MUX2_X1 U15581 ( .A(n14181), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14186), .Z(
        P2_U3544) );
  MUX2_X1 U15582 ( .A(n14182), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14186), .Z(
        P2_U3543) );
  MUX2_X1 U15583 ( .A(n14183), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14186), .Z(
        P2_U3542) );
  MUX2_X1 U15584 ( .A(n14184), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14186), .Z(
        P2_U3541) );
  MUX2_X1 U15585 ( .A(n14185), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14186), .Z(
        P2_U3540) );
  MUX2_X1 U15586 ( .A(n14187), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14186), .Z(
        P2_U3539) );
  MUX2_X1 U15587 ( .A(n14188), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14186), .Z(
        P2_U3538) );
  MUX2_X1 U15588 ( .A(n14189), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14186), .Z(
        P2_U3537) );
  MUX2_X1 U15589 ( .A(n14190), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14186), .Z(
        P2_U3536) );
  MUX2_X1 U15590 ( .A(n14191), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14186), .Z(
        P2_U3535) );
  MUX2_X1 U15591 ( .A(n14192), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14186), .Z(
        P2_U3534) );
  MUX2_X1 U15592 ( .A(n14193), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14186), .Z(
        P2_U3533) );
  MUX2_X1 U15593 ( .A(n10348), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14186), .Z(
        P2_U3532) );
  MUX2_X1 U15594 ( .A(n14194), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14186), .Z(
        P2_U3531) );
  AOI211_X1 U15595 ( .C1(n14197), .C2(n14196), .A(n14195), .B(n15368), .ZN(
        n14198) );
  INV_X1 U15596 ( .A(n14198), .ZN(n14206) );
  AOI22_X1 U15597 ( .A1(n15271), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14205) );
  NAND2_X1 U15598 ( .A1(n15374), .A2(n14199), .ZN(n14204) );
  OAI211_X1 U15599 ( .C1(n14202), .C2(n14201), .A(n15333), .B(n14200), .ZN(
        n14203) );
  NAND4_X1 U15600 ( .A1(n14206), .A2(n14205), .A3(n14204), .A4(n14203), .ZN(
        P2_U3216) );
  NOR2_X1 U15601 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14207), .ZN(n14209) );
  INV_X1 U15602 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15448) );
  NOR2_X1 U15603 ( .A1(n15377), .A2(n15448), .ZN(n14208) );
  AOI211_X1 U15604 ( .C1(n15374), .C2(n14210), .A(n14209), .B(n14208), .ZN(
        n14220) );
  AOI211_X1 U15605 ( .C1(n14213), .C2(n14212), .A(n14211), .B(n15368), .ZN(
        n14214) );
  INV_X1 U15606 ( .A(n14214), .ZN(n14219) );
  OAI211_X1 U15607 ( .C1(n14217), .C2(n14216), .A(n15333), .B(n14215), .ZN(
        n14218) );
  NAND3_X1 U15608 ( .A1(n14220), .A2(n14219), .A3(n14218), .ZN(P2_U3217) );
  AOI211_X1 U15609 ( .C1(n14222), .C2(n14221), .A(n15368), .B(n7239), .ZN(
        n14223) );
  INV_X1 U15610 ( .A(n14223), .ZN(n14232) );
  AND2_X1 U15611 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14225) );
  INV_X1 U15612 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15491) );
  NOR2_X1 U15613 ( .A1(n15377), .A2(n15491), .ZN(n14224) );
  AOI211_X1 U15614 ( .C1(n15374), .C2(n14226), .A(n14225), .B(n14224), .ZN(
        n14231) );
  OAI211_X1 U15615 ( .C1(n14229), .C2(n14228), .A(n15333), .B(n14227), .ZN(
        n14230) );
  NAND3_X1 U15616 ( .A1(n14232), .A2(n14231), .A3(n14230), .ZN(P2_U3221) );
  AOI211_X1 U15617 ( .C1(n14235), .C2(n14234), .A(n15368), .B(n14233), .ZN(
        n14236) );
  INV_X1 U15618 ( .A(n14236), .ZN(n14245) );
  OAI21_X1 U15619 ( .B1(n15322), .B2(n14238), .A(n14237), .ZN(n14239) );
  AOI21_X1 U15620 ( .B1(n15271), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n14239), .ZN(
        n14244) );
  OAI211_X1 U15621 ( .C1(n14242), .C2(n14241), .A(n15333), .B(n14240), .ZN(
        n14243) );
  NAND3_X1 U15622 ( .A1(n14245), .A2(n14244), .A3(n14243), .ZN(P2_U3222) );
  NAND2_X1 U15623 ( .A1(n14246), .A2(n7209), .ZN(n14435) );
  NAND2_X1 U15624 ( .A1(n14248), .A2(n14247), .ZN(n14438) );
  NOR2_X1 U15625 ( .A1(n15947), .A2(n14438), .ZN(n14256) );
  NOR2_X1 U15626 ( .A1(n7653), .A2(n15940), .ZN(n14249) );
  AOI211_X1 U15627 ( .C1(n15947), .C2(P2_REG2_REG_31__SCAN_IN), .A(n14256), 
        .B(n14249), .ZN(n14250) );
  OAI21_X1 U15628 ( .B1(n15717), .B2(n14435), .A(n14250), .ZN(P2_U3234) );
  NAND2_X1 U15629 ( .A1(n14524), .A2(n14251), .ZN(n14252) );
  NAND2_X1 U15630 ( .A1(n14252), .A2(n7209), .ZN(n14253) );
  NOR2_X1 U15631 ( .A1(n15721), .A2(n14255), .ZN(n14257) );
  AOI211_X1 U15632 ( .C1(n14524), .C2(n15917), .A(n14257), .B(n14256), .ZN(
        n14258) );
  OAI21_X1 U15633 ( .B1(n14439), .B2(n15717), .A(n14258), .ZN(P2_U3235) );
  INV_X1 U15634 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n14259) );
  OAI22_X1 U15635 ( .A1(n14260), .A2(n15714), .B1(n14259), .B2(n15721), .ZN(
        n14261) );
  AOI21_X1 U15636 ( .B1(n14262), .B2(n15917), .A(n14261), .ZN(n14263) );
  OAI21_X1 U15637 ( .B1(n14264), .B2(n15717), .A(n14263), .ZN(n14265) );
  AOI21_X1 U15638 ( .B1(n14266), .B2(n15807), .A(n14265), .ZN(n14267) );
  OAI21_X1 U15639 ( .B1(n14268), .B2(n15947), .A(n14267), .ZN(P2_U3236) );
  AOI21_X1 U15640 ( .B1(n14269), .B2(n14274), .A(n15702), .ZN(n14272) );
  INV_X1 U15641 ( .A(n14295), .ZN(n14278) );
  INV_X1 U15642 ( .A(n14276), .ZN(n14277) );
  AOI211_X1 U15643 ( .C1(n14444), .C2(n14278), .A(n14360), .B(n14277), .ZN(
        n14443) );
  NAND2_X1 U15644 ( .A1(n14443), .A2(n15934), .ZN(n14282) );
  INV_X1 U15645 ( .A(n14279), .ZN(n14280) );
  AOI22_X1 U15646 ( .A1(n14280), .A2(n15936), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n15947), .ZN(n14281) );
  OAI211_X1 U15647 ( .C1(n14283), .C2(n15940), .A(n14282), .B(n14281), .ZN(
        n14284) );
  AOI21_X1 U15648 ( .B1(n14442), .B2(n15807), .A(n14284), .ZN(n14285) );
  OAI21_X1 U15649 ( .B1(n15947), .B2(n14446), .A(n14285), .ZN(P2_U3237) );
  XNOR2_X1 U15650 ( .A(n14286), .B(n14289), .ZN(n14288) );
  AOI21_X1 U15651 ( .B1(n14288), .B2(n15797), .A(n14287), .ZN(n14452) );
  NAND2_X1 U15652 ( .A1(n14290), .A2(n14289), .ZN(n14291) );
  NAND2_X1 U15653 ( .A1(n14292), .A2(n14291), .ZN(n14453) );
  INV_X1 U15654 ( .A(n14453), .ZN(n14300) );
  NAND2_X1 U15655 ( .A1(n14309), .A2(n14448), .ZN(n14293) );
  NAND2_X1 U15656 ( .A1(n14293), .A2(n7209), .ZN(n14294) );
  OR2_X1 U15657 ( .A1(n14295), .A2(n14294), .ZN(n14450) );
  AOI22_X1 U15658 ( .A1(n14296), .A2(n15936), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15947), .ZN(n14298) );
  NAND2_X1 U15659 ( .A1(n14448), .A2(n15917), .ZN(n14297) );
  OAI211_X1 U15660 ( .C1(n14450), .C2(n15717), .A(n14298), .B(n14297), .ZN(
        n14299) );
  AOI21_X1 U15661 ( .B1(n14300), .B2(n15807), .A(n14299), .ZN(n14301) );
  OAI21_X1 U15662 ( .B1(n15947), .B2(n14452), .A(n14301), .ZN(P2_U3238) );
  XNOR2_X1 U15663 ( .A(n14302), .B(n14303), .ZN(n14305) );
  OAI21_X1 U15664 ( .B1(n14305), .B2(n15702), .A(n14304), .ZN(n14454) );
  INV_X1 U15665 ( .A(n14454), .ZN(n14316) );
  XNOR2_X1 U15666 ( .A(n14307), .B(n14306), .ZN(n14456) );
  OR2_X1 U15667 ( .A1(n14322), .A2(n14531), .ZN(n14310) );
  AND3_X1 U15668 ( .A1(n14310), .A2(n14309), .A3(n14308), .ZN(n14455) );
  NAND2_X1 U15669 ( .A1(n14455), .A2(n15934), .ZN(n14313) );
  AOI22_X1 U15670 ( .A1(n14311), .A2(n15936), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15947), .ZN(n14312) );
  OAI211_X1 U15671 ( .C1(n14531), .C2(n15940), .A(n14313), .B(n14312), .ZN(
        n14314) );
  AOI21_X1 U15672 ( .B1(n14456), .B2(n15807), .A(n14314), .ZN(n14315) );
  OAI21_X1 U15673 ( .B1(n14316), .B2(n15947), .A(n14315), .ZN(P2_U3239) );
  XNOR2_X1 U15674 ( .A(n14317), .B(n14320), .ZN(n14319) );
  OAI21_X1 U15675 ( .B1(n14319), .B2(n15702), .A(n14318), .ZN(n14459) );
  INV_X1 U15676 ( .A(n14459), .ZN(n14329) );
  XNOR2_X1 U15677 ( .A(n14321), .B(n14320), .ZN(n14461) );
  AOI211_X1 U15678 ( .C1(n14323), .C2(n7639), .A(n14360), .B(n14322), .ZN(
        n14460) );
  NAND2_X1 U15679 ( .A1(n14460), .A2(n15934), .ZN(n14326) );
  AOI22_X1 U15680 ( .A1(n14324), .A2(n15936), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n15947), .ZN(n14325) );
  OAI211_X1 U15681 ( .C1(n14535), .C2(n15940), .A(n14326), .B(n14325), .ZN(
        n14327) );
  AOI21_X1 U15682 ( .B1(n15807), .B2(n14461), .A(n14327), .ZN(n14328) );
  OAI21_X1 U15683 ( .B1(n15947), .B2(n14329), .A(n14328), .ZN(P2_U3240) );
  XNOR2_X1 U15684 ( .A(n14330), .B(n14332), .ZN(n14468) );
  AOI21_X1 U15685 ( .B1(n14332), .B2(n14331), .A(n7271), .ZN(n14334) );
  OAI21_X1 U15686 ( .B1(n14334), .B2(n15702), .A(n14333), .ZN(n14464) );
  NAND2_X1 U15687 ( .A1(n7240), .A2(n14466), .ZN(n14335) );
  NAND2_X1 U15688 ( .A1(n14335), .A2(n7209), .ZN(n14336) );
  NOR2_X1 U15689 ( .A1(n7635), .A2(n14336), .ZN(n14465) );
  NAND2_X1 U15690 ( .A1(n14465), .A2(n15934), .ZN(n14339) );
  AOI22_X1 U15691 ( .A1(n14337), .A2(n15936), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n15947), .ZN(n14338) );
  OAI211_X1 U15692 ( .C1(n7638), .C2(n15940), .A(n14339), .B(n14338), .ZN(
        n14340) );
  AOI21_X1 U15693 ( .B1(n14464), .B2(n15721), .A(n14340), .ZN(n14341) );
  OAI21_X1 U15694 ( .B1(n14369), .B2(n14468), .A(n14341), .ZN(P2_U3241) );
  INV_X1 U15695 ( .A(n14346), .ZN(n14342) );
  XNOR2_X1 U15696 ( .A(n14343), .B(n14342), .ZN(n14345) );
  AOI21_X1 U15697 ( .B1(n14345), .B2(n15797), .A(n14344), .ZN(n14475) );
  XNOR2_X1 U15698 ( .A(n14347), .B(n14346), .ZN(n14473) );
  AOI21_X1 U15699 ( .B1(n14361), .B2(n14469), .A(n14360), .ZN(n14348) );
  NAND2_X1 U15700 ( .A1(n14348), .A2(n7240), .ZN(n14471) );
  INV_X1 U15701 ( .A(n14349), .ZN(n14350) );
  AOI22_X1 U15702 ( .A1(n14350), .A2(n15936), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n15947), .ZN(n14352) );
  NAND2_X1 U15703 ( .A1(n14469), .A2(n15917), .ZN(n14351) );
  OAI211_X1 U15704 ( .C1(n14471), .C2(n15717), .A(n14352), .B(n14351), .ZN(
        n14353) );
  AOI21_X1 U15705 ( .B1(n14473), .B2(n15807), .A(n14353), .ZN(n14354) );
  OAI21_X1 U15706 ( .B1(n14475), .B2(n15947), .A(n14354), .ZN(P2_U3242) );
  XNOR2_X1 U15707 ( .A(n7252), .B(n14357), .ZN(n14478) );
  OAI211_X1 U15708 ( .C1(n14357), .C2(n14356), .A(n14355), .B(n15797), .ZN(
        n14359) );
  AND2_X1 U15709 ( .A1(n14359), .A2(n14358), .ZN(n14477) );
  INV_X1 U15710 ( .A(n14477), .ZN(n14367) );
  AOI21_X1 U15711 ( .B1(n14540), .B2(n14372), .A(n14360), .ZN(n14362) );
  NAND2_X1 U15712 ( .A1(n14362), .A2(n14361), .ZN(n14476) );
  AOI22_X1 U15713 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(n15947), .B1(n14363), 
        .B2(n15936), .ZN(n14365) );
  NAND2_X1 U15714 ( .A1(n14540), .A2(n15917), .ZN(n14364) );
  OAI211_X1 U15715 ( .C1(n14476), .C2(n15717), .A(n14365), .B(n14364), .ZN(
        n14366) );
  AOI21_X1 U15716 ( .B1(n14367), .B2(n15721), .A(n14366), .ZN(n14368) );
  OAI21_X1 U15717 ( .B1(n14478), .B2(n14369), .A(n14368), .ZN(P2_U3243) );
  XNOR2_X1 U15718 ( .A(n14371), .B(n14370), .ZN(n14481) );
  OAI211_X1 U15719 ( .C1(n14545), .C2(n14391), .A(n7209), .B(n14372), .ZN(
        n14482) );
  INV_X1 U15720 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n14374) );
  OAI22_X1 U15721 ( .A1(n15721), .A2(n14374), .B1(n14373), .B2(n15714), .ZN(
        n14375) );
  AOI21_X1 U15722 ( .B1(n14376), .B2(n15917), .A(n14375), .ZN(n14377) );
  OAI21_X1 U15723 ( .B1(n14482), .B2(n15717), .A(n14377), .ZN(n14384) );
  OAI211_X1 U15724 ( .C1(n14380), .C2(n14379), .A(n14378), .B(n15797), .ZN(
        n14382) );
  AND2_X1 U15725 ( .A1(n14382), .A2(n14381), .ZN(n14483) );
  NOR2_X1 U15726 ( .A1(n14483), .A2(n15947), .ZN(n14383) );
  AOI211_X1 U15727 ( .C1(n15807), .C2(n14481), .A(n14384), .B(n14383), .ZN(
        n14385) );
  INV_X1 U15728 ( .A(n14385), .ZN(P2_U3244) );
  XNOR2_X1 U15729 ( .A(n14389), .B(n14386), .ZN(n14388) );
  OAI21_X1 U15730 ( .B1(n14388), .B2(n15702), .A(n14387), .ZN(n14487) );
  INV_X1 U15731 ( .A(n14487), .ZN(n14398) );
  XOR2_X1 U15732 ( .A(n7397), .B(n14389), .Z(n14489) );
  AOI211_X1 U15733 ( .C1(n14392), .C2(n14403), .A(n14360), .B(n14391), .ZN(
        n14488) );
  NAND2_X1 U15734 ( .A1(n14488), .A2(n15934), .ZN(n14395) );
  AOI22_X1 U15735 ( .A1(n15947), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14393), 
        .B2(n15936), .ZN(n14394) );
  OAI211_X1 U15736 ( .C1(n14549), .C2(n15940), .A(n14395), .B(n14394), .ZN(
        n14396) );
  AOI21_X1 U15737 ( .B1(n15807), .B2(n14489), .A(n14396), .ZN(n14397) );
  OAI21_X1 U15738 ( .B1(n15947), .B2(n14398), .A(n14397), .ZN(P2_U3245) );
  INV_X1 U15739 ( .A(n14411), .ZN(n14400) );
  NAND2_X1 U15740 ( .A1(n14400), .A2(n14399), .ZN(n14401) );
  NAND2_X1 U15741 ( .A1(n14402), .A2(n14401), .ZN(n14492) );
  INV_X1 U15742 ( .A(n14403), .ZN(n14404) );
  AOI211_X1 U15743 ( .C1(n14405), .C2(n14427), .A(n14360), .B(n14404), .ZN(
        n14494) );
  NOR2_X1 U15744 ( .A1(n7640), .A2(n15940), .ZN(n14409) );
  OAI22_X1 U15745 ( .A1(n15721), .A2(n14407), .B1(n14406), .B2(n15714), .ZN(
        n14408) );
  AOI211_X1 U15746 ( .C1(n14494), .C2(n15934), .A(n14409), .B(n14408), .ZN(
        n14416) );
  XNOR2_X1 U15747 ( .A(n14411), .B(n14410), .ZN(n14412) );
  NAND2_X1 U15748 ( .A1(n14412), .A2(n15797), .ZN(n14413) );
  OAI211_X1 U15749 ( .C1(n14492), .C2(n14423), .A(n14414), .B(n14413), .ZN(
        n14493) );
  NAND2_X1 U15750 ( .A1(n14493), .A2(n15721), .ZN(n14415) );
  OAI211_X1 U15751 ( .C1(n14492), .C2(n14431), .A(n14416), .B(n14415), .ZN(
        P2_U3246) );
  XNOR2_X1 U15752 ( .A(n14417), .B(n14420), .ZN(n14425) );
  INV_X1 U15753 ( .A(n14418), .ZN(n14419) );
  AOI21_X1 U15754 ( .B1(n14421), .B2(n14420), .A(n14419), .ZN(n14503) );
  OAI21_X1 U15755 ( .B1(n14503), .B2(n14423), .A(n14422), .ZN(n14424) );
  AOI21_X1 U15756 ( .B1(n14425), .B2(n15797), .A(n14424), .ZN(n14502) );
  INV_X1 U15757 ( .A(n14427), .ZN(n14428) );
  AOI211_X1 U15758 ( .C1(n14500), .C2(n7644), .A(n14360), .B(n14428), .ZN(
        n14499) );
  AOI22_X1 U15759 ( .A1(n15947), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14429), 
        .B2(n15936), .ZN(n14430) );
  OAI21_X1 U15760 ( .B1(n7838), .B2(n15940), .A(n14430), .ZN(n14433) );
  NOR2_X1 U15761 ( .A1(n14503), .A2(n14431), .ZN(n14432) );
  AOI211_X1 U15762 ( .C1(n14499), .C2(n15934), .A(n14433), .B(n14432), .ZN(
        n14434) );
  OAI21_X1 U15763 ( .B1(n15947), .B2(n14502), .A(n14434), .ZN(P2_U3247) );
  AND2_X1 U15764 ( .A1(n14435), .A2(n14438), .ZN(n14519) );
  MUX2_X1 U15765 ( .A(n14436), .B(n14519), .S(n15970), .Z(n14437) );
  OAI21_X1 U15766 ( .B1(n7653), .B2(n14498), .A(n14437), .ZN(P2_U3530) );
  NAND2_X1 U15767 ( .A1(n14439), .A2(n14438), .ZN(n14522) );
  MUX2_X1 U15768 ( .A(n14522), .B(P2_REG1_REG_30__SCAN_IN), .S(n15968), .Z(
        n14440) );
  AOI21_X1 U15769 ( .B1(n14510), .B2(n14524), .A(n14440), .ZN(n14441) );
  INV_X1 U15770 ( .A(n14441), .ZN(P2_U3529) );
  INV_X1 U15771 ( .A(n14442), .ZN(n14447) );
  AOI21_X1 U15772 ( .B1(n15959), .B2(n14444), .A(n14443), .ZN(n14445) );
  OAI211_X1 U15773 ( .C1(n14447), .C2(n15834), .A(n14446), .B(n14445), .ZN(
        n14526) );
  MUX2_X1 U15774 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14526), .S(n15970), .Z(
        P2_U3527) );
  NAND2_X1 U15775 ( .A1(n14448), .A2(n15959), .ZN(n14449) );
  AND2_X1 U15776 ( .A1(n14450), .A2(n14449), .ZN(n14451) );
  OAI211_X1 U15777 ( .C1(n15834), .C2(n14453), .A(n14452), .B(n14451), .ZN(
        n14527) );
  MUX2_X1 U15778 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14527), .S(n15970), .Z(
        P2_U3526) );
  AOI211_X1 U15779 ( .C1(n15964), .C2(n14456), .A(n14455), .B(n14454), .ZN(
        n14528) );
  MUX2_X1 U15780 ( .A(n14457), .B(n14528), .S(n15970), .Z(n14458) );
  OAI21_X1 U15781 ( .B1(n14531), .B2(n14498), .A(n14458), .ZN(P2_U3525) );
  AOI211_X1 U15782 ( .C1(n14461), .C2(n15964), .A(n14460), .B(n14459), .ZN(
        n14532) );
  MUX2_X1 U15783 ( .A(n14462), .B(n14532), .S(n15970), .Z(n14463) );
  OAI21_X1 U15784 ( .B1(n14535), .B2(n14498), .A(n14463), .ZN(P2_U3524) );
  AOI211_X1 U15785 ( .C1(n15959), .C2(n14466), .A(n14465), .B(n14464), .ZN(
        n14467) );
  OAI21_X1 U15786 ( .B1(n15834), .B2(n14468), .A(n14467), .ZN(n14536) );
  MUX2_X1 U15787 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14536), .S(n15970), .Z(
        P2_U3523) );
  NAND2_X1 U15788 ( .A1(n14469), .A2(n15959), .ZN(n14470) );
  NAND2_X1 U15789 ( .A1(n14471), .A2(n14470), .ZN(n14472) );
  AOI21_X1 U15790 ( .B1(n14473), .B2(n15964), .A(n14472), .ZN(n14474) );
  NAND2_X1 U15791 ( .A1(n14475), .A2(n14474), .ZN(n14537) );
  MUX2_X1 U15792 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14537), .S(n15970), .Z(
        P2_U3522) );
  OAI211_X1 U15793 ( .C1(n14478), .C2(n15834), .A(n14477), .B(n14476), .ZN(
        n14538) );
  MUX2_X1 U15794 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14538), .S(n15970), .Z(
        n14479) );
  AOI21_X1 U15795 ( .B1(n14510), .B2(n14540), .A(n14479), .ZN(n14480) );
  INV_X1 U15796 ( .A(n14480), .ZN(P2_U3521) );
  NAND2_X1 U15797 ( .A1(n14481), .A2(n15964), .ZN(n14484) );
  MUX2_X1 U15798 ( .A(n14543), .B(n14485), .S(n15968), .Z(n14486) );
  OAI21_X1 U15799 ( .B1(n14545), .B2(n14498), .A(n14486), .ZN(P2_U3520) );
  AOI211_X1 U15800 ( .C1(n15964), .C2(n14489), .A(n14488), .B(n14487), .ZN(
        n14546) );
  MUX2_X1 U15801 ( .A(n14490), .B(n14546), .S(n15970), .Z(n14491) );
  OAI21_X1 U15802 ( .B1(n14549), .B2(n14498), .A(n14491), .ZN(P2_U3519) );
  INV_X1 U15803 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14496) );
  INV_X1 U15804 ( .A(n14492), .ZN(n14495) );
  AOI211_X1 U15805 ( .C1(n14495), .C2(n15758), .A(n14494), .B(n14493), .ZN(
        n14550) );
  MUX2_X1 U15806 ( .A(n14496), .B(n14550), .S(n15970), .Z(n14497) );
  OAI21_X1 U15807 ( .B1(n7640), .B2(n14498), .A(n14497), .ZN(P2_U3518) );
  AOI21_X1 U15808 ( .B1(n15959), .B2(n14500), .A(n14499), .ZN(n14501) );
  OAI211_X1 U15809 ( .C1(n14503), .C2(n9421), .A(n14502), .B(n14501), .ZN(
        n14554) );
  MUX2_X1 U15810 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14554), .S(n15970), .Z(
        P2_U3517) );
  NOR2_X1 U15811 ( .A1(n14505), .A2(n14504), .ZN(n14508) );
  NAND2_X1 U15812 ( .A1(n14506), .A2(n15964), .ZN(n14507) );
  NAND2_X1 U15813 ( .A1(n14508), .A2(n14507), .ZN(n14555) );
  MUX2_X1 U15814 ( .A(n14555), .B(P2_REG1_REG_17__SCAN_IN), .S(n15968), .Z(
        n14509) );
  AOI21_X1 U15815 ( .B1(n14510), .B2(n14557), .A(n14509), .ZN(n14511) );
  INV_X1 U15816 ( .A(n14511), .ZN(P2_U3516) );
  NAND2_X1 U15817 ( .A1(n14512), .A2(n15959), .ZN(n14514) );
  OAI211_X1 U15818 ( .C1(n14515), .C2(n9421), .A(n14514), .B(n14513), .ZN(
        n14516) );
  OR2_X1 U15819 ( .A1(n14517), .A2(n14516), .ZN(n14560) );
  MUX2_X1 U15820 ( .A(n14560), .B(P2_REG1_REG_16__SCAN_IN), .S(n15968), .Z(
        P2_U3515) );
  MUX2_X1 U15821 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14518), .S(n15970), .Z(
        P2_U3510) );
  INV_X1 U15822 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14520) );
  MUX2_X1 U15823 ( .A(n14520), .B(n14519), .S(n15973), .Z(n14521) );
  OAI21_X1 U15824 ( .B1(n7653), .B2(n14553), .A(n14521), .ZN(P2_U3498) );
  MUX2_X1 U15825 ( .A(n14522), .B(P2_REG0_REG_30__SCAN_IN), .S(n15971), .Z(
        n14523) );
  AOI21_X1 U15826 ( .B1(n14558), .B2(n14524), .A(n14523), .ZN(n14525) );
  INV_X1 U15827 ( .A(n14525), .ZN(P2_U3497) );
  MUX2_X1 U15828 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14526), .S(n15973), .Z(
        P2_U3495) );
  MUX2_X1 U15829 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14527), .S(n15973), .Z(
        P2_U3494) );
  INV_X1 U15830 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14529) );
  MUX2_X1 U15831 ( .A(n14529), .B(n14528), .S(n15973), .Z(n14530) );
  OAI21_X1 U15832 ( .B1(n14531), .B2(n14553), .A(n14530), .ZN(P2_U3493) );
  INV_X1 U15833 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14533) );
  MUX2_X1 U15834 ( .A(n14533), .B(n14532), .S(n15973), .Z(n14534) );
  OAI21_X1 U15835 ( .B1(n14535), .B2(n14553), .A(n14534), .ZN(P2_U3492) );
  MUX2_X1 U15836 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14536), .S(n15973), .Z(
        P2_U3491) );
  MUX2_X1 U15837 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14537), .S(n15973), .Z(
        P2_U3490) );
  MUX2_X1 U15838 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14538), .S(n15973), .Z(
        n14539) );
  AOI21_X1 U15839 ( .B1(n14558), .B2(n14540), .A(n14539), .ZN(n14541) );
  INV_X1 U15840 ( .A(n14541), .ZN(P2_U3489) );
  INV_X1 U15841 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14542) );
  MUX2_X1 U15842 ( .A(n14543), .B(n14542), .S(n15971), .Z(n14544) );
  OAI21_X1 U15843 ( .B1(n14545), .B2(n14553), .A(n14544), .ZN(P2_U3488) );
  INV_X1 U15844 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n14547) );
  MUX2_X1 U15845 ( .A(n14547), .B(n14546), .S(n15973), .Z(n14548) );
  OAI21_X1 U15846 ( .B1(n14549), .B2(n14553), .A(n14548), .ZN(P2_U3487) );
  INV_X1 U15847 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14551) );
  MUX2_X1 U15848 ( .A(n14551), .B(n14550), .S(n15973), .Z(n14552) );
  OAI21_X1 U15849 ( .B1(n7640), .B2(n14553), .A(n14552), .ZN(P2_U3486) );
  MUX2_X1 U15850 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14554), .S(n15973), .Z(
        P2_U3484) );
  MUX2_X1 U15851 ( .A(n14555), .B(P2_REG0_REG_17__SCAN_IN), .S(n15971), .Z(
        n14556) );
  AOI21_X1 U15852 ( .B1(n14558), .B2(n14557), .A(n14556), .ZN(n14559) );
  INV_X1 U15853 ( .A(n14559), .ZN(P2_U3481) );
  MUX2_X1 U15854 ( .A(n14560), .B(P2_REG0_REG_16__SCAN_IN), .S(n15971), .Z(
        P2_U3478) );
  INV_X1 U15855 ( .A(n14561), .ZN(n15214) );
  INV_X1 U15856 ( .A(n14562), .ZN(n14564) );
  NOR4_X1 U15857 ( .A1(n14564), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14563), .A4(
        P2_U3088), .ZN(n14565) );
  AOI21_X1 U15858 ( .B1(n14576), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14565), 
        .ZN(n14566) );
  OAI21_X1 U15859 ( .B1(n15214), .B2(n14578), .A(n14566), .ZN(P2_U3296) );
  INV_X1 U15860 ( .A(n14567), .ZN(n15216) );
  INV_X1 U15861 ( .A(n14568), .ZN(n14570) );
  INV_X1 U15862 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14569) );
  OAI222_X1 U15863 ( .A1(n14578), .A2(n15216), .B1(P2_U3088), .B2(n14570), 
        .C1(n14569), .C2(n14592), .ZN(P2_U3297) );
  INV_X1 U15864 ( .A(n14571), .ZN(n15219) );
  INV_X1 U15865 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14572) );
  OAI222_X1 U15866 ( .A1(P2_U3088), .A2(n14573), .B1(n14578), .B2(n15219), 
        .C1(n14572), .C2(n14592), .ZN(P2_U3298) );
  INV_X1 U15867 ( .A(n14574), .ZN(n15222) );
  AOI21_X1 U15868 ( .B1(n14576), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14575), 
        .ZN(n14577) );
  OAI21_X1 U15869 ( .B1(n15222), .B2(n14578), .A(n14577), .ZN(P2_U3299) );
  INV_X1 U15870 ( .A(n14579), .ZN(n15226) );
  OAI222_X1 U15871 ( .A1(n14592), .A2(n14581), .B1(n14578), .B2(n15226), .C1(
        n14580), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15872 ( .A(n14582), .ZN(n15229) );
  OAI222_X1 U15873 ( .A1(P2_U3088), .A2(n14584), .B1(n14578), .B2(n15229), 
        .C1(n14583), .C2(n14592), .ZN(P2_U3301) );
  OAI222_X1 U15874 ( .A1(n14592), .A2(n14588), .B1(n14578), .B2(n14587), .C1(
        P2_U3088), .C2(n14586), .ZN(P2_U3302) );
  INV_X1 U15875 ( .A(n14589), .ZN(n15232) );
  OAI222_X1 U15876 ( .A1(n14592), .A2(n14591), .B1(n14578), .B2(n15232), .C1(
        P2_U3088), .C2(n14590), .ZN(P2_U3303) );
  INV_X1 U15877 ( .A(n14593), .ZN(n14594) );
  MUX2_X1 U15878 ( .A(n14594), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NOR2_X1 U15879 ( .A1(n16031), .A2(n14889), .ZN(n14598) );
  AOI22_X1 U15880 ( .A1(n15978), .A2(n14727), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14596) );
  OAI21_X1 U15881 ( .B1(n14888), .B2(n16016), .A(n14596), .ZN(n14597) );
  AOI211_X1 U15882 ( .C1(n15114), .C2(n16027), .A(n14598), .B(n14597), .ZN(
        n14599) );
  OAI21_X1 U15883 ( .B1(n14600), .B2(n16022), .A(n14599), .ZN(P1_U3214) );
  INV_X1 U15884 ( .A(n14601), .ZN(n14602) );
  AOI21_X1 U15885 ( .B1(n14604), .B2(n14603), .A(n14602), .ZN(n14612) );
  OAI21_X1 U15886 ( .B1(n16019), .B2(n14606), .A(n14605), .ZN(n14607) );
  AOI21_X1 U15887 ( .B1(n15980), .B2(n14734), .A(n14607), .ZN(n14608) );
  OAI21_X1 U15888 ( .B1(n14609), .B2(n16031), .A(n14608), .ZN(n14610) );
  AOI21_X1 U15889 ( .B1(n15950), .B2(n16027), .A(n14610), .ZN(n14611) );
  OAI21_X1 U15890 ( .B1(n14612), .B2(n16022), .A(n14611), .ZN(P1_U3215) );
  OAI21_X1 U15891 ( .B1(n14614), .B2(n14613), .A(n14664), .ZN(n14615) );
  NAND2_X1 U15892 ( .A1(n14615), .A2(n16010), .ZN(n14619) );
  OAI22_X1 U15893 ( .A1(n7794), .A2(n15042), .B1(n14972), .B2(n15041), .ZN(
        n15140) );
  OAI22_X1 U15894 ( .A1(n14945), .A2(n16031), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14616), .ZN(n14617) );
  AOI21_X1 U15895 ( .B1(n15140), .B2(n16011), .A(n14617), .ZN(n14618) );
  OAI211_X1 U15896 ( .C1(n14949), .C2(n15982), .A(n14619), .B(n14618), .ZN(
        P1_U3216) );
  OAI211_X1 U15897 ( .C1(n14620), .C2(n14622), .A(n14621), .B(n16010), .ZN(
        n14628) );
  AOI22_X1 U15898 ( .A1(n15978), .A2(n14741), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14627) );
  INV_X1 U15899 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14623) );
  AOI22_X1 U15900 ( .A1(n16027), .A2(n14624), .B1(n14721), .B2(n14623), .ZN(
        n14626) );
  NAND2_X1 U15901 ( .A1(n15980), .A2(n14743), .ZN(n14625) );
  NAND4_X1 U15902 ( .A1(n14628), .A2(n14627), .A3(n14626), .A4(n14625), .ZN(
        P1_U3218) );
  XOR2_X1 U15903 ( .A(n14630), .B(n14629), .Z(n14635) );
  NAND2_X1 U15904 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14820)
         );
  OAI21_X1 U15905 ( .B1(n16016), .B2(n16018), .A(n14820), .ZN(n14631) );
  AOI21_X1 U15906 ( .B1(n14733), .B2(n15978), .A(n14631), .ZN(n14632) );
  OAI21_X1 U15907 ( .B1(n15004), .B2(n16031), .A(n14632), .ZN(n14633) );
  AOI21_X1 U15908 ( .B1(n15170), .B2(n16027), .A(n14633), .ZN(n14634) );
  OAI21_X1 U15909 ( .B1(n14635), .B2(n16022), .A(n14634), .ZN(P1_U3219) );
  INV_X1 U15910 ( .A(n14636), .ZN(n14637) );
  AOI21_X1 U15911 ( .B1(n14639), .B2(n14638), .A(n14637), .ZN(n14644) );
  AOI22_X1 U15912 ( .A1(n14733), .A2(n15980), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14641) );
  NAND2_X1 U15913 ( .A1(n14721), .A2(n14971), .ZN(n14640) );
  OAI211_X1 U15914 ( .C1(n14972), .C2(n16019), .A(n14641), .B(n14640), .ZN(
        n14642) );
  AOI21_X1 U15915 ( .B1(n15154), .B2(n16027), .A(n14642), .ZN(n14643) );
  OAI21_X1 U15916 ( .B1(n14644), .B2(n16022), .A(n14643), .ZN(P1_U3223) );
  OAI211_X1 U15917 ( .C1(n7326), .C2(n14646), .A(n14645), .B(n16010), .ZN(
        n14653) );
  NOR2_X1 U15918 ( .A1(n16031), .A2(n14647), .ZN(n14651) );
  OAI21_X1 U15919 ( .B1(n16019), .B2(n14649), .A(n14648), .ZN(n14650) );
  AOI211_X1 U15920 ( .C1(n15980), .C2(n14736), .A(n14651), .B(n14650), .ZN(
        n14652) );
  OAI211_X1 U15921 ( .C1(n7584), .C2(n15982), .A(n14653), .B(n14652), .ZN(
        P1_U3224) );
  OAI21_X1 U15922 ( .B1(n14656), .B2(n14655), .A(n14654), .ZN(n14657) );
  NAND2_X1 U15923 ( .A1(n14657), .A2(n16010), .ZN(n14663) );
  NAND2_X1 U15924 ( .A1(n14731), .A2(n15075), .ZN(n14659) );
  OR2_X1 U15925 ( .A1(n14888), .A2(n15042), .ZN(n14658) );
  NAND2_X1 U15926 ( .A1(n14659), .A2(n14658), .ZN(n15125) );
  INV_X1 U15927 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14660) );
  OAI22_X1 U15928 ( .A1(n16031), .A2(n14916), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14660), .ZN(n14661) );
  AOI21_X1 U15929 ( .B1(n15125), .B2(n16011), .A(n14661), .ZN(n14662) );
  OAI211_X1 U15930 ( .C1(n15128), .C2(n15982), .A(n14663), .B(n14662), .ZN(
        P1_U3225) );
  INV_X1 U15931 ( .A(n14664), .ZN(n14667) );
  NOR3_X1 U15932 ( .A1(n14667), .A2(n14666), .A3(n14665), .ZN(n14670) );
  INV_X1 U15933 ( .A(n14668), .ZN(n14669) );
  OAI21_X1 U15934 ( .B1(n14670), .B2(n14669), .A(n16010), .ZN(n14675) );
  INV_X1 U15935 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14671) );
  OAI22_X1 U15936 ( .A1(n16019), .A2(n14926), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14671), .ZN(n14673) );
  NOR2_X1 U15937 ( .A1(n14927), .A2(n16016), .ZN(n14672) );
  AOI211_X1 U15938 ( .C1(n14721), .C2(n14933), .A(n14673), .B(n14672), .ZN(
        n14674) );
  OAI211_X1 U15939 ( .C1(n14936), .C2(n15982), .A(n14675), .B(n14674), .ZN(
        P1_U3229) );
  AOI21_X1 U15940 ( .B1(n14677), .B2(n14676), .A(n16022), .ZN(n14679) );
  NAND2_X1 U15941 ( .A1(n14679), .A2(n14678), .ZN(n14683) );
  AOI22_X1 U15942 ( .A1(n14984), .A2(n15978), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14680) );
  OAI21_X1 U15943 ( .B1(n8101), .B2(n16016), .A(n14680), .ZN(n14681) );
  AOI21_X1 U15944 ( .B1(n14985), .B2(n14721), .A(n14681), .ZN(n14682) );
  OAI211_X1 U15945 ( .C1(n15161), .C2(n15982), .A(n14683), .B(n14682), .ZN(
        P1_U3233) );
  OAI211_X1 U15946 ( .C1(n14686), .C2(n14685), .A(n14684), .B(n16010), .ZN(
        n14693) );
  INV_X1 U15947 ( .A(n14687), .ZN(n14691) );
  INV_X1 U15948 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n14688) );
  OAI22_X1 U15949 ( .A1(n14689), .A2(n15924), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14688), .ZN(n14690) );
  AOI21_X1 U15950 ( .B1(n14691), .B2(n14721), .A(n14690), .ZN(n14692) );
  OAI211_X1 U15951 ( .C1(n15926), .C2(n15982), .A(n14693), .B(n14692), .ZN(
        P1_U3234) );
  NAND2_X1 U15952 ( .A1(n14695), .A2(n14694), .ZN(n14696) );
  XNOR2_X1 U15953 ( .A(n14697), .B(n14696), .ZN(n14704) );
  OAI22_X1 U15954 ( .A1(n14699), .A2(n16016), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14698), .ZN(n14700) );
  AOI21_X1 U15955 ( .B1(n14960), .B2(n14721), .A(n14700), .ZN(n14701) );
  OAI21_X1 U15956 ( .B1(n14927), .B2(n16019), .A(n14701), .ZN(n14702) );
  AOI21_X1 U15957 ( .B1(n14959), .B2(n16027), .A(n14702), .ZN(n14703) );
  OAI21_X1 U15958 ( .B1(n14704), .B2(n16022), .A(n14703), .ZN(P1_U3235) );
  XOR2_X1 U15959 ( .A(n14706), .B(n14705), .Z(n14711) );
  NAND2_X1 U15960 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15405)
         );
  OAI21_X1 U15961 ( .B1(n16019), .B2(n8101), .A(n15405), .ZN(n14707) );
  AOI21_X1 U15962 ( .B1(n15980), .B2(n15057), .A(n14707), .ZN(n14708) );
  OAI21_X1 U15963 ( .B1(n15019), .B2(n16031), .A(n14708), .ZN(n14709) );
  AOI21_X1 U15964 ( .B1(n15175), .B2(n16027), .A(n14709), .ZN(n14710) );
  OAI21_X1 U15965 ( .B1(n14711), .B2(n16022), .A(n14710), .ZN(P1_U3238) );
  NOR2_X1 U15966 ( .A1(n14712), .A2(n7556), .ZN(n14717) );
  AOI21_X1 U15967 ( .B1(n14715), .B2(n14714), .A(n14713), .ZN(n14716) );
  OAI21_X1 U15968 ( .B1(n14717), .B2(n14716), .A(n16010), .ZN(n14723) );
  INV_X1 U15969 ( .A(n14718), .ZN(n14905) );
  AOI22_X1 U15970 ( .A1(n15978), .A2(n14728), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14719) );
  OAI21_X1 U15971 ( .B1(n14926), .B2(n16016), .A(n14719), .ZN(n14720) );
  AOI21_X1 U15972 ( .B1(n14905), .B2(n14721), .A(n14720), .ZN(n14722) );
  OAI211_X1 U15973 ( .C1(n14724), .C2(n15982), .A(n14723), .B(n14722), .ZN(
        P1_U3240) );
  MUX2_X1 U15974 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14855), .S(n14745), .Z(
        P1_U3591) );
  MUX2_X1 U15975 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14725), .S(n14745), .Z(
        P1_U3590) );
  MUX2_X1 U15976 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14726), .S(n14745), .Z(
        P1_U3589) );
  MUX2_X1 U15977 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14727), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15978 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14728), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15979 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14729), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15980 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14730), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15981 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14731), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15982 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14958), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15983 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14732), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15984 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14984), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15985 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14733), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15986 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15031), .S(n14745), .Z(
        P1_U3579) );
  MUX2_X1 U15987 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15001), .S(n14745), .Z(
        P1_U3578) );
  MUX2_X1 U15988 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15057), .S(n14745), .Z(
        P1_U3577) );
  MUX2_X1 U15989 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15977), .S(n14745), .Z(
        P1_U3576) );
  MUX2_X1 U15990 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15058), .S(n14745), .Z(
        P1_U3575) );
  MUX2_X1 U15991 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15979), .S(n14745), .Z(
        P1_U3574) );
  MUX2_X1 U15992 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14734), .S(n14745), .Z(
        P1_U3573) );
  MUX2_X1 U15993 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14735), .S(n14745), .Z(
        P1_U3572) );
  MUX2_X1 U15994 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14736), .S(n14745), .Z(
        P1_U3571) );
  MUX2_X1 U15995 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14737), .S(n14745), .Z(
        P1_U3569) );
  MUX2_X1 U15996 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14738), .S(n14745), .Z(
        P1_U3568) );
  MUX2_X1 U15997 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14739), .S(n14745), .Z(
        P1_U3567) );
  MUX2_X1 U15998 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14740), .S(n14745), .Z(
        P1_U3565) );
  MUX2_X1 U15999 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14741), .S(n14745), .Z(
        P1_U3564) );
  MUX2_X1 U16000 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14742), .S(n14745), .Z(
        P1_U3563) );
  MUX2_X1 U16001 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14743), .S(n14745), .Z(
        P1_U3562) );
  MUX2_X1 U16002 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14744), .S(n14745), .Z(
        P1_U3561) );
  MUX2_X1 U16003 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14746), .S(n14745), .Z(
        P1_U3560) );
  OAI211_X1 U16004 ( .C1(n14749), .C2(n14748), .A(n15426), .B(n14747), .ZN(
        n14757) );
  OAI211_X1 U16005 ( .C1(n14752), .C2(n14751), .A(n15427), .B(n14750), .ZN(
        n14756) );
  AOI22_X1 U16006 ( .A1(n15381), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14755) );
  NAND2_X1 U16007 ( .A1(n15423), .A2(n14753), .ZN(n14754) );
  NAND4_X1 U16008 ( .A1(n14757), .A2(n14756), .A3(n14755), .A4(n14754), .ZN(
        P1_U3244) );
  NAND2_X1 U16009 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n14758) );
  OAI21_X1 U16010 ( .B1(n15430), .B2(n15451), .A(n14758), .ZN(n14759) );
  AOI21_X1 U16011 ( .B1(n14760), .B2(n15423), .A(n14759), .ZN(n14769) );
  OAI211_X1 U16012 ( .C1(n14763), .C2(n14762), .A(n15427), .B(n14761), .ZN(
        n14768) );
  OAI211_X1 U16013 ( .C1(n14766), .C2(n14765), .A(n15426), .B(n14764), .ZN(
        n14767) );
  NAND3_X1 U16014 ( .A1(n14769), .A2(n14768), .A3(n14767), .ZN(P1_U3246) );
  OAI21_X1 U16015 ( .B1(n15430), .B2(n15480), .A(n14770), .ZN(n14771) );
  AOI21_X1 U16016 ( .B1(n14772), .B2(n15423), .A(n14771), .ZN(n14781) );
  OAI211_X1 U16017 ( .C1(n14775), .C2(n14774), .A(n15426), .B(n14773), .ZN(
        n14780) );
  OAI211_X1 U16018 ( .C1(n14778), .C2(n14777), .A(n15427), .B(n14776), .ZN(
        n14779) );
  NAND3_X1 U16019 ( .A1(n14781), .A2(n14780), .A3(n14779), .ZN(P1_U3249) );
  INV_X1 U16020 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15483) );
  OAI21_X1 U16021 ( .B1(n15430), .B2(n15483), .A(n14782), .ZN(n14783) );
  AOI21_X1 U16022 ( .B1(n14784), .B2(n15423), .A(n14783), .ZN(n14793) );
  OAI211_X1 U16023 ( .C1(n14787), .C2(n14786), .A(n15426), .B(n14785), .ZN(
        n14792) );
  OAI211_X1 U16024 ( .C1(n14790), .C2(n14789), .A(n14788), .B(n15427), .ZN(
        n14791) );
  NAND3_X1 U16025 ( .A1(n14793), .A2(n14792), .A3(n14791), .ZN(P1_U3250) );
  OAI211_X1 U16026 ( .C1(n14796), .C2(n14795), .A(n14794), .B(n15427), .ZN(
        n14805) );
  INV_X1 U16027 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15519) );
  OAI21_X1 U16028 ( .B1(n15430), .B2(n15519), .A(n14797), .ZN(n14798) );
  AOI21_X1 U16029 ( .B1(n14799), .B2(n15423), .A(n14798), .ZN(n14804) );
  OAI211_X1 U16030 ( .C1(n14802), .C2(n14801), .A(n14800), .B(n15426), .ZN(
        n14803) );
  NAND3_X1 U16031 ( .A1(n14805), .A2(n14804), .A3(n14803), .ZN(P1_U3253) );
  OAI211_X1 U16032 ( .C1(n14808), .C2(n14807), .A(n14806), .B(n15427), .ZN(
        n14819) );
  NAND2_X1 U16033 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14810)
         );
  NAND2_X1 U16034 ( .A1(n15381), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14809) );
  OAI211_X1 U16035 ( .C1(n14812), .C2(n14811), .A(n14810), .B(n14809), .ZN(
        n14813) );
  INV_X1 U16036 ( .A(n14813), .ZN(n14818) );
  OAI211_X1 U16037 ( .C1(n14816), .C2(n14815), .A(n14814), .B(n15426), .ZN(
        n14817) );
  NAND3_X1 U16038 ( .A1(n14819), .A2(n14818), .A3(n14817), .ZN(P1_U3256) );
  INV_X1 U16039 ( .A(n14820), .ZN(n14851) );
  NAND2_X1 U16040 ( .A1(n14825), .A2(n14824), .ZN(n14826) );
  INV_X1 U16041 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n16000) );
  XNOR2_X1 U16042 ( .A(n14827), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n15409) );
  NAND2_X1 U16043 ( .A1(n15410), .A2(n15409), .ZN(n15408) );
  NAND2_X1 U16044 ( .A1(n15418), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n14828) );
  NAND2_X1 U16045 ( .A1(n15408), .A2(n14828), .ZN(n15387) );
  INV_X1 U16046 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14829) );
  XNOR2_X1 U16047 ( .A(n15394), .B(n14829), .ZN(n15386) );
  NAND2_X1 U16048 ( .A1(n15387), .A2(n15386), .ZN(n15385) );
  NAND2_X1 U16049 ( .A1(n15394), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n14830) );
  NAND2_X1 U16050 ( .A1(n15385), .A2(n14830), .ZN(n14831) );
  NOR2_X1 U16051 ( .A1(n14831), .A2(n15404), .ZN(n14832) );
  INV_X1 U16052 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15399) );
  XOR2_X1 U16053 ( .A(n14834), .B(n14833), .Z(n14848) );
  INV_X1 U16054 ( .A(n14848), .ZN(n14845) );
  OAI21_X1 U16055 ( .B1(n14837), .B2(n14836), .A(n14835), .ZN(n14838) );
  XNOR2_X1 U16056 ( .A(n14838), .B(n15424), .ZN(n15422) );
  OAI22_X1 U16057 ( .A1(n15422), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n15424), 
        .B2(n14838), .ZN(n15414) );
  XNOR2_X1 U16058 ( .A(n15418), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n15415) );
  NOR2_X1 U16059 ( .A1(n15414), .A2(n15415), .ZN(n15412) );
  AOI21_X1 U16060 ( .B1(n15418), .B2(P1_REG2_REG_16__SCAN_IN), .A(n15412), 
        .ZN(n15391) );
  NAND2_X1 U16061 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n15394), .ZN(n14839) );
  OAI21_X1 U16062 ( .B1(n15394), .B2(P1_REG2_REG_17__SCAN_IN), .A(n14839), 
        .ZN(n15390) );
  NOR2_X1 U16063 ( .A1(n15391), .A2(n15390), .ZN(n15389) );
  AOI21_X1 U16064 ( .B1(n15394), .B2(P1_REG2_REG_17__SCAN_IN), .A(n15389), 
        .ZN(n14841) );
  NOR2_X1 U16065 ( .A1(n14841), .A2(n14840), .ZN(n14843) );
  AOI21_X1 U16066 ( .B1(n14841), .B2(n14840), .A(n14843), .ZN(n14842) );
  INV_X1 U16067 ( .A(n14842), .ZN(n15401) );
  NOR2_X1 U16068 ( .A1(n15401), .A2(n15020), .ZN(n15400) );
  NOR2_X1 U16069 ( .A1(n14843), .A2(n15400), .ZN(n14844) );
  XOR2_X1 U16070 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14844), .Z(n14846) );
  AOI21_X1 U16071 ( .B1(n14846), .B2(n15426), .A(n15423), .ZN(n14847) );
  OAI21_X1 U16072 ( .B1(n14848), .B2(n15397), .A(n14847), .ZN(n14850) );
  INV_X1 U16073 ( .A(n14852), .ZN(n14859) );
  NAND2_X1 U16074 ( .A1(n14859), .A2(n15094), .ZN(n14858) );
  XNOR2_X1 U16075 ( .A(n15091), .B(n14858), .ZN(n14853) );
  NAND2_X1 U16076 ( .A1(n14853), .A2(n15071), .ZN(n15090) );
  NAND2_X1 U16077 ( .A1(n14855), .A2(n14854), .ZN(n15092) );
  NOR2_X1 U16078 ( .A1(n15667), .A2(n15092), .ZN(n14861) );
  NOR2_X1 U16079 ( .A1(n15091), .A2(n15078), .ZN(n14856) );
  AOI211_X1 U16080 ( .C1(n15667), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14861), 
        .B(n14856), .ZN(n14857) );
  OAI21_X1 U16081 ( .B1(n15090), .B2(n15086), .A(n14857), .ZN(P1_U3263) );
  OAI211_X1 U16082 ( .C1(n14859), .C2(n15094), .A(n15071), .B(n14858), .ZN(
        n15093) );
  NOR2_X1 U16083 ( .A1(n15094), .A2(n15078), .ZN(n14860) );
  AOI211_X1 U16084 ( .C1(n15667), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14861), 
        .B(n14860), .ZN(n14862) );
  OAI21_X1 U16085 ( .B1(n15086), .B2(n15093), .A(n14862), .ZN(P1_U3264) );
  INV_X1 U16086 ( .A(n14863), .ZN(n14864) );
  AOI21_X1 U16087 ( .B1(n14864), .B2(n14871), .A(n15747), .ZN(n14867) );
  AOI21_X1 U16088 ( .B1(n14867), .B2(n14866), .A(n14865), .ZN(n15110) );
  OAI21_X1 U16089 ( .B1(n14886), .B2(n14868), .A(n15071), .ZN(n14870) );
  NOR2_X1 U16090 ( .A1(n14870), .A2(n14869), .ZN(n15104) );
  INV_X1 U16091 ( .A(n15104), .ZN(n14878) );
  OR2_X1 U16092 ( .A1(n14872), .A2(n14871), .ZN(n15107) );
  NAND3_X1 U16093 ( .A1(n15107), .A2(n15106), .A3(n15088), .ZN(n14877) );
  OAI22_X1 U16094 ( .A1(n15021), .A2(n14874), .B1(n14873), .B2(n15660), .ZN(
        n14875) );
  AOI21_X1 U16095 ( .B1(n15105), .B2(n15066), .A(n14875), .ZN(n14876) );
  OAI211_X1 U16096 ( .C1(n14878), .C2(n15086), .A(n14877), .B(n14876), .ZN(
        n14879) );
  INV_X1 U16097 ( .A(n14879), .ZN(n14880) );
  OAI21_X1 U16098 ( .B1(n15110), .B2(n15667), .A(n14880), .ZN(P1_U3265) );
  AOI21_X1 U16099 ( .B1(n8234), .B2(n14882), .A(n14881), .ZN(n15117) );
  XNOR2_X1 U16100 ( .A(n14883), .B(n8234), .ZN(n15111) );
  NAND2_X1 U16101 ( .A1(n15111), .A2(n15083), .ZN(n14896) );
  NAND2_X1 U16102 ( .A1(n14902), .A2(n15114), .ZN(n14884) );
  NAND2_X1 U16103 ( .A1(n14884), .A2(n15071), .ZN(n14885) );
  NOR2_X1 U16104 ( .A1(n14886), .A2(n14885), .ZN(n15112) );
  NAND2_X1 U16105 ( .A1(n15114), .A2(n15066), .ZN(n14892) );
  OAI22_X1 U16106 ( .A1(n14888), .A2(n15041), .B1(n14887), .B2(n15042), .ZN(
        n15113) );
  INV_X1 U16107 ( .A(n14889), .ZN(n14890) );
  AOI22_X1 U16108 ( .A1(n15021), .A2(n15113), .B1(n15043), .B2(n14890), .ZN(
        n14891) );
  OAI211_X1 U16109 ( .C1(n15021), .C2(n14893), .A(n14892), .B(n14891), .ZN(
        n14894) );
  AOI21_X1 U16110 ( .B1(n15112), .B2(n15049), .A(n14894), .ZN(n14895) );
  OAI211_X1 U16111 ( .C1(n15117), .C2(n14897), .A(n14896), .B(n14895), .ZN(
        P1_U3266) );
  OAI21_X1 U16112 ( .B1(n14899), .B2(n14900), .A(n14898), .ZN(n15124) );
  XOR2_X1 U16113 ( .A(n14901), .B(n14900), .Z(n15118) );
  NAND2_X1 U16114 ( .A1(n15118), .A2(n15083), .ZN(n14911) );
  AOI21_X1 U16115 ( .B1(n14915), .B2(n15121), .A(n15731), .ZN(n14903) );
  AND2_X1 U16116 ( .A1(n14903), .A2(n14902), .ZN(n15119) );
  NAND2_X1 U16117 ( .A1(n15121), .A2(n15066), .ZN(n14907) );
  OAI22_X1 U16118 ( .A1(n14926), .A2(n15041), .B1(n14904), .B2(n15042), .ZN(
        n15120) );
  AOI22_X1 U16119 ( .A1(n15021), .A2(n15120), .B1(n14905), .B2(n15043), .ZN(
        n14906) );
  OAI211_X1 U16120 ( .C1(n15021), .C2(n14908), .A(n14907), .B(n14906), .ZN(
        n14909) );
  AOI21_X1 U16121 ( .B1(n15119), .B2(n15049), .A(n14909), .ZN(n14910) );
  OAI211_X1 U16122 ( .C1(n15124), .C2(n15069), .A(n14911), .B(n14910), .ZN(
        P1_U3267) );
  XNOR2_X1 U16123 ( .A(n14912), .B(n14914), .ZN(n15132) );
  OAI21_X1 U16124 ( .B1(n7309), .B2(n14914), .A(n14913), .ZN(n15130) );
  OAI211_X1 U16125 ( .C1(n14932), .C2(n15128), .A(n15071), .B(n14915), .ZN(
        n15127) );
  OAI22_X1 U16126 ( .A1(n15021), .A2(n14917), .B1(n14916), .B2(n15660), .ZN(
        n14918) );
  AOI21_X1 U16127 ( .B1(n15125), .B2(n15021), .A(n14918), .ZN(n14921) );
  NAND2_X1 U16128 ( .A1(n14919), .A2(n15066), .ZN(n14920) );
  OAI211_X1 U16129 ( .C1(n15127), .C2(n15086), .A(n14921), .B(n14920), .ZN(
        n14922) );
  AOI21_X1 U16130 ( .B1(n15130), .B2(n15083), .A(n14922), .ZN(n14923) );
  OAI21_X1 U16131 ( .B1(n15069), .B2(n15132), .A(n14923), .ZN(P1_U3268) );
  OAI21_X1 U16132 ( .B1(n14925), .B2(n14929), .A(n14924), .ZN(n15133) );
  OAI22_X1 U16133 ( .A1(n14927), .A2(n15041), .B1(n14926), .B2(n15042), .ZN(
        n14931) );
  AOI211_X1 U16134 ( .C1(n14929), .C2(n14928), .A(n15747), .B(n7412), .ZN(
        n14930) );
  AOI211_X1 U16135 ( .C1(n15025), .C2(n15133), .A(n14931), .B(n14930), .ZN(
        n15137) );
  AOI211_X1 U16136 ( .C1(n15135), .C2(n7592), .A(n15731), .B(n14932), .ZN(
        n15134) );
  NAND2_X1 U16137 ( .A1(n15134), .A2(n15049), .ZN(n14935) );
  AOI22_X1 U16138 ( .A1(n14933), .A2(n15043), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15667), .ZN(n14934) );
  OAI211_X1 U16139 ( .C1(n14936), .C2(n15078), .A(n14935), .B(n14934), .ZN(
        n14937) );
  AOI21_X1 U16140 ( .B1(n15034), .B2(n15133), .A(n14937), .ZN(n14938) );
  OAI21_X1 U16141 ( .B1(n15137), .B2(n15667), .A(n14938), .ZN(P1_U3269) );
  XNOR2_X1 U16142 ( .A(n14940), .B(n14939), .ZN(n15145) );
  OAI21_X1 U16143 ( .B1(n14943), .B2(n14942), .A(n14941), .ZN(n15142) );
  NAND2_X1 U16144 ( .A1(n15142), .A2(n15083), .ZN(n14952) );
  AOI211_X1 U16145 ( .C1(n15141), .C2(n7593), .A(n15731), .B(n14944), .ZN(
        n15139) );
  INV_X1 U16146 ( .A(n14945), .ZN(n14946) );
  AOI22_X1 U16147 ( .A1(n14946), .A2(n15043), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15667), .ZN(n14948) );
  NAND2_X1 U16148 ( .A1(n15140), .A2(n15021), .ZN(n14947) );
  OAI211_X1 U16149 ( .C1(n14949), .C2(n15078), .A(n14948), .B(n14947), .ZN(
        n14950) );
  AOI21_X1 U16150 ( .B1(n15139), .B2(n15049), .A(n14950), .ZN(n14951) );
  OAI211_X1 U16151 ( .C1(n15145), .C2(n15069), .A(n14952), .B(n14951), .ZN(
        P1_U3270) );
  XNOR2_X1 U16152 ( .A(n14954), .B(n14953), .ZN(n15151) );
  NAND2_X1 U16153 ( .A1(n14959), .A2(n7247), .ZN(n14955) );
  NAND2_X1 U16154 ( .A1(n14955), .A2(n15071), .ZN(n14956) );
  NOR2_X1 U16155 ( .A1(n14957), .A2(n14956), .ZN(n15147) );
  AOI22_X1 U16156 ( .A1(n14958), .A2(n15076), .B1(n15075), .B2(n14984), .ZN(
        n15146) );
  NAND2_X1 U16157 ( .A1(n14959), .A2(n15066), .ZN(n14962) );
  AOI22_X1 U16158 ( .A1(n14960), .A2(n15043), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15667), .ZN(n14961) );
  OAI211_X1 U16159 ( .C1(n15667), .C2(n15146), .A(n14962), .B(n14961), .ZN(
        n14963) );
  AOI21_X1 U16160 ( .B1(n15147), .B2(n15049), .A(n14963), .ZN(n14967) );
  XNOR2_X1 U16161 ( .A(n14964), .B(n14965), .ZN(n15149) );
  NAND2_X1 U16162 ( .A1(n15149), .A2(n15088), .ZN(n14966) );
  OAI211_X1 U16163 ( .C1(n15151), .C2(n15052), .A(n14967), .B(n14966), .ZN(
        P1_U3271) );
  XNOR2_X1 U16164 ( .A(n14968), .B(n9599), .ZN(n15158) );
  OAI21_X1 U16165 ( .B1(n7320), .B2(n9599), .A(n14969), .ZN(n15155) );
  AOI21_X1 U16166 ( .B1(n14981), .B2(n15154), .A(n15731), .ZN(n14970) );
  AND2_X1 U16167 ( .A1(n14970), .A2(n7247), .ZN(n15152) );
  NAND2_X1 U16168 ( .A1(n15152), .A2(n15049), .ZN(n14976) );
  AOI22_X1 U16169 ( .A1(n14971), .A2(n15043), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15667), .ZN(n14975) );
  NAND2_X1 U16170 ( .A1(n15154), .A2(n15066), .ZN(n14974) );
  OAI22_X1 U16171 ( .A1(n14972), .A2(n15042), .B1(n15000), .B2(n15041), .ZN(
        n15153) );
  NAND2_X1 U16172 ( .A1(n15153), .A2(n15021), .ZN(n14973) );
  NAND4_X1 U16173 ( .A1(n14976), .A2(n14975), .A3(n14974), .A4(n14973), .ZN(
        n14977) );
  AOI21_X1 U16174 ( .B1(n15155), .B2(n15088), .A(n14977), .ZN(n14978) );
  OAI21_X1 U16175 ( .B1(n15158), .B2(n15052), .A(n14978), .ZN(P1_U3272) );
  AOI21_X1 U16176 ( .B1(n14990), .B2(n14979), .A(n7327), .ZN(n15166) );
  INV_X1 U16177 ( .A(n14999), .ZN(n14980) );
  AOI21_X1 U16178 ( .B1(n14980), .B2(n14988), .A(n15731), .ZN(n14982) );
  NAND2_X1 U16179 ( .A1(n14982), .A2(n14981), .ZN(n15160) );
  AND2_X1 U16180 ( .A1(n15031), .A2(n15075), .ZN(n14983) );
  AOI21_X1 U16181 ( .B1(n14984), .B2(n15076), .A(n14983), .ZN(n15159) );
  AOI22_X1 U16182 ( .A1(n14985), .A2(n15043), .B1(n15667), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14986) );
  OAI21_X1 U16183 ( .B1(n15159), .B2(n15667), .A(n14986), .ZN(n14987) );
  AOI21_X1 U16184 ( .B1(n14988), .B2(n15066), .A(n14987), .ZN(n14989) );
  OAI21_X1 U16185 ( .B1(n15160), .B2(n15086), .A(n14989), .ZN(n14993) );
  NOR2_X1 U16186 ( .A1(n14991), .A2(n14990), .ZN(n15163) );
  NOR3_X1 U16187 ( .A1(n15163), .A2(n15162), .A3(n15069), .ZN(n14992) );
  AOI211_X1 U16188 ( .C1(n15166), .C2(n15083), .A(n14993), .B(n14992), .ZN(
        n14994) );
  INV_X1 U16189 ( .A(n14994), .ZN(P1_U3273) );
  XNOR2_X1 U16190 ( .A(n14996), .B(n14995), .ZN(n15171) );
  NAND2_X1 U16191 ( .A1(n15170), .A2(n15017), .ZN(n14997) );
  NAND2_X1 U16192 ( .A1(n14997), .A2(n15071), .ZN(n14998) );
  NOR2_X1 U16193 ( .A1(n14999), .A2(n14998), .ZN(n15168) );
  NAND2_X1 U16194 ( .A1(n15168), .A2(n15049), .ZN(n15008) );
  OR2_X1 U16195 ( .A1(n15000), .A2(n15042), .ZN(n15003) );
  NAND2_X1 U16196 ( .A1(n15001), .A2(n15075), .ZN(n15002) );
  NAND2_X1 U16197 ( .A1(n15003), .A2(n15002), .ZN(n15169) );
  INV_X1 U16198 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15005) );
  OAI22_X1 U16199 ( .A1(n15021), .A2(n15005), .B1(n15004), .B2(n15660), .ZN(
        n15006) );
  AOI21_X1 U16200 ( .B1(n15169), .B2(n15021), .A(n15006), .ZN(n15007) );
  OAI211_X1 U16201 ( .C1(n15009), .C2(n15078), .A(n15008), .B(n15007), .ZN(
        n15012) );
  XNOR2_X1 U16202 ( .A(n15010), .B(n7937), .ZN(n15174) );
  NOR2_X1 U16203 ( .A1(n15174), .A2(n15069), .ZN(n15011) );
  AOI211_X1 U16204 ( .C1(n15171), .C2(n15083), .A(n15012), .B(n15011), .ZN(
        n15013) );
  INV_X1 U16205 ( .A(n15013), .ZN(P1_U3274) );
  NAND2_X1 U16206 ( .A1(n15026), .A2(n15014), .ZN(n15015) );
  NAND2_X1 U16207 ( .A1(n15016), .A2(n15015), .ZN(n15180) );
  OAI211_X1 U16208 ( .C1(n15018), .C2(n15040), .A(n15071), .B(n15017), .ZN(
        n15178) );
  OAI22_X1 U16209 ( .A1(n15021), .A2(n15020), .B1(n15019), .B2(n15660), .ZN(
        n15022) );
  AOI21_X1 U16210 ( .B1(n15175), .B2(n15066), .A(n15022), .ZN(n15023) );
  OAI21_X1 U16211 ( .B1(n15178), .B2(n15086), .A(n15023), .ZN(n15033) );
  AND2_X1 U16212 ( .A1(n15057), .A2(n15075), .ZN(n15024) );
  AOI21_X1 U16213 ( .B1(n15180), .B2(n15025), .A(n15024), .ZN(n15030) );
  XNOR2_X1 U16214 ( .A(n15027), .B(n15026), .ZN(n15028) );
  NAND2_X1 U16215 ( .A1(n15028), .A2(n15993), .ZN(n15029) );
  NAND2_X1 U16216 ( .A1(n15031), .A2(n15076), .ZN(n15177) );
  AOI21_X1 U16217 ( .B1(n15182), .B2(n15177), .A(n15667), .ZN(n15032) );
  AOI211_X1 U16218 ( .C1(n15034), .C2(n15180), .A(n15033), .B(n15032), .ZN(
        n15035) );
  INV_X1 U16219 ( .A(n15035), .ZN(P1_U3275) );
  XNOR2_X1 U16220 ( .A(n7189), .B(n15039), .ZN(n15188) );
  INV_X1 U16221 ( .A(n15036), .ZN(n15037) );
  AOI21_X1 U16222 ( .B1(n15039), .B2(n15038), .A(n15037), .ZN(n15185) );
  NAND2_X1 U16223 ( .A1(n15185), .A2(n15088), .ZN(n15051) );
  AOI211_X1 U16224 ( .C1(n16026), .C2(n15062), .A(n15731), .B(n15040), .ZN(
        n15183) );
  INV_X1 U16225 ( .A(n16026), .ZN(n15047) );
  OAI22_X1 U16226 ( .A1(n16018), .A2(n15042), .B1(n16017), .B2(n15041), .ZN(
        n15184) );
  INV_X1 U16227 ( .A(n16030), .ZN(n15044) );
  AOI22_X1 U16228 ( .A1(n15184), .A2(n15021), .B1(n15044), .B2(n15043), .ZN(
        n15046) );
  NAND2_X1 U16229 ( .A1(n15667), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n15045) );
  OAI211_X1 U16230 ( .C1(n15047), .C2(n15078), .A(n15046), .B(n15045), .ZN(
        n15048) );
  AOI21_X1 U16231 ( .B1(n15183), .B2(n15049), .A(n15048), .ZN(n15050) );
  OAI211_X1 U16232 ( .C1(n15188), .C2(n15052), .A(n15051), .B(n15050), .ZN(
        P1_U3276) );
  XNOR2_X1 U16233 ( .A(n15053), .B(n15055), .ZN(n15194) );
  OAI21_X1 U16234 ( .B1(n15056), .B2(n15055), .A(n15054), .ZN(n15061) );
  NAND2_X1 U16235 ( .A1(n15057), .A2(n15076), .ZN(n15060) );
  NAND2_X1 U16236 ( .A1(n15058), .A2(n15075), .ZN(n15059) );
  NAND2_X1 U16237 ( .A1(n15060), .A2(n15059), .ZN(n16012) );
  AOI21_X1 U16238 ( .B1(n15061), .B2(n15993), .A(n16012), .ZN(n15193) );
  INV_X1 U16239 ( .A(n15193), .ZN(n15065) );
  OAI21_X1 U16240 ( .B1(n15189), .B2(n15074), .A(n15062), .ZN(n15190) );
  OAI22_X1 U16241 ( .A1(n15190), .A2(n15063), .B1(n16015), .B2(n15660), .ZN(
        n15064) );
  OAI21_X1 U16242 ( .B1(n15065), .B2(n15064), .A(n15021), .ZN(n15068) );
  AOI22_X1 U16243 ( .A1(n16008), .A2(n15066), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n15667), .ZN(n15067) );
  OAI211_X1 U16244 ( .C1(n15194), .C2(n15069), .A(n15068), .B(n15067), .ZN(
        P1_U3277) );
  OAI21_X1 U16245 ( .B1(n7233), .B2(n15081), .A(n7324), .ZN(n15997) );
  NAND2_X1 U16246 ( .A1(n15077), .A2(n15070), .ZN(n15072) );
  NAND2_X1 U16247 ( .A1(n15072), .A2(n15071), .ZN(n15073) );
  OR2_X1 U16248 ( .A1(n15074), .A2(n15073), .ZN(n15989) );
  AOI22_X1 U16249 ( .A1(n15977), .A2(n15076), .B1(n15075), .B2(n15979), .ZN(
        n15988) );
  OAI22_X1 U16250 ( .A1(n15667), .A2(n15988), .B1(n15987), .B2(n15660), .ZN(
        n15080) );
  INV_X1 U16251 ( .A(n15077), .ZN(n15991) );
  NOR2_X1 U16252 ( .A1(n15991), .A2(n15078), .ZN(n15079) );
  AOI211_X1 U16253 ( .C1(n15667), .C2(P1_REG2_REG_15__SCAN_IN), .A(n15080), 
        .B(n15079), .ZN(n15085) );
  NAND2_X1 U16254 ( .A1(n15082), .A2(n15081), .ZN(n15992) );
  NAND3_X1 U16255 ( .A1(n15994), .A2(n15992), .A3(n15083), .ZN(n15084) );
  OAI211_X1 U16256 ( .C1(n15989), .C2(n15086), .A(n15085), .B(n15084), .ZN(
        n15087) );
  AOI21_X1 U16257 ( .B1(n15088), .B2(n15997), .A(n15087), .ZN(n15089) );
  INV_X1 U16258 ( .A(n15089), .ZN(P1_U3278) );
  OAI211_X1 U16259 ( .C1(n15091), .C2(n15990), .A(n15090), .B(n15092), .ZN(
        n15195) );
  MUX2_X1 U16260 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15195), .S(n16001), .Z(
        P1_U3559) );
  OAI211_X1 U16261 ( .C1(n15094), .C2(n15990), .A(n15093), .B(n15092), .ZN(
        n15196) );
  MUX2_X1 U16262 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15196), .S(n16001), .Z(
        P1_U3558) );
  NOR2_X1 U16263 ( .A1(n15096), .A2(n15731), .ZN(n15101) );
  OAI211_X1 U16264 ( .C1(n15099), .C2(n15990), .A(n15098), .B(n15097), .ZN(
        n15100) );
  AOI21_X1 U16265 ( .B1(n15949), .B2(n15105), .A(n15104), .ZN(n15109) );
  NAND3_X1 U16266 ( .A1(n15107), .A2(n15106), .A3(n15998), .ZN(n15108) );
  NAND3_X1 U16267 ( .A1(n15110), .A2(n15109), .A3(n15108), .ZN(n15197) );
  MUX2_X1 U16268 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15197), .S(n16001), .Z(
        P1_U3556) );
  NAND2_X1 U16269 ( .A1(n15111), .A2(n15993), .ZN(n15116) );
  AOI211_X1 U16270 ( .C1(n15949), .C2(n15114), .A(n15113), .B(n15112), .ZN(
        n15115) );
  OAI211_X1 U16271 ( .C1(n15953), .C2(n15117), .A(n15116), .B(n15115), .ZN(
        n15198) );
  MUX2_X1 U16272 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15198), .S(n16001), .Z(
        P1_U3555) );
  NAND2_X1 U16273 ( .A1(n15118), .A2(n15993), .ZN(n15123) );
  AOI211_X1 U16274 ( .C1(n15949), .C2(n15121), .A(n15120), .B(n15119), .ZN(
        n15122) );
  OAI211_X1 U16275 ( .C1(n15953), .C2(n15124), .A(n15123), .B(n15122), .ZN(
        n15199) );
  MUX2_X1 U16276 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15199), .S(n16001), .Z(
        P1_U3554) );
  INV_X1 U16277 ( .A(n15125), .ZN(n15126) );
  OAI211_X1 U16278 ( .C1(n15128), .C2(n15990), .A(n15127), .B(n15126), .ZN(
        n15129) );
  AOI21_X1 U16279 ( .B1(n15130), .B2(n15993), .A(n15129), .ZN(n15131) );
  OAI21_X1 U16280 ( .B1(n15953), .B2(n15132), .A(n15131), .ZN(n15200) );
  MUX2_X1 U16281 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15200), .S(n16001), .Z(
        P1_U3553) );
  INV_X1 U16282 ( .A(n15133), .ZN(n15138) );
  AOI21_X1 U16283 ( .B1(n15949), .B2(n15135), .A(n15134), .ZN(n15136) );
  OAI211_X1 U16284 ( .C1(n15138), .C2(n15773), .A(n15137), .B(n15136), .ZN(
        n15201) );
  MUX2_X1 U16285 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15201), .S(n16001), .Z(
        P1_U3552) );
  AOI211_X1 U16286 ( .C1(n15949), .C2(n15141), .A(n15140), .B(n15139), .ZN(
        n15144) );
  NAND2_X1 U16287 ( .A1(n15142), .A2(n15993), .ZN(n15143) );
  OAI211_X1 U16288 ( .C1(n15953), .C2(n15145), .A(n15144), .B(n15143), .ZN(
        n15202) );
  MUX2_X1 U16289 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15202), .S(n16001), .Z(
        P1_U3551) );
  OAI21_X1 U16290 ( .B1(n7591), .B2(n15990), .A(n15146), .ZN(n15148) );
  AOI211_X1 U16291 ( .C1(n15149), .C2(n15998), .A(n15148), .B(n15147), .ZN(
        n15150) );
  OAI21_X1 U16292 ( .B1(n15151), .B2(n15747), .A(n15150), .ZN(n15203) );
  MUX2_X1 U16293 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15203), .S(n16001), .Z(
        P1_U3550) );
  AOI211_X1 U16294 ( .C1(n15949), .C2(n15154), .A(n15153), .B(n15152), .ZN(
        n15157) );
  NAND2_X1 U16295 ( .A1(n15155), .A2(n15998), .ZN(n15156) );
  OAI211_X1 U16296 ( .C1(n15158), .C2(n15747), .A(n15157), .B(n15156), .ZN(
        n15204) );
  MUX2_X1 U16297 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15204), .S(n16001), .Z(
        P1_U3549) );
  OAI211_X1 U16298 ( .C1(n15161), .C2(n15990), .A(n15160), .B(n15159), .ZN(
        n15165) );
  NOR3_X1 U16299 ( .A1(n15163), .A2(n15162), .A3(n15953), .ZN(n15164) );
  AOI211_X1 U16300 ( .C1(n15166), .C2(n15993), .A(n15165), .B(n15164), .ZN(
        n15167) );
  INV_X1 U16301 ( .A(n15167), .ZN(n15205) );
  MUX2_X1 U16302 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15205), .S(n16001), .Z(
        P1_U3548) );
  AOI211_X1 U16303 ( .C1(n15949), .C2(n15170), .A(n15169), .B(n15168), .ZN(
        n15173) );
  NAND2_X1 U16304 ( .A1(n15171), .A2(n15993), .ZN(n15172) );
  OAI211_X1 U16305 ( .C1(n15953), .C2(n15174), .A(n15173), .B(n15172), .ZN(
        n15206) );
  MUX2_X1 U16306 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15206), .S(n16001), .Z(
        P1_U3547) );
  NAND2_X1 U16307 ( .A1(n15175), .A2(n15949), .ZN(n15176) );
  NAND3_X1 U16308 ( .A1(n15178), .A2(n15177), .A3(n15176), .ZN(n15179) );
  AOI21_X1 U16309 ( .B1(n15180), .B2(n15912), .A(n15179), .ZN(n15181) );
  NAND2_X1 U16310 ( .A1(n15182), .A2(n15181), .ZN(n15207) );
  MUX2_X1 U16311 ( .A(n15207), .B(P1_REG1_REG_18__SCAN_IN), .S(n15999), .Z(
        P1_U3546) );
  AOI211_X1 U16312 ( .C1(n15949), .C2(n16026), .A(n15184), .B(n15183), .ZN(
        n15187) );
  NAND2_X1 U16313 ( .A1(n15185), .A2(n15998), .ZN(n15186) );
  OAI211_X1 U16314 ( .C1(n15747), .C2(n15188), .A(n15187), .B(n15186), .ZN(
        n15208) );
  MUX2_X1 U16315 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15208), .S(n16001), .Z(
        P1_U3545) );
  OAI22_X1 U16316 ( .A1(n15190), .A2(n15731), .B1(n15189), .B2(n15990), .ZN(
        n15191) );
  INV_X1 U16317 ( .A(n15191), .ZN(n15192) );
  OAI211_X1 U16318 ( .C1(n15953), .C2(n15194), .A(n15193), .B(n15192), .ZN(
        n15209) );
  MUX2_X1 U16319 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15209), .S(n16001), .Z(
        P1_U3544) );
  MUX2_X1 U16320 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15195), .S(n16005), .Z(
        P1_U3527) );
  MUX2_X1 U16321 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15196), .S(n16005), .Z(
        P1_U3526) );
  MUX2_X1 U16322 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15197), .S(n16005), .Z(
        P1_U3524) );
  MUX2_X1 U16323 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15198), .S(n16005), .Z(
        P1_U3523) );
  MUX2_X1 U16324 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15199), .S(n16005), .Z(
        P1_U3522) );
  MUX2_X1 U16325 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15200), .S(n16005), .Z(
        P1_U3521) );
  MUX2_X1 U16326 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15201), .S(n16005), .Z(
        P1_U3520) );
  MUX2_X1 U16327 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15202), .S(n16005), .Z(
        P1_U3519) );
  MUX2_X1 U16328 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15203), .S(n16005), .Z(
        P1_U3518) );
  MUX2_X1 U16329 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15204), .S(n16005), .Z(
        P1_U3517) );
  MUX2_X1 U16330 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15205), .S(n16005), .Z(
        P1_U3516) );
  MUX2_X1 U16331 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15206), .S(n16005), .Z(
        P1_U3515) );
  MUX2_X1 U16332 ( .A(n15207), .B(P1_REG0_REG_18__SCAN_IN), .S(n16002), .Z(
        P1_U3513) );
  MUX2_X1 U16333 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15208), .S(n16005), .Z(
        P1_U3510) );
  MUX2_X1 U16334 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15209), .S(n16005), .Z(
        P1_U3507) );
  NOR4_X1 U16335 ( .A1(n15210), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9537), .A4(
        P1_U3086), .ZN(n15211) );
  AOI21_X1 U16336 ( .B1(n15212), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15211), 
        .ZN(n15213) );
  OAI21_X1 U16337 ( .B1(n15214), .B2(n15233), .A(n15213), .ZN(P1_U3324) );
  OAI222_X1 U16338 ( .A1(n15235), .A2(n15217), .B1(n15233), .B2(n15216), .C1(
        n15215), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U16339 ( .A1(n15220), .A2(P1_U3086), .B1(n15233), .B2(n15219), 
        .C1(n15218), .C2(n15235), .ZN(P1_U3326) );
  OAI222_X1 U16340 ( .A1(P1_U3086), .A2(n15227), .B1(n15233), .B2(n15226), 
        .C1(n15225), .C2(n15224), .ZN(P1_U3328) );
  OAI222_X1 U16341 ( .A1(n15235), .A2(n15230), .B1(n15233), .B2(n15229), .C1(
        P1_U3086), .C2(n15228), .ZN(P1_U3329) );
  OAI222_X1 U16342 ( .A1(n15235), .A2(n15234), .B1(n15233), .B2(n15232), .C1(
        n15231), .C2(P1_U3086), .ZN(P1_U3331) );
  MUX2_X1 U16343 ( .A(n15237), .B(n15236), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16344 ( .A(n15238), .ZN(n15239) );
  MUX2_X1 U16345 ( .A(n15239), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U16346 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15240), .ZN(P1_U3323) );
  AND2_X1 U16347 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15240), .ZN(P1_U3322) );
  AND2_X1 U16348 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15240), .ZN(P1_U3321) );
  AND2_X1 U16349 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15240), .ZN(P1_U3320) );
  AND2_X1 U16350 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15240), .ZN(P1_U3319) );
  AND2_X1 U16351 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15240), .ZN(P1_U3318) );
  AND2_X1 U16352 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15240), .ZN(P1_U3317) );
  AND2_X1 U16353 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15240), .ZN(P1_U3316) );
  AND2_X1 U16354 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15240), .ZN(P1_U3315) );
  AND2_X1 U16355 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15240), .ZN(P1_U3314) );
  AND2_X1 U16356 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15240), .ZN(P1_U3313) );
  AND2_X1 U16357 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15240), .ZN(P1_U3312) );
  AND2_X1 U16358 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15240), .ZN(P1_U3311) );
  AND2_X1 U16359 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15240), .ZN(P1_U3310) );
  AND2_X1 U16360 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15240), .ZN(P1_U3309) );
  AND2_X1 U16361 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15240), .ZN(P1_U3308) );
  AND2_X1 U16362 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15240), .ZN(P1_U3307) );
  AND2_X1 U16363 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15240), .ZN(P1_U3306) );
  AND2_X1 U16364 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15240), .ZN(P1_U3305) );
  AND2_X1 U16365 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15240), .ZN(P1_U3304) );
  AND2_X1 U16366 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15240), .ZN(P1_U3303) );
  AND2_X1 U16367 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15240), .ZN(P1_U3302) );
  AND2_X1 U16368 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15240), .ZN(P1_U3301) );
  AND2_X1 U16369 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15240), .ZN(P1_U3300) );
  AND2_X1 U16370 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15240), .ZN(P1_U3299) );
  AND2_X1 U16371 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15240), .ZN(P1_U3298) );
  AND2_X1 U16372 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15240), .ZN(P1_U3297) );
  AND2_X1 U16373 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15240), .ZN(P1_U3296) );
  AND2_X1 U16374 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15240), .ZN(P1_U3295) );
  AND2_X1 U16375 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15240), .ZN(P1_U3294) );
  INV_X1 U16376 ( .A(n15241), .ZN(n15242) );
  AOI21_X1 U16377 ( .B1(n15243), .B2(n15247), .A(n15242), .ZN(P2_U3417) );
  AND2_X1 U16378 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15245), .ZN(P2_U3295) );
  AND2_X1 U16379 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15245), .ZN(P2_U3294) );
  AND2_X1 U16380 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15245), .ZN(P2_U3293) );
  AND2_X1 U16381 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15245), .ZN(P2_U3292) );
  AND2_X1 U16382 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15245), .ZN(P2_U3291) );
  AND2_X1 U16383 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15245), .ZN(P2_U3290) );
  AND2_X1 U16384 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15245), .ZN(P2_U3289) );
  AND2_X1 U16385 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15245), .ZN(P2_U3288) );
  AND2_X1 U16386 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15245), .ZN(P2_U3287) );
  AND2_X1 U16387 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15245), .ZN(P2_U3286) );
  AND2_X1 U16388 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15245), .ZN(P2_U3285) );
  AND2_X1 U16389 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15245), .ZN(P2_U3284) );
  AND2_X1 U16390 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15245), .ZN(P2_U3283) );
  AND2_X1 U16391 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15245), .ZN(P2_U3282) );
  AND2_X1 U16392 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15245), .ZN(P2_U3281) );
  AND2_X1 U16393 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15245), .ZN(P2_U3280) );
  AND2_X1 U16394 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15245), .ZN(P2_U3279) );
  AND2_X1 U16395 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15245), .ZN(P2_U3278) );
  AND2_X1 U16396 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15245), .ZN(P2_U3277) );
  AND2_X1 U16397 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15245), .ZN(P2_U3276) );
  AND2_X1 U16398 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15245), .ZN(P2_U3275) );
  AND2_X1 U16399 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15245), .ZN(P2_U3274) );
  AND2_X1 U16400 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15245), .ZN(P2_U3273) );
  AND2_X1 U16401 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15245), .ZN(P2_U3272) );
  AND2_X1 U16402 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15245), .ZN(P2_U3271) );
  AND2_X1 U16403 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15245), .ZN(P2_U3270) );
  AND2_X1 U16404 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15245), .ZN(P2_U3269) );
  AND2_X1 U16405 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15245), .ZN(P2_U3268) );
  AND2_X1 U16406 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15245), .ZN(P2_U3267) );
  AND2_X1 U16407 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15245), .ZN(P2_U3266) );
  NOR2_X1 U16408 ( .A1(n15271), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16409 ( .A1(P3_U3897), .A2(n15246), .ZN(P3_U3150) );
  INV_X1 U16410 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15248) );
  AOI22_X1 U16411 ( .A1(n15250), .A2(n15249), .B1(n15248), .B2(n15247), .ZN(
        P2_U3416) );
  AOI22_X1 U16412 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15333), .B1(n15251), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15256) );
  OAI22_X1 U16413 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15364), .B1(n15368), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15252) );
  NOR2_X1 U16414 ( .A1(n15374), .A2(n15252), .ZN(n15254) );
  AOI22_X1 U16415 ( .A1(n15271), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15253) );
  OAI221_X1 U16416 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n15256), .C1(n15255), .C2(
        n15254), .A(n15253), .ZN(P2_U3214) );
  AOI22_X1 U16417 ( .A1(n15271), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(n15374), 
        .B2(n15257), .ZN(n15269) );
  AOI211_X1 U16418 ( .C1(n15260), .C2(n15259), .A(n15258), .B(n15368), .ZN(
        n15267) );
  INV_X1 U16419 ( .A(n15261), .ZN(n15264) );
  INV_X1 U16420 ( .A(n15262), .ZN(n15263) );
  AOI211_X1 U16421 ( .C1(n15265), .C2(n15264), .A(n15263), .B(n15364), .ZN(
        n15266) );
  AOI211_X1 U16422 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(P2_U3088), .A(n15267), 
        .B(n15266), .ZN(n15268) );
  NAND2_X1 U16423 ( .A1(n15269), .A2(n15268), .ZN(P2_U3215) );
  AOI22_X1 U16424 ( .A1(n15271), .A2(P2_ADDR_REG_6__SCAN_IN), .B1(n15374), 
        .B2(n15270), .ZN(n15282) );
  AOI211_X1 U16425 ( .C1(n15274), .C2(n15273), .A(n15368), .B(n15272), .ZN(
        n15280) );
  OAI211_X1 U16426 ( .C1(n15277), .C2(n15276), .A(n15333), .B(n15275), .ZN(
        n15278) );
  INV_X1 U16427 ( .A(n15278), .ZN(n15279) );
  AOI211_X1 U16428 ( .C1(P2_REG3_REG_6__SCAN_IN), .C2(P2_U3088), .A(n15280), 
        .B(n15279), .ZN(n15281) );
  NAND2_X1 U16429 ( .A1(n15282), .A2(n15281), .ZN(P2_U3220) );
  INV_X1 U16430 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15299) );
  NOR2_X1 U16431 ( .A1(n15283), .A2(n15289), .ZN(n15285) );
  XNOR2_X1 U16432 ( .A(n15308), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15286) );
  AOI211_X1 U16433 ( .C1(n15287), .C2(n15286), .A(n15300), .B(n15368), .ZN(
        n15296) );
  NOR2_X1 U16434 ( .A1(n15289), .A2(n15288), .ZN(n15291) );
  NOR2_X1 U16435 ( .A1(n15291), .A2(n15290), .ZN(n15294) );
  NAND2_X1 U16436 ( .A1(n15308), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n15292) );
  OAI21_X1 U16437 ( .B1(n15308), .B2(P2_REG2_REG_16__SCAN_IN), .A(n15292), 
        .ZN(n15293) );
  NOR2_X1 U16438 ( .A1(n15294), .A2(n15293), .ZN(n15307) );
  AOI211_X1 U16439 ( .C1(n15294), .C2(n15293), .A(n15307), .B(n15364), .ZN(
        n15295) );
  AOI211_X1 U16440 ( .C1(n15308), .C2(n15374), .A(n15296), .B(n15295), .ZN(
        n15298) );
  OAI211_X1 U16441 ( .C1(n15299), .C2(n15377), .A(n15298), .B(n15297), .ZN(
        P2_U3230) );
  INV_X1 U16442 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15318) );
  NAND2_X1 U16443 ( .A1(n15308), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n15301) );
  INV_X1 U16444 ( .A(n15303), .ZN(n15306) );
  XNOR2_X1 U16445 ( .A(n15323), .B(n15302), .ZN(n15304) );
  INV_X1 U16446 ( .A(n15304), .ZN(n15305) );
  AOI211_X1 U16447 ( .C1(n15306), .C2(n15305), .A(n15325), .B(n15368), .ZN(
        n15315) );
  AOI21_X1 U16448 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n15308), .A(n15307), 
        .ZN(n15313) );
  INV_X1 U16449 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n15309) );
  XNOR2_X1 U16450 ( .A(n15323), .B(n15309), .ZN(n15311) );
  INV_X1 U16451 ( .A(n15311), .ZN(n15312) );
  INV_X1 U16452 ( .A(n15313), .ZN(n15310) );
  AOI211_X1 U16453 ( .C1(n15313), .C2(n15312), .A(n15320), .B(n15364), .ZN(
        n15314) );
  AOI211_X1 U16454 ( .C1(n15374), .C2(n15323), .A(n15315), .B(n15314), .ZN(
        n15317) );
  OAI211_X1 U16455 ( .C1(n15318), .C2(n15377), .A(n15317), .B(n15316), .ZN(
        P2_U3231) );
  INV_X1 U16456 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15336) );
  AND2_X1 U16457 ( .A1(n15323), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n15319) );
  NOR2_X1 U16458 ( .A1(n15320), .A2(n15319), .ZN(n15344) );
  XNOR2_X1 U16459 ( .A(n15344), .B(n15326), .ZN(n15321) );
  NAND2_X1 U16460 ( .A1(n15321), .A2(n8938), .ZN(n15341) );
  OAI21_X1 U16461 ( .B1(n15321), .B2(n8938), .A(n15341), .ZN(n15332) );
  NOR2_X1 U16462 ( .A1(n15322), .A2(n15343), .ZN(n15331) );
  INV_X1 U16463 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15329) );
  AND2_X1 U16464 ( .A1(n15323), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n15324) );
  NAND2_X1 U16465 ( .A1(n15327), .A2(n15326), .ZN(n15337) );
  OAI21_X1 U16466 ( .B1(n15327), .B2(n15326), .A(n15337), .ZN(n15328) );
  AOI211_X1 U16467 ( .C1(n15329), .C2(n15328), .A(n15338), .B(n15368), .ZN(
        n15330) );
  AOI211_X1 U16468 ( .C1(n15333), .C2(n15332), .A(n15331), .B(n15330), .ZN(
        n15335) );
  OAI211_X1 U16469 ( .C1(n15336), .C2(n15377), .A(n15335), .B(n15334), .ZN(
        P2_U3232) );
  NAND2_X1 U16470 ( .A1(n15374), .A2(n15339), .ZN(n15340) );
  INV_X1 U16471 ( .A(n15341), .ZN(n15342) );
  AOI21_X1 U16472 ( .B1(n15344), .B2(n15343), .A(n15342), .ZN(n15346) );
  MUX2_X1 U16473 ( .A(n14407), .B(P2_REG2_REG_19__SCAN_IN), .S(n9420), .Z(
        n15345) );
  XNOR2_X1 U16474 ( .A(n15346), .B(n15345), .ZN(n15347) );
  INV_X1 U16475 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15361) );
  INV_X1 U16476 ( .A(n15349), .ZN(n15350) );
  AOI211_X1 U16477 ( .C1(n15352), .C2(n15351), .A(n15364), .B(n15350), .ZN(
        n15357) );
  AOI211_X1 U16478 ( .C1(n15355), .C2(n15354), .A(n15368), .B(n15353), .ZN(
        n15356) );
  AOI211_X1 U16479 ( .C1(n15374), .C2(n15358), .A(n15357), .B(n15356), .ZN(
        n15360) );
  NAND2_X1 U16480 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n15359)
         );
  OAI211_X1 U16481 ( .C1(n15361), .C2(n15377), .A(n15360), .B(n15359), .ZN(
        P2_U3227) );
  INV_X1 U16482 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15515) );
  INV_X1 U16483 ( .A(n15362), .ZN(n15363) );
  AOI211_X1 U16484 ( .C1(n15366), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        n15372) );
  AOI211_X1 U16485 ( .C1(n15370), .C2(n15369), .A(n15368), .B(n15367), .ZN(
        n15371) );
  AOI211_X1 U16486 ( .C1(n15374), .C2(n15373), .A(n15372), .B(n15371), .ZN(
        n15376) );
  NAND2_X1 U16487 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n15375)
         );
  OAI211_X1 U16488 ( .C1(n15515), .C2(n15377), .A(n15376), .B(n15375), .ZN(
        P2_U3224) );
  OAI21_X1 U16489 ( .B1(n15379), .B2(P1_REG1_REG_0__SCAN_IN), .A(n15378), .ZN(
        n15380) );
  XNOR2_X1 U16490 ( .A(n15380), .B(n7345), .ZN(n15384) );
  AOI22_X1 U16491 ( .A1(n15381), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15382) );
  OAI21_X1 U16492 ( .B1(n15384), .B2(n15383), .A(n15382), .ZN(P1_U3243) );
  INV_X1 U16493 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15586) );
  OAI211_X1 U16494 ( .C1(n15387), .C2(n15386), .A(n15385), .B(n15427), .ZN(
        n15388) );
  INV_X1 U16495 ( .A(n15388), .ZN(n15393) );
  AOI211_X1 U16496 ( .C1(n15391), .C2(n15390), .A(n15413), .B(n15389), .ZN(
        n15392) );
  AOI211_X1 U16497 ( .C1(n15423), .C2(n15394), .A(n15393), .B(n15392), .ZN(
        n15395) );
  NAND2_X1 U16498 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3086), .ZN(n16028)
         );
  OAI211_X1 U16499 ( .C1(n15586), .C2(n15430), .A(n15395), .B(n16028), .ZN(
        P1_U3260) );
  INV_X1 U16500 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15407) );
  AOI211_X1 U16501 ( .C1(n15399), .C2(n15398), .A(n15397), .B(n15396), .ZN(
        n15403) );
  AOI211_X1 U16502 ( .C1(n15020), .C2(n15401), .A(n15413), .B(n15400), .ZN(
        n15402) );
  AOI211_X1 U16503 ( .C1(n15423), .C2(n15404), .A(n15403), .B(n15402), .ZN(
        n15406) );
  OAI211_X1 U16504 ( .C1(n15407), .C2(n15430), .A(n15406), .B(n15405), .ZN(
        P1_U3261) );
  INV_X1 U16505 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15573) );
  OAI211_X1 U16506 ( .C1(n15410), .C2(n15409), .A(n15408), .B(n15427), .ZN(
        n15411) );
  INV_X1 U16507 ( .A(n15411), .ZN(n15417) );
  AOI211_X1 U16508 ( .C1(n15415), .C2(n15414), .A(n15413), .B(n15412), .ZN(
        n15416) );
  AOI211_X1 U16509 ( .C1(n15423), .C2(n15418), .A(n15417), .B(n15416), .ZN(
        n15419) );
  NAND2_X1 U16510 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n16013)
         );
  OAI211_X1 U16511 ( .C1(n15573), .C2(n15430), .A(n15419), .B(n16013), .ZN(
        P1_U3259) );
  INV_X1 U16512 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15431) );
  OAI21_X1 U16513 ( .B1(n15421), .B2(n16000), .A(n15420), .ZN(n15428) );
  XNOR2_X1 U16514 ( .A(n15422), .B(P1_REG2_REG_15__SCAN_IN), .ZN(n15425) );
  AOI222_X1 U16515 ( .A1(n15428), .A2(n15427), .B1(n15426), .B2(n15425), .C1(
        n15424), .C2(n15423), .ZN(n15429) );
  NAND2_X1 U16516 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15985)
         );
  OAI211_X1 U16517 ( .C1(n15431), .C2(n15430), .A(n15429), .B(n15985), .ZN(
        P1_U3258) );
  XOR2_X1 U16518 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15437), .Z(SUB_1596_U53) );
  INV_X1 U16519 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15434) );
  NAND2_X1 U16520 ( .A1(n15436), .A2(n15435), .ZN(n15433) );
  OAI21_X1 U16521 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n15434), .A(n15433), .ZN(
        n15444) );
  XNOR2_X1 U16522 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n15445) );
  XOR2_X1 U16523 ( .A(n15444), .B(n15445), .Z(n15441) );
  NAND2_X1 U16524 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15437), .ZN(n15607) );
  NAND2_X1 U16525 ( .A1(n15608), .A2(n15607), .ZN(n15438) );
  NOR2_X1 U16526 ( .A1(n15608), .A2(n15607), .ZN(n15606) );
  NAND2_X1 U16527 ( .A1(n15441), .A2(n15440), .ZN(n15442) );
  OAI21_X1 U16528 ( .B1(n15441), .B2(n15440), .A(n15442), .ZN(n15439) );
  XNOR2_X1 U16529 ( .A(n15439), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  NOR2_X1 U16530 ( .A1(n15441), .A2(n15440), .ZN(n15443) );
  OAI21_X1 U16531 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n15443), .A(n15442), .ZN(
        n15456) );
  NAND2_X1 U16532 ( .A1(n15445), .A2(n15444), .ZN(n15446) );
  XNOR2_X1 U16533 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n15452), .ZN(n15457) );
  XOR2_X1 U16534 ( .A(n15456), .B(n15457), .Z(n15449) );
  NAND2_X1 U16535 ( .A1(n15449), .A2(n15448), .ZN(n15458) );
  OAI21_X1 U16536 ( .B1(n15449), .B2(n15448), .A(n15458), .ZN(SUB_1596_U60) );
  NAND2_X1 U16537 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15450), .ZN(n15454) );
  NAND2_X1 U16538 ( .A1(n15452), .A2(n15451), .ZN(n15453) );
  NAND2_X1 U16539 ( .A1(n15454), .A2(n15453), .ZN(n15463) );
  XNOR2_X1 U16540 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P3_ADDR_REG_4__SCAN_IN), 
        .ZN(n15455) );
  XOR2_X1 U16541 ( .A(n15463), .B(n15455), .Z(n15466) );
  XNOR2_X1 U16542 ( .A(n15466), .B(n15465), .ZN(n15461) );
  NAND2_X1 U16543 ( .A1(n15457), .A2(n15456), .ZN(n15459) );
  NAND2_X1 U16544 ( .A1(n15459), .A2(n15458), .ZN(n15460) );
  NOR2_X1 U16545 ( .A1(n15461), .A2(n15460), .ZN(n15467) );
  AOI21_X1 U16546 ( .B1(n15461), .B2(n15460), .A(n15467), .ZN(SUB_1596_U59) );
  XNOR2_X1 U16547 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n15464) );
  XNOR2_X1 U16548 ( .A(n15464), .B(n15478), .ZN(n15471) );
  NOR2_X1 U16549 ( .A1(n15466), .A2(n15465), .ZN(n15468) );
  XNOR2_X1 U16550 ( .A(n15471), .B(n15472), .ZN(n15470) );
  NOR2_X1 U16551 ( .A1(n15470), .A2(n15469), .ZN(n15473) );
  AOI21_X1 U16552 ( .B1(n15470), .B2(n15469), .A(n15473), .ZN(SUB_1596_U58) );
  NOR2_X1 U16553 ( .A1(n15472), .A2(n15471), .ZN(n15474) );
  XNOR2_X1 U16554 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n15479) );
  NAND2_X1 U16555 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n15475), .ZN(n15477) );
  XOR2_X1 U16556 ( .A(n15479), .B(n15481), .Z(n15603) );
  NAND2_X1 U16557 ( .A1(n15604), .A2(n15603), .ZN(n15602) );
  AND2_X1 U16558 ( .A1(n15480), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n15482) );
  XOR2_X1 U16559 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n15486), .Z(n15487) );
  XNOR2_X1 U16560 ( .A(n15483), .B(n15487), .ZN(n15484) );
  NAND2_X1 U16561 ( .A1(n15485), .A2(n15484), .ZN(n15492) );
  OAI21_X1 U16562 ( .B1(n15485), .B2(n15484), .A(n15492), .ZN(SUB_1596_U56) );
  XNOR2_X1 U16563 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n15496) );
  INV_X1 U16564 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15628) );
  NOR2_X1 U16565 ( .A1(n15628), .A2(n15486), .ZN(n15489) );
  NOR2_X1 U16566 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n15487), .ZN(n15488) );
  XNOR2_X1 U16567 ( .A(n15496), .B(n15495), .ZN(n15500) );
  NAND2_X1 U16568 ( .A1(n15491), .A2(n15490), .ZN(n15493) );
  NAND2_X1 U16569 ( .A1(n15493), .A2(n15492), .ZN(n15499) );
  NAND2_X1 U16570 ( .A1(n15500), .A2(n15499), .ZN(n15501) );
  OAI21_X1 U16571 ( .B1(n15500), .B2(n15499), .A(n15501), .ZN(n15494) );
  XNOR2_X1 U16572 ( .A(n15494), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  NAND2_X1 U16573 ( .A1(n15496), .A2(n15495), .ZN(n15497) );
  XOR2_X1 U16574 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n15510), .Z(n15508) );
  XNOR2_X1 U16575 ( .A(n15507), .B(n15508), .ZN(n15505) );
  NOR2_X1 U16576 ( .A1(n15500), .A2(n15499), .ZN(n15502) );
  OAI21_X1 U16577 ( .B1(n15505), .B2(n15504), .A(n15506), .ZN(n15503) );
  XNOR2_X1 U16578 ( .A(n15503), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  NAND2_X1 U16579 ( .A1(n15508), .A2(n15507), .ZN(n15509) );
  XOR2_X1 U16580 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n15516) );
  XNOR2_X1 U16581 ( .A(n15517), .B(n15516), .ZN(n15512) );
  NAND2_X1 U16582 ( .A1(n15511), .A2(n15512), .ZN(n15514) );
  INV_X1 U16583 ( .A(n15513), .ZN(n15522) );
  NAND2_X1 U16584 ( .A1(n15515), .A2(n15514), .ZN(n15521) );
  OAI222_X1 U16585 ( .A1(n15515), .A2(n15514), .B1(n15515), .B2(n15522), .C1(
        n15513), .C2(n15521), .ZN(SUB_1596_U70) );
  XNOR2_X1 U16586 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n15520) );
  XNOR2_X1 U16587 ( .A(n15520), .B(n15531), .ZN(n15525) );
  NAND2_X1 U16588 ( .A1(n15522), .A2(n15521), .ZN(n15524) );
  NOR2_X1 U16589 ( .A1(n15525), .A2(n15524), .ZN(n15526) );
  AOI21_X1 U16590 ( .B1(n15525), .B2(n15524), .A(n15526), .ZN(n15523) );
  XOR2_X1 U16591 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15523), .Z(SUB_1596_U69)
         );
  NAND2_X1 U16592 ( .A1(n15525), .A2(n15524), .ZN(n15527) );
  XNOR2_X1 U16593 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n15540) );
  NAND2_X1 U16594 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n15528), .ZN(n15530) );
  INV_X1 U16595 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15529) );
  XOR2_X1 U16596 ( .A(n15540), .B(n15539), .Z(n15534) );
  INV_X1 U16597 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15532) );
  OAI21_X1 U16598 ( .B1(n15533), .B2(n15532), .A(n15536), .ZN(SUB_1596_U68) );
  NAND2_X1 U16599 ( .A1(n15535), .A2(n15534), .ZN(n15537) );
  INV_X1 U16600 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15551) );
  INV_X1 U16601 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15538) );
  XOR2_X1 U16602 ( .A(n15551), .B(n15538), .Z(n15549) );
  INV_X1 U16603 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15542) );
  NAND2_X1 U16604 ( .A1(n15540), .A2(n15539), .ZN(n15541) );
  XNOR2_X1 U16605 ( .A(n15549), .B(n15548), .ZN(n15544) );
  NAND2_X1 U16606 ( .A1(n15545), .A2(n15544), .ZN(n15546) );
  OAI21_X1 U16607 ( .B1(n15545), .B2(n15544), .A(n15546), .ZN(n15543) );
  XNOR2_X1 U16608 ( .A(n15543), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  NOR2_X1 U16609 ( .A1(n15545), .A2(n15544), .ZN(n15547) );
  NOR2_X1 U16610 ( .A1(n15549), .A2(n15548), .ZN(n15550) );
  AOI21_X1 U16611 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n15551), .A(n15550), 
        .ZN(n15558) );
  XOR2_X1 U16612 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n15557) );
  XNOR2_X1 U16613 ( .A(n15558), .B(n15557), .ZN(n15553) );
  OAI21_X1 U16614 ( .B1(n15554), .B2(n15553), .A(n15555), .ZN(n15552) );
  XNOR2_X1 U16615 ( .A(n15552), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  INV_X1 U16616 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15565) );
  INV_X1 U16617 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15571) );
  NOR2_X1 U16618 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15571), .ZN(n15556) );
  AOI21_X1 U16619 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15571), .A(n15556), 
        .ZN(n15569) );
  INV_X1 U16620 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15560) );
  NOR2_X1 U16621 ( .A1(n15558), .A2(n15557), .ZN(n15559) );
  AOI21_X1 U16622 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n15560), .A(n15559), 
        .ZN(n15568) );
  XNOR2_X1 U16623 ( .A(n15569), .B(n15568), .ZN(n15562) );
  NAND2_X1 U16624 ( .A1(n15561), .A2(n15562), .ZN(n15564) );
  INV_X1 U16625 ( .A(n15563), .ZN(n15567) );
  NAND2_X1 U16626 ( .A1(n15565), .A2(n15564), .ZN(n15566) );
  OAI222_X1 U16627 ( .A1(n15565), .A2(n15564), .B1(n15565), .B2(n15567), .C1(
        n15563), .C2(n15566), .ZN(SUB_1596_U65) );
  NAND2_X1 U16628 ( .A1(n15569), .A2(n15568), .ZN(n15570) );
  XOR2_X1 U16629 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n15574), .Z(n15575) );
  XNOR2_X1 U16630 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n15575), .ZN(n15578) );
  NAND2_X1 U16631 ( .A1(n15579), .A2(n15578), .ZN(n15580) );
  OAI21_X1 U16632 ( .B1(n15579), .B2(n15578), .A(n15580), .ZN(n15572) );
  XNOR2_X1 U16633 ( .A(n15572), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NOR2_X1 U16634 ( .A1(n15574), .A2(n15573), .ZN(n15577) );
  NOR2_X1 U16635 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15575), .ZN(n15576) );
  NOR2_X1 U16636 ( .A1(n15577), .A2(n15576), .ZN(n15587) );
  XNOR2_X1 U16637 ( .A(n15586), .B(n15587), .ZN(n15588) );
  XOR2_X1 U16638 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n15588), .Z(n15583) );
  XNOR2_X1 U16639 ( .A(n15583), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(n15582) );
  AOI21_X1 U16640 ( .B1(n15582), .B2(n15581), .A(n15584), .ZN(SUB_1596_U63) );
  AND2_X1 U16641 ( .A1(n15583), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n15585) );
  NOR2_X1 U16642 ( .A1(n15587), .A2(n15586), .ZN(n15590) );
  NOR2_X1 U16643 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n15588), .ZN(n15589) );
  NOR2_X1 U16644 ( .A1(n15590), .A2(n15589), .ZN(n15598) );
  NAND2_X1 U16645 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15600), .ZN(n15591) );
  OAI21_X1 U16646 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15600), .A(n15591), 
        .ZN(n15597) );
  XNOR2_X1 U16647 ( .A(n15598), .B(n15597), .ZN(n15593) );
  NOR2_X1 U16648 ( .A1(n15594), .A2(n15593), .ZN(n15595) );
  AOI21_X1 U16649 ( .B1(n15594), .B2(n15593), .A(n15595), .ZN(n15592) );
  XOR2_X1 U16650 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n15592), .Z(SUB_1596_U62)
         );
  NAND2_X1 U16651 ( .A1(n15594), .A2(n15593), .ZN(n15596) );
  NOR2_X1 U16652 ( .A1(n15598), .A2(n15597), .ZN(n15599) );
  AOI21_X1 U16653 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15600), .A(n15599), 
        .ZN(n15601) );
  OAI21_X1 U16654 ( .B1(n15604), .B2(n15603), .A(n15602), .ZN(n15605) );
  XNOR2_X1 U16655 ( .A(n15605), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(SUB_1596_U57)
         );
  AOI21_X1 U16656 ( .B1(n15608), .B2(n15607), .A(n15606), .ZN(n15609) );
  XOR2_X1 U16657 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n15609), .Z(SUB_1596_U5) );
  AOI21_X1 U16658 ( .B1(n15612), .B2(n15611), .A(n15610), .ZN(n15620) );
  OAI21_X1 U16659 ( .B1(n15615), .B2(n15614), .A(n15613), .ZN(n15616) );
  AOI22_X1 U16660 ( .A1(n15618), .A2(n15617), .B1(n15616), .B2(n15638), .ZN(
        n15619) );
  OAI21_X1 U16661 ( .B1(n15620), .B2(n15636), .A(n15619), .ZN(n15625) );
  AOI21_X1 U16662 ( .B1(n15822), .B2(n15622), .A(n15621), .ZN(n15623) );
  NOR2_X1 U16663 ( .A1(n15623), .A2(n15631), .ZN(n15624) );
  NOR2_X1 U16664 ( .A1(n15625), .A2(n15624), .ZN(n15627) );
  OAI211_X1 U16665 ( .C1(n15628), .C2(n15651), .A(n15627), .B(n15626), .ZN(
        P3_U3189) );
  INV_X1 U16666 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15652) );
  AOI21_X1 U16667 ( .B1(n12162), .B2(n15630), .A(n15629), .ZN(n15632) );
  NOR2_X1 U16668 ( .A1(n15632), .A2(n15631), .ZN(n15647) );
  AOI21_X1 U16669 ( .B1(n15635), .B2(n15634), .A(n15633), .ZN(n15637) );
  NOR2_X1 U16670 ( .A1(n15637), .A2(n15636), .ZN(n15646) );
  OAI21_X1 U16671 ( .B1(n15640), .B2(n15639), .A(n15638), .ZN(n15644) );
  OAI22_X1 U16672 ( .A1(n15644), .A2(n15643), .B1(n15642), .B2(n15641), .ZN(
        n15645) );
  NOR3_X1 U16673 ( .A1(n15647), .A2(n15646), .A3(n15645), .ZN(n15650) );
  INV_X1 U16674 ( .A(n15648), .ZN(n15649) );
  OAI211_X1 U16675 ( .C1(n15652), .C2(n15651), .A(n15650), .B(n15649), .ZN(
        P3_U3191) );
  OAI221_X1 U16677 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n7677), .C2(n8274), .A(n15653), .ZN(U29) );
  AOI22_X1 U16678 ( .A1(n16005), .A2(n15655), .B1(n9716), .B2(n16002), .ZN(
        P1_U3459) );
  INV_X1 U16679 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n15659) );
  NAND2_X1 U16680 ( .A1(n15657), .A2(n15656), .ZN(n15658) );
  OAI21_X1 U16681 ( .B1(n15660), .B2(n15659), .A(n15658), .ZN(n15662) );
  AOI211_X1 U16682 ( .C1(n15664), .C2(n15663), .A(n15662), .B(n15661), .ZN(
        n15665) );
  AOI22_X1 U16683 ( .A1(n15667), .A2(n15666), .B1(n15665), .B2(n15021), .ZN(
        P1_U3293) );
  OAI211_X1 U16684 ( .C1(n15670), .C2(n15990), .A(n15669), .B(n15668), .ZN(
        n15674) );
  NOR2_X1 U16685 ( .A1(n15672), .A2(n15671), .ZN(n15673) );
  AOI211_X1 U16686 ( .C1(n15912), .C2(n15675), .A(n15674), .B(n15673), .ZN(
        n15677) );
  AOI22_X1 U16687 ( .A1(n16001), .A2(n15677), .B1(n15676), .B2(n15999), .ZN(
        P1_U3529) );
  AOI22_X1 U16688 ( .A1(n16005), .A2(n15677), .B1(n9701), .B2(n16002), .ZN(
        P1_U3462) );
  OAI22_X1 U16689 ( .A1(n15679), .A2(n15858), .B1(n15886), .B2(n15678), .ZN(
        n15680) );
  NOR2_X1 U16690 ( .A1(n15681), .A2(n15680), .ZN(n15684) );
  AOI22_X1 U16691 ( .A1(n15894), .A2(n15684), .B1(n15682), .B2(n15892), .ZN(
        P3_U3461) );
  INV_X1 U16692 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15683) );
  AOI22_X1 U16693 ( .A1(n15898), .A2(n15684), .B1(n15683), .B2(n15895), .ZN(
        P3_U3396) );
  OAI21_X1 U16694 ( .B1(n15686), .B2(n15990), .A(n15685), .ZN(n15687) );
  AOI21_X1 U16695 ( .B1(n15688), .B2(n15912), .A(n15687), .ZN(n15689) );
  AND2_X1 U16696 ( .A1(n15690), .A2(n15689), .ZN(n15691) );
  AOI22_X1 U16697 ( .A1(n16001), .A2(n15691), .B1(n10863), .B2(n15999), .ZN(
        P1_U3530) );
  AOI22_X1 U16698 ( .A1(n16005), .A2(n15691), .B1(n9724), .B2(n16002), .ZN(
        P1_U3465) );
  OAI21_X1 U16699 ( .B1(n15698), .B2(n15693), .A(n15692), .ZN(n15712) );
  INV_X1 U16700 ( .A(n15959), .ZN(n15851) );
  OAI211_X1 U16701 ( .C1(n15708), .C2(n15695), .A(n7209), .B(n15694), .ZN(
        n15716) );
  OAI21_X1 U16702 ( .B1(n15708), .B2(n15851), .A(n15716), .ZN(n15704) );
  NAND3_X1 U16703 ( .A1(n15698), .A2(n15697), .A3(n15696), .ZN(n15700) );
  AND2_X1 U16704 ( .A1(n15700), .A2(n15699), .ZN(n15703) );
  OAI21_X1 U16705 ( .B1(n15703), .B2(n15702), .A(n15701), .ZN(n15710) );
  AOI211_X1 U16706 ( .C1(n15964), .C2(n15712), .A(n15704), .B(n15710), .ZN(
        n15706) );
  AOI22_X1 U16707 ( .A1(n15970), .A2(n15706), .B1(n10764), .B2(n15968), .ZN(
        P2_U3501) );
  INV_X1 U16708 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15705) );
  AOI22_X1 U16709 ( .A1(n15973), .A2(n15706), .B1(n15705), .B2(n15971), .ZN(
        P2_U3436) );
  INV_X1 U16710 ( .A(n15707), .ZN(n15709) );
  NOR2_X1 U16711 ( .A1(n15709), .A2(n15708), .ZN(n15711) );
  AOI211_X1 U16712 ( .C1(n15713), .C2(n15712), .A(n15711), .B(n15710), .ZN(
        n15722) );
  OAI22_X1 U16713 ( .A1(n15717), .A2(n15716), .B1(n15715), .B2(n15714), .ZN(
        n15718) );
  INV_X1 U16714 ( .A(n15718), .ZN(n15719) );
  OAI221_X1 U16715 ( .B1(n15947), .B2(n15722), .C1(n15721), .C2(n15720), .A(
        n15719), .ZN(P2_U3263) );
  NOR2_X1 U16716 ( .A1(n15723), .A2(n15886), .ZN(n15725) );
  AOI211_X1 U16717 ( .C1(n15873), .C2(n15726), .A(n15725), .B(n15724), .ZN(
        n15729) );
  AOI22_X1 U16718 ( .A1(n15894), .A2(n15729), .B1(n15727), .B2(n15892), .ZN(
        P3_U3462) );
  INV_X1 U16719 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15728) );
  AOI22_X1 U16720 ( .A1(n15898), .A2(n15729), .B1(n15728), .B2(n15895), .ZN(
        P3_U3399) );
  OAI22_X1 U16721 ( .A1(n15732), .A2(n15731), .B1(n15730), .B2(n15990), .ZN(
        n15734) );
  AOI211_X1 U16722 ( .C1(n15735), .C2(n15998), .A(n15734), .B(n15733), .ZN(
        n15736) );
  AOI22_X1 U16723 ( .A1(n16001), .A2(n15736), .B1(n10864), .B2(n15999), .ZN(
        P1_U3531) );
  AOI22_X1 U16724 ( .A1(n16005), .A2(n15736), .B1(n9696), .B2(n16002), .ZN(
        P1_U3468) );
  OAI22_X1 U16725 ( .A1(n15738), .A2(n15858), .B1(n15886), .B2(n15737), .ZN(
        n15740) );
  NOR2_X1 U16726 ( .A1(n15740), .A2(n15739), .ZN(n15743) );
  AOI22_X1 U16727 ( .A1(n15894), .A2(n15743), .B1(n15741), .B2(n15892), .ZN(
        P3_U3463) );
  INV_X1 U16728 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15742) );
  AOI22_X1 U16729 ( .A1(n15898), .A2(n15743), .B1(n15742), .B2(n15895), .ZN(
        P3_U3402) );
  OAI211_X1 U16730 ( .C1(n15746), .C2(n15990), .A(n15745), .B(n15744), .ZN(
        n15750) );
  NOR2_X1 U16731 ( .A1(n15748), .A2(n15747), .ZN(n15749) );
  AOI211_X1 U16732 ( .C1(n15751), .C2(n15998), .A(n15750), .B(n15749), .ZN(
        n15752) );
  AOI22_X1 U16733 ( .A1(n16001), .A2(n15752), .B1(n10865), .B2(n15999), .ZN(
        P1_U3532) );
  AOI22_X1 U16734 ( .A1(n16005), .A2(n15752), .B1(n9749), .B2(n16002), .ZN(
        P1_U3471) );
  OAI21_X1 U16735 ( .B1(n15754), .B2(n15851), .A(n15753), .ZN(n15756) );
  AOI211_X1 U16736 ( .C1(n15758), .C2(n15757), .A(n15756), .B(n15755), .ZN(
        n15760) );
  AOI22_X1 U16737 ( .A1(n15970), .A2(n15760), .B1(n10766), .B2(n15968), .ZN(
        P2_U3503) );
  INV_X1 U16738 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15759) );
  AOI22_X1 U16739 ( .A1(n15973), .A2(n15760), .B1(n15759), .B2(n15971), .ZN(
        P2_U3442) );
  AOI21_X1 U16740 ( .B1(n15872), .B2(n15762), .A(n15761), .ZN(n15763) );
  OAI21_X1 U16741 ( .B1(n15764), .B2(n15765), .A(n15763), .ZN(n15769) );
  INV_X1 U16742 ( .A(n15765), .ZN(n15770) );
  AOI22_X1 U16743 ( .A1(n15769), .A2(n15894), .B1(n15766), .B2(n15770), .ZN(
        n15767) );
  OAI21_X1 U16744 ( .B1(n15894), .B2(n15768), .A(n15767), .ZN(P3_U3464) );
  AOI21_X1 U16745 ( .B1(n15873), .B2(n15770), .A(n15769), .ZN(n15772) );
  INV_X1 U16746 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15771) );
  AOI22_X1 U16747 ( .A1(n15898), .A2(n15772), .B1(n15771), .B2(n15895), .ZN(
        P3_U3405) );
  NOR2_X1 U16748 ( .A1(n15774), .A2(n15773), .ZN(n15778) );
  NOR4_X1 U16749 ( .A1(n15778), .A2(n15777), .A3(n15776), .A4(n15775), .ZN(
        n15780) );
  AOI22_X1 U16750 ( .A1(n16001), .A2(n15780), .B1(n10866), .B2(n15999), .ZN(
        P1_U3533) );
  INV_X1 U16751 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15779) );
  AOI22_X1 U16752 ( .A1(n16005), .A2(n15780), .B1(n15779), .B2(n16002), .ZN(
        P1_U3474) );
  AOI22_X1 U16753 ( .A1(n15782), .A2(n15873), .B1(n15872), .B2(n15781), .ZN(
        n15783) );
  AND2_X1 U16754 ( .A1(n15784), .A2(n15783), .ZN(n15787) );
  AOI22_X1 U16755 ( .A1(n15894), .A2(n15787), .B1(n15785), .B2(n15892), .ZN(
        P3_U3465) );
  INV_X1 U16756 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15786) );
  AOI22_X1 U16757 ( .A1(n15898), .A2(n15787), .B1(n15786), .B2(n15895), .ZN(
        P3_U3408) );
  NAND2_X1 U16758 ( .A1(n15789), .A2(n15788), .ZN(n15791) );
  AOI211_X1 U16759 ( .C1(n15912), .C2(n15792), .A(n15791), .B(n15790), .ZN(
        n15793) );
  AOI22_X1 U16760 ( .A1(n16001), .A2(n15793), .B1(n10867), .B2(n15999), .ZN(
        P1_U3534) );
  AOI22_X1 U16761 ( .A1(n16005), .A2(n15793), .B1(n9687), .B2(n16002), .ZN(
        P1_U3477) );
  XNOR2_X1 U16762 ( .A(n15794), .B(n15795), .ZN(n15798) );
  AOI21_X1 U16763 ( .B1(n15798), .B2(n15797), .A(n15796), .ZN(n15812) );
  INV_X1 U16764 ( .A(n15799), .ZN(n15800) );
  AOI222_X1 U16765 ( .A1(n15801), .A2(n15917), .B1(P2_REG2_REG_6__SCAN_IN), 
        .B2(n15947), .C1(n15936), .C2(n15800), .ZN(n15809) );
  XNOR2_X1 U16766 ( .A(n15802), .B(n15803), .ZN(n15815) );
  OAI211_X1 U16767 ( .C1(n15805), .C2(n15811), .A(n7209), .B(n15804), .ZN(
        n15810) );
  INV_X1 U16768 ( .A(n15810), .ZN(n15806) );
  AOI22_X1 U16769 ( .A1(n15815), .A2(n15807), .B1(n15934), .B2(n15806), .ZN(
        n15808) );
  OAI211_X1 U16770 ( .C1(n15947), .C2(n15812), .A(n15809), .B(n15808), .ZN(
        P2_U3259) );
  OAI21_X1 U16771 ( .B1(n15811), .B2(n15851), .A(n15810), .ZN(n15814) );
  INV_X1 U16772 ( .A(n15812), .ZN(n15813) );
  AOI211_X1 U16773 ( .C1(n15815), .C2(n15964), .A(n15814), .B(n15813), .ZN(
        n15817) );
  AOI22_X1 U16774 ( .A1(n15970), .A2(n15817), .B1(n11264), .B2(n15968), .ZN(
        P2_U3505) );
  INV_X1 U16775 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15816) );
  AOI22_X1 U16776 ( .A1(n15973), .A2(n15817), .B1(n15816), .B2(n15971), .ZN(
        P2_U3448) );
  NOR2_X1 U16777 ( .A1(n15818), .A2(n15886), .ZN(n15820) );
  AOI211_X1 U16778 ( .C1(n15873), .C2(n15821), .A(n15820), .B(n15819), .ZN(
        n15824) );
  AOI22_X1 U16779 ( .A1(n15894), .A2(n15824), .B1(n15822), .B2(n15892), .ZN(
        P3_U3466) );
  INV_X1 U16780 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15823) );
  AOI22_X1 U16781 ( .A1(n15898), .A2(n15824), .B1(n15823), .B2(n15895), .ZN(
        P3_U3411) );
  OAI21_X1 U16782 ( .B1(n7583), .B2(n15990), .A(n15825), .ZN(n15827) );
  AOI211_X1 U16783 ( .C1(n15912), .C2(n15828), .A(n15827), .B(n15826), .ZN(
        n15830) );
  AOI22_X1 U16784 ( .A1(n16001), .A2(n15830), .B1(n10868), .B2(n15999), .ZN(
        P1_U3535) );
  INV_X1 U16785 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15829) );
  AOI22_X1 U16786 ( .A1(n16005), .A2(n15830), .B1(n15829), .B2(n16002), .ZN(
        P1_U3480) );
  AND2_X1 U16787 ( .A1(n15831), .A2(n15959), .ZN(n15832) );
  NOR2_X1 U16788 ( .A1(n15833), .A2(n15832), .ZN(n15837) );
  OR2_X1 U16789 ( .A1(n15835), .A2(n15834), .ZN(n15836) );
  AND3_X1 U16790 ( .A1(n15838), .A2(n15837), .A3(n15836), .ZN(n15840) );
  AOI22_X1 U16791 ( .A1(n15970), .A2(n15840), .B1(n11265), .B2(n15968), .ZN(
        P2_U3506) );
  INV_X1 U16792 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15839) );
  AOI22_X1 U16793 ( .A1(n15973), .A2(n15840), .B1(n15839), .B2(n15971), .ZN(
        P2_U3451) );
  AOI22_X1 U16794 ( .A1(n15842), .A2(n15873), .B1(n15872), .B2(n15841), .ZN(
        n15843) );
  AND2_X1 U16795 ( .A1(n15844), .A2(n15843), .ZN(n15846) );
  AOI22_X1 U16796 ( .A1(n15894), .A2(n15846), .B1(n11772), .B2(n15892), .ZN(
        P3_U3467) );
  INV_X1 U16797 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15845) );
  AOI22_X1 U16798 ( .A1(n15898), .A2(n15846), .B1(n15845), .B2(n15895), .ZN(
        P3_U3414) );
  NAND3_X1 U16799 ( .A1(n15848), .A2(n15847), .A3(n15964), .ZN(n15850) );
  OAI211_X1 U16800 ( .C1(n15852), .C2(n15851), .A(n15850), .B(n15849), .ZN(
        n15853) );
  NOR2_X1 U16801 ( .A1(n15854), .A2(n15853), .ZN(n15856) );
  AOI22_X1 U16802 ( .A1(n15970), .A2(n15856), .B1(n11266), .B2(n15968), .ZN(
        P2_U3507) );
  INV_X1 U16803 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15855) );
  AOI22_X1 U16804 ( .A1(n15973), .A2(n15856), .B1(n15855), .B2(n15971), .ZN(
        P2_U3454) );
  OAI22_X1 U16805 ( .A1(n15859), .A2(n15858), .B1(n15886), .B2(n15857), .ZN(
        n15860) );
  NOR2_X1 U16806 ( .A1(n15861), .A2(n15860), .ZN(n15863) );
  AOI22_X1 U16807 ( .A1(n15894), .A2(n15863), .B1(n12162), .B2(n15892), .ZN(
        P3_U3468) );
  INV_X1 U16808 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15862) );
  AOI22_X1 U16809 ( .A1(n15898), .A2(n15863), .B1(n15862), .B2(n15895), .ZN(
        P3_U3417) );
  OAI21_X1 U16810 ( .B1(n15865), .B2(n15990), .A(n15864), .ZN(n15867) );
  AOI211_X1 U16811 ( .C1(n15912), .C2(n15868), .A(n15867), .B(n15866), .ZN(
        n15870) );
  AOI22_X1 U16812 ( .A1(n16001), .A2(n15870), .B1(n10969), .B2(n15999), .ZN(
        P1_U3537) );
  INV_X1 U16813 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15869) );
  AOI22_X1 U16814 ( .A1(n16005), .A2(n15870), .B1(n15869), .B2(n16002), .ZN(
        P1_U3486) );
  AOI22_X1 U16815 ( .A1(n15874), .A2(n15873), .B1(n15872), .B2(n15871), .ZN(
        n15875) );
  AOI22_X1 U16816 ( .A1(n15894), .A2(n15878), .B1(n12180), .B2(n15892), .ZN(
        P3_U3469) );
  INV_X1 U16817 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15877) );
  AOI22_X1 U16818 ( .A1(n15898), .A2(n15878), .B1(n15877), .B2(n15895), .ZN(
        P3_U3420) );
  OAI21_X1 U16819 ( .B1(n15880), .B2(n15990), .A(n15879), .ZN(n15882) );
  AOI211_X1 U16820 ( .C1(n15998), .C2(n15883), .A(n15882), .B(n15881), .ZN(
        n15885) );
  AOI22_X1 U16821 ( .A1(n16001), .A2(n15885), .B1(n10970), .B2(n15999), .ZN(
        P1_U3538) );
  INV_X1 U16822 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15884) );
  AOI22_X1 U16823 ( .A1(n16005), .A2(n15885), .B1(n15884), .B2(n16002), .ZN(
        P1_U3489) );
  NOR2_X1 U16824 ( .A1(n15887), .A2(n15886), .ZN(n15889) );
  AOI211_X1 U16825 ( .C1(n15891), .C2(n15890), .A(n15889), .B(n15888), .ZN(
        n15897) );
  AOI22_X1 U16826 ( .A1(n15894), .A2(n15897), .B1(n15893), .B2(n15892), .ZN(
        P3_U3470) );
  INV_X1 U16827 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15896) );
  AOI22_X1 U16828 ( .A1(n15898), .A2(n15897), .B1(n15896), .B2(n15895), .ZN(
        P3_U3423) );
  AOI21_X1 U16829 ( .B1(n15949), .B2(n15900), .A(n15899), .ZN(n15901) );
  OAI211_X1 U16830 ( .C1(n15953), .C2(n15903), .A(n15902), .B(n15901), .ZN(
        n15904) );
  INV_X1 U16831 ( .A(n15904), .ZN(n15906) );
  AOI22_X1 U16832 ( .A1(n16001), .A2(n15906), .B1(n11456), .B2(n15999), .ZN(
        P1_U3539) );
  INV_X1 U16833 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15905) );
  AOI22_X1 U16834 ( .A1(n16005), .A2(n15906), .B1(n15905), .B2(n16002), .ZN(
        P1_U3492) );
  INV_X1 U16835 ( .A(n15907), .ZN(n15911) );
  OAI21_X1 U16836 ( .B1(n7584), .B2(n15990), .A(n15908), .ZN(n15910) );
  AOI211_X1 U16837 ( .C1(n15912), .C2(n15911), .A(n15910), .B(n15909), .ZN(
        n15914) );
  AOI22_X1 U16838 ( .A1(n16001), .A2(n15914), .B1(n11885), .B2(n15999), .ZN(
        P1_U3540) );
  INV_X1 U16839 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n15913) );
  AOI22_X1 U16840 ( .A1(n16005), .A2(n15914), .B1(n15913), .B2(n16002), .ZN(
        P1_U3495) );
  INV_X1 U16841 ( .A(n15915), .ZN(n15916) );
  AOI222_X1 U16842 ( .A1(n15918), .A2(n15917), .B1(P2_REG2_REG_12__SCAN_IN), 
        .B2(n15947), .C1(n15936), .C2(n15916), .ZN(n15922) );
  AOI22_X1 U16843 ( .A1(n15920), .A2(n15934), .B1(n15944), .B2(n15919), .ZN(
        n15921) );
  OAI211_X1 U16844 ( .C1(n15947), .C2(n15923), .A(n15922), .B(n15921), .ZN(
        P2_U3253) );
  OAI211_X1 U16845 ( .C1(n15926), .C2(n15990), .A(n15925), .B(n15924), .ZN(
        n15929) );
  NOR2_X1 U16846 ( .A1(n15927), .A2(n15953), .ZN(n15928) );
  AOI211_X1 U16847 ( .C1(n15930), .C2(n15993), .A(n15929), .B(n15928), .ZN(
        n15933) );
  AOI22_X1 U16848 ( .A1(n16001), .A2(n15933), .B1(n15931), .B2(n15999), .ZN(
        P1_U3541) );
  INV_X1 U16849 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15932) );
  AOI22_X1 U16850 ( .A1(n16005), .A2(n15933), .B1(n15932), .B2(n16002), .ZN(
        P1_U3498) );
  NAND2_X1 U16851 ( .A1(n15935), .A2(n15934), .ZN(n15939) );
  AOI22_X1 U16852 ( .A1(n15947), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n15937), 
        .B2(n15936), .ZN(n15938) );
  OAI211_X1 U16853 ( .C1(n15941), .C2(n15940), .A(n15939), .B(n15938), .ZN(
        n15942) );
  AOI21_X1 U16854 ( .B1(n15944), .B2(n15943), .A(n15942), .ZN(n15945) );
  OAI21_X1 U16855 ( .B1(n15947), .B2(n15946), .A(n15945), .ZN(P2_U3252) );
  AOI21_X1 U16856 ( .B1(n15950), .B2(n15949), .A(n15948), .ZN(n15952) );
  OAI211_X1 U16857 ( .C1(n15954), .C2(n15953), .A(n15952), .B(n15951), .ZN(
        n15955) );
  AOI21_X1 U16858 ( .B1(n15956), .B2(n15993), .A(n15955), .ZN(n15958) );
  AOI22_X1 U16859 ( .A1(n16001), .A2(n15958), .B1(n9787), .B2(n15999), .ZN(
        P1_U3542) );
  INV_X1 U16860 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15957) );
  AOI22_X1 U16861 ( .A1(n16005), .A2(n15958), .B1(n15957), .B2(n16002), .ZN(
        P1_U3501) );
  NAND2_X1 U16862 ( .A1(n15960), .A2(n15959), .ZN(n15961) );
  NAND2_X1 U16863 ( .A1(n15962), .A2(n15961), .ZN(n15963) );
  AOI21_X1 U16864 ( .B1(n15965), .B2(n15964), .A(n15963), .ZN(n15966) );
  AOI22_X1 U16865 ( .A1(n15970), .A2(n15972), .B1(n15969), .B2(n15968), .ZN(
        P2_U3514) );
  AOI22_X1 U16866 ( .A1(n15973), .A2(n15972), .B1(n9186), .B2(n15971), .ZN(
        P2_U3475) );
  OAI21_X1 U16867 ( .B1(n15976), .B2(n15975), .A(n15974), .ZN(n15984) );
  AOI22_X1 U16868 ( .A1(n15980), .A2(n15979), .B1(n15978), .B2(n15977), .ZN(
        n15981) );
  OAI21_X1 U16869 ( .B1(n15991), .B2(n15982), .A(n15981), .ZN(n15983) );
  AOI21_X1 U16870 ( .B1(n15984), .B2(n16010), .A(n15983), .ZN(n15986) );
  OAI211_X1 U16871 ( .C1(n16031), .C2(n15987), .A(n15986), .B(n15985), .ZN(
        P1_U3241) );
  OAI211_X1 U16872 ( .C1(n15991), .C2(n15990), .A(n15989), .B(n15988), .ZN(
        n15996) );
  AND3_X1 U16873 ( .A1(n15994), .A2(n15993), .A3(n15992), .ZN(n15995) );
  AOI211_X1 U16874 ( .C1(n15998), .C2(n15997), .A(n15996), .B(n15995), .ZN(
        n16004) );
  AOI22_X1 U16875 ( .A1(n16001), .A2(n16004), .B1(n16000), .B2(n15999), .ZN(
        P1_U3543) );
  INV_X1 U16876 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n16003) );
  AOI22_X1 U16877 ( .A1(n16005), .A2(n16004), .B1(n16003), .B2(n16002), .ZN(
        P1_U3504) );
  XNOR2_X1 U16878 ( .A(n16006), .B(n16007), .ZN(n16009) );
  AOI222_X1 U16879 ( .A1(n16012), .A2(n16011), .B1(n16010), .B2(n16009), .C1(
        n16008), .C2(n16027), .ZN(n16014) );
  OAI211_X1 U16880 ( .C1(n16031), .C2(n16015), .A(n16014), .B(n16013), .ZN(
        P1_U3226) );
  OAI22_X1 U16881 ( .A1(n16019), .A2(n16018), .B1(n16017), .B2(n16016), .ZN(
        n16025) );
  XOR2_X1 U16882 ( .A(n16021), .B(n16020), .Z(n16023) );
  NOR2_X1 U16883 ( .A1(n16023), .A2(n16022), .ZN(n16024) );
  AOI211_X1 U16884 ( .C1(n16027), .C2(n16026), .A(n16025), .B(n16024), .ZN(
        n16029) );
  OAI211_X1 U16885 ( .C1(n16031), .C2(n16030), .A(n16029), .B(n16028), .ZN(
        P1_U3228) );
  AOI21_X1 U16886 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16032) );
  OAI21_X1 U16887 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16032), 
        .ZN(U28) );
  CLKBUF_X2 U7323 ( .A(n9003), .Z(n7168) );
  BUF_X2 U9865 ( .A(n12999), .Z(n13019) );
  INV_X1 U7277 ( .A(n14192), .ZN(n11104) );
  CLKBUF_X1 U7285 ( .A(n13789), .Z(n7166) );
  CLKBUF_X2 U7296 ( .A(n9003), .Z(n7169) );
  CLKBUF_X1 U7347 ( .A(n10770), .Z(n7526) );
endmodule

