

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1,
         READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786,
         n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
         n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
         n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
         n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
         n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
         n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
         n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
         n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
         n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882,
         n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
         n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954,
         n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
         n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
         n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
         n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
         n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
         n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002,
         n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010,
         n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
         n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026,
         n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
         n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
         n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
         n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
         n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066,
         n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074,
         n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
         n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
         n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098,
         n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122,
         n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
         n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138,
         n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146,
         n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
         n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
         n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170,
         n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
         n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
         n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194,
         n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
         n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
         n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
         n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
         n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
         n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242,
         n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
         n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
         n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266,
         n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
         n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
         n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
         n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
         n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
         n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314,
         n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
         n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
         n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338,
         n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
         n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
         n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
         n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
         n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
         n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386,
         n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
         n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
         n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
         n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
         n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
         n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
         n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
         n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
         n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
         n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
         n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
         n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
         n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
         n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
         n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
         n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
         n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
         n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
         n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
         n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
         n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
         n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
         n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
         n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
         n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602,
         n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
         n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
         n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626,
         n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
         n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
         n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
         n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658,
         n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
         n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
         n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
         n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
         n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698,
         n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
         n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714,
         n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722,
         n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
         n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
         n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746,
         n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754,
         n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
         n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770,
         n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778,
         n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786,
         n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794,
         n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
         n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
         n22811, n22812, n22813, n22814;

  OR2_X1 U11264 ( .A1(n17316), .A2(n11497), .ZN(n17516) );
  NOR2_X1 U11265 ( .A1(n18638), .A2(n18639), .ZN(n18607) );
  INV_X2 U11266 ( .A(n18832), .ZN(n18820) );
  NOR2_X1 U11267 ( .A1(n21792), .A2(n20639), .ZN(n20682) );
  OAI21_X1 U11268 ( .B1(n15285), .B2(n12203), .A(n12199), .ZN(n14889) );
  INV_X1 U11269 ( .A(n18640), .ZN(n21649) );
  AND4_X1 U11270 ( .A1(n14096), .A2(n14097), .A3(n14095), .A4(n14112), .ZN(
        n11480) );
  XNOR2_X1 U11271 ( .A(n12164), .B(n12163), .ZN(n12854) );
  AND2_X1 U11272 ( .A1(n14109), .A2(n14108), .ZN(n14164) );
  AND2_X1 U11273 ( .A1(n14109), .A2(n14105), .ZN(n14160) );
  NAND2_X1 U11274 ( .A1(n19589), .A2(n21179), .ZN(n15992) );
  INV_X2 U11275 ( .A(n21219), .ZN(n21179) );
  BUF_X1 U11276 ( .A(n14986), .Z(n18048) );
  CLKBUF_X1 U11277 ( .A(n15058), .Z(n11175) );
  CLKBUF_X2 U11278 ( .A(n12032), .Z(n12627) );
  CLKBUF_X1 U11279 ( .A(n12048), .Z(n12637) );
  CLKBUF_X2 U11280 ( .A(n16234), .Z(n11159) );
  INV_X1 U11281 ( .A(n11852), .ZN(n18347) );
  INV_X1 U11282 ( .A(n18099), .ZN(n18371) );
  AND2_X2 U11283 ( .A1(n16397), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16211) );
  BUF_X2 U11284 ( .A(n14985), .Z(n18320) );
  INV_X1 U11285 ( .A(n18099), .ZN(n18323) );
  BUF_X2 U11286 ( .A(n14986), .Z(n11170) );
  AND2_X1 U11287 ( .A1(n16249), .A2(n13329), .ZN(n16240) );
  AND2_X1 U11288 ( .A1(n13328), .A2(n16249), .ZN(n16242) );
  CLKBUF_X2 U11289 ( .A(n13064), .Z(n14878) );
  INV_X1 U11290 ( .A(n14405), .ZN(n14257) );
  INV_X1 U11291 ( .A(n13104), .ZN(n13114) );
  AND2_X1 U11292 ( .A1(n15090), .A2(n16896), .ZN(n12015) );
  AND2_X1 U11293 ( .A1(n11801), .A2(n16896), .ZN(n12067) );
  AND2_X1 U11294 ( .A1(n11866), .A2(n15098), .ZN(n12048) );
  AND2_X1 U11295 ( .A1(n11866), .A2(n11868), .ZN(n11907) );
  AND2_X1 U11296 ( .A1(n11775), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15090) );
  AND2_X1 U11297 ( .A1(n14797), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11866) );
  NAND3_X1 U11298 ( .A1(n14219), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16374) );
  INV_X2 U11299 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14219) );
  CLKBUF_X1 U11300 ( .A(n20982), .Z(n11157) );
  NOR4_X1 U11301 ( .A1(n21537), .A2(n20682), .A3(n21056), .A4(n21837), .ZN(
        n20982) );
  AND2_X1 U11302 ( .A1(n13328), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11162) );
  NOR2_X2 U11303 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11868) );
  NAND2_X1 U11304 ( .A1(n11560), .A2(n20178), .ZN(n11559) );
  INV_X1 U11305 ( .A(n14178), .ZN(n14203) );
  INV_X1 U11306 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15226) );
  AND2_X1 U11307 ( .A1(n15090), .A2(n15076), .ZN(n12032) );
  AND2_X2 U11308 ( .A1(n13328), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13042) );
  CLKBUF_X3 U11309 ( .A(n16400), .Z(n16384) );
  AND2_X1 U11310 ( .A1(n13330), .A2(n16249), .ZN(n13368) );
  OAI21_X1 U11311 ( .B1(n11583), .B2(n11582), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U11313 ( .A1(n21342), .A2(n21361), .ZN(n14966) );
  AND2_X1 U11314 ( .A1(n11964), .A2(n14540), .ZN(n14558) );
  XNOR2_X1 U11316 ( .A(n11988), .B(n12003), .ZN(n12030) );
  NAND2_X1 U11317 ( .A1(n12076), .A2(n12075), .ZN(n12177) );
  NAND2_X1 U11318 ( .A1(n11581), .A2(n11579), .ZN(n13104) );
  INV_X1 U11319 ( .A(n13619), .ZN(n13624) );
  OR2_X1 U11320 ( .A1(n13158), .A2(n13157), .ZN(n13160) );
  AND2_X1 U11321 ( .A1(n14109), .A2(n14103), .ZN(n14161) );
  NAND2_X2 U11322 ( .A1(n21324), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14967) );
  OR2_X2 U11323 ( .A1(n11884), .A2(n11883), .ZN(n16595) );
  INV_X2 U11324 ( .A(n11861), .ZN(n20552) );
  INV_X1 U11325 ( .A(n12752), .ZN(n15304) );
  INV_X2 U11326 ( .A(n16595), .ZN(n15592) );
  OR2_X1 U11328 ( .A1(n16366), .A2(n16365), .ZN(n11225) );
  AND2_X1 U11329 ( .A1(n13160), .A2(n13159), .ZN(n14086) );
  INV_X1 U11331 ( .A(n18346), .ZN(n17979) );
  AOI221_X1 U11332 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18524), 
        .C1(n21706), .C2(n18523), .A(n18522), .ZN(n18525) );
  INV_X1 U11333 ( .A(n22203), .ZN(n22187) );
  INV_X2 U11334 ( .A(n14764), .ZN(n15391) );
  OR2_X1 U11335 ( .A1(n15416), .A2(n15417), .ZN(n15702) );
  NAND2_X1 U11336 ( .A1(n15772), .A2(n15771), .ZN(n15870) );
  INV_X1 U11337 ( .A(n13110), .ZN(n13358) );
  OAI21_X1 U11338 ( .B1(n17285), .B2(n17283), .A(n17284), .ZN(n17275) );
  INV_X1 U11339 ( .A(n20980), .ZN(n20996) );
  NAND2_X1 U11340 ( .A1(n18639), .A2(n11598), .ZN(n21664) );
  AND2_X1 U11341 ( .A1(n21628), .A2(n20684), .ZN(n21788) );
  INV_X1 U11342 ( .A(n14808), .ZN(n14686) );
  INV_X1 U11343 ( .A(n18745), .ZN(n18682) );
  NAND2_X1 U11344 ( .A1(n20684), .A2(n21850), .ZN(n18832) );
  INV_X1 U11345 ( .A(n13109), .ZN(n19175) );
  AND2_X1 U11346 ( .A1(n11906), .A2(n11905), .ZN(n11158) );
  XNOR2_X1 U11347 ( .A(n14093), .B(n14092), .ZN(n15239) );
  INV_X2 U11348 ( .A(n17205), .ZN(n11477) );
  NOR2_X4 U11349 ( .A1(n15298), .A2(n15297), .ZN(n15299) );
  NAND2_X2 U11350 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21341) );
  NOR3_X2 U11352 ( .A1(n15982), .A2(n15981), .A3(n15980), .ZN(n15983) );
  NAND2_X2 U11353 ( .A1(n15990), .A2(n18395), .ZN(n15982) );
  AND4_X2 U11354 ( .A1(n14118), .A2(n14126), .A3(n14117), .A4(n14120), .ZN(
        n11482) );
  AND4_X2 U11355 ( .A1(n14113), .A2(n14111), .A3(n14094), .A4(n14110), .ZN(
        n11479) );
  AND2_X4 U11356 ( .A1(n13326), .A2(n15226), .ZN(n13027) );
  OAI22_X2 U11357 ( .A1(n17027), .A2(n17021), .B1(n11178), .B2(n16285), .ZN(
        n17015) );
  AND2_X2 U11358 ( .A1(n14107), .A2(n14106), .ZN(n19796) );
  AND2_X1 U11359 ( .A1(n16384), .A2(n15200), .ZN(n16234) );
  OR2_X2 U11360 ( .A1(n20687), .A2(n14966), .ZN(n18099) );
  AND2_X2 U11361 ( .A1(n14107), .A2(n14108), .ZN(n14149) );
  AND2_X2 U11362 ( .A1(n14099), .A2(n14105), .ZN(n14146) );
  INV_X2 U11363 ( .A(n14116), .ZN(n14163) );
  NOR2_X1 U11364 ( .A1(n14965), .A2(n14964), .ZN(n11160) );
  NOR2_X1 U11365 ( .A1(n14965), .A2(n14964), .ZN(n11161) );
  XNOR2_X2 U11366 ( .A(n12177), .B(n12176), .ZN(n15112) );
  BUF_X4 U11367 ( .A(n17979), .Z(n20722) );
  NOR2_X2 U11369 ( .A1(n14460), .A2(n17199), .ZN(n14484) );
  AOI21_X2 U11370 ( .B1(n17212), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14460) );
  BUF_X4 U11371 ( .A(n14984), .Z(n18366) );
  AOI211_X4 U11372 ( .C1(n20684), .C2(n15985), .A(n20638), .B(n17680), .ZN(
        n21318) );
  INV_X1 U11373 ( .A(n14710), .ZN(n13338) );
  AND2_X1 U11374 ( .A1(n14410), .A2(n14710), .ZN(n11566) );
  AND2_X2 U11375 ( .A1(n16041), .A2(n17295), .ZN(n17285) );
  OAI211_X2 U11376 ( .C1(n11769), .C2(n11766), .A(n17178), .B(n11765), .ZN(
        n17168) );
  AOI21_X1 U11377 ( .B1(n15754), .B2(n14200), .A(n14201), .ZN(n14202) );
  NAND2_X1 U11378 ( .A1(n18575), .A2(n21694), .ZN(n18574) );
  INV_X1 U11379 ( .A(n18813), .ZN(n18821) );
  INV_X4 U11380 ( .A(n18815), .ZN(n18828) );
  AND2_X1 U11381 ( .A1(n14109), .A2(n14106), .ZN(n14151) );
  INV_X1 U11382 ( .A(n21748), .ZN(n21628) );
  NAND2_X1 U11383 ( .A1(n11501), .A2(n12013), .ZN(n15101) );
  NOR2_X1 U11384 ( .A1(n15882), .A2(n15881), .ZN(n15921) );
  NAND2_X1 U11385 ( .A1(n20493), .A2(n15309), .ZN(n20483) );
  OR2_X1 U11386 ( .A1(n21337), .A2(n21339), .ZN(n11519) );
  INV_X4 U11387 ( .A(n21054), .ZN(n21080) );
  NOR2_X1 U11388 ( .A1(n18632), .A2(n20693), .ZN(n18656) );
  INV_X4 U11389 ( .A(n16060), .ZN(n14287) );
  CLKBUF_X3 U11390 ( .A(n13114), .Z(n19982) );
  NAND4_X2 U11391 ( .A1(n14550), .A2(n12943), .A3(n15592), .A4(n15529), .ZN(
        n14785) );
  INV_X2 U11392 ( .A(n14410), .ZN(n20079) );
  AND2_X1 U11393 ( .A1(n18674), .A2(n11288), .ZN(n18499) );
  NOR2_X1 U11394 ( .A1(n18451), .A2(n18461), .ZN(n18674) );
  BUF_X1 U11395 ( .A(n11182), .Z(n11174) );
  CLKBUF_X2 U11396 ( .A(n13027), .Z(n16398) );
  INV_X4 U11397 ( .A(n14959), .ZN(n18348) );
  BUF_X1 U11398 ( .A(n11181), .Z(n11173) );
  CLKBUF_X2 U11399 ( .A(n11907), .Z(n12581) );
  CLKBUF_X2 U11400 ( .A(n12015), .Z(n12588) );
  BUF_X4 U11401 ( .A(n15006), .Z(n11163) );
  CLKBUF_X2 U11402 ( .A(n11959), .Z(n12635) );
  NOR2_X4 U11403 ( .A1(n14966), .A2(n14964), .ZN(n18324) );
  INV_X2 U11405 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21342) );
  NAND2_X1 U11406 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21344) );
  NOR2_X1 U11408 ( .A1(n17154), .A2(n17153), .ZN(n17371) );
  AND2_X1 U11409 ( .A1(n16174), .A2(n16175), .ZN(n11755) );
  MUX2_X1 U11410 ( .A(n17152), .B(n17162), .S(n17151), .Z(n17154) );
  OR2_X1 U11411 ( .A1(n16590), .A2(n11832), .ZN(n16594) );
  INV_X1 U11412 ( .A(n11496), .ZN(n17212) );
  XNOR2_X1 U11413 ( .A(n16142), .B(n11430), .ZN(n16124) );
  NAND2_X1 U11414 ( .A1(n16432), .A2(n13651), .ZN(n16450) );
  AND2_X1 U11415 ( .A1(n17139), .A2(n11561), .ZN(n16142) );
  NAND2_X1 U11416 ( .A1(n11359), .A2(n11358), .ZN(n11496) );
  AND2_X1 U11417 ( .A1(n17127), .A2(n17128), .ZN(n17130) );
  AOI21_X1 U11418 ( .B1(n17216), .B2(n16046), .A(n14467), .ZN(n17206) );
  NOR2_X1 U11419 ( .A1(n17177), .A2(n16078), .ZN(n17139) );
  OR2_X1 U11420 ( .A1(n17177), .A2(n11331), .ZN(n16143) );
  XNOR2_X1 U11421 ( .A(n16329), .B(n11837), .ZN(n17004) );
  NAND2_X1 U11422 ( .A1(n17008), .A2(n11831), .ZN(n16329) );
  OR2_X1 U11423 ( .A1(n16702), .A2(n11788), .ZN(n12929) );
  XNOR2_X1 U11424 ( .A(n16151), .B(n16150), .ZN(n16169) );
  XNOR2_X1 U11425 ( .A(n16145), .B(n11732), .ZN(n16414) );
  OR2_X1 U11426 ( .A1(n16986), .A2(n16997), .ZN(n19150) );
  NAND2_X1 U11427 ( .A1(n11472), .A2(n11245), .ZN(n17193) );
  OAI21_X1 U11428 ( .B1(n14529), .B2(n11328), .A(n11861), .ZN(n20544) );
  NAND2_X1 U11429 ( .A1(n18601), .A2(n21665), .ZN(n21647) );
  NAND2_X1 U11430 ( .A1(n15902), .A2(n11310), .ZN(n17027) );
  CLKBUF_X1 U11431 ( .A(n14529), .Z(n16734) );
  XNOR2_X1 U11432 ( .A(n18659), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21621) );
  NAND2_X1 U11433 ( .A1(n18606), .A2(n21666), .ZN(n18601) );
  NAND2_X1 U11434 ( .A1(n18607), .A2(n18640), .ZN(n18606) );
  AND2_X1 U11435 ( .A1(n16067), .A2(n11463), .ZN(n11462) );
  NAND2_X1 U11436 ( .A1(n18658), .A2(n21664), .ZN(n18659) );
  AND2_X1 U11437 ( .A1(n17151), .A2(n17163), .ZN(n16067) );
  AND2_X1 U11438 ( .A1(n16063), .A2(n16075), .ZN(n17151) );
  NAND2_X1 U11439 ( .A1(n14315), .A2(n18984), .ZN(n14316) );
  AND2_X1 U11440 ( .A1(n14311), .A2(n14310), .ZN(n17611) );
  NOR2_X1 U11441 ( .A1(n16074), .A2(n17377), .ZN(n17162) );
  OR2_X1 U11442 ( .A1(n11762), .A2(n17180), .ZN(n11765) );
  NAND2_X1 U11443 ( .A1(n11467), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11466) );
  AND2_X1 U11444 ( .A1(n18613), .A2(n11388), .ZN(n18598) );
  AND2_X1 U11445 ( .A1(n15419), .A2(n15443), .ZN(n11835) );
  OR2_X1 U11446 ( .A1(n16069), .A2(n16068), .ZN(n16072) );
  AND2_X1 U11447 ( .A1(n18574), .A2(n11592), .ZN(n18614) );
  NAND2_X1 U11448 ( .A1(n18574), .A2(n21649), .ZN(n18613) );
  OR2_X1 U11449 ( .A1(n17180), .A2(n11767), .ZN(n11766) );
  AND2_X1 U11450 ( .A1(n18563), .A2(n18564), .ZN(n18575) );
  INV_X1 U11451 ( .A(n16056), .ZN(n13636) );
  AND2_X1 U11452 ( .A1(n11593), .A2(n11325), .ZN(n11592) );
  OR2_X1 U11453 ( .A1(n17067), .A2(n17058), .ZN(n17060) );
  AND2_X1 U11454 ( .A1(n14171), .A2(n14170), .ZN(n14174) );
  OR2_X1 U11455 ( .A1(n16051), .A2(n16050), .ZN(n16056) );
  NAND2_X1 U11456 ( .A1(n14192), .A2(n14191), .ZN(n14204) );
  NOR2_X1 U11457 ( .A1(n18668), .A2(n18640), .ZN(n18522) );
  OR2_X1 U11458 ( .A1(n14189), .A2(n14188), .ZN(n14192) );
  NAND2_X1 U11459 ( .A1(n11230), .A2(n12212), .ZN(n14953) );
  NOR2_X1 U11460 ( .A1(n15499), .A2(n15455), .ZN(n22783) );
  AND2_X2 U11461 ( .A1(n12890), .A2(n12908), .ZN(n11861) );
  NOR2_X2 U11462 ( .A1(n18827), .A2(n18815), .ZN(n18671) );
  NOR2_X2 U11463 ( .A1(n21655), .A2(n18831), .ZN(n18745) );
  OR2_X1 U11464 ( .A1(n14359), .A2(n14357), .ZN(n14374) );
  AND2_X1 U11465 ( .A1(n18437), .A2(n11848), .ZN(n11859) );
  NAND2_X1 U11466 ( .A1(n21370), .A2(n21850), .ZN(n18831) );
  AND2_X1 U11467 ( .A1(n14870), .A2(n14868), .ZN(n12190) );
  CLKBUF_X1 U11468 ( .A(n12854), .Z(n15172) );
  NAND2_X1 U11469 ( .A1(n11513), .A2(n11511), .ZN(n12202) );
  INV_X1 U11470 ( .A(n21489), .ZN(n21721) );
  NAND2_X1 U11471 ( .A1(n14816), .A2(n14815), .ZN(n14857) );
  AND2_X1 U11472 ( .A1(n14844), .A2(n14686), .ZN(n14104) );
  OR2_X1 U11473 ( .A1(n18436), .A2(n21743), .ZN(n18437) );
  NOR2_X1 U11474 ( .A1(n18708), .A2(n21731), .ZN(n18436) );
  AND2_X1 U11475 ( .A1(n16575), .A2(n16518), .ZN(n16567) );
  NAND2_X1 U11476 ( .A1(n18698), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n21489) );
  AND2_X1 U11477 ( .A1(n18426), .A2(n11260), .ZN(n11541) );
  NAND2_X1 U11478 ( .A1(n11577), .A2(n13160), .ZN(n11552) );
  OR2_X1 U11479 ( .A1(n14705), .A2(n14704), .ZN(n14821) );
  AND2_X1 U11480 ( .A1(n17634), .A2(n19183), .ZN(n14108) );
  AND2_X1 U11481 ( .A1(n15239), .A2(n19183), .ZN(n14105) );
  NAND2_X2 U11482 ( .A1(n16659), .A2(n14896), .ZN(n16667) );
  AND2_X1 U11483 ( .A1(n18748), .A2(n18392), .ZN(n18737) );
  XNOR2_X1 U11484 ( .A(n14819), .B(n14818), .ZN(n14705) );
  NAND2_X1 U11485 ( .A1(n18762), .A2(n18421), .ZN(n18756) );
  OAI21_X1 U11486 ( .B1(n19183), .B2(n17692), .A(n14699), .ZN(n14819) );
  NAND2_X1 U11487 ( .A1(n12084), .A2(n12058), .ZN(n12170) );
  OR2_X1 U11488 ( .A1(n14799), .A2(n12184), .ZN(n12185) );
  NAND2_X1 U11489 ( .A1(n18764), .A2(n18388), .ZN(n18453) );
  NAND2_X1 U11490 ( .A1(n13173), .A2(n13172), .ZN(n14085) );
  NAND2_X4 U11491 ( .A1(n21775), .A2(n21768), .ZN(n21748) );
  CLKBUF_X1 U11492 ( .A(n15134), .Z(n22430) );
  NOR2_X1 U11493 ( .A1(n21122), .A2(n21121), .ZN(n21302) );
  NOR2_X2 U11494 ( .A1(n20077), .A2(n20234), .ZN(n20078) );
  NOR2_X2 U11495 ( .A1(n20028), .A2(n20234), .ZN(n20029) );
  NOR2_X2 U11496 ( .A1(n19980), .A2(n20234), .ZN(n19981) );
  NOR2_X2 U11497 ( .A1(n19932), .A2(n20234), .ZN(n19933) );
  NOR2_X2 U11498 ( .A1(n19721), .A2(n20234), .ZN(n19722) );
  INV_X2 U11499 ( .A(n17044), .ZN(n15444) );
  AND2_X1 U11500 ( .A1(n13628), .A2(n13627), .ZN(n14321) );
  INV_X1 U11501 ( .A(n11519), .ZN(n21327) );
  OAI221_X2 U11502 ( .B1(n18396), .B2(n21320), .C1(n18396), .C2(n21319), .A(
        n21348), .ZN(n21606) );
  CLKBUF_X1 U11503 ( .A(n13176), .Z(n13294) );
  AOI21_X1 U11504 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13176), .A(
        n13167), .ZN(n13169) );
  NAND2_X1 U11505 ( .A1(n14281), .A2(n14282), .ZN(n14314) );
  AND2_X1 U11506 ( .A1(n14288), .A2(n14300), .ZN(n14281) );
  AOI21_X1 U11507 ( .B1(n19455), .B2(n15992), .A(n15991), .ZN(n21348) );
  AND2_X1 U11508 ( .A1(n14289), .A2(n14290), .ZN(n14288) );
  NAND2_X1 U11509 ( .A1(n18795), .A2(n18381), .ZN(n18787) );
  AND2_X1 U11510 ( .A1(n21367), .A2(n15983), .ZN(n20638) );
  AND2_X1 U11511 ( .A1(n11987), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12003) );
  NOR2_X1 U11512 ( .A1(n14297), .A2(n14298), .ZN(n14289) );
  AND2_X1 U11513 ( .A1(n13129), .A2(n13128), .ZN(n11803) );
  NOR2_X2 U11514 ( .A1(n21655), .A2(n18389), .ZN(n18640) );
  OR2_X1 U11515 ( .A1(n14388), .A2(n14216), .ZN(n13142) );
  AOI21_X1 U11516 ( .B1(n14535), .B2(n14789), .A(n11980), .ZN(n11981) );
  CLKBUF_X1 U11517 ( .A(n12662), .Z(n15103) );
  INV_X2 U11518 ( .A(n13532), .ZN(n13394) );
  INV_X1 U11519 ( .A(n14249), .ZN(n15280) );
  NOR2_X1 U11520 ( .A1(n21165), .A2(n18408), .ZN(n18359) );
  NAND2_X1 U11521 ( .A1(n11562), .A2(n11566), .ZN(n14378) );
  INV_X1 U11522 ( .A(n21115), .ZN(n19589) );
  AND3_X1 U11523 ( .A1(n11566), .A2(n11258), .A3(n11563), .ZN(n14383) );
  NOR2_X1 U11524 ( .A1(n18362), .A2(n18363), .ZN(n18365) );
  AND2_X1 U11525 ( .A1(n11565), .A2(n13112), .ZN(n11562) );
  NOR2_X1 U11526 ( .A1(n15979), .A2(n21180), .ZN(n21363) );
  NAND2_X1 U11527 ( .A1(n11232), .A2(n11411), .ZN(n21115) );
  CLKBUF_X1 U11528 ( .A(n19175), .Z(n11178) );
  AND2_X1 U11529 ( .A1(n13468), .A2(n13467), .ZN(n16060) );
  OR2_X1 U11530 ( .A1(n14895), .A2(n11979), .ZN(n14789) );
  AND2_X1 U11531 ( .A1(n15406), .A2(n12820), .ZN(n14730) );
  AND2_X1 U11532 ( .A1(n18361), .A2(n18412), .ZN(n18362) );
  AND3_X1 U11533 ( .A1(n14878), .A2(n20030), .A3(n13114), .ZN(n11427) );
  NAND2_X1 U11534 ( .A1(n14700), .A2(n13114), .ZN(n13123) );
  NAND2_X1 U11535 ( .A1(n15981), .A2(n21180), .ZN(n21122) );
  NAND2_X1 U11536 ( .A1(n14550), .A2(n16595), .ZN(n14559) );
  OR2_X1 U11537 ( .A1(n13354), .A2(n13353), .ZN(n14264) );
  NAND2_X1 U11538 ( .A1(n11204), .A2(n11235), .ZN(n21366) );
  AND2_X1 U11539 ( .A1(n12842), .A2(n11158), .ZN(n12943) );
  OR2_X1 U11540 ( .A1(n13420), .A2(n13419), .ZN(n14140) );
  OR2_X1 U11541 ( .A1(n13406), .A2(n13405), .ZN(n14127) );
  INV_X1 U11542 ( .A(n20684), .ZN(n21370) );
  OAI21_X2 U11543 ( .B1(n22630), .B2(n20605), .A(n15590), .ZN(n15591) );
  OAI21_X2 U11544 ( .B1(n22630), .B2(n20613), .A(n15389), .ZN(n15390) );
  OAI21_X2 U11545 ( .B1(n22630), .B2(n20617), .A(n15381), .ZN(n15382) );
  NOR2_X2 U11546 ( .A1(n14983), .A2(n14982), .ZN(n20684) );
  INV_X1 U11547 ( .A(n15127), .ZN(n22414) );
  NOR2_X2 U11548 ( .A1(n14973), .A2(n14972), .ZN(n21219) );
  NAND2_X1 U11549 ( .A1(n13017), .A2(n13016), .ZN(n13064) );
  NAND2_X1 U11550 ( .A1(n13103), .A2(n13102), .ZN(n14405) );
  INV_X4 U11551 ( .A(n13113), .ZN(n20237) );
  OAI21_X2 U11552 ( .B1(n22630), .B2(n20623), .A(n15527), .ZN(n15528) );
  OAI21_X2 U11553 ( .B1(n22630), .B2(n20610), .A(n15141), .ZN(n15142) );
  NAND2_X2 U11554 ( .A1(n14764), .A2(n11177), .ZN(n12752) );
  NAND2_X1 U11555 ( .A1(n11922), .A2(n15309), .ZN(n16591) );
  NAND2_X1 U11556 ( .A1(n11228), .A2(n11894), .ZN(n11921) );
  AND4_X1 U11557 ( .A1(n13070), .A2(n13069), .A3(n13068), .A4(n13067), .ZN(
        n13071) );
  NAND2_X2 U11558 ( .A1(U214), .A2(n20565), .ZN(n20626) );
  INV_X2 U11559 ( .A(U214), .ZN(n20615) );
  AND2_X2 U11560 ( .A1(n11192), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13446) );
  BUF_X2 U11561 ( .A(n14985), .Z(n18335) );
  INV_X2 U11562 ( .A(n18728), .ZN(n11165) );
  AND2_X1 U11563 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11410) );
  AND4_X1 U11564 ( .A1(n11941), .A2(n11940), .A3(n11939), .A4(n11938), .ZN(
        n11952) );
  AND4_X1 U11565 ( .A1(n11949), .A2(n11948), .A3(n11947), .A4(n11946), .ZN(
        n11950) );
  AND4_X1 U11566 ( .A1(n11893), .A2(n11892), .A3(n11891), .A4(n11890), .ZN(
        n11894) );
  AND2_X1 U11567 ( .A1(n18715), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18750) );
  NAND2_X2 U11568 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17907), .ZN(n17900) );
  INV_X2 U11569 ( .A(n11852), .ZN(n11180) );
  BUF_X2 U11570 ( .A(n18324), .Z(n18254) );
  INV_X1 U11571 ( .A(n11187), .ZN(n11191) );
  BUF_X2 U11572 ( .A(n12107), .Z(n12348) );
  AND2_X2 U11573 ( .A1(n16399), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13460) );
  BUF_X2 U11574 ( .A(n12107), .Z(n12626) );
  INV_X2 U11575 ( .A(n19581), .ZN(U215) );
  OR2_X2 U11576 ( .A1(n22805), .A2(n17750), .ZN(n17710) );
  NAND2_X1 U11577 ( .A1(n20710), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n18346) );
  BUF_X2 U11578 ( .A(n11937), .Z(n12630) );
  NOR2_X4 U11579 ( .A1(n21355), .A2(n14967), .ZN(n14984) );
  INV_X2 U11580 ( .A(n20347), .ZN(n20372) );
  BUF_X4 U11581 ( .A(n18223), .Z(n11167) );
  INV_X2 U11582 ( .A(n20428), .ZN(n11168) );
  INV_X2 U11583 ( .A(n20426), .ZN(n11169) );
  AND2_X1 U11584 ( .A1(n11866), .A2(n11801), .ZN(n12107) );
  NOR2_X2 U11585 ( .A1(n21811), .A2(n19314), .ZN(n19576) );
  BUF_X4 U11586 ( .A(n14988), .Z(n11171) );
  BUF_X4 U11587 ( .A(n18321), .Z(n11172) );
  AND2_X1 U11588 ( .A1(n15088), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11801) );
  AND2_X2 U11589 ( .A1(n14243), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13321) );
  NOR2_X1 U11590 ( .A1(n14422), .A2(n17461), .ZN(n11358) );
  AND2_X1 U11591 ( .A1(n11983), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11867) );
  AND2_X1 U11592 ( .A1(n21342), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n21345) );
  NAND2_X1 U11593 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21361), .ZN(
        n21355) );
  NOR2_X1 U11594 ( .A1(n21341), .A2(n21310), .ZN(n20710) );
  NAND2_X1 U11595 ( .A1(n21310), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n21347) );
  INV_X2 U11596 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21310) );
  INV_X1 U11597 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21324) );
  INV_X2 U11598 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21855) );
  AND2_X2 U11599 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14243) );
  AND2_X1 U11600 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13330) );
  AND2_X1 U11601 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15098) );
  AND2_X2 U11602 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15076) );
  AOI22_X1 U11603 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19796), .B1(
        n14164), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14110) );
  NOR3_X1 U11604 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n21347), .ZN(n15058) );
  NAND2_X2 U11605 ( .A1(n14882), .A2(n14881), .ZN(n15330) );
  OAI211_X1 U11606 ( .C1(n13150), .C2(n17752), .A(n13149), .B(n13148), .ZN(
        n14089) );
  NOR2_X4 U11607 ( .A1(n16473), .A2(n16474), .ZN(n16460) );
  NAND4_X1 U11608 ( .A1(n11953), .A2(n11952), .A3(n11951), .A4(n11950), .ZN(
        n11176) );
  NAND4_X1 U11609 ( .A1(n11953), .A2(n11952), .A3(n11951), .A4(n11950), .ZN(
        n11177) );
  AOI21_X1 U11610 ( .B1(n13161), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13162), .ZN(n13168) );
  INV_X1 U11611 ( .A(n14764), .ZN(n11179) );
  NAND2_X2 U11612 ( .A1(n14700), .A2(n11183), .ZN(n13110) );
  NAND3_X2 U11613 ( .A1(n11431), .A2(n11553), .A3(n11555), .ZN(n15556) );
  INV_X2 U11614 ( .A(n11210), .ZN(n12786) );
  NAND2_X1 U11615 ( .A1(n14087), .A2(n14086), .ZN(n11577) );
  INV_X4 U11616 ( .A(n16374), .ZN(n16400) );
  AOI21_X2 U11617 ( .B1(n16433), .B2(n16432), .A(n16431), .ZN(n16678) );
  NOR3_X1 U11618 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n21347), .ZN(n11181) );
  NOR3_X1 U11619 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n21347), .ZN(n11182) );
  NAND2_X1 U11620 ( .A1(n11581), .A2(n11579), .ZN(n11183) );
  XNOR2_X2 U11621 ( .A(n11800), .B(n14143), .ZN(n15649) );
  NAND2_X2 U11622 ( .A1(n15556), .A2(n14139), .ZN(n11800) );
  AOI21_X2 U11623 ( .B1(n17227), .B2(n16039), .A(n14371), .ZN(n17216) );
  NOR2_X2 U11624 ( .A1(n15346), .A2(n15345), .ZN(n15419) );
  NOR2_X2 U11625 ( .A1(n11425), .A2(n17616), .ZN(n17612) );
  NOR2_X2 U11626 ( .A1(n14199), .A2(n14198), .ZN(n11425) );
  NOR2_X4 U11627 ( .A1(n16923), .A2(n17000), .ZN(n16995) );
  NAND2_X2 U11628 ( .A1(n17030), .A2(n11315), .ZN(n16923) );
  NOR2_X2 U11629 ( .A1(n15704), .A2(n15705), .ZN(n15685) );
  AND2_X1 U11630 ( .A1(n14844), .A2(n14808), .ZN(n14099) );
  AND2_X1 U11631 ( .A1(n14243), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11184) );
  AND2_X2 U11632 ( .A1(n14243), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11185) );
  INV_X2 U11633 ( .A(n16259), .ZN(n11186) );
  INV_X1 U11634 ( .A(n16259), .ZN(n11187) );
  INV_X1 U11635 ( .A(n16259), .ZN(n11188) );
  INV_X1 U11636 ( .A(n11186), .ZN(n11189) );
  INV_X1 U11637 ( .A(n11186), .ZN(n11190) );
  INV_X1 U11638 ( .A(n11187), .ZN(n11192) );
  INV_X1 U11639 ( .A(n11187), .ZN(n11193) );
  INV_X1 U11640 ( .A(n11188), .ZN(n11194) );
  INV_X1 U11641 ( .A(n11188), .ZN(n11195) );
  INV_X1 U11642 ( .A(n11188), .ZN(n11196) );
  AND2_X2 U11643 ( .A1(n15192), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16259) );
  BUF_X4 U11646 ( .A(n13021), .Z(n16399) );
  NAND2_X1 U11647 ( .A1(n14580), .A2(n15127), .ZN(n12014) );
  AND2_X1 U11648 ( .A1(n14701), .A2(n14700), .ZN(n16347) );
  NAND2_X1 U11649 ( .A1(n14851), .A2(n14850), .ZN(n14853) );
  NAND2_X1 U11650 ( .A1(n14864), .A2(n14812), .ZN(n14851) );
  OR2_X1 U11651 ( .A1(n21860), .A2(n12726), .ZN(n14075) );
  NOR2_X1 U11652 ( .A1(n17060), .A2(n11589), .ZN(n11591) );
  NAND2_X1 U11653 ( .A1(n11590), .A2(n13608), .ZN(n11589) );
  INV_X1 U11654 ( .A(n14447), .ZN(n11590) );
  AND2_X1 U11655 ( .A1(n14567), .A2(n11976), .ZN(n11993) );
  NOR2_X1 U11656 ( .A1(n11477), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11476) );
  INV_X1 U11657 ( .A(n14312), .ZN(n14201) );
  NAND2_X1 U11658 ( .A1(n11428), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11487) );
  NAND2_X1 U11659 ( .A1(n21172), .A2(n11536), .ZN(n18407) );
  NAND2_X1 U11660 ( .A1(n11540), .A2(n18412), .ZN(n11536) );
  AND2_X1 U11661 ( .A1(n11273), .A2(n16512), .ZN(n11826) );
  NAND3_X1 U11662 ( .A1(n11514), .A2(n11367), .A3(n11246), .ZN(n14529) );
  NAND2_X1 U11663 ( .A1(n11236), .A2(n11792), .ZN(n11514) );
  XNOR2_X1 U11664 ( .A(n12890), .B(n12148), .ZN(n12898) );
  INV_X1 U11665 ( .A(n16503), .ZN(n11749) );
  NAND2_X1 U11666 ( .A1(n11580), .A2(n15200), .ZN(n11579) );
  INV_X1 U11667 ( .A(n17101), .ZN(n11624) );
  INV_X1 U11668 ( .A(n15187), .ZN(n11735) );
  NAND2_X1 U11669 ( .A1(n17129), .A2(n17141), .ZN(n11757) );
  INV_X1 U11670 ( .A(n13164), .ZN(n13287) );
  NOR2_X1 U11671 ( .A1(n11607), .A2(n15839), .ZN(n11606) );
  INV_X1 U11672 ( .A(n11610), .ZN(n11607) );
  OAI22_X1 U11673 ( .A1(n11270), .A2(n11441), .B1(n18973), .B2(n11444), .ZN(
        n11440) );
  NOR2_X1 U11674 ( .A1(n13336), .A2(n13335), .ZN(n14190) );
  INV_X1 U11675 ( .A(n13572), .ZN(n13534) );
  OR2_X1 U11676 ( .A1(n14757), .A2(n13380), .ZN(n13391) );
  NAND2_X1 U11677 ( .A1(n14853), .A2(n14852), .ZN(n14880) );
  NAND2_X1 U11678 ( .A1(n13314), .A2(n13119), .ZN(n14382) );
  NAND2_X1 U11679 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21310), .ZN(
        n14964) );
  INV_X1 U11680 ( .A(n21345), .ZN(n14965) );
  NAND2_X1 U11681 ( .A1(n18614), .A2(n18596), .ZN(n18599) );
  INV_X1 U11682 ( .A(n18597), .ZN(n11388) );
  INV_X1 U11683 ( .A(n18362), .ZN(n18408) );
  NAND2_X1 U11684 ( .A1(n16465), .A2(n16452), .ZN(n16451) );
  AND2_X1 U11685 ( .A1(n16669), .A2(n16672), .ZN(n13652) );
  AND2_X1 U11686 ( .A1(n16478), .A2(n16463), .ZN(n16465) );
  AND2_X1 U11687 ( .A1(n16488), .A2(n16476), .ZN(n16478) );
  AND2_X1 U11688 ( .A1(n14547), .A2(n22809), .ZN(n14583) );
  AND2_X1 U11689 ( .A1(n14755), .A2(n14754), .ZN(n14757) );
  NOR2_X1 U11690 ( .A1(n15688), .A2(n15773), .ZN(n11739) );
  NAND2_X1 U11691 ( .A1(n11739), .A2(n11738), .ZN(n15889) );
  INV_X1 U11692 ( .A(n14381), .ZN(n11738) );
  INV_X1 U11693 ( .A(n11466), .ZN(n11465) );
  NAND2_X1 U11694 ( .A1(n11464), .A2(n11466), .ZN(n11463) );
  INV_X1 U11695 ( .A(n11433), .ZN(n11432) );
  OAI21_X1 U11696 ( .B1(n14317), .B2(n11434), .A(n11773), .ZN(n11433) );
  AOI21_X1 U11697 ( .B1(n11201), .B2(n11774), .A(n11282), .ZN(n11773) );
  NAND2_X1 U11698 ( .A1(n14209), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14210) );
  NAND2_X1 U11699 ( .A1(n21649), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U11700 ( .A1(n11374), .A2(n11238), .ZN(n11373) );
  INV_X1 U11701 ( .A(n14770), .ZN(n11374) );
  NAND2_X1 U11702 ( .A1(n16115), .A2(n19189), .ZN(n16119) );
  XNOR2_X1 U11703 ( .A(n13661), .B(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n13664) );
  XNOR2_X1 U11704 ( .A(n13662), .B(DATAI_31_), .ZN(n13663) );
  INV_X1 U11705 ( .A(keyinput_0), .ZN(n13661) );
  INV_X1 U11706 ( .A(keyinput_4), .ZN(n13668) );
  AOI21_X1 U11707 ( .B1(n11720), .B2(n11719), .A(n11718), .ZN(n13681) );
  NAND2_X1 U11708 ( .A1(n20459), .A2(keyinput_48), .ZN(n11713) );
  AOI21_X1 U11709 ( .B1(n11689), .B2(n11686), .A(n13768), .ZN(n11685) );
  AND2_X1 U11710 ( .A1(n11688), .A2(n11687), .ZN(n11686) );
  OR2_X1 U11711 ( .A1(n13764), .A2(n11690), .ZN(n11689) );
  NAND2_X1 U11712 ( .A1(n11698), .A2(n13810), .ZN(n11697) );
  OAI21_X1 U11713 ( .B1(n13798), .B2(n11700), .A(n11699), .ZN(n11698) );
  AOI21_X1 U11714 ( .B1(n12581), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n11280), .ZN(n12045) );
  NAND2_X1 U11715 ( .A1(n13382), .A2(n13381), .ZN(n11630) );
  NAND2_X1 U11716 ( .A1(n14895), .A2(n12842), .ZN(n11995) );
  CLKBUF_X1 U11717 ( .A(n12107), .Z(n12610) );
  CLKBUF_X2 U11718 ( .A(n11885), .Z(n12587) );
  CLKBUF_X2 U11719 ( .A(n12067), .Z(n12560) );
  OR2_X1 U11720 ( .A1(n12014), .A2(n22225), .ZN(n12695) );
  NAND2_X1 U11721 ( .A1(n13161), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11802) );
  NAND2_X1 U11722 ( .A1(n13163), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11804) );
  AND2_X1 U11723 ( .A1(n11554), .A2(n14140), .ZN(n11770) );
  NOR2_X1 U11724 ( .A1(n13301), .A2(n13305), .ZN(n13302) );
  INV_X1 U11725 ( .A(n13306), .ZN(n13301) );
  NAND2_X1 U11726 ( .A1(n21368), .A2(n15979), .ZN(n15999) );
  AND2_X1 U11727 ( .A1(n12687), .A2(n12718), .ZN(n12721) );
  NAND2_X1 U11728 ( .A1(n11992), .A2(n11991), .ZN(n12061) );
  NOR2_X1 U11729 ( .A1(n12435), .A2(n11828), .ZN(n11827) );
  INV_X1 U11730 ( .A(n16647), .ZN(n11828) );
  NAND2_X1 U11731 ( .A1(n11215), .A2(n11278), .ZN(n11818) );
  INV_X1 U11732 ( .A(n15885), .ZN(n11820) );
  INV_X1 U11733 ( .A(n12264), .ZN(n12652) );
  AND2_X1 U11734 ( .A1(n15427), .A2(n15562), .ZN(n11821) );
  AND2_X1 U11735 ( .A1(n12216), .A2(n12158), .ZN(n12880) );
  INV_X1 U11736 ( .A(n12650), .ZN(n12657) );
  INV_X1 U11737 ( .A(n17711), .ZN(n12650) );
  NAND2_X1 U11738 ( .A1(n16549), .A2(n11744), .ZN(n11743) );
  INV_X1 U11739 ( .A(n14578), .ZN(n11744) );
  INV_X1 U11740 ( .A(n12915), .ZN(n11797) );
  NAND2_X1 U11741 ( .A1(n11502), .A2(n12915), .ZN(n11794) );
  INV_X1 U11742 ( .A(n15777), .ZN(n11502) );
  NOR2_X1 U11743 ( .A1(n12215), .A2(n12157), .ZN(n11812) );
  NOR2_X1 U11744 ( .A1(n11786), .A2(n11783), .ZN(n11782) );
  INV_X1 U11745 ( .A(n15605), .ZN(n11783) );
  INV_X1 U11746 ( .A(n15716), .ZN(n11786) );
  NAND2_X1 U11747 ( .A1(n11210), .A2(n12752), .ZN(n12794) );
  AND2_X1 U11748 ( .A1(n12848), .A2(n11365), .ZN(n12851) );
  INV_X1 U11749 ( .A(n11366), .ZN(n11365) );
  OAI21_X1 U11750 ( .B1(n12850), .B2(n12849), .A(n12847), .ZN(n11366) );
  INV_X1 U11751 ( .A(n12695), .ZN(n12720) );
  NOR2_X1 U11752 ( .A1(n12704), .A2(n12686), .ZN(n12723) );
  NAND2_X1 U11753 ( .A1(n22225), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11378) );
  NOR2_X1 U11754 ( .A1(n16064), .A2(n11651), .ZN(n11650) );
  INV_X1 U11755 ( .A(n16055), .ZN(n11651) );
  NOR2_X1 U11756 ( .A1(n11682), .A2(n11681), .ZN(n11680) );
  NAND2_X1 U11757 ( .A1(n13631), .A2(n14329), .ZN(n14337) );
  INV_X1 U11758 ( .A(n14331), .ZN(n13631) );
  NAND2_X1 U11759 ( .A1(n14321), .A2(n11644), .ZN(n14331) );
  AND2_X1 U11760 ( .A1(n11231), .A2(n11645), .ZN(n11644) );
  INV_X1 U11761 ( .A(n14325), .ZN(n11645) );
  OAI211_X1 U11762 ( .C1(n13143), .C2(n13621), .A(n13156), .B(n13155), .ZN(
        n13157) );
  NOR2_X1 U11763 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16249) );
  NOR2_X1 U11764 ( .A1(n12955), .A2(n12956), .ZN(n12954) );
  INV_X1 U11765 ( .A(n12982), .ZN(n11723) );
  INV_X1 U11766 ( .A(n16925), .ZN(n11736) );
  NOR2_X1 U11767 ( .A1(n14392), .A2(n11612), .ZN(n17411) );
  NAND2_X1 U11768 ( .A1(n11218), .A2(n17111), .ZN(n11612) );
  NAND2_X1 U11769 ( .A1(n17411), .A2(n17410), .ZN(n17409) );
  INV_X1 U11770 ( .A(n11476), .ZN(n11473) );
  NAND2_X1 U11771 ( .A1(n11470), .A2(n16040), .ZN(n11469) );
  NOR2_X1 U11772 ( .A1(n11244), .A2(n11475), .ZN(n11474) );
  AND2_X1 U11773 ( .A1(n11477), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11475) );
  INV_X1 U11774 ( .A(n15334), .ZN(n11734) );
  NAND2_X1 U11775 ( .A1(n11618), .A2(n17509), .ZN(n11617) );
  INV_X1 U11776 ( .A(n11620), .ZN(n11618) );
  NAND2_X1 U11777 ( .A1(n14340), .A2(n14339), .ZN(n16041) );
  NOR2_X1 U11778 ( .A1(n13455), .A2(n13454), .ZN(n13468) );
  AOI21_X1 U11779 ( .B1(n17620), .B2(n11263), .A(n11611), .ZN(n11610) );
  INV_X1 U11780 ( .A(n17601), .ZN(n11611) );
  AND3_X1 U11781 ( .A1(n13423), .A2(n13422), .A3(n13421), .ZN(n15326) );
  NAND2_X1 U11782 ( .A1(n13139), .A2(n20237), .ZN(n11740) );
  NOR2_X1 U11783 ( .A1(n13134), .A2(n11485), .ZN(n11484) );
  INV_X1 U11784 ( .A(n13142), .ZN(n11485) );
  OAI21_X1 U11785 ( .B1(n13101), .B2(n13100), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13102) );
  NOR2_X1 U11786 ( .A1(n21344), .A2(n14966), .ZN(n18122) );
  OR2_X1 U11787 ( .A1(n14967), .A2(n11384), .ZN(n14959) );
  NAND2_X1 U11788 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11384) );
  INV_X1 U11789 ( .A(n14994), .ZN(n11415) );
  NAND2_X1 U11790 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11413) );
  INV_X1 U11791 ( .A(n14993), .ZN(n11414) );
  AND2_X1 U11792 ( .A1(n11659), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11658) );
  NAND3_X1 U11793 ( .A1(n18423), .A2(n11541), .A3(n11545), .ZN(n11544) );
  INV_X1 U11794 ( .A(n18383), .ZN(n11588) );
  NOR2_X1 U11795 ( .A1(n11588), .A2(n11383), .ZN(n11382) );
  NAND2_X1 U11796 ( .A1(n21122), .A2(n11408), .ZN(n16005) );
  OR2_X1 U11797 ( .A1(n21115), .A2(n21366), .ZN(n11408) );
  NOR2_X1 U11798 ( .A1(n21219), .A2(n19455), .ZN(n18395) );
  OR2_X1 U11799 ( .A1(n15999), .A2(n21320), .ZN(n15978) );
  NAND2_X1 U11800 ( .A1(n21318), .A2(n21348), .ZN(n21337) );
  AND2_X1 U11801 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12207), .ZN(
        n12209) );
  AND4_X1 U11802 ( .A1(n11945), .A2(n11944), .A3(n11943), .A4(n11942), .ZN(
        n11951) );
  AND4_X1 U11803 ( .A1(n11936), .A2(n11935), .A3(n11934), .A4(n11933), .ZN(
        n11953) );
  AND2_X1 U11804 ( .A1(n11823), .A2(n12604), .ZN(n11822) );
  NOR2_X1 U11805 ( .A1(n16433), .A2(n11824), .ZN(n11823) );
  INV_X1 U11806 ( .A(n13650), .ZN(n11824) );
  NAND2_X1 U11807 ( .A1(n12925), .A2(n20552), .ZN(n16708) );
  NAND2_X1 U11808 ( .A1(n12315), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12329) );
  NAND2_X1 U11809 ( .A1(n12209), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12217) );
  INV_X1 U11810 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12220) );
  NOR2_X1 U11811 ( .A1(n12217), .A2(n12220), .ZN(n12218) );
  AOI21_X1 U11812 ( .B1(n11509), .B2(n11272), .A(n11507), .ZN(n11506) );
  INV_X1 U11813 ( .A(n12937), .ZN(n11507) );
  OAI21_X1 U11814 ( .B1(n20545), .B2(n11779), .A(n11776), .ZN(n16693) );
  NAND2_X1 U11815 ( .A1(n20544), .A2(n11780), .ZN(n11779) );
  AOI21_X1 U11816 ( .B1(n20544), .B2(n11777), .A(n20552), .ZN(n11776) );
  AND2_X1 U11817 ( .A1(n11780), .A2(n11778), .ZN(n11777) );
  AND2_X1 U11818 ( .A1(n16567), .A2(n11314), .ZN(n16488) );
  INV_X1 U11819 ( .A(n16489), .ZN(n11748) );
  NAND2_X1 U11820 ( .A1(n11398), .A2(n11397), .ZN(n16872) );
  NAND2_X1 U11821 ( .A1(n15776), .A2(n20552), .ZN(n11397) );
  NAND2_X1 U11822 ( .A1(n16767), .A2(n11861), .ZN(n11398) );
  NOR2_X1 U11823 ( .A1(n16872), .A2(n16879), .ZN(n16873) );
  NAND2_X1 U11824 ( .A1(n11368), .A2(n12914), .ZN(n15778) );
  NAND2_X1 U11825 ( .A1(n15778), .A2(n15777), .ZN(n15776) );
  AOI21_X1 U11826 ( .B1(n15515), .B2(n11361), .A(n11248), .ZN(n11360) );
  INV_X1 U11827 ( .A(n15515), .ZN(n11362) );
  INV_X1 U11828 ( .A(n12879), .ZN(n11361) );
  AOI21_X1 U11829 ( .B1(n16184), .B2(n15304), .A(n12741), .ZN(n14907) );
  OR3_X1 U11830 ( .A1(n14892), .A2(n14780), .A3(n14779), .ZN(n15104) );
  INV_X1 U11831 ( .A(n22626), .ZN(n22411) );
  AND2_X1 U11832 ( .A1(n15172), .A2(n11512), .ZN(n15436) );
  INV_X1 U11833 ( .A(n11677), .ZN(n11675) );
  AOI21_X1 U11834 ( .B1(n19032), .B2(n11679), .A(n11678), .ZN(n11677) );
  INV_X1 U11835 ( .A(n19148), .ZN(n11679) );
  INV_X1 U11836 ( .A(n19169), .ZN(n11678) );
  NAND2_X1 U11837 ( .A1(n11202), .A2(n15321), .ZN(n15327) );
  OAI211_X1 U11838 ( .C1(n13572), .C2(n13360), .A(n13359), .B(n13389), .ZN(
        n14754) );
  OAI21_X1 U11839 ( .B1(n13532), .B2(n13343), .A(n13342), .ZN(n14755) );
  AND2_X1 U11840 ( .A1(n13242), .A2(n13241), .ZN(n14381) );
  INV_X1 U11841 ( .A(n11569), .ZN(n11568) );
  OAI21_X1 U11842 ( .B1(n11573), .B2(n11570), .A(n16977), .ZN(n11569) );
  INV_X1 U11843 ( .A(n11571), .ZN(n11570) );
  AOI21_X1 U11844 ( .B1(n16365), .B2(n11574), .A(n11572), .ZN(n11571) );
  INV_X1 U11845 ( .A(n16984), .ZN(n11572) );
  OR2_X1 U11846 ( .A1(n16365), .A2(n11574), .ZN(n11573) );
  AND2_X1 U11847 ( .A1(n11625), .A2(n11623), .ZN(n11622) );
  INV_X1 U11848 ( .A(n17065), .ZN(n11623) );
  AND3_X1 U11849 ( .A1(n13483), .A2(n13482), .A3(n13481), .ZN(n15839) );
  AND2_X1 U11850 ( .A1(n12954), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13002) );
  AND2_X1 U11851 ( .A1(n13236), .A2(n13235), .ZN(n15773) );
  AND2_X1 U11852 ( .A1(n16995), .A2(n11220), .ZN(n16145) );
  NAND2_X1 U11853 ( .A1(n17131), .A2(n11758), .ZN(n11634) );
  AND2_X1 U11854 ( .A1(n17128), .A2(n17345), .ZN(n11758) );
  OR2_X1 U11855 ( .A1(n17129), .A2(n17141), .ZN(n11458) );
  OR2_X1 U11856 ( .A1(n19107), .A2(n16054), .ZN(n17178) );
  NAND2_X1 U11857 ( .A1(n11769), .A2(n11226), .ZN(n11768) );
  NAND2_X1 U11858 ( .A1(n11496), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11493) );
  AOI21_X1 U11859 ( .B1(n17337), .B2(n11199), .A(n17572), .ZN(n11813) );
  NAND2_X1 U11860 ( .A1(n11557), .A2(n11199), .ZN(n11556) );
  NAND2_X1 U11861 ( .A1(n11608), .A2(n11610), .ZN(n17600) );
  INV_X1 U11862 ( .A(n11440), .ZN(n11439) );
  AND2_X1 U11863 ( .A1(n11269), .A2(n15748), .ZN(n11599) );
  NAND2_X1 U11864 ( .A1(n11481), .A2(n11478), .ZN(n11431) );
  NAND2_X1 U11865 ( .A1(n11772), .A2(n14129), .ZN(n11481) );
  NAND2_X1 U11866 ( .A1(n11771), .A2(n14115), .ZN(n11478) );
  OR2_X1 U11867 ( .A1(n14823), .A2(n14822), .ZN(n14858) );
  NAND2_X1 U11868 ( .A1(n11584), .A2(n13393), .ZN(n11587) );
  AND2_X1 U11869 ( .A1(n14880), .A2(n14856), .ZN(n14862) );
  INV_X1 U11870 ( .A(n14853), .ZN(n14855) );
  NAND2_X1 U11871 ( .A1(n14858), .A2(n14857), .ZN(n14861) );
  NAND2_X1 U11872 ( .A1(n14862), .A2(n14861), .ZN(n14882) );
  NOR2_X1 U11873 ( .A1(n19863), .A2(n17805), .ZN(n19824) );
  AND2_X1 U11874 ( .A1(n19863), .A2(n17805), .ZN(n19790) );
  OR2_X1 U11875 ( .A1(n19745), .A2(n19743), .ZN(n19835) );
  NAND2_X1 U11876 ( .A1(n19211), .A2(n17752), .ZN(n17694) );
  NAND2_X1 U11877 ( .A1(n19863), .A2(n19845), .ZN(n19746) );
  AND2_X1 U11878 ( .A1(n15212), .A2(n15211), .ZN(n17645) );
  AOI21_X1 U11879 ( .B1(n18399), .B2(n15996), .A(n15995), .ZN(n21793) );
  NOR2_X1 U11880 ( .A1(n11539), .A2(n11538), .ZN(n11537) );
  AOI211_X1 U11881 ( .C1(n11180), .C2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n18330), .B(n18329), .ZN(n18331) );
  INV_X1 U11882 ( .A(n18333), .ZN(n11538) );
  NOR2_X1 U11883 ( .A1(n21050), .A2(n11647), .ZN(n11646) );
  NOR2_X1 U11884 ( .A1(n18534), .A2(n20986), .ZN(n18555) );
  NOR2_X1 U11885 ( .A1(n18831), .A2(n11529), .ZN(n11528) );
  NAND2_X1 U11886 ( .A1(n21721), .A2(n21655), .ZN(n11529) );
  AOI21_X1 U11887 ( .B1(n18392), .B2(n21479), .A(n18736), .ZN(n11389) );
  INV_X1 U11888 ( .A(n18392), .ZN(n11390) );
  AND2_X1 U11889 ( .A1(n11544), .A2(n11543), .ZN(n21491) );
  NAND2_X1 U11890 ( .A1(n18422), .A2(n11546), .ZN(n11545) );
  INV_X1 U11891 ( .A(n18425), .ZN(n11546) );
  NAND2_X1 U11892 ( .A1(n21648), .A2(n21655), .ZN(n21720) );
  INV_X1 U11893 ( .A(n21795), .ZN(n21648) );
  NOR3_X1 U11894 ( .A1(n16509), .A2(n12734), .A3(n12735), .ZN(n16455) );
  NAND2_X1 U11895 ( .A1(n22215), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16509) );
  AND2_X1 U11896 ( .A1(n14073), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12729) );
  NOR2_X1 U11897 ( .A1(n15410), .A2(n12831), .ZN(n22165) );
  OR2_X1 U11898 ( .A1(n22034), .A2(n22030), .ZN(n22200) );
  OR2_X1 U11899 ( .A1(n13649), .A2(n13650), .ZN(n13651) );
  AND2_X1 U11900 ( .A1(n20506), .A2(n14804), .ZN(n20520) );
  OR2_X1 U11901 ( .A1(n13652), .A2(n11505), .ZN(n11504) );
  INV_X1 U11902 ( .A(n11509), .ZN(n11505) );
  NOR2_X1 U11903 ( .A1(n12938), .A2(n11272), .ZN(n11508) );
  MUX2_X1 U11904 ( .A(n12830), .B(n12829), .S(n12828), .Z(n16804) );
  MUX2_X1 U11905 ( .A(n16440), .B(n12820), .S(n16451), .Z(n12830) );
  AND2_X1 U11906 ( .A1(n14583), .A2(n14582), .ZN(n21993) );
  NOR2_X1 U11907 ( .A1(n15270), .A2(n19219), .ZN(n18968) );
  INV_X1 U11908 ( .A(n19732), .ZN(n19743) );
  NAND2_X1 U11909 ( .A1(n19222), .A2(n14475), .ZN(n17762) );
  OR2_X1 U11910 ( .A1(n16162), .A2(n16161), .ZN(n16163) );
  XNOR2_X1 U11911 ( .A(n16154), .B(n16153), .ZN(n19687) );
  INV_X1 U11912 ( .A(n11591), .ZN(n16154) );
  INV_X1 U11913 ( .A(n19193), .ZN(n17628) );
  AND2_X1 U11914 ( .A1(n14421), .A2(n14386), .ZN(n17633) );
  AND2_X1 U11915 ( .A1(n14421), .A2(n14391), .ZN(n19189) );
  CLKBUF_X1 U11916 ( .A(n13314), .Z(n13315) );
  AOI21_X1 U11917 ( .B1(n21100), .B2(n21099), .A(n21098), .ZN(n11655) );
  INV_X1 U11918 ( .A(n21103), .ZN(n11656) );
  INV_X1 U11919 ( .A(n21023), .ZN(n21096) );
  AOI21_X1 U11920 ( .B1(n21235), .B2(n11405), .A(n11404), .ZN(n11403) );
  INV_X1 U11921 ( .A(P3_EAX_REG_31__SCAN_IN), .ZN(n11404) );
  OR2_X1 U11922 ( .A1(n21306), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n11405) );
  NOR2_X1 U11923 ( .A1(n21253), .A2(n21230), .ZN(n11406) );
  NAND2_X1 U11924 ( .A1(n21238), .A2(n21290), .ZN(n21235) );
  INV_X1 U11925 ( .A(n21242), .ZN(n21239) );
  NOR2_X1 U11926 ( .A1(n21264), .A2(n21263), .ZN(n21262) );
  NOR2_X1 U11927 ( .A1(n21283), .A2(n21282), .ZN(n21281) );
  NAND2_X1 U11928 ( .A1(n21179), .A2(n21305), .ZN(n21290) );
  NOR2_X1 U11929 ( .A1(n21121), .A2(n11417), .ZN(n21294) );
  INV_X1 U11930 ( .A(n11419), .ZN(n11417) );
  NAND2_X1 U11931 ( .A1(n11534), .A2(n11533), .ZN(n11532) );
  NAND2_X1 U11932 ( .A1(n18672), .A2(n21094), .ZN(n11533) );
  NAND2_X1 U11933 ( .A1(n18652), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11534) );
  OAI22_X1 U11934 ( .A1(n21664), .A2(n11597), .B1(n18658), .B2(n11596), .ZN(
        n18641) );
  NAND2_X1 U11935 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U11936 ( .A1(n21630), .A2(n21618), .ZN(n11596) );
  INV_X1 U11937 ( .A(keyinput_1), .ZN(n13662) );
  INV_X1 U11938 ( .A(n13676), .ZN(n11719) );
  AND3_X1 U11939 ( .A1(n13673), .A2(n13672), .A3(n13671), .ZN(n13674) );
  XNOR2_X1 U11940 ( .A(n22413), .B(keyinput_8), .ZN(n11718) );
  OAI21_X1 U11941 ( .B1(n11840), .B2(n13685), .A(n13684), .ZN(n13686) );
  NOR2_X1 U11942 ( .A1(DATAI_22_), .A2(keyinput_10), .ZN(n13685) );
  OR3_X1 U11943 ( .A1(n11846), .A2(n11849), .A3(n13696), .ZN(n13700) );
  OAI21_X1 U11944 ( .B1(n13723), .B2(n13722), .A(n13721), .ZN(n13727) );
  OR2_X1 U11945 ( .A1(n13747), .A2(n11711), .ZN(n11710) );
  NAND2_X1 U11946 ( .A1(n11713), .A2(n11712), .ZN(n11711) );
  NAND2_X1 U11947 ( .A1(n13748), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n11712) );
  INV_X1 U11948 ( .A(n13750), .ZN(n11709) );
  NAND2_X1 U11949 ( .A1(n13752), .A2(n13751), .ZN(n11705) );
  NAND2_X1 U11950 ( .A1(keyinput_52), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n11704) );
  INV_X1 U11951 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n11707) );
  AOI21_X1 U11952 ( .B1(n11708), .B2(n11706), .A(n11703), .ZN(n13759) );
  XNOR2_X1 U11953 ( .A(n11707), .B(keyinput_51), .ZN(n11706) );
  NAND2_X1 U11954 ( .A1(n11705), .A2(n11704), .ZN(n11703) );
  NAND2_X1 U11955 ( .A1(n11710), .A2(n11709), .ZN(n11708) );
  NAND2_X1 U11956 ( .A1(n11692), .A2(n11691), .ZN(n11690) );
  NAND2_X1 U11957 ( .A1(n13765), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n11691) );
  NAND2_X1 U11958 ( .A1(n22191), .A2(keyinput_60), .ZN(n11692) );
  NAND2_X1 U11959 ( .A1(n16526), .A2(keyinput_61), .ZN(n11688) );
  NAND2_X1 U11960 ( .A1(n13766), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n11687) );
  OAI21_X1 U11961 ( .B1(n16548), .B2(keyinput_64), .A(n13767), .ZN(n11684) );
  AOI21_X1 U11962 ( .B1(n11683), .B2(n13775), .A(n13774), .ZN(n13777) );
  OR2_X1 U11963 ( .A1(n11685), .A2(n11684), .ZN(n11683) );
  INV_X1 U11964 ( .A(n11671), .ZN(n11670) );
  OAI21_X1 U11965 ( .B1(n13781), .B2(n13784), .A(n13787), .ZN(n11671) );
  AOI21_X1 U11966 ( .B1(n11670), .B2(n13784), .A(n11329), .ZN(n11669) );
  INV_X1 U11967 ( .A(n13809), .ZN(n11699) );
  NAND2_X1 U11968 ( .A1(n11702), .A2(n11701), .ZN(n11700) );
  NAND2_X1 U11969 ( .A1(n13799), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n11701) );
  NAND2_X1 U11970 ( .A1(n22082), .A2(keyinput_77), .ZN(n11702) );
  AND2_X1 U11971 ( .A1(n13813), .A2(n11695), .ZN(n11694) );
  NOR2_X1 U11972 ( .A1(n13808), .A2(n11696), .ZN(n11695) );
  NOR2_X1 U11973 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_88), .ZN(n11696)
         );
  NAND2_X1 U11974 ( .A1(n11693), .A2(n13826), .ZN(n13831) );
  NAND2_X1 U11975 ( .A1(n11697), .A2(n11694), .ZN(n11693) );
  AOI21_X1 U11976 ( .B1(n12581), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n11303), .ZN(n12542) );
  AOI21_X1 U11977 ( .B1(n12610), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n11320), .ZN(n12613) );
  AOI21_X1 U11978 ( .B1(n12605), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n11317), .ZN(n12562) );
  AOI21_X1 U11979 ( .B1(n12581), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n11300), .ZN(n12477) );
  AOI21_X1 U11980 ( .B1(n12610), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n11297), .ZN(n12485) );
  AOI21_X1 U11981 ( .B1(n12581), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n11268), .ZN(n12135) );
  NAND2_X1 U11982 ( .A1(n11978), .A2(n14895), .ZN(n14535) );
  OAI21_X1 U11983 ( .B1(n12695), .B2(n12703), .A(n12694), .ZN(n12702) );
  NOR2_X1 U11984 ( .A1(n14548), .A2(n12689), .ZN(n12711) );
  AOI22_X1 U11985 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13031) );
  OR2_X1 U11986 ( .A1(n15050), .A2(n15051), .ZN(n15046) );
  NAND2_X1 U11987 ( .A1(n22402), .A2(keyinput_117), .ZN(n11728) );
  NAND2_X1 U11988 ( .A1(n13855), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11727) );
  AOI21_X1 U11989 ( .B1(n12610), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n11296), .ZN(n12227) );
  AOI21_X1 U11990 ( .B1(n12581), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n11301), .ZN(n12502) );
  AOI21_X1 U11991 ( .B1(n12610), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n11319), .ZN(n12453) );
  AOI21_X1 U11992 ( .B1(n12610), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n11298), .ZN(n12401) );
  AOI21_X1 U11993 ( .B1(n12581), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n11302), .ZN(n12424) );
  AOI21_X1 U11994 ( .B1(n12636), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n11304), .ZN(n12382) );
  NOR2_X1 U11995 ( .A1(n11791), .A2(n11793), .ZN(n11790) );
  INV_X1 U11996 ( .A(n12918), .ZN(n11791) );
  INV_X1 U11997 ( .A(n11793), .ZN(n11792) );
  AOI21_X1 U11998 ( .B1(n12610), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n11318), .ZN(n12366) );
  AND2_X1 U11999 ( .A1(n11372), .A2(n11371), .ZN(n12335) );
  AOI21_X1 U12000 ( .B1(n12581), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n11299), .ZN(n12301) );
  CLKBUF_X1 U12001 ( .A(n11908), .Z(n12628) );
  CLKBUF_X1 U12002 ( .A(n12456), .Z(n12636) );
  AOI21_X1 U12003 ( .B1(n12581), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n11281), .ZN(n12096) );
  OR2_X1 U12004 ( .A1(n12118), .A2(n12117), .ZN(n12881) );
  OR2_X1 U12005 ( .A1(n12054), .A2(n12053), .ZN(n12855) );
  INV_X1 U12006 ( .A(n12027), .ZN(n12028) );
  NAND2_X1 U12007 ( .A1(n15074), .A2(n22225), .ZN(n12029) );
  INV_X1 U12008 ( .A(n12705), .ZN(n12696) );
  AOI22_X1 U12009 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11887) );
  NOR2_X1 U12010 ( .A1(n12705), .A2(n12688), .ZN(n12715) );
  AOI22_X1 U12011 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13019) );
  INV_X1 U12012 ( .A(n13022), .ZN(n11582) );
  INV_X1 U12013 ( .A(n14486), .ZN(n11613) );
  INV_X1 U12014 ( .A(n17118), .ZN(n13582) );
  INV_X1 U12015 ( .A(n14392), .ZN(n11614) );
  NAND2_X1 U12016 ( .A1(n14203), .A2(n14205), .ZN(n14208) );
  NOR2_X1 U12017 ( .A1(n14116), .A2(n14100), .ZN(n14101) );
  INV_X1 U12018 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14121) );
  NOR2_X1 U12019 ( .A1(n13388), .A2(n11630), .ZN(n11629) );
  AOI21_X1 U12020 ( .B1(n16211), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n11632), .ZN(n11631) );
  NAND2_X1 U12021 ( .A1(n15280), .A2(n18958), .ZN(n13126) );
  NOR2_X1 U12022 ( .A1(n14404), .A2(n17752), .ZN(n11437) );
  AND2_X1 U12023 ( .A1(n20178), .A2(n19876), .ZN(n13337) );
  NOR2_X1 U12024 ( .A1(n20178), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13357) );
  AOI22_X1 U12025 ( .A1(n16399), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11195), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U12026 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13081) );
  INV_X1 U12027 ( .A(n13099), .ZN(n13100) );
  AOI22_X1 U12028 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13036) );
  AND2_X1 U12029 ( .A1(n19891), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14218) );
  NOR2_X1 U12030 ( .A1(n21156), .A2(n18358), .ZN(n18386) );
  INV_X1 U12031 ( .A(n18407), .ZN(n18405) );
  NAND2_X1 U12032 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11521) );
  INV_X1 U12033 ( .A(n15023), .ZN(n11522) );
  NAND2_X1 U12034 ( .A1(n11979), .A2(n16591), .ZN(n11401) );
  NAND2_X1 U12035 ( .A1(n11253), .A2(n14540), .ZN(n11399) );
  NAND2_X1 U12036 ( .A1(n14559), .A2(n14776), .ZN(n11400) );
  AOI21_X1 U12037 ( .B1(n11730), .B2(n11729), .A(n11726), .ZN(n13856) );
  AOI22_X1 U12038 ( .A1(n13854), .A2(n13853), .B1(keyinput_116), .B2(
        P1_EAX_REG_31__SCAN_IN), .ZN(n11729) );
  NAND2_X1 U12039 ( .A1(n11728), .A2(n11727), .ZN(n11726) );
  NOR2_X1 U12040 ( .A1(n14764), .A2(n15127), .ZN(n14548) );
  INV_X1 U12041 ( .A(n12943), .ZN(n14554) );
  AOI21_X1 U12042 ( .B1(n11959), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n11251), .ZN(n11917) );
  NAND2_X1 U12043 ( .A1(n11913), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11942) );
  AOI21_X1 U12044 ( .B1(n12635), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n11305), .ZN(n12273) );
  NOR2_X1 U12045 ( .A1(n16682), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11780) );
  INV_X1 U12046 ( .A(n20476), .ZN(n11750) );
  NAND2_X1 U12047 ( .A1(n20545), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12925) );
  INV_X1 U12048 ( .A(n16848), .ZN(n11752) );
  NOR2_X1 U12049 ( .A1(n15941), .A2(n11754), .ZN(n11753) );
  INV_X1 U12050 ( .A(n15920), .ZN(n11754) );
  OR2_X1 U12051 ( .A1(n20552), .A2(n12920), .ZN(n16768) );
  OR2_X1 U12052 ( .A1(n20552), .A2(n21889), .ZN(n16771) );
  NAND2_X1 U12053 ( .A1(n11747), .A2(n15479), .ZN(n11746) );
  INV_X1 U12054 ( .A(n15358), .ZN(n11747) );
  NAND2_X1 U12055 ( .A1(n15304), .A2(n12820), .ZN(n12819) );
  INV_X1 U12056 ( .A(n12906), .ZN(n14533) );
  OR2_X1 U12057 ( .A1(n12073), .A2(n12072), .ZN(n12856) );
  INV_X1 U12058 ( .A(n12909), .ZN(n12146) );
  NAND2_X1 U12059 ( .A1(n12082), .A2(n12907), .ZN(n12168) );
  NAND2_X1 U12060 ( .A1(n11513), .A2(n11512), .ZN(n12200) );
  OAI21_X1 U12061 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12004), .A(
        n12003), .ZN(n12005) );
  AOI21_X1 U12062 ( .B1(n21858), .B2(n22224), .A(n22228), .ZN(n15143) );
  NOR2_X1 U12063 ( .A1(n11661), .A2(n11664), .ZN(n11660) );
  INV_X1 U12064 ( .A(n16048), .ZN(n11664) );
  INV_X1 U12065 ( .A(n11662), .ZN(n11661) );
  NOR2_X1 U12066 ( .A1(n11663), .A2(n16032), .ZN(n11662) );
  AND2_X1 U12067 ( .A1(n14352), .A2(n14353), .ZN(n14361) );
  AND2_X1 U12068 ( .A1(n14344), .A2(n14345), .ZN(n14352) );
  NOR2_X1 U12069 ( .A1(n14350), .A2(n14348), .ZN(n14344) );
  NOR2_X1 U12070 ( .A1(n14337), .A2(n14336), .ZN(n11652) );
  NAND2_X1 U12071 ( .A1(n13154), .A2(n13153), .ZN(n13158) );
  NOR2_X1 U12072 ( .A1(n14710), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13355) );
  NOR2_X2 U12073 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13329) );
  NAND2_X1 U12074 ( .A1(n11803), .A2(n11804), .ZN(n13130) );
  NAND2_X1 U12075 ( .A1(n11802), .A2(n13121), .ZN(n13131) );
  AOI22_X1 U12076 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n13042), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13050) );
  INV_X1 U12077 ( .A(n16994), .ZN(n11574) );
  NOR2_X1 U12078 ( .A1(n11627), .A2(n11626), .ZN(n11625) );
  INV_X1 U12079 ( .A(n17077), .ZN(n11626) );
  NAND2_X1 U12080 ( .A1(n11628), .A2(n16928), .ZN(n11627) );
  INV_X1 U12081 ( .A(n17091), .ZN(n11628) );
  INV_X1 U12082 ( .A(n17038), .ZN(n11578) );
  AND2_X1 U12083 ( .A1(n13109), .A2(n20237), .ZN(n14412) );
  INV_X1 U12084 ( .A(n16347), .ZN(n16324) );
  AND2_X1 U12085 ( .A1(n19175), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14701) );
  NOR2_X1 U12086 ( .A1(n17158), .A2(n11716), .ZN(n11715) );
  INV_X1 U12087 ( .A(n14445), .ZN(n11731) );
  NAND2_X1 U12088 ( .A1(n17141), .A2(n17345), .ZN(n11761) );
  INV_X1 U12089 ( .A(n11468), .ZN(n11464) );
  NAND2_X1 U12090 ( .A1(n17169), .A2(n16057), .ZN(n11468) );
  INV_X1 U12091 ( .A(n17169), .ZN(n11467) );
  AND2_X1 U12092 ( .A1(n17022), .A2(n17017), .ZN(n11737) );
  INV_X1 U12093 ( .A(n11226), .ZN(n11763) );
  NAND2_X1 U12094 ( .A1(n11614), .A2(n13582), .ZN(n17120) );
  NAND2_X1 U12095 ( .A1(n11621), .A2(n15908), .ZN(n11620) );
  INV_X1 U12096 ( .A(n15924), .ZN(n11621) );
  INV_X1 U12097 ( .A(n15812), .ZN(n11619) );
  AND2_X1 U12098 ( .A1(n11311), .A2(n14328), .ZN(n11774) );
  INV_X1 U12099 ( .A(n11774), .ZN(n11434) );
  OR2_X1 U12100 ( .A1(n15911), .A2(n16060), .ZN(n14341) );
  NOR2_X1 U12101 ( .A1(n14208), .A2(n16060), .ZN(n14209) );
  XNOR2_X1 U12102 ( .A(n14208), .B(n16060), .ZN(n14206) );
  NAND2_X1 U12103 ( .A1(n17611), .A2(n17610), .ZN(n11435) );
  INV_X1 U12104 ( .A(n11445), .ZN(n11444) );
  NAND2_X1 U12105 ( .A1(n11357), .A2(n14141), .ZN(n14142) );
  NAND2_X1 U12106 ( .A1(n13164), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13146) );
  NAND2_X1 U12107 ( .A1(n13143), .A2(n14219), .ZN(n11488) );
  AND2_X1 U12109 ( .A1(n13115), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U12110 ( .A1(n11564), .A2(n14249), .ZN(n14388) );
  NAND2_X1 U12111 ( .A1(n11247), .A2(n14378), .ZN(n11564) );
  NOR2_X1 U12112 ( .A1(n13375), .A2(n13374), .ZN(n14133) );
  AOI21_X1 U12113 ( .B1(n14808), .B2(n14812), .A(n14811), .ZN(n14813) );
  INV_X1 U12114 ( .A(n14404), .ZN(n13115) );
  NAND2_X1 U12115 ( .A1(n13108), .A2(n20237), .ZN(n14416) );
  AOI22_X1 U12116 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13070) );
  AOI22_X1 U12117 ( .A1(n11193), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16400), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U12118 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13073) );
  NOR2_X1 U12119 ( .A1(n14844), .A2(n14808), .ZN(n14107) );
  AND2_X1 U12120 ( .A1(n15963), .A2(n14093), .ZN(n14106) );
  AND2_X1 U12121 ( .A1(n15963), .A2(n14088), .ZN(n14103) );
  NOR2_X1 U12122 ( .A1(n14966), .A2(n14967), .ZN(n14986) );
  INV_X1 U12123 ( .A(n21341), .ZN(n11517) );
  OR3_X1 U12124 ( .A1(n21342), .A2(n21361), .A3(n20687), .ZN(n11852) );
  INV_X1 U12125 ( .A(n18332), .ZN(n11539) );
  NOR2_X1 U12126 ( .A1(n18428), .A2(n11638), .ZN(n11637) );
  INV_X1 U12127 ( .A(n20845), .ZN(n11657) );
  AND2_X1 U12128 ( .A1(n18739), .A2(n11287), .ZN(n11659) );
  NAND2_X1 U12129 ( .A1(n18708), .A2(n18431), .ZN(n18475) );
  NAND2_X1 U12130 ( .A1(n18773), .A2(n18418), .ZN(n18420) );
  NOR2_X1 U12131 ( .A1(n15031), .A2(n11410), .ZN(n11409) );
  INV_X1 U12132 ( .A(n21122), .ZN(n21307) );
  NAND2_X1 U12133 ( .A1(n11519), .A2(n11424), .ZN(n21117) );
  INV_X1 U12134 ( .A(n20638), .ZN(n11424) );
  INV_X1 U12135 ( .A(n11973), .ZN(n11972) );
  INV_X1 U12136 ( .A(n14785), .ZN(n11966) );
  INV_X1 U12137 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n22037) );
  INV_X1 U12138 ( .A(n12059), .ZN(n12060) );
  NAND2_X1 U12139 ( .A1(n14558), .A2(n11805), .ZN(n14783) );
  AND2_X1 U12140 ( .A1(n15592), .A2(n11179), .ZN(n11805) );
  AOI21_X1 U12141 ( .B1(n15126), .B2(n22405), .A(n17713), .ZN(n20381) );
  INV_X1 U12142 ( .A(n22813), .ZN(n14766) );
  AND2_X1 U12143 ( .A1(n12656), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12727) );
  OR2_X1 U12144 ( .A1(n12603), .A2(n12602), .ZN(n16462) );
  CLKBUF_X1 U12145 ( .A(n16473), .Z(n16486) );
  AND2_X1 U12146 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n12555), .ZN(
        n12556) );
  AND2_X1 U12147 ( .A1(n12657), .A2(n16715), .ZN(n12536) );
  NOR2_X1 U12148 ( .A1(n12515), .A2(n16719), .ZN(n12516) );
  NOR2_X1 U12149 ( .A1(n12467), .A2(n16730), .ZN(n12468) );
  NAND2_X1 U12150 ( .A1(n12468), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12515) );
  AND2_X1 U12151 ( .A1(n12471), .A2(n12470), .ZN(n16512) );
  NOR2_X1 U12152 ( .A1(n12432), .A2(n16737), .ZN(n12414) );
  AND2_X1 U12153 ( .A1(n12399), .A2(n12398), .ZN(n16647) );
  NOR2_X1 U12154 ( .A1(n12359), .A2(n16762), .ZN(n12360) );
  NAND2_X1 U12155 ( .A1(n12360), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12395) );
  OR2_X1 U12156 ( .A1(n12329), .A2(n22123), .ZN(n12359) );
  NOR2_X1 U12157 ( .A1(n11818), .A2(n11817), .ZN(n11816) );
  INV_X1 U12158 ( .A(n15879), .ZN(n11817) );
  NOR2_X1 U12159 ( .A1(n12311), .A2(n12310), .ZN(n12315) );
  NOR2_X1 U12160 ( .A1(n12282), .A2(n14072), .ZN(n12283) );
  NAND2_X1 U12161 ( .A1(n12253), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12282) );
  NOR2_X1 U12162 ( .A1(n12239), .A2(n15488), .ZN(n12253) );
  CLKBUF_X1 U12163 ( .A(n14062), .Z(n14063) );
  INV_X1 U12164 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15488) );
  NAND2_X1 U12165 ( .A1(n12218), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12239) );
  NAND2_X1 U12166 ( .A1(n12155), .A2(n12154), .ZN(n15424) );
  NOR2_X1 U12167 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  AOI21_X1 U12168 ( .B1(n12891), .B2(n12338), .A(n12224), .ZN(n15297) );
  AOI21_X1 U12169 ( .B1(n12880), .B2(n12338), .A(n12161), .ZN(n15130) );
  NAND2_X1 U12170 ( .A1(n12214), .A2(n12213), .ZN(n15298) );
  INV_X1 U12171 ( .A(n15130), .ZN(n12214) );
  INV_X1 U12172 ( .A(n14952), .ZN(n12213) );
  OR2_X1 U12173 ( .A1(n17669), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12947) );
  INV_X1 U12174 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11788) );
  NAND2_X1 U12175 ( .A1(n16567), .A2(n11294), .ZN(n16505) );
  NAND2_X1 U12176 ( .A1(n16567), .A2(n11292), .ZN(n20479) );
  NAND2_X1 U12177 ( .A1(n16567), .A2(n16566), .ZN(n20477) );
  NOR3_X1 U12178 ( .A1(n16583), .A2(n11295), .A3(n11743), .ZN(n16575) );
  NOR2_X1 U12179 ( .A1(n16583), .A2(n14578), .ZN(n16550) );
  NAND2_X1 U12180 ( .A1(n11795), .A2(n11796), .ZN(n16748) );
  OR2_X1 U12181 ( .A1(n15778), .A2(n11797), .ZN(n11795) );
  OR2_X1 U12182 ( .A1(n16580), .A2(n16581), .ZN(n16583) );
  OR2_X1 U12183 ( .A1(n20552), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n20526) );
  AND2_X1 U12184 ( .A1(n15921), .A2(n11751), .ZN(n20467) );
  AND2_X1 U12185 ( .A1(n11211), .A2(n12782), .ZN(n11751) );
  NAND2_X1 U12186 ( .A1(n15921), .A2(n11211), .ZN(n16845) );
  NAND2_X1 U12187 ( .A1(n15921), .A2(n11753), .ZN(n16847) );
  AND2_X1 U12188 ( .A1(n12771), .A2(n12770), .ZN(n15881) );
  OR2_X1 U12189 ( .A1(n14069), .A2(n14070), .ZN(n15882) );
  NOR2_X1 U12190 ( .A1(n15525), .A2(n15487), .ZN(n15580) );
  AOI21_X1 U12191 ( .B1(n15716), .B2(n11785), .A(n11249), .ZN(n11784) );
  INV_X1 U12192 ( .A(n12897), .ZN(n11785) );
  OR2_X1 U12193 ( .A1(n15523), .A2(n11850), .ZN(n15525) );
  OR2_X1 U12194 ( .A1(n15359), .A2(n11746), .ZN(n15478) );
  NOR2_X1 U12195 ( .A1(n15359), .A2(n15358), .ZN(n15480) );
  NAND2_X1 U12196 ( .A1(n12750), .A2(n12749), .ZN(n15359) );
  INV_X1 U12197 ( .A(n15353), .ZN(n12750) );
  AND2_X1 U12198 ( .A1(n14573), .A2(n14572), .ZN(n21920) );
  NAND2_X1 U12199 ( .A1(n14907), .A2(n14906), .ZN(n15353) );
  NOR2_X1 U12200 ( .A1(n22015), .A2(n14900), .ZN(n21922) );
  XNOR2_X1 U12201 ( .A(n12740), .B(n12741), .ZN(n16184) );
  INV_X1 U12202 ( .A(n14803), .ZN(n11364) );
  XNOR2_X1 U12203 ( .A(n15101), .B(n15133), .ZN(n15080) );
  AND2_X1 U12204 ( .A1(n14558), .A2(n15391), .ZN(n11806) );
  OR2_X1 U12205 ( .A1(n16178), .A2(n15287), .ZN(n15461) );
  NOR2_X1 U12206 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15143), .ZN(n22626) );
  AND2_X1 U12207 ( .A1(n16178), .A2(n15112), .ZN(n22427) );
  OR3_X1 U12208 ( .A1(n22464), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n15143), 
        .ZN(n22629) );
  AND2_X1 U12209 ( .A1(n15100), .A2(n15099), .ZN(n17739) );
  NAND2_X1 U12210 ( .A1(n11376), .A2(n11276), .ZN(n16422) );
  INV_X1 U12211 ( .A(n11377), .ZN(n11376) );
  AOI21_X1 U12212 ( .B1(n12722), .B2(n11378), .A(n12723), .ZN(n11377) );
  NOR2_X1 U12213 ( .A1(n11649), .A2(n16058), .ZN(n11648) );
  INV_X1 U12214 ( .A(n11650), .ZN(n11649) );
  NOR2_X1 U12215 ( .A1(n15851), .A2(n15850), .ZN(n15852) );
  NAND2_X1 U12216 ( .A1(n12988), .A2(n11212), .ZN(n12992) );
  NAND2_X1 U12217 ( .A1(n11652), .A2(n11306), .ZN(n14350) );
  NAND2_X1 U12218 ( .A1(n12978), .A2(n11208), .ZN(n12987) );
  INV_X1 U12219 ( .A(n11652), .ZN(n14342) );
  NAND2_X1 U12220 ( .A1(n12978), .A2(n11680), .ZN(n12974) );
  INV_X1 U12221 ( .A(n14314), .ZN(n13628) );
  NAND2_X1 U12222 ( .A1(n14321), .A2(n11231), .ZN(n14326) );
  INV_X1 U12223 ( .A(n14088), .ZN(n14093) );
  NAND2_X1 U12224 ( .A1(n11624), .A2(n11625), .ZN(n17064) );
  XNOR2_X1 U12225 ( .A(n17013), .B(n16305), .ZN(n17010) );
  NAND2_X1 U12226 ( .A1(n17015), .A2(n17014), .ZN(n17013) );
  NAND2_X1 U12227 ( .A1(n15902), .A2(n11293), .ZN(n17042) );
  AND2_X1 U12228 ( .A1(n19982), .A2(n14710), .ZN(n14747) );
  NOR2_X1 U12229 ( .A1(n11617), .A2(n11616), .ZN(n11615) );
  INV_X1 U12230 ( .A(n15805), .ZN(n11616) );
  AND2_X1 U12231 ( .A1(n14880), .A2(n14879), .ZN(n14881) );
  AND2_X1 U12232 ( .A1(n14734), .A2(n18957), .ZN(n17823) );
  XNOR2_X1 U12233 ( .A(n11665), .B(n12959), .ZN(n16172) );
  NAND2_X1 U12234 ( .A1(n13002), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11665) );
  AND2_X1 U12235 ( .A1(n11219), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11714) );
  INV_X1 U12236 ( .A(n12954), .ZN(n12958) );
  NAND2_X1 U12237 ( .A1(n12996), .A2(n11715), .ZN(n12998) );
  NOR2_X1 U12238 ( .A1(n12965), .A2(n17183), .ZN(n12996) );
  INV_X1 U12239 ( .A(n12966), .ZN(n11667) );
  NAND2_X1 U12240 ( .A1(n11666), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12965) );
  AND2_X1 U12241 ( .A1(n13247), .A2(n13246), .ZN(n15888) );
  INV_X1 U12242 ( .A(n11810), .ZN(n11809) );
  AND2_X1 U12243 ( .A1(n13229), .A2(n13228), .ZN(n15701) );
  AND2_X1 U12244 ( .A1(n12988), .A2(n11271), .ZN(n12990) );
  NOR2_X1 U12245 ( .A1(n12987), .A2(n17277), .ZN(n12988) );
  AND2_X1 U12246 ( .A1(n13214), .A2(n13213), .ZN(n15334) );
  AND2_X1 U12247 ( .A1(n15178), .A2(n11237), .ZN(n15446) );
  NAND2_X1 U12248 ( .A1(n15178), .A2(n11227), .ZN(n15335) );
  NAND2_X1 U12249 ( .A1(n15178), .A2(n15177), .ZN(n15188) );
  INV_X1 U12250 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17318) );
  NAND2_X1 U12251 ( .A1(n13194), .A2(n13193), .ZN(n15118) );
  AND2_X1 U12252 ( .A1(n13199), .A2(n13198), .ZN(n15117) );
  NOR2_X1 U12253 ( .A1(n15755), .A2(n11722), .ZN(n11721) );
  NOR2_X1 U12254 ( .A1(n16112), .A2(n17141), .ZN(n11561) );
  NAND2_X1 U12255 ( .A1(n13592), .A2(n13591), .ZN(n17101) );
  INV_X1 U12256 ( .A(n17409), .ZN(n13592) );
  NOR2_X1 U12257 ( .A1(n17101), .A2(n17091), .ZN(n17090) );
  OR3_X1 U12258 ( .A1(n17563), .A2(n17428), .A3(n17422), .ZN(n17413) );
  AND2_X1 U12259 ( .A1(n13260), .A2(n13259), .ZN(n17029) );
  NAND2_X1 U12260 ( .A1(n16041), .A2(n11240), .ZN(n11472) );
  NAND2_X1 U12261 ( .A1(n14472), .A2(n14473), .ZN(n17036) );
  NOR2_X1 U12262 ( .A1(n17316), .A2(n17422), .ZN(n17199) );
  OR2_X1 U12263 ( .A1(n15787), .A2(n15788), .ZN(n15851) );
  AND2_X1 U12264 ( .A1(n13223), .A2(n13222), .ZN(n15417) );
  AND2_X1 U12265 ( .A1(n11237), .A2(n15445), .ZN(n11733) );
  NAND2_X1 U12266 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11810) );
  NAND2_X1 U12267 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11498) );
  NOR2_X1 U12268 ( .A1(n11605), .A2(n11604), .ZN(n11603) );
  INV_X1 U12269 ( .A(n17558), .ZN(n11604) );
  INV_X1 U12270 ( .A(n11606), .ZN(n11605) );
  OR2_X1 U12271 ( .A1(n17332), .A2(n11201), .ZN(n17321) );
  OR2_X1 U12272 ( .A1(n19005), .A2(n14335), .ZN(n17322) );
  NAND2_X1 U12273 ( .A1(n17321), .A2(n14328), .ZN(n17327) );
  NOR2_X1 U12274 ( .A1(n17316), .A2(n17532), .ZN(n17315) );
  XOR2_X1 U12275 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n14206), .Z(
        n17337) );
  AND2_X1 U12276 ( .A1(n14197), .A2(n14196), .ZN(n14198) );
  AND2_X1 U12277 ( .A1(n14434), .A2(n14433), .ZN(n17614) );
  INV_X1 U12278 ( .A(n15326), .ZN(n11600) );
  INV_X1 U12279 ( .A(n14826), .ZN(n11586) );
  AND2_X1 U12280 ( .A1(n13183), .A2(n13182), .ZN(n15740) );
  NAND2_X1 U12281 ( .A1(n11352), .A2(n14280), .ZN(n11351) );
  NAND2_X1 U12282 ( .A1(n14309), .A2(n18973), .ZN(n15736) );
  NAND2_X1 U12283 ( .A1(n11205), .A2(n11242), .ZN(n11446) );
  NAND2_X1 U12284 ( .A1(n14287), .A2(n15729), .ZN(n11447) );
  OAI21_X1 U12285 ( .B1(n14286), .B2(n14287), .A(n15729), .ZN(n15644) );
  XNOR2_X1 U12286 ( .A(n14757), .B(n13363), .ZN(n14943) );
  CLKBUF_X1 U12287 ( .A(n13326), .Z(n13327) );
  OR2_X1 U12288 ( .A1(n14240), .A2(n14238), .ZN(n17641) );
  NOR2_X1 U12289 ( .A1(n13116), .A2(n13113), .ZN(n13117) );
  INV_X1 U12290 ( .A(n19865), .ZN(n19910) );
  NAND3_X1 U12291 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19717), .A3(n19910), 
        .ZN(n20081) );
  NAND3_X1 U12292 ( .A1(n19718), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19910), 
        .ZN(n20080) );
  OR2_X1 U12293 ( .A1(n20234), .A2(n19908), .ZN(n19865) );
  NAND2_X1 U12294 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19914), .ZN(n20236) );
  INV_X1 U12295 ( .A(n20081), .ZN(n20240) );
  INV_X1 U12296 ( .A(n20080), .ZN(n20241) );
  INV_X1 U12297 ( .A(n19801), .ZN(n19846) );
  NOR3_X1 U12298 ( .A1(n17680), .A2(n20638), .A3(n21327), .ZN(n21792) );
  NAND2_X1 U12299 ( .A1(n20953), .A2(n20952), .ZN(n20968) );
  NAND2_X1 U12300 ( .A1(n11641), .A2(n20925), .ZN(n11640) );
  NOR2_X1 U12301 ( .A1(n21248), .A2(n18906), .ZN(n11416) );
  NOR2_X1 U12302 ( .A1(n11387), .A2(n11386), .ZN(n11385) );
  INV_X1 U12303 ( .A(n18318), .ZN(n11386) );
  NOR2_X1 U12304 ( .A1(n21296), .A2(n11420), .ZN(n11419) );
  NOR2_X1 U12305 ( .A1(n11415), .A2(n11412), .ZN(n11411) );
  NOR2_X1 U12306 ( .A1(n20639), .A2(n17679), .ZN(n18888) );
  NAND2_X1 U12307 ( .A1(n18589), .A2(n11213), .ZN(n18632) );
  NAND2_X1 U12308 ( .A1(n18589), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18593) );
  NOR2_X1 U12309 ( .A1(n21694), .A2(n18552), .ZN(n18588) );
  NAND2_X1 U12310 ( .A1(n21389), .A2(n18544), .ZN(n18552) );
  NAND2_X1 U12311 ( .A1(n18499), .A2(n11853), .ZN(n18534) );
  AND2_X1 U12312 ( .A1(n11637), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11636) );
  NAND2_X1 U12313 ( .A1(n18674), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18429) );
  AND3_X1 U12314 ( .A1(n18750), .A2(n11658), .A3(n11657), .ZN(n18687) );
  NAND2_X1 U12315 ( .A1(n18750), .A2(n11658), .ZN(n18472) );
  AND2_X1 U12316 ( .A1(n18750), .A2(n11659), .ZN(n20835) );
  XNOR2_X1 U12317 ( .A(n18420), .B(n11535), .ZN(n18763) );
  INV_X1 U12318 ( .A(n18419), .ZN(n11535) );
  NAND2_X1 U12319 ( .A1(n18763), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18762) );
  AND2_X1 U12320 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18792) );
  NOR2_X1 U12321 ( .A1(n11595), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11594) );
  INV_X1 U12322 ( .A(n18637), .ZN(n11595) );
  INV_X1 U12323 ( .A(n18552), .ZN(n21676) );
  NAND2_X1 U12324 ( .A1(n18438), .A2(n11859), .ZN(n18669) );
  NOR2_X1 U12325 ( .A1(n18435), .A2(n18436), .ZN(n18492) );
  NAND2_X1 U12326 ( .A1(n11544), .A2(n11542), .ZN(n18683) );
  AND2_X1 U12327 ( .A1(n11543), .A2(n21518), .ZN(n11542) );
  NOR2_X1 U12328 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21649), .ZN(
        n18736) );
  XNOR2_X1 U12329 ( .A(n18453), .B(n18390), .ZN(n18749) );
  NAND2_X1 U12330 ( .A1(n18749), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18748) );
  NAND2_X1 U12331 ( .A1(n11229), .A2(n11381), .ZN(n18778) );
  NAND2_X1 U12332 ( .A1(n18786), .A2(n11382), .ZN(n11381) );
  NAND2_X1 U12333 ( .A1(n11588), .A2(n11383), .ZN(n11379) );
  INV_X1 U12334 ( .A(n21793), .ZN(n21797) );
  AOI211_X1 U12335 ( .C1(n15056), .C2(n15055), .A(n18399), .B(n15995), .ZN(
        n21790) );
  NAND2_X1 U12336 ( .A1(n21310), .A2(n21324), .ZN(n20687) );
  NOR2_X1 U12337 ( .A1(n15992), .A2(n15978), .ZN(n15985) );
  NAND2_X1 U12338 ( .A1(n18394), .A2(n18393), .ZN(n21728) );
  NOR2_X1 U12339 ( .A1(n15043), .A2(n15042), .ZN(n19455) );
  AND2_X1 U12340 ( .A1(n11516), .A2(n11515), .ZN(n21787) );
  NAND2_X1 U12341 ( .A1(n21788), .A2(n21790), .ZN(n11515) );
  NAND2_X1 U12342 ( .A1(n21648), .A2(n21794), .ZN(n11516) );
  CLKBUF_X1 U12343 ( .A(n14712), .Z(n19718) );
  AND2_X1 U12344 ( .A1(n11972), .A2(n11954), .ZN(n22810) );
  AND2_X1 U12345 ( .A1(n22199), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n22215) );
  NAND2_X1 U12346 ( .A1(n16527), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n22190) );
  NOR2_X1 U12347 ( .A1(n22191), .A2(n22190), .ZN(n22199) );
  NOR2_X1 U12348 ( .A1(n22181), .A2(n16729), .ZN(n16527) );
  NAND2_X1 U12349 ( .A1(n22121), .A2(n16515), .ZN(n22181) );
  NOR2_X1 U12350 ( .A1(n22103), .A2(n16516), .ZN(n22121) );
  NAND2_X1 U12351 ( .A1(n14075), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22152) );
  INV_X1 U12352 ( .A(n22200), .ZN(n22189) );
  INV_X1 U12353 ( .A(n22209), .ZN(n22172) );
  NAND2_X1 U12354 ( .A1(n14075), .A2(n14074), .ZN(n22203) );
  NOR2_X1 U12355 ( .A1(n22055), .A2(n22056), .ZN(n22072) );
  AND2_X1 U12356 ( .A1(n21860), .A2(n11284), .ZN(n22034) );
  INV_X1 U12357 ( .A(n14075), .ZN(n22030) );
  XNOR2_X1 U12359 ( .A(n16442), .B(n16441), .ZN(n16815) );
  INV_X1 U12360 ( .A(n20483), .ZN(n20489) );
  INV_X1 U12361 ( .A(n20480), .ZN(n20488) );
  INV_X1 U12362 ( .A(DATAI_24_), .ZN(n22413) );
  AND2_X1 U12363 ( .A1(n16659), .A2(n14897), .ZN(n15948) );
  INV_X1 U12364 ( .A(n15948), .ZN(n15954) );
  CLKBUF_X1 U12365 ( .A(n20393), .Z(n20399) );
  CLKBUF_X1 U12366 ( .A(n20390), .Z(n21862) );
  XNOR2_X1 U12367 ( .A(n11825), .B(n12661), .ZN(n16590) );
  INV_X1 U12368 ( .A(n11825), .ZN(n16431) );
  OR2_X1 U12369 ( .A1(n16618), .A2(n16499), .ZN(n22210) );
  AOI21_X1 U12370 ( .B1(n20551), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20514), .ZN(n11394) );
  OR2_X1 U12371 ( .A1(n16465), .A2(n16464), .ZN(n21984) );
  XNOR2_X1 U12372 ( .A(n16866), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20513) );
  NAND2_X1 U12373 ( .A1(n15776), .A2(n11396), .ZN(n21879) );
  OR2_X1 U12374 ( .A1(n15778), .A2(n15777), .ZN(n11396) );
  NAND2_X1 U12375 ( .A1(n11787), .A2(n12897), .ZN(n15717) );
  NAND2_X1 U12376 ( .A1(n15606), .A2(n15605), .ZN(n11787) );
  OR2_X1 U12377 ( .A1(n15285), .A2(n15172), .ZN(n15499) );
  CLKBUF_X1 U12378 ( .A(n15080), .Z(n22041) );
  AND2_X1 U12379 ( .A1(n22428), .A2(n22427), .ZN(n22749) );
  OAI21_X1 U12380 ( .B1(n15290), .B2(n22698), .A(n22509), .ZN(n22700) );
  NOR2_X1 U12381 ( .A1(n22411), .A2(n22410), .ZN(n22522) );
  INV_X1 U12382 ( .A(n22550), .ZN(n22552) );
  INV_X1 U12383 ( .A(n22585), .ZN(n22593) );
  INV_X1 U12384 ( .A(n22620), .ZN(n22622) );
  INV_X1 U12385 ( .A(n22660), .ZN(n22667) );
  INV_X1 U12386 ( .A(n22685), .ZN(n15638) );
  INV_X1 U12387 ( .A(n22804), .ZN(n15639) );
  INV_X1 U12388 ( .A(n22728), .ZN(n22732) );
  AND2_X1 U12389 ( .A1(n15436), .A2(n15379), .ZN(n22800) );
  INV_X1 U12390 ( .A(n22787), .ZN(n22799) );
  NOR2_X1 U12391 ( .A1(n16422), .A2(n22464), .ZN(n22228) );
  NAND2_X1 U12392 ( .A1(n11672), .A2(n11673), .ZN(n16914) );
  AOI21_X1 U12393 ( .B1(n11674), .B2(n19134), .A(n19134), .ZN(n11673) );
  NAND2_X1 U12394 ( .A1(n11676), .A2(n11677), .ZN(n19166) );
  OR2_X1 U12395 ( .A1(n19147), .A2(n19134), .ZN(n11676) );
  NAND2_X1 U12396 ( .A1(n19146), .A2(n19032), .ZN(n19168) );
  NAND2_X1 U12397 ( .A1(n16949), .A2(n11724), .ZN(n19065) );
  NAND2_X1 U12398 ( .A1(n12963), .A2(n11725), .ZN(n11724) );
  INV_X1 U12399 ( .A(n16960), .ZN(n11725) );
  INV_X1 U12400 ( .A(n19131), .ZN(n19163) );
  AND2_X1 U12401 ( .A1(n13644), .A2(n13643), .ZN(n19156) );
  INV_X1 U12402 ( .A(n19158), .ZN(n19108) );
  INV_X1 U12403 ( .A(n19183), .ZN(n15963) );
  AND2_X1 U12404 ( .A1(n13644), .A2(n13642), .ZN(n19131) );
  INV_X1 U12405 ( .A(n11739), .ZN(n14380) );
  NAND2_X1 U12406 ( .A1(n11835), .A2(n15421), .ZN(n15704) );
  NAND2_X1 U12407 ( .A1(n15330), .A2(n15329), .ZN(n16011) );
  AND2_X1 U12408 ( .A1(n14709), .A2(n18966), .ZN(n17044) );
  NOR2_X1 U12409 ( .A1(n11857), .A2(n11591), .ZN(n16115) );
  NAND2_X1 U12410 ( .A1(n11576), .A2(n11575), .ZN(n16409) );
  NAND2_X1 U12411 ( .A1(n11567), .A2(n11571), .ZN(n16979) );
  AND2_X1 U12412 ( .A1(n17060), .A2(n17059), .ZN(n19160) );
  INV_X1 U12413 ( .A(n20223), .ZN(n17123) );
  AND2_X1 U12414 ( .A1(n15849), .A2(n19718), .ZN(n20225) );
  AND2_X1 U12415 ( .A1(n15849), .A2(n19717), .ZN(n20224) );
  NOR2_X1 U12416 ( .A1(n20123), .A2(n20169), .ZN(n19979) );
  INV_X1 U12417 ( .A(n20228), .ZN(n20123) );
  AND2_X1 U12418 ( .A1(n19929), .A2(n13338), .ZN(n20169) );
  INV_X1 U12419 ( .A(n19929), .ZN(n20221) );
  NOR2_X1 U12420 ( .A1(n17823), .A2(n17851), .ZN(n17836) );
  CLKBUF_X1 U12422 ( .A(n17841), .Z(n17851) );
  CLKBUF_X1 U12423 ( .A(n14678), .Z(n14682) );
  NAND2_X1 U12424 ( .A1(n11356), .A2(n11493), .ZN(n11355) );
  NAND2_X1 U12425 ( .A1(n11809), .A2(n11326), .ZN(n11807) );
  INV_X1 U12426 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17338) );
  INV_X1 U12427 ( .A(n17770), .ZN(n17782) );
  CLKBUF_X1 U12428 ( .A(n19040), .Z(n19047) );
  AND2_X1 U12429 ( .A1(n17762), .A2(n14476), .ZN(n17784) );
  AND2_X1 U12430 ( .A1(n17762), .A2(n14626), .ZN(n17754) );
  INV_X1 U12431 ( .A(n17774), .ZN(n17785) );
  INV_X1 U12432 ( .A(n17784), .ZN(n17773) );
  XNOR2_X1 U12433 ( .A(n11633), .B(n16077), .ZN(n16104) );
  OAI21_X1 U12434 ( .B1(n11200), .B2(n11457), .A(n11456), .ZN(n11455) );
  AND2_X1 U12435 ( .A1(n11459), .A2(n11458), .ZN(n11457) );
  NAND2_X1 U12436 ( .A1(n11200), .A2(n11458), .ZN(n11456) );
  NAND2_X1 U12437 ( .A1(n11449), .A2(n11207), .ZN(n11448) );
  INV_X1 U12438 ( .A(n17130), .ZN(n11449) );
  NAND2_X1 U12439 ( .A1(n17130), .A2(n11453), .ZN(n11451) );
  NOR2_X1 U12440 ( .A1(n11200), .A2(n11454), .ZN(n11453) );
  INV_X1 U12441 ( .A(n11458), .ZN(n11454) );
  NAND2_X1 U12442 ( .A1(n17130), .A2(n17129), .ZN(n17137) );
  NAND2_X1 U12443 ( .A1(n11768), .A2(n11764), .ZN(n17182) );
  INV_X1 U12444 ( .A(n11493), .ZN(n11491) );
  OR2_X1 U12445 ( .A1(n11498), .A2(n11810), .ZN(n11497) );
  NAND2_X1 U12446 ( .A1(n11609), .A2(n11263), .ZN(n17602) );
  OR2_X1 U12447 ( .A1(n17621), .A2(n17620), .ZN(n11609) );
  INV_X1 U12448 ( .A(n15557), .ZN(n11555) );
  INV_X1 U12449 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19891) );
  INV_X1 U12450 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19889) );
  INV_X1 U12451 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19766) );
  AND2_X1 U12452 ( .A1(n14858), .A2(n14824), .ZN(n19845) );
  NAND2_X1 U12453 ( .A1(n11587), .A2(n11836), .ZN(n14827) );
  AND2_X1 U12454 ( .A1(n14863), .A2(n14882), .ZN(n19863) );
  INV_X1 U12455 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19777) );
  OR2_X1 U12456 ( .A1(n14819), .A2(n14753), .ZN(n19732) );
  INV_X1 U12457 ( .A(n17659), .ZN(n19211) );
  NAND2_X1 U12458 ( .A1(n14821), .A2(n14706), .ZN(n19745) );
  NOR2_X1 U12459 ( .A1(n19895), .A2(n19846), .ZN(n20315) );
  OAI21_X1 U12460 ( .B1(n19857), .B2(n19854), .A(n19853), .ZN(n20310) );
  NOR2_X2 U12461 ( .A1(n19836), .A2(n19835), .ZN(n20308) );
  INV_X1 U12462 ( .A(n19803), .ZN(n20284) );
  INV_X1 U12463 ( .A(n20193), .ZN(n20272) );
  INV_X1 U12464 ( .A(n20327), .ZN(n20337) );
  INV_X1 U12465 ( .A(n19964), .ZN(n19968) );
  AND2_X1 U12466 ( .A1(n15278), .A2(n15277), .ZN(n19218) );
  NOR2_X2 U12467 ( .A1(n21787), .A2(n21847), .ZN(n21850) );
  AND2_X1 U12468 ( .A1(n20968), .A2(n21054), .ZN(n20969) );
  AND2_X1 U12469 ( .A1(n11643), .A2(n11642), .ZN(n20951) );
  NOR2_X1 U12470 ( .A1(n20926), .A2(n20927), .ZN(n20941) );
  NOR2_X1 U12471 ( .A1(n21080), .A2(n20925), .ZN(n20926) );
  NOR2_X1 U12472 ( .A1(n20989), .A2(n18188), .ZN(n18194) );
  INV_X1 U12473 ( .A(n18246), .ZN(n18219) );
  NOR2_X1 U12474 ( .A1(n18234), .A2(n18233), .ZN(n18247) );
  BUF_X1 U12475 ( .A(n18248), .Z(n18268) );
  NAND2_X1 U12476 ( .A1(n21225), .A2(n11222), .ZN(n21242) );
  NAND2_X1 U12477 ( .A1(n21225), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n21247) );
  NOR2_X1 U12478 ( .A1(n21256), .A2(n21220), .ZN(n21225) );
  OR2_X1 U12479 ( .A1(n21254), .A2(n21255), .ZN(n21256) );
  NAND2_X1 U12480 ( .A1(n11423), .A2(n11327), .ZN(n21264) );
  INV_X1 U12481 ( .A(n21217), .ZN(n11422) );
  INV_X1 U12482 ( .A(n21218), .ZN(n11421) );
  INV_X1 U12483 ( .A(n21275), .ZN(n21266) );
  NOR2_X1 U12484 ( .A1(n21289), .A2(n21177), .ZN(n21178) );
  NAND2_X1 U12485 ( .A1(n21305), .A2(n11418), .ZN(n21289) );
  AND2_X1 U12486 ( .A1(n21176), .A2(n11419), .ZN(n11418) );
  NOR2_X1 U12487 ( .A1(n18309), .A2(n18308), .ZN(n21165) );
  INV_X1 U12488 ( .A(n21303), .ZN(n21175) );
  NOR2_X1 U12489 ( .A1(n21314), .A2(n18827), .ZN(n18901) );
  CLKBUF_X1 U12490 ( .A(n18901), .Z(n21785) );
  CLKBUF_X1 U12491 ( .A(n18903), .Z(n18911) );
  INV_X1 U12492 ( .A(n20680), .ZN(n20670) );
  NOR2_X1 U12493 ( .A1(n20678), .A2(n20670), .ZN(n20669) );
  INV_X1 U12494 ( .A(n20672), .ZN(n20678) );
  NOR2_X1 U12496 ( .A1(n18650), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11531) );
  NAND2_X1 U12497 ( .A1(n18589), .A2(n11646), .ZN(n18667) );
  INV_X1 U12498 ( .A(n21389), .ZN(n18548) );
  NAND2_X1 U12499 ( .A1(n18674), .A2(n11636), .ZN(n18515) );
  NOR2_X1 U12500 ( .A1(n21539), .A2(n21545), .ZN(n11526) );
  OR2_X1 U12501 ( .A1(n11528), .A2(n21491), .ZN(n11524) );
  OR2_X1 U12502 ( .A1(n11528), .A2(n18820), .ZN(n11523) );
  NOR2_X1 U12503 ( .A1(n11525), .A2(n11528), .ZN(n18733) );
  AND2_X1 U12504 ( .A1(n18820), .A2(n21491), .ZN(n11525) );
  NAND2_X1 U12505 ( .A1(n18792), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18776) );
  INV_X1 U12506 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20745) );
  INV_X1 U12507 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n21314) );
  OAI21_X1 U12508 ( .B1(n21643), .B2(n21720), .A(n11279), .ZN(n11550) );
  NAND2_X1 U12509 ( .A1(n21638), .A2(n21639), .ZN(n11551) );
  AND2_X1 U12510 ( .A1(n18640), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11598) );
  INV_X1 U12511 ( .A(n18638), .ZN(n21666) );
  NAND2_X1 U12512 ( .A1(n18735), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18734) );
  INV_X1 U12513 ( .A(n21788), .ZN(n21675) );
  INV_X1 U12514 ( .A(n21766), .ZN(n21601) );
  INV_X1 U12515 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21806) );
  INV_X1 U12516 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21809) );
  INV_X1 U12517 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19534) );
  CLKBUF_X1 U12518 ( .A(n19247), .Z(n19581) );
  NOR2_X1 U12519 ( .A1(n16456), .A2(n16455), .ZN(n16457) );
  NOR2_X1 U12520 ( .A1(n13656), .A2(n11799), .ZN(n11798) );
  INV_X1 U12521 ( .A(n13655), .ZN(n11799) );
  OAI21_X1 U12522 ( .B1(n20513), .B2(n22216), .A(n11392), .ZN(P1_U2988) );
  AOI21_X1 U12523 ( .B1(n11395), .B2(n20557), .A(n11393), .ZN(n11392) );
  OAI21_X1 U12524 ( .B1(n20561), .B2(n22108), .A(n11394), .ZN(n11393) );
  INV_X1 U12525 ( .A(n22104), .ZN(n11395) );
  NAND2_X1 U12526 ( .A1(n11363), .A2(n16805), .ZN(P1_U3000) );
  AOI21_X1 U12527 ( .B1(n19687), .B2(n19189), .A(n16163), .ZN(n16164) );
  AOI211_X1 U12528 ( .C1(n16414), .C2(n17633), .A(n16121), .B(n16120), .ZN(
        n16122) );
  OAI21_X1 U12529 ( .B1(n21105), .B2(n21104), .A(n11655), .ZN(n11654) );
  AOI211_X1 U12530 ( .C1(n21082), .C2(n21076), .A(n21075), .B(n21074), .ZN(
        n21077) );
  INV_X1 U12531 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20718) );
  NAND2_X1 U12532 ( .A1(n11407), .A2(n11402), .ZN(P3_U2704) );
  NAND2_X1 U12533 ( .A1(n21229), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n11407) );
  NOR2_X1 U12534 ( .A1(n11406), .A2(n11403), .ZN(n11402) );
  NAND2_X1 U12535 ( .A1(n21305), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n21297) );
  AND2_X1 U12536 ( .A1(n21604), .A2(n11531), .ZN(n11530) );
  OAI21_X1 U12537 ( .B1(n11549), .B2(n21764), .A(n11547), .ZN(P3_U2831) );
  AOI21_X1 U12538 ( .B1(n21644), .B2(n21779), .A(n11548), .ZN(n11547) );
  AOI21_X1 U12539 ( .B1(n21640), .B2(n21788), .A(n11550), .ZN(n11549) );
  OAI21_X1 U12540 ( .B1(n21755), .B2(n21646), .A(n21645), .ZN(n11548) );
  NOR2_X1 U12541 ( .A1(n14964), .A2(n21355), .ZN(n14988) );
  INV_X1 U12542 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17763) );
  NAND2_X1 U12543 ( .A1(n11431), .A2(n11553), .ZN(n14286) );
  NAND2_X1 U12544 ( .A1(n11819), .A2(n11324), .ZN(n15875) );
  INV_X2 U12545 ( .A(n22278), .ZN(n17907) );
  NAND2_X1 U12546 ( .A1(n14207), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11199) );
  INV_X1 U12547 ( .A(n11158), .ZN(n14776) );
  XOR2_X1 U12548 ( .A(n17131), .B(n17345), .Z(n11200) );
  NAND2_X1 U12549 ( .A1(n17575), .A2(n17573), .ZN(n11201) );
  CLKBUF_X1 U12550 ( .A(n13042), .Z(n16390) );
  OR2_X1 U12551 ( .A1(n17316), .A2(n11321), .ZN(n17188) );
  AND2_X1 U12552 ( .A1(n15902), .A2(n11308), .ZN(n17026) );
  AND2_X1 U12553 ( .A1(n11585), .A2(n11587), .ZN(n11202) );
  NAND2_X1 U12554 ( .A1(n16584), .A2(n11273), .ZN(n11203) );
  INV_X1 U12555 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n17752) );
  NAND2_X1 U12556 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12982) );
  AND4_X1 U12557 ( .A1(n15030), .A2(n15029), .A3(n15028), .A4(n15027), .ZN(
        n11204) );
  AND2_X1 U12558 ( .A1(n14307), .A2(n14306), .ZN(n11205) );
  AND3_X1 U12559 ( .A1(n14200), .A2(n11351), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11206) );
  NOR2_X1 U12560 ( .A1(n15016), .A2(n15015), .ZN(n21180) );
  INV_X1 U12561 ( .A(n13123), .ZN(n11563) );
  AND2_X1 U12562 ( .A1(n11200), .A2(n11460), .ZN(n11207) );
  AND2_X1 U12563 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n11680), .ZN(
        n11208) );
  NAND2_X1 U12564 ( .A1(n12968), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12966) );
  NAND2_X1 U12565 ( .A1(n12970), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12969) );
  NOR2_X1 U12566 ( .A1(n14061), .A2(n11818), .ZN(n15877) );
  NOR2_X1 U12567 ( .A1(n11619), .A2(n11620), .ZN(n15923) );
  AND4_X1 U12568 ( .A1(n11723), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11209) );
  AND2_X1 U12569 ( .A1(n15383), .A2(n15127), .ZN(n11210) );
  AND2_X1 U12570 ( .A1(n11753), .A2(n11752), .ZN(n11211) );
  AND2_X1 U12571 ( .A1(n11271), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11212) );
  NAND2_X1 U12572 ( .A1(n14413), .A2(n13624), .ZN(n14419) );
  NOR2_X1 U12573 ( .A1(n11619), .A2(n11617), .ZN(n15804) );
  NAND2_X1 U12574 ( .A1(n21281), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n21271) );
  INV_X1 U12575 ( .A(n21271), .ZN(n11423) );
  AND2_X1 U12576 ( .A1(n11646), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11213) );
  AND2_X1 U12577 ( .A1(n15329), .A2(n11322), .ZN(n11214) );
  OR2_X1 U12578 ( .A1(n11324), .A2(n11820), .ZN(n11215) );
  AND2_X1 U12579 ( .A1(n11506), .A2(n22004), .ZN(n11216) );
  AND2_X1 U12580 ( .A1(n11506), .A2(n20556), .ZN(n11217) );
  NAND2_X1 U12581 ( .A1(n11608), .A2(n11603), .ZN(n15811) );
  AND2_X1 U12582 ( .A1(n13582), .A2(n11613), .ZN(n11218) );
  AND2_X1 U12583 ( .A1(n11715), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11219) );
  AND2_X1 U12584 ( .A1(n11307), .A2(n11731), .ZN(n11220) );
  OR3_X1 U12585 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n22463), .ZN(n11221) );
  AND2_X1 U12586 ( .A1(n11416), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n11222) );
  NAND2_X2 U12587 ( .A1(n17907), .A2(n22289), .ZN(n17904) );
  OR2_X1 U12588 ( .A1(n17036), .A2(n17035), .ZN(n11223) );
  INV_X1 U12589 ( .A(n13344), .ZN(n13443) );
  NOR2_X1 U12590 ( .A1(n20687), .A2(n21355), .ZN(n18223) );
  NAND2_X1 U12591 ( .A1(n14107), .A2(n14103), .ZN(n14147) );
  OR2_X1 U12592 ( .A1(n18522), .A2(n18442), .ZN(n11593) );
  AND4_X1 U12593 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11224) );
  INV_X2 U12594 ( .A(n16149), .ZN(n13176) );
  NAND2_X1 U12595 ( .A1(n16584), .A2(n16647), .ZN(n16529) );
  NAND2_X1 U12596 ( .A1(n12925), .A2(n20544), .ZN(n16680) );
  NAND2_X1 U12597 ( .A1(n11435), .A2(n14317), .ZN(n17332) );
  OR2_X1 U12598 ( .A1(n17191), .A2(n16080), .ZN(n11226) );
  OR2_X1 U12599 ( .A1(n17336), .A2(n17337), .ZN(n11814) );
  NAND2_X1 U12600 ( .A1(n11518), .A2(n11517), .ZN(n18010) );
  NAND2_X1 U12601 ( .A1(n11487), .A2(n13142), .ZN(n13161) );
  AND2_X1 U12602 ( .A1(n11735), .A2(n15177), .ZN(n11227) );
  NAND2_X1 U12603 ( .A1(n15776), .A2(n12915), .ZN(n16767) );
  AND4_X1 U12604 ( .A1(n11889), .A2(n11888), .A3(n11887), .A4(n11886), .ZN(
        n11228) );
  NAND2_X1 U12605 ( .A1(n13649), .A2(n13650), .ZN(n16432) );
  AND2_X1 U12606 ( .A1(n16584), .A2(n11827), .ZN(n16531) );
  AND2_X1 U12607 ( .A1(n11380), .A2(n11379), .ZN(n11229) );
  OR2_X1 U12608 ( .A1(n12873), .A2(n12203), .ZN(n11230) );
  NOR2_X1 U12609 ( .A1(n18377), .A2(n18376), .ZN(n18826) );
  INV_X1 U12610 ( .A(n18826), .ZN(n11540) );
  AND2_X1 U12611 ( .A1(n14322), .A2(n14318), .ZN(n11231) );
  INV_X1 U12612 ( .A(n21318), .ZN(n18396) );
  AND4_X1 U12613 ( .A1(n14992), .A2(n14991), .A3(n14990), .A4(n14989), .ZN(
        n11232) );
  AND4_X1 U12614 ( .A1(n13074), .A2(n15200), .A3(n13073), .A4(n13072), .ZN(
        n11233) );
  OAI21_X1 U12615 ( .B1(n17168), .B2(n11465), .A(n11462), .ZN(n17127) );
  AND2_X1 U12616 ( .A1(n18788), .A2(n11588), .ZN(n11234) );
  AND3_X1 U12617 ( .A1(n15033), .A2(n11409), .A3(n15032), .ZN(n11235) );
  AND2_X1 U12618 ( .A1(n15234), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13328) );
  NAND3_X1 U12619 ( .A1(n13110), .A2(n13109), .A3(n11426), .ZN(n13139) );
  AND2_X1 U12620 ( .A1(n12918), .A2(n11797), .ZN(n11236) );
  AND2_X1 U12621 ( .A1(n11227), .A2(n11734), .ZN(n11237) );
  OR2_X1 U12622 ( .A1(n16890), .A2(n16422), .ZN(n11238) );
  NOR2_X1 U12623 ( .A1(n17304), .A2(n11807), .ZN(n11239) );
  INV_X1 U12624 ( .A(n11375), .ZN(n16482) );
  NOR2_X1 U12625 ( .A1(n16509), .A2(n12734), .ZN(n11375) );
  AND2_X1 U12626 ( .A1(n16040), .A2(n11473), .ZN(n11240) );
  NAND2_X1 U12627 ( .A1(n11461), .A2(n11466), .ZN(n17150) );
  OR2_X1 U12628 ( .A1(n17130), .A2(n17129), .ZN(n11241) );
  INV_X1 U12629 ( .A(n14061), .ZN(n11819) );
  NAND2_X1 U12630 ( .A1(n14308), .A2(n11447), .ZN(n11242) );
  OR2_X1 U12631 ( .A1(n14443), .A2(n14442), .ZN(n11243) );
  NAND4_X1 U12632 ( .A1(n17203), .A2(n16046), .A3(n16045), .A4(n16044), .ZN(
        n11244) );
  AND2_X1 U12633 ( .A1(n11474), .A2(n11469), .ZN(n11245) );
  NOR2_X1 U12634 ( .A1(n16747), .A2(n12922), .ZN(n11246) );
  INV_X1 U12635 ( .A(n11460), .ZN(n11459) );
  NAND2_X1 U12636 ( .A1(n17129), .A2(n17141), .ZN(n11460) );
  OR2_X1 U12637 ( .A1(n17304), .A2(n11808), .ZN(n17448) );
  INV_X1 U12638 ( .A(n17448), .ZN(n11359) );
  AND2_X1 U12639 ( .A1(n19175), .A2(n14257), .ZN(n11247) );
  AND2_X1 U12640 ( .A1(n12889), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11248) );
  AND2_X1 U12641 ( .A1(n12905), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11249) );
  NAND2_X1 U12642 ( .A1(n14321), .A2(n14322), .ZN(n11250) );
  INV_X1 U12643 ( .A(n11811), .ZN(n17287) );
  OR2_X1 U12644 ( .A1(n17304), .A2(n17533), .ZN(n11811) );
  AND2_X1 U12645 ( .A1(n11913), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11251) );
  NOR2_X1 U12646 ( .A1(n18733), .A2(n21539), .ZN(n11252) );
  AND2_X1 U12647 ( .A1(n11922), .A2(n16595), .ZN(n11253) );
  NOR2_X1 U12648 ( .A1(n18755), .A2(n21479), .ZN(n18422) );
  MUX2_X1 U12649 ( .A(n13063), .B(n13062), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14410) );
  INV_X1 U12650 ( .A(n15981), .ZN(n15979) );
  OR2_X1 U12651 ( .A1(n15022), .A2(n11520), .ZN(n15981) );
  NAND2_X1 U12652 ( .A1(n17030), .A2(n11737), .ZN(n16924) );
  AND2_X1 U12653 ( .A1(n17030), .A2(n17022), .ZN(n17016) );
  NAND2_X1 U12654 ( .A1(n11437), .A2(n11436), .ZN(n13143) );
  AND2_X1 U12655 ( .A1(n11954), .A2(n15391), .ZN(n11254) );
  AND2_X1 U12656 ( .A1(n14416), .A2(n11740), .ZN(n11255) );
  AND2_X1 U12657 ( .A1(n11499), .A2(n12005), .ZN(n11256) );
  AND2_X1 U12658 ( .A1(n11814), .A2(n11199), .ZN(n11257) );
  AND2_X1 U12659 ( .A1(n13113), .A2(n11565), .ZN(n11258) );
  NAND2_X1 U12660 ( .A1(n14441), .A2(n14440), .ZN(n11259) );
  NAND2_X1 U12661 ( .A1(n14382), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13127) );
  NAND2_X1 U12662 ( .A1(n18757), .A2(n18756), .ZN(n11260) );
  NAND2_X1 U12663 ( .A1(n20526), .A2(n14577), .ZN(n11261) );
  INV_X1 U12664 ( .A(n11495), .ZN(n11494) );
  NAND2_X1 U12665 ( .A1(n11496), .A2(n14427), .ZN(n11495) );
  OR2_X1 U12666 ( .A1(n18653), .A2(n11532), .ZN(n11262) );
  AND2_X2 U12667 ( .A1(n11801), .A2(n15076), .ZN(n11913) );
  NAND2_X1 U12668 ( .A1(n14747), .A2(n13337), .ZN(n13532) );
  OR2_X1 U12669 ( .A1(n16060), .A2(n13572), .ZN(n11263) );
  NAND2_X1 U12670 ( .A1(n14888), .A2(n14953), .ZN(n14952) );
  NOR2_X1 U12671 ( .A1(n12979), .A2(n17338), .ZN(n12980) );
  NOR2_X1 U12672 ( .A1(n12982), .A2(n17763), .ZN(n12983) );
  NAND2_X1 U12673 ( .A1(n12978), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12975) );
  OR2_X1 U12674 ( .A1(n16583), .A2(n11743), .ZN(n11264) );
  INV_X1 U12675 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11983) );
  AND2_X1 U12676 ( .A1(n21225), .A2(n11416), .ZN(n11265) );
  AND2_X1 U12677 ( .A1(n18674), .A2(n11637), .ZN(n11266) );
  NOR2_X1 U12678 ( .A1(n12977), .A2(n17318), .ZN(n12978) );
  AND2_X1 U12679 ( .A1(n12988), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12971) );
  NAND2_X1 U12680 ( .A1(n13122), .A2(n13619), .ZN(n14403) );
  AND2_X1 U12681 ( .A1(n11614), .A2(n11218), .ZN(n11267) );
  AND2_X1 U12682 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11268) );
  AND2_X1 U12683 ( .A1(n11600), .A2(n15321), .ZN(n11269) );
  OAI21_X1 U12684 ( .B1(n11435), .B2(n11434), .A(n11432), .ZN(n17294) );
  AND2_X1 U12685 ( .A1(n11205), .A2(n15729), .ZN(n11270) );
  NAND2_X1 U12686 ( .A1(n11391), .A2(n12879), .ZN(n15514) );
  AND2_X1 U12687 ( .A1(n15812), .A2(n11615), .ZN(n15803) );
  AND2_X1 U12688 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11271) );
  AND2_X1 U12689 ( .A1(n15902), .A2(n15901), .ZN(n16201) );
  AND2_X1 U12690 ( .A1(n20552), .A2(n16823), .ZN(n11272) );
  AND2_X1 U12691 ( .A1(n11827), .A2(n16573), .ZN(n11273) );
  AND2_X1 U12692 ( .A1(n15299), .A2(n15424), .ZN(n11274) );
  INV_X1 U12693 ( .A(n21121), .ZN(n21305) );
  AOI21_X1 U12694 ( .B1(n21117), .B2(n21118), .A(n21116), .ZN(n21121) );
  AND3_X1 U12695 ( .A1(n15299), .A2(n15424), .A3(n15427), .ZN(n11275) );
  OR2_X1 U12696 ( .A1(n12705), .A2(n12686), .ZN(n11276) );
  AND2_X1 U12697 ( .A1(n12106), .A2(n12105), .ZN(n15171) );
  INV_X1 U12698 ( .A(n15171), .ZN(n11512) );
  OR3_X1 U12699 ( .A1(n16583), .A2(n11743), .A3(n16537), .ZN(n11277) );
  AND2_X1 U12700 ( .A1(n15937), .A2(n15936), .ZN(n11278) );
  AND2_X1 U12701 ( .A1(n17191), .A2(n16080), .ZN(n11767) );
  INV_X1 U12702 ( .A(n11767), .ZN(n11764) );
  INV_X1 U12703 ( .A(n11639), .ZN(n19142) );
  NAND2_X1 U12704 ( .A1(n16072), .A2(n16070), .ZN(n11639) );
  AND2_X1 U12705 ( .A1(n12145), .A2(n12144), .ZN(n12215) );
  AND2_X1 U12706 ( .A1(n21642), .A2(n11551), .ZN(n11279) );
  AND2_X1 U12707 ( .A1(n11913), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11280) );
  AND2_X1 U12708 ( .A1(n11913), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11281) );
  NAND2_X1 U12709 ( .A1(n17305), .A2(n17322), .ZN(n11282) );
  NOR2_X1 U12710 ( .A1(n15889), .A2(n15888), .ZN(n14472) );
  NOR2_X1 U12711 ( .A1(n15702), .A2(n15701), .ZN(n15689) );
  NOR2_X1 U12712 ( .A1(n17101), .A2(n11627), .ZN(n16927) );
  AND2_X1 U12713 ( .A1(n14710), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11283) );
  NOR2_X1 U12714 ( .A1(n12832), .A2(n22414), .ZN(n11284) );
  AND2_X1 U12715 ( .A1(n12120), .A2(n12119), .ZN(n11285) );
  NOR2_X1 U12716 ( .A1(n11746), .A2(n15356), .ZN(n11286) );
  AND2_X1 U12717 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11287) );
  NOR2_X1 U12718 ( .A1(n11675), .A2(n16099), .ZN(n11674) );
  AND2_X1 U12719 ( .A1(n11636), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11288) );
  AND2_X1 U12720 ( .A1(n11212), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11289) );
  NAND2_X1 U12721 ( .A1(keyinput_3), .A2(DATAI_29_), .ZN(n11290) );
  AND2_X1 U12722 ( .A1(n11214), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11291) );
  INV_X1 U12723 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15755) );
  INV_X1 U12724 ( .A(n13321), .ZN(n15214) );
  INV_X1 U12725 ( .A(n19182), .ZN(n17636) );
  INV_X1 U12726 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U12727 ( .A1(n17621), .A2(n11263), .ZN(n11608) );
  NOR2_X1 U12728 ( .A1(n18585), .A2(n18617), .ZN(n18589) );
  AND2_X1 U12729 ( .A1(n15330), .A2(n11214), .ZN(n15120) );
  AND2_X1 U12730 ( .A1(n12988), .A2(n11289), .ZN(n12970) );
  NOR2_X1 U12731 ( .A1(n12969), .A2(n17221), .ZN(n12968) );
  NOR2_X1 U12732 ( .A1(n15811), .A2(n15813), .ZN(n15812) );
  NAND2_X1 U12733 ( .A1(n18555), .A2(n11854), .ZN(n18585) );
  AND2_X1 U12734 ( .A1(n11608), .A2(n11606), .ZN(n15838) );
  NAND2_X1 U12735 ( .A1(n12996), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12960) );
  NAND2_X1 U12736 ( .A1(n15921), .A2(n15920), .ZN(n15919) );
  NAND2_X1 U12737 ( .A1(n14583), .A2(n14553), .ZN(n22010) );
  NOR2_X1 U12738 ( .A1(n15739), .A2(n15740), .ZN(n14937) );
  INV_X1 U12739 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11638) );
  NAND2_X1 U12740 ( .A1(n15580), .A2(n15579), .ZN(n14069) );
  AND2_X1 U12741 ( .A1(n16566), .A2(n11750), .ZN(n11292) );
  AND2_X1 U12742 ( .A1(n15901), .A2(n17043), .ZN(n11293) );
  AND2_X1 U12743 ( .A1(n11292), .A2(n11749), .ZN(n11294) );
  NAND2_X1 U12744 ( .A1(n14403), .A2(n11756), .ZN(n14387) );
  OR2_X1 U12745 ( .A1(n16537), .A2(n16574), .ZN(n11295) );
  AND2_X1 U12746 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11296) );
  AND2_X1 U12747 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11297) );
  AND2_X1 U12748 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11298) );
  AND2_X1 U12749 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11299) );
  AND2_X1 U12750 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11300) );
  AND2_X1 U12751 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11301) );
  AND2_X1 U12752 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11302) );
  AND2_X1 U12753 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11303) );
  AND2_X1 U12754 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11304) );
  AND2_X1 U12755 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11305) );
  OR2_X1 U12756 ( .A1(n16136), .A2(n13633), .ZN(n11306) );
  INV_X1 U12757 ( .A(n11921), .ZN(n14550) );
  AND2_X1 U12758 ( .A1(n16987), .A2(n16996), .ZN(n11307) );
  AND2_X1 U12759 ( .A1(n11293), .A2(n11578), .ZN(n11308) );
  AND2_X1 U12760 ( .A1(n12996), .A2(n11219), .ZN(n11309) );
  INV_X1 U12761 ( .A(n14469), .ZN(n11663) );
  NAND2_X1 U12762 ( .A1(n12963), .A2(n12995), .ZN(n16949) );
  INV_X1 U12763 ( .A(n20556), .ZN(n22216) );
  NAND2_X1 U12764 ( .A1(n20467), .A2(n20466), .ZN(n16580) );
  INV_X1 U12765 ( .A(n16144), .ZN(n11732) );
  INV_X1 U12766 ( .A(n17283), .ZN(n11471) );
  NAND2_X1 U12767 ( .A1(n11667), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12967) );
  INV_X1 U12768 ( .A(n12967), .ZN(n11666) );
  AND2_X1 U12769 ( .A1(n11308), .A2(n17028), .ZN(n11310) );
  INV_X1 U12770 ( .A(n21860), .ZN(n15410) );
  AND2_X1 U12771 ( .A1(n11373), .A2(n22809), .ZN(n21860) );
  NAND2_X1 U12772 ( .A1(n14333), .A2(n17547), .ZN(n11311) );
  OR2_X1 U12773 ( .A1(n21092), .A2(n21094), .ZN(n11312) );
  AND2_X1 U12774 ( .A1(n11202), .A2(n11269), .ZN(n11313) );
  AND2_X1 U12775 ( .A1(n11294), .A2(n11748), .ZN(n11314) );
  AND2_X1 U12776 ( .A1(n11737), .A2(n11736), .ZN(n11315) );
  AND2_X1 U12777 ( .A1(n11220), .A2(n16144), .ZN(n11316) );
  INV_X1 U12778 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14797) );
  AND2_X1 U12779 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11317) );
  AND2_X1 U12780 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11318) );
  AND2_X1 U12781 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11319) );
  AND2_X1 U12782 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11320) );
  OR2_X1 U12783 ( .A1(n17422), .A2(n17428), .ZN(n11321) );
  AND2_X1 U12784 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11322) );
  OR2_X1 U12785 ( .A1(n11321), .A2(n16080), .ZN(n11323) );
  NAND2_X1 U12786 ( .A1(n12285), .A2(n12284), .ZN(n11324) );
  NOR2_X1 U12787 ( .A1(n18567), .A2(n18566), .ZN(n11325) );
  INV_X1 U12788 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18798) );
  NAND4_X1 U12789 ( .A1(n18750), .A2(n11658), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A4(n11657), .ZN(n18451) );
  INV_X1 U12790 ( .A(n20538), .ZN(n20557) );
  INV_X1 U12791 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11647) );
  INV_X1 U12792 ( .A(n20927), .ZN(n11641) );
  INV_X1 U12793 ( .A(n20943), .ZN(n11642) );
  NOR2_X1 U12794 ( .A1(n18776), .A2(n20745), .ZN(n18715) );
  NOR2_X1 U12795 ( .A1(n14211), .A2(n17504), .ZN(n11326) );
  AND4_X1 U12796 ( .A1(n11422), .A2(n11421), .A3(P3_EAX_REG_22__SCAN_IN), .A4(
        P3_EAX_REG_19__SCAN_IN), .ZN(n11327) );
  INV_X1 U12797 ( .A(n21539), .ZN(n11527) );
  INV_X1 U12798 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15234) );
  OR3_X1 U12799 ( .A1(n12924), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11328) );
  XOR2_X1 U12800 ( .A(n22113), .B(keyinput_71), .Z(n11329) );
  INV_X1 U12801 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11716) );
  INV_X1 U12802 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11717) );
  NAND2_X1 U12803 ( .A1(n11561), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11330) );
  OR2_X1 U12804 ( .A1(n16078), .A2(n11330), .ZN(n11331) );
  OR2_X1 U12805 ( .A1(n16078), .A2(n17141), .ZN(n11332) );
  INV_X1 U12806 ( .A(DATAI_29_), .ZN(n13670) );
  INV_X1 U12807 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n11420) );
  INV_X1 U12808 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11681) );
  INV_X1 U12809 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11503) );
  INV_X1 U12810 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11778) );
  AND2_X1 U12811 ( .A1(n12927), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11333) );
  INV_X1 U12812 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11430) );
  NAND2_X1 U12813 ( .A1(keyinput_115), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11334)
         );
  NOR2_X1 U12814 ( .A1(n21785), .A2(n18888), .ZN(n18903) );
  NOR2_X1 U12815 ( .A1(n20381), .A2(n21862), .ZN(n20393) );
  INV_X1 U12816 ( .A(n16592), .ZN(n16588) );
  NAND2_X1 U12817 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11371) );
  OAI22_X2 U12818 ( .A1(n22422), .A2(n22632), .B1(n22421), .B2(n22630), .ZN(
        n22523) );
  OR2_X1 U12819 ( .A1(n16592), .A2(n20538), .ZN(n22630) );
  INV_X1 U12820 ( .A(n22668), .ZN(n11335) );
  INV_X1 U12821 ( .A(n11335), .ZN(n11336) );
  OAI22_X2 U12822 ( .A1(n22558), .A2(n22632), .B1(n22557), .B2(n22630), .ZN(
        n22594) );
  INV_X1 U12823 ( .A(n22725), .ZN(n11337) );
  INV_X1 U12824 ( .A(n11337), .ZN(n11338) );
  INV_X1 U12825 ( .A(n22617), .ZN(n11339) );
  INV_X1 U12826 ( .A(n11339), .ZN(n11340) );
  INV_X1 U12827 ( .A(n22547), .ZN(n11341) );
  INV_X1 U12828 ( .A(n11341), .ZN(n11342) );
  INV_X1 U12829 ( .A(n11221), .ZN(n11343) );
  INV_X1 U12830 ( .A(n22782), .ZN(n11344) );
  INV_X1 U12831 ( .A(n11344), .ZN(n11345) );
  INV_X1 U12832 ( .A(n22588), .ZN(n11346) );
  INV_X1 U12833 ( .A(n11346), .ZN(n11347) );
  INV_X1 U12834 ( .A(n22663), .ZN(n11348) );
  INV_X1 U12835 ( .A(n11348), .ZN(n11349) );
  NAND2_X1 U12836 ( .A1(n21653), .A2(n21648), .ZN(n21476) );
  INV_X1 U12837 ( .A(n21653), .ZN(n21764) );
  NOR2_X2 U12838 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19725), .ZN(n19911) );
  NOR3_X2 U12839 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12668), .A3(
        n22463), .ZN(n22729) );
  NOR2_X2 U12840 ( .A1(n19275), .A2(n19298), .ZN(n19622) );
  OAI22_X2 U12841 ( .A1(n22413), .A2(n22632), .B1(n22412), .B2(n22630), .ZN(
        n22517) );
  NAND2_X1 U12842 ( .A1(n19142), .A2(n14287), .ZN(n17129) );
  OR2_X1 U12843 ( .A1(n14280), .A2(n14287), .ZN(n14309) );
  AOI21_X1 U12844 ( .B1(n18973), .B2(n14287), .A(n15742), .ZN(n11445) );
  OR3_X1 U12845 ( .A1(n16653), .A2(n16592), .A3(n16591), .ZN(n16662) );
  INV_X1 U12846 ( .A(n16662), .ZN(n11350) );
  INV_X1 U12847 ( .A(n16659), .ZN(n16653) );
  NAND2_X1 U12848 ( .A1(n14200), .A2(n11351), .ZN(n11353) );
  INV_X1 U12849 ( .A(n14193), .ZN(n11352) );
  NAND2_X1 U12850 ( .A1(n11353), .A2(n15742), .ZN(n15753) );
  NAND3_X1 U12851 ( .A1(n11566), .A2(n11563), .A3(n11565), .ZN(n14249) );
  AND2_X2 U12852 ( .A1(n14383), .A2(n14701), .ZN(n13164) );
  NAND2_X1 U12853 ( .A1(n11354), .A2(n14505), .ZN(P2_U2996) );
  NAND2_X1 U12854 ( .A1(n11355), .A2(n17782), .ZN(n11354) );
  NAND2_X1 U12855 ( .A1(n11494), .A2(n17250), .ZN(n11356) );
  NAND3_X1 U12856 ( .A1(n11771), .A2(n11772), .A3(n11554), .ZN(n11357) );
  NAND2_X2 U12857 ( .A1(n11482), .A2(n11483), .ZN(n11772) );
  NAND2_X2 U12858 ( .A1(n11480), .A2(n11479), .ZN(n11771) );
  OR2_X2 U12859 ( .A1(n17316), .A2(n11498), .ZN(n17304) );
  OAI21_X2 U12860 ( .B1(n11391), .B2(n11362), .A(n11360), .ZN(n15606) );
  NAND2_X1 U12861 ( .A1(n15606), .A2(n11782), .ZN(n11781) );
  NAND3_X1 U12862 ( .A1(n11510), .A2(n11216), .A3(n11504), .ZN(n11363) );
  XNOR2_X1 U12863 ( .A(n12851), .B(n11364), .ZN(n14838) );
  NAND2_X1 U12864 ( .A1(n11790), .A2(n15778), .ZN(n11367) );
  NAND2_X1 U12865 ( .A1(n15694), .A2(n15695), .ZN(n11368) );
  NAND2_X4 U12866 ( .A1(n11224), .A2(n11860), .ZN(n14764) );
  NAND3_X1 U12867 ( .A1(n16693), .A2(n16681), .A3(n16708), .ZN(n16702) );
  NAND2_X1 U12868 ( .A1(n11369), .A2(n12005), .ZN(n11501) );
  NAND2_X1 U12869 ( .A1(n11369), .A2(n11256), .ZN(n11500) );
  NAND2_X1 U12870 ( .A1(n15397), .A2(n11369), .ZN(n15134) );
  OR2_X2 U12871 ( .A1(n12031), .A2(n12030), .ZN(n11369) );
  CLKBUF_X1 U12872 ( .A(n11913), .Z(n11370) );
  NAND2_X1 U12873 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11372) );
  NAND2_X1 U12874 ( .A1(n18787), .A2(n18788), .ZN(n18786) );
  NAND2_X1 U12875 ( .A1(n18787), .A2(n11234), .ZN(n11380) );
  NAND2_X1 U12876 ( .A1(n18786), .A2(n18382), .ZN(n18384) );
  NAND2_X1 U12877 ( .A1(n18778), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18777) );
  INV_X1 U12878 ( .A(n18382), .ZN(n11383) );
  INV_X2 U12879 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21361) );
  NAND2_X2 U12880 ( .A1(n18331), .A2(n11537), .ZN(n18412) );
  NAND2_X1 U12881 ( .A1(n18317), .A2(n11385), .ZN(n18361) );
  INV_X1 U12882 ( .A(n18319), .ZN(n11387) );
  INV_X1 U12883 ( .A(n18412), .ZN(n21301) );
  INV_X1 U12884 ( .A(n18361), .ZN(n21172) );
  OAI21_X1 U12885 ( .B1(n18749), .B2(n11390), .A(n11389), .ZN(n11602) );
  AND2_X2 U12886 ( .A1(n11602), .A2(n11601), .ZN(n18708) );
  NOR2_X4 U12887 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16896) );
  NAND2_X1 U12888 ( .A1(n15161), .A2(n15160), .ZN(n11391) );
  OAI21_X1 U12889 ( .B1(n15112), .B2(n12906), .A(n12844), .ZN(n14801) );
  NAND4_X1 U12890 ( .A1(n11401), .A2(n11995), .A3(n11400), .A4(n11399), .ZN(
        n11973) );
  NAND3_X1 U12891 ( .A1(n21321), .A2(n15999), .A3(n16005), .ZN(n15986) );
  NAND3_X1 U12892 ( .A1(n11414), .A2(n14995), .A3(n11413), .ZN(n11412) );
  AND2_X1 U12893 ( .A1(n11425), .A2(n17616), .ZN(n17771) );
  NAND2_X1 U12894 ( .A1(n11426), .A2(n20079), .ZN(n13065) );
  NOR2_X1 U12895 ( .A1(n11426), .A2(n14404), .ZN(n14413) );
  NOR2_X1 U12896 ( .A1(n11426), .A2(n13619), .ZN(n11436) );
  NAND2_X2 U12897 ( .A1(n11427), .A2(n13338), .ZN(n11426) );
  NAND2_X1 U12898 ( .A1(n11255), .A2(n11429), .ZN(n11428) );
  NAND2_X1 U12899 ( .A1(n13140), .A2(n13624), .ZN(n11429) );
  NOR2_X2 U12900 ( .A1(n17316), .A2(n11323), .ZN(n17176) );
  AND2_X2 U12901 ( .A1(n17569), .A2(n14210), .ZN(n17316) );
  NAND2_X1 U12902 ( .A1(n11438), .A2(n11446), .ZN(n15738) );
  NAND2_X1 U12903 ( .A1(n14286), .A2(n11270), .ZN(n11438) );
  OAI211_X1 U12904 ( .C1(n14280), .C2(n11444), .A(n11442), .B(n11439), .ZN(
        n14311) );
  INV_X1 U12905 ( .A(n11446), .ZN(n11441) );
  NAND2_X1 U12906 ( .A1(n11443), .A2(n11446), .ZN(n11442) );
  INV_X1 U12907 ( .A(n14286), .ZN(n11443) );
  NAND3_X1 U12908 ( .A1(n11451), .A2(n11455), .A3(n11448), .ZN(n17353) );
  NAND3_X1 U12909 ( .A1(n11451), .A2(n11450), .A3(n11448), .ZN(n11452) );
  AND2_X1 U12910 ( .A1(n11455), .A2(n17636), .ZN(n11450) );
  NAND2_X1 U12911 ( .A1(n17352), .A2(n11452), .ZN(P2_U3018) );
  NAND2_X1 U12912 ( .A1(n17168), .A2(n11468), .ZN(n11461) );
  NOR2_X1 U12913 ( .A1(n11476), .A2(n11471), .ZN(n11470) );
  NAND3_X1 U12914 ( .A1(n11772), .A2(n11771), .A3(n11554), .ZN(n11553) );
  NAND2_X1 U12915 ( .A1(n11487), .A2(n11484), .ZN(n11486) );
  NAND2_X1 U12916 ( .A1(n11486), .A2(n11488), .ZN(n13138) );
  INV_X1 U12917 ( .A(n13143), .ZN(n16146) );
  NAND2_X1 U12918 ( .A1(n13066), .A2(n13065), .ZN(n13140) );
  OAI21_X1 U12919 ( .B1(n11495), .B2(n11492), .A(n11490), .ZN(P2_U3028) );
  AOI21_X1 U12920 ( .B1(n11491), .B2(n17628), .A(n11259), .ZN(n11490) );
  NAND2_X1 U12921 ( .A1(n17250), .A2(n17628), .ZN(n11492) );
  NAND2_X1 U12922 ( .A1(n17250), .A2(n14427), .ZN(n17233) );
  INV_X1 U12923 ( .A(n12013), .ZN(n11499) );
  AND2_X2 U12924 ( .A1(n15101), .A2(n11500), .ZN(n15074) );
  XNOR2_X1 U12925 ( .A(n11861), .B(n11503), .ZN(n15777) );
  NAND3_X1 U12926 ( .A1(n11504), .A2(n11510), .A3(n11217), .ZN(n12952) );
  NAND2_X1 U12927 ( .A1(n13652), .A2(n11508), .ZN(n11510) );
  AND2_X1 U12928 ( .A1(n12936), .A2(n12935), .ZN(n11509) );
  INV_X1 U12929 ( .A(n12202), .ZN(n12133) );
  NOR2_X1 U12930 ( .A1(n15171), .A2(n11285), .ZN(n11511) );
  INV_X1 U12931 ( .A(n12191), .ZN(n11513) );
  INV_X1 U12932 ( .A(n21347), .ZN(n11518) );
  NOR2_X2 U12933 ( .A1(n21766), .A2(n21789), .ZN(n21768) );
  NAND2_X2 U12934 ( .A1(n11519), .A2(n21318), .ZN(n21766) );
  NAND4_X1 U12935 ( .A1(n11522), .A2(n15024), .A3(n15025), .A4(n11521), .ZN(
        n11520) );
  NAND3_X1 U12936 ( .A1(n11524), .A2(n11523), .A3(n11526), .ZN(n18493) );
  NOR2_X2 U12937 ( .A1(n18831), .A2(n18400), .ZN(n18746) );
  AOI21_X1 U12938 ( .B1(n18624), .B2(n11530), .A(n11262), .ZN(n18654) );
  NAND2_X1 U12939 ( .A1(n18624), .A2(n21604), .ZN(n18649) );
  NOR2_X2 U12940 ( .A1(n18495), .A2(n18496), .ZN(n21389) );
  NAND2_X1 U12941 ( .A1(n18426), .A2(n21477), .ZN(n11543) );
  NAND3_X1 U12942 ( .A1(n11545), .A2(n11260), .A3(n18423), .ZN(n18735) );
  AOI21_X1 U12943 ( .B1(n13175), .B2(n11552), .A(n13174), .ZN(n15655) );
  XNOR2_X2 U12944 ( .A(n11552), .B(n14085), .ZN(n14844) );
  AND2_X1 U12945 ( .A1(n14115), .A2(n14129), .ZN(n11554) );
  NOR2_X1 U12946 ( .A1(n17612), .A2(n14202), .ZN(n17336) );
  OAI21_X1 U12947 ( .B1(n17612), .B2(n11556), .A(n11813), .ZN(n17569) );
  INV_X1 U12948 ( .A(n14202), .ZN(n11557) );
  INV_X1 U12949 ( .A(n13126), .ZN(n11560) );
  NAND3_X1 U12950 ( .A1(n14403), .A2(n11558), .A3(n11756), .ZN(n13136) );
  NAND3_X1 U12951 ( .A1(n11756), .A2(n14403), .A3(n13115), .ZN(n14384) );
  NAND3_X2 U12952 ( .A1(n13136), .A2(n13127), .A3(n11559), .ZN(n13163) );
  OR2_X1 U12953 ( .A1(n17177), .A2(n11332), .ZN(n17132) );
  AND2_X2 U12954 ( .A1(n15685), .A2(n15686), .ZN(n15772) );
  NOR2_X2 U12955 ( .A1(n14405), .A2(n13111), .ZN(n11565) );
  NAND2_X1 U12956 ( .A1(n16366), .A2(n11573), .ZN(n11567) );
  NAND2_X1 U12957 ( .A1(n16366), .A2(n16365), .ZN(n16992) );
  OAI21_X1 U12958 ( .B1(n16366), .B2(n11570), .A(n11568), .ZN(n11576) );
  INV_X1 U12959 ( .A(n16976), .ZN(n11575) );
  NAND2_X1 U12960 ( .A1(n15330), .A2(n11291), .ZN(n15346) );
  NOR2_X4 U12961 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15192) );
  NAND4_X1 U12962 ( .A1(n13026), .A2(n13023), .A3(n13024), .A4(n13025), .ZN(
        n11580) );
  NAND3_X1 U12963 ( .A1(n13020), .A2(n13018), .A3(n13019), .ZN(n11583) );
  NAND2_X1 U12964 ( .A1(n14947), .A2(n13391), .ZN(n11584) );
  NAND2_X1 U12965 ( .A1(n11836), .A2(n11586), .ZN(n11585) );
  NOR2_X1 U12966 ( .A1(n17060), .A2(n14447), .ZN(n14449) );
  AND2_X1 U12967 ( .A1(n18600), .A2(n21598), .ZN(n18638) );
  NAND2_X1 U12968 ( .A1(n18600), .A2(n11594), .ZN(n18658) );
  NOR2_X2 U12969 ( .A1(n18600), .A2(n21598), .ZN(n18639) );
  NAND2_X1 U12970 ( .A1(n11202), .A2(n11599), .ZN(n15747) );
  INV_X1 U12971 ( .A(n15747), .ZN(n13436) );
  INV_X1 U12972 ( .A(n11602), .ZN(n18476) );
  NAND2_X1 U12973 ( .A1(n15812), .A2(n15908), .ZN(n15907) );
  NAND2_X1 U12974 ( .A1(n11624), .A2(n11622), .ZN(n17067) );
  NAND3_X1 U12975 ( .A1(n13337), .A2(n11283), .A3(n19982), .ZN(n13361) );
  NAND3_X1 U12976 ( .A1(n11631), .A2(n13383), .A3(n11629), .ZN(n14132) );
  NAND2_X1 U12977 ( .A1(n14132), .A2(n13624), .ZN(n13620) );
  AND2_X1 U12978 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11632) );
  INV_X1 U12979 ( .A(n16106), .ZN(n11633) );
  AND2_X2 U12980 ( .A1(n11635), .A2(n11634), .ZN(n16106) );
  NAND3_X1 U12981 ( .A1(n11760), .A2(n11759), .A3(n17128), .ZN(n11635) );
  NAND2_X1 U12982 ( .A1(n21054), .A2(n11640), .ZN(n11643) );
  INV_X1 U12983 ( .A(n11643), .ZN(n20942) );
  INV_X1 U12984 ( .A(n18632), .ZN(n18631) );
  NAND2_X1 U12985 ( .A1(n13636), .A2(n11650), .ZN(n16059) );
  NAND2_X1 U12986 ( .A1(n13636), .A2(n11648), .ZN(n16069) );
  NAND2_X1 U12987 ( .A1(n13636), .A2(n16055), .ZN(n16066) );
  OAI21_X1 U12988 ( .B1(n21093), .B2(n11312), .A(n11653), .ZN(P3_U2640) );
  NOR2_X1 U12989 ( .A1(n11656), .A2(n11654), .ZN(n11653) );
  NOR2_X1 U12990 ( .A1(n21081), .A2(n21080), .ZN(n21093) );
  NAND2_X1 U12991 ( .A1(n14468), .A2(n11662), .ZN(n16049) );
  NAND2_X1 U12992 ( .A1(n14468), .A2(n11660), .ZN(n16051) );
  NAND2_X1 U12993 ( .A1(n14468), .A2(n14469), .ZN(n16033) );
  NAND2_X1 U12994 ( .A1(n13782), .A2(n11670), .ZN(n11668) );
  NAND2_X1 U12995 ( .A1(n11668), .A2(n11669), .ZN(n13797) );
  NAND2_X1 U12996 ( .A1(n19147), .A2(n11674), .ZN(n11672) );
  NAND2_X1 U12997 ( .A1(n19147), .A2(n19148), .ZN(n19146) );
  NAND2_X1 U12998 ( .A1(n12996), .A2(n11714), .ZN(n12955) );
  NAND3_X1 U12999 ( .A1(n13674), .A2(n13675), .A3(n11290), .ZN(n11720) );
  NAND2_X1 U13000 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11722) );
  NAND3_X1 U13001 ( .A1(n11723), .A2(n11721), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12979) );
  NAND3_X1 U13002 ( .A1(n11723), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12981) );
  INV_X2 U13003 ( .A(n12963), .ZN(n19134) );
  NAND3_X1 U13004 ( .A1(n13852), .A2(n13851), .A3(n11334), .ZN(n11730) );
  NAND2_X1 U13005 ( .A1(n16995), .A2(n11316), .ZN(n16151) );
  NAND2_X1 U13006 ( .A1(n16995), .A2(n11307), .ZN(n16989) );
  AND2_X1 U13007 ( .A1(n16995), .A2(n16996), .ZN(n16986) );
  NAND2_X1 U13008 ( .A1(n15178), .A2(n11733), .ZN(n15416) );
  NAND2_X1 U13009 ( .A1(n12739), .A2(n11741), .ZN(n12741) );
  NAND3_X1 U13010 ( .A1(n15304), .A2(n12820), .A3(n11742), .ZN(n11741) );
  INV_X1 U13011 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n11742) );
  INV_X1 U13012 ( .A(n15359), .ZN(n11745) );
  NAND2_X1 U13013 ( .A1(n11745), .A2(n11286), .ZN(n15523) );
  OAI21_X1 U13014 ( .B1(n16176), .B2(n17774), .A(n11755), .ZN(P2_U2983) );
  NOR2_X1 U13015 ( .A1(n13125), .A2(n13124), .ZN(n11756) );
  NAND3_X1 U13016 ( .A1(n11757), .A2(n17150), .A3(n16067), .ZN(n11760) );
  NAND2_X1 U13017 ( .A1(n16073), .A2(n11761), .ZN(n11759) );
  NAND2_X1 U13018 ( .A1(n19157), .A2(n14287), .ZN(n17131) );
  INV_X1 U13019 ( .A(n17193), .ZN(n11769) );
  NAND2_X1 U13020 ( .A1(n11764), .A2(n11763), .ZN(n11762) );
  NAND3_X1 U13021 ( .A1(n11772), .A2(n11771), .A3(n11770), .ZN(n14173) );
  INV_X1 U13022 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11775) );
  NAND2_X1 U13023 ( .A1(n11972), .A2(n11254), .ZN(n12662) );
  NAND2_X1 U13024 ( .A1(n11781), .A2(n11784), .ZN(n15694) );
  NAND2_X1 U13025 ( .A1(n11789), .A2(n11333), .ZN(n12928) );
  INV_X1 U13026 ( .A(n16702), .ZN(n11789) );
  AND2_X1 U13027 ( .A1(n12918), .A2(n11794), .ZN(n11796) );
  NAND2_X1 U13028 ( .A1(n11261), .A2(n11794), .ZN(n11793) );
  OAI21_X1 U13029 ( .B1(n16828), .B2(n22216), .A(n11798), .ZN(P1_U2970) );
  XNOR2_X1 U13030 ( .A(n13652), .B(n16670), .ZN(n16828) );
  NOR2_X1 U13031 ( .A1(n14144), .A2(n11800), .ZN(n14145) );
  AND2_X2 U13032 ( .A1(n11867), .A2(n11801), .ZN(n11959) );
  AND2_X2 U13033 ( .A1(n13330), .A2(n15226), .ZN(n13320) );
  NAND4_X1 U13034 ( .A1(n11802), .A2(n11803), .A3(n13121), .A4(n11804), .ZN(
        n13151) );
  NAND2_X1 U13035 ( .A1(n16888), .A2(n11806), .ZN(n15092) );
  NAND3_X1 U13036 ( .A1(n11809), .A2(n11326), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11808) );
  NAND2_X1 U13037 ( .A1(n12133), .A2(n12156), .ZN(n12216) );
  NAND2_X1 U13038 ( .A1(n12133), .A2(n11812), .ZN(n12890) );
  INV_X1 U13039 ( .A(n14061), .ZN(n11815) );
  NAND2_X1 U13040 ( .A1(n11815), .A2(n11816), .ZN(n15878) );
  NAND3_X1 U13041 ( .A1(n15299), .A2(n15424), .A3(n11821), .ZN(n14062) );
  AND2_X2 U13042 ( .A1(n16460), .A2(n12604), .ZN(n13649) );
  NAND2_X1 U13043 ( .A1(n16460), .A2(n11822), .ZN(n11825) );
  NAND2_X1 U13044 ( .A1(n16584), .A2(n11826), .ZN(n16513) );
  NAND2_X1 U13045 ( .A1(n12980), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12977) );
  CLKBUF_X1 U13046 ( .A(n12963), .Z(n19032) );
  INV_X1 U13047 ( .A(n14938), .ZN(n13194) );
  OAI21_X1 U13048 ( .B1(n15239), .B2(n17692), .A(n14703), .ZN(n14704) );
  INV_X1 U13049 ( .A(n15239), .ZN(n17634) );
  INV_X1 U13050 ( .A(n16423), .ZN(n14762) );
  AND2_X1 U13051 ( .A1(n13147), .A2(n13146), .ZN(n13149) );
  OAI21_X1 U13052 ( .B1(n14147), .B2(n14098), .A(n11178), .ZN(n14102) );
  NAND2_X1 U13053 ( .A1(n12929), .A2(n12930), .ZN(n16669) );
  NAND2_X1 U13054 ( .A1(n13116), .A2(n13106), .ZN(n13107) );
  INV_X1 U13055 ( .A(n12162), .ZN(n12164) );
  CLKBUF_X1 U13056 ( .A(n17569), .Z(n17570) );
  NAND2_X1 U13057 ( .A1(n12270), .A2(n12269), .ZN(n14061) );
  INV_X1 U13058 ( .A(n14062), .ZN(n12270) );
  AOI22_X1 U13059 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U13060 ( .A1(n11162), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13018) );
  NOR2_X1 U13061 ( .A1(n12842), .A2(n11176), .ZN(n11964) );
  CLKBUF_X1 U13062 ( .A(n15132), .Z(n16178) );
  NAND2_X1 U13063 ( .A1(n12898), .A2(n12338), .ZN(n12155) );
  NAND4_X1 U13064 ( .A1(n20030), .A2(n14710), .A3(n14405), .A4(n13104), .ZN(
        n13116) );
  AND2_X1 U13065 ( .A1(n13111), .A2(n14710), .ZN(n13088) );
  AND2_X1 U13066 ( .A1(n14457), .A2(n14456), .ZN(n11829) );
  AND3_X1 U13067 ( .A1(n13647), .A2(n13646), .A3(n13645), .ZN(n11830) );
  OR2_X1 U13068 ( .A1(n17013), .A2(n16307), .ZN(n11831) );
  NAND2_X1 U13069 ( .A1(n16659), .A2(n16596), .ZN(n11832) );
  AND2_X1 U13070 ( .A1(n17694), .A2(n19725), .ZN(n20234) );
  AND2_X1 U13071 ( .A1(n14482), .A2(n14481), .ZN(n11833) );
  AND2_X1 U13072 ( .A1(n14497), .A2(n14496), .ZN(n11834) );
  NAND3_X1 U13073 ( .A1(n14947), .A2(n13391), .A3(n13392), .ZN(n11836) );
  INV_X1 U13074 ( .A(n13357), .ZN(n13470) );
  INV_X1 U13075 ( .A(n13355), .ZN(n13469) );
  AND2_X1 U13076 ( .A1(n16326), .A2(n16346), .ZN(n11837) );
  OR2_X1 U13077 ( .A1(n13714), .A2(n13713), .ZN(n11838) );
  NOR2_X1 U13078 ( .A1(n21908), .A2(n13776), .ZN(n11839) );
  OR2_X1 U13079 ( .A1(n13681), .A2(n13680), .ZN(n11840) );
  AND4_X1 U13080 ( .A1(n14157), .A2(n14156), .A3(n14155), .A4(n14154), .ZN(
        n11841) );
  AND2_X1 U13081 ( .A1(n13731), .A2(n13730), .ZN(n11842) );
  AND2_X1 U13082 ( .A1(n14058), .A2(n14057), .ZN(n11843) );
  OR2_X1 U13083 ( .A1(n21080), .A2(n21066), .ZN(n11844) );
  INV_X1 U13084 ( .A(n12749), .ZN(n15352) );
  AND2_X1 U13085 ( .A1(n14059), .A2(n11843), .ZN(n11845) );
  NOR2_X1 U13086 ( .A1(DATAI_14_), .A2(n13659), .ZN(n11846) );
  AND4_X1 U13087 ( .A1(n14168), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        n11847) );
  OR2_X1 U13088 ( .A1(n21649), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11848) );
  NOR2_X1 U13089 ( .A1(n13897), .A2(keyinput_18), .ZN(n11849) );
  INV_X1 U13090 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12665) );
  INV_X1 U13091 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12953) );
  INV_X1 U13092 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18364) );
  AND2_X1 U13093 ( .A1(n12759), .A2(n12758), .ZN(n11850) );
  OR2_X1 U13094 ( .A1(n14764), .A2(n12732), .ZN(n11851) );
  AND2_X1 U13095 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11853) );
  AND2_X1 U13096 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11854) );
  NOR2_X1 U13097 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_67), .ZN(n11855)
         );
  AND2_X1 U13098 ( .A1(n16132), .A2(n16131), .ZN(n11856) );
  AOI21_X1 U13099 ( .B1(n14073), .B2(n20520), .A(n12949), .ZN(n12950) );
  INV_X1 U13100 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18432) );
  AOI22_X1 U13101 ( .A1(n16172), .A2(n17752), .B1(n16155), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n12963) );
  NOR2_X1 U13102 ( .A1(n14449), .A2(n13608), .ZN(n11857) );
  AND2_X1 U13103 ( .A1(n12660), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11858) );
  INV_X1 U13104 ( .A(n13105), .ZN(n13112) );
  AND2_X2 U13105 ( .A1(n14099), .A2(n14106), .ZN(n14152) );
  AND2_X2 U13106 ( .A1(n14104), .A2(n14106), .ZN(n14158) );
  AND2_X2 U13107 ( .A1(n14104), .A2(n14103), .ZN(n14150) );
  AND4_X1 U13108 ( .A1(n11958), .A2(n11957), .A3(n11956), .A4(n11955), .ZN(
        n11860) );
  CLKBUF_X3 U13109 ( .A(n12745), .Z(n12820) );
  INV_X1 U13110 ( .A(n12180), .ZN(n12264) );
  INV_X1 U13111 ( .A(keyinput_3), .ZN(n13669) );
  NAND2_X1 U13112 ( .A1(n13670), .A2(n13669), .ZN(n13671) );
  OAI22_X1 U13113 ( .A1(n22633), .A2(n13682), .B1(DATAI_20_), .B2(keyinput_12), 
        .ZN(n13683) );
  INV_X1 U13114 ( .A(n13683), .ZN(n13684) );
  OAI22_X1 U13115 ( .A1(n22558), .A2(keyinput_14), .B1(n13688), .B2(DATAI_18_), 
        .ZN(n13689) );
  INV_X1 U13116 ( .A(n13689), .ZN(n13690) );
  XNOR2_X1 U13117 ( .A(keyinput_17), .B(DATAI_15_), .ZN(n13693) );
  OAI22_X1 U13118 ( .A1(n13902), .A2(keyinput_20), .B1(n13701), .B2(DATAI_12_), 
        .ZN(n13702) );
  OAI22_X1 U13119 ( .A1(n17708), .A2(n13728), .B1(BS16), .B2(keyinput_35), 
        .ZN(n13729) );
  INV_X1 U13120 ( .A(keyinput_38), .ZN(n13733) );
  XNOR2_X1 U13121 ( .A(n13733), .B(P1_READREQUEST_REG_SCAN_IN), .ZN(n13734) );
  NAND2_X1 U13122 ( .A1(n13735), .A2(n13734), .ZN(n13736) );
  NOR2_X1 U13123 ( .A1(n11842), .A2(n13736), .ZN(n13739) );
  AOI211_X1 U13124 ( .C1(n13746), .C2(n13745), .A(n13744), .B(n13743), .ZN(
        n13747) );
  OAI22_X1 U13125 ( .A1(n16547), .A2(keyinput_65), .B1(n13769), .B2(
        P1_REIP_REG_18__SCAN_IN), .ZN(n13770) );
  NAND2_X1 U13126 ( .A1(n13773), .A2(n13772), .ZN(n13774) );
  OAI22_X1 U13127 ( .A1(n16849), .A2(n13783), .B1(P1_REIP_REG_14__SCAN_IN), 
        .B2(keyinput_69), .ZN(n13784) );
  OAI22_X1 U13128 ( .A1(n15940), .A2(n13785), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(keyinput_70), .ZN(n13786) );
  INV_X1 U13129 ( .A(n13786), .ZN(n13787) );
  NAND2_X1 U13130 ( .A1(n13792), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n13793) );
  NAND2_X1 U13131 ( .A1(n13794), .A2(n13793), .ZN(n13795) );
  XNOR2_X1 U13132 ( .A(n22122), .B(keyinput_101), .ZN(n13828) );
  NOR2_X1 U13133 ( .A1(n13829), .A2(n13828), .ZN(n13830) );
  INV_X1 U13134 ( .A(keyinput_110), .ZN(n13839) );
  XNOR2_X1 U13135 ( .A(n13839), .B(P1_EBX_REG_5__SCAN_IN), .ZN(n13840) );
  INV_X1 U13136 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13849) );
  NAND2_X1 U13137 ( .A1(n13850), .A2(n13849), .ZN(n13851) );
  NAND2_X1 U13138 ( .A1(n16423), .A2(n11851), .ZN(n11969) );
  NAND2_X1 U13139 ( .A1(n13123), .A2(n13105), .ZN(n14252) );
  NAND2_X1 U13140 ( .A1(n13105), .A2(n14257), .ZN(n13106) );
  INV_X1 U13141 ( .A(n12700), .ZN(n12679) );
  AND4_X1 U13142 ( .A1(n11898), .A2(n11897), .A3(n11896), .A4(n11895), .ZN(
        n11906) );
  AOI22_X1 U13143 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13098) );
  OR2_X1 U13144 ( .A1(n12043), .A2(n12042), .ZN(n12909) );
  AND2_X1 U13145 ( .A1(n12057), .A2(n12056), .ZN(n12085) );
  NAND2_X1 U13146 ( .A1(n13311), .A2(n13300), .ZN(n13306) );
  NAND2_X1 U13147 ( .A1(n13639), .A2(n16071), .ZN(n14453) );
  INV_X1 U13148 ( .A(n14204), .ZN(n14205) );
  AOI22_X1 U13149 ( .A1(n11162), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13085) );
  OR2_X1 U13150 ( .A1(n12682), .A2(n12681), .ZN(n12684) );
  NAND2_X1 U13151 ( .A1(n12014), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12705) );
  OR2_X1 U13152 ( .A1(n16530), .A2(n16546), .ZN(n12435) );
  NOR2_X1 U13153 ( .A1(n12599), .A2(n16698), .ZN(n12600) );
  INV_X1 U13154 ( .A(n16658), .ZN(n12364) );
  INV_X1 U13155 ( .A(n15342), .ZN(n15343) );
  AND2_X1 U13156 ( .A1(n16329), .A2(n11837), .ZN(n16330) );
  NAND2_X1 U13157 ( .A1(n15852), .A2(n14393), .ZN(n14392) );
  NOR2_X1 U13158 ( .A1(n13433), .A2(n13432), .ZN(n14169) );
  OR2_X1 U13159 ( .A1(n16948), .A2(n16060), .ZN(n17205) );
  AND3_X1 U13160 ( .A1(n17230), .A2(n17243), .A3(n17226), .ZN(n16039) );
  NAND2_X1 U13161 ( .A1(n14178), .A2(n14176), .ZN(n14280) );
  INV_X1 U13162 ( .A(n20956), .ZN(n20952) );
  INV_X1 U13163 ( .A(n21180), .ZN(n21368) );
  NAND2_X1 U13164 ( .A1(n12684), .A2(n12683), .ZN(n12686) );
  NAND2_X1 U13165 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12193) );
  INV_X1 U13166 ( .A(n12654), .ZN(n12619) );
  NAND2_X1 U13167 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11936) );
  AND2_X1 U13168 ( .A1(n12600), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12656) );
  NAND2_X1 U13169 ( .A1(n12556), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12599) );
  NOR2_X1 U13170 ( .A1(n12395), .A2(n22153), .ZN(n12396) );
  AND2_X1 U13171 ( .A1(n21855), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12660) );
  OR2_X1 U13172 ( .A1(n12104), .A2(n12103), .ZN(n12868) );
  INV_X1 U13173 ( .A(n16788), .ZN(n21918) );
  AND2_X1 U13174 ( .A1(n12744), .A2(n12743), .ZN(n14906) );
  AND2_X1 U13175 ( .A1(n14583), .A2(n14570), .ZN(n14900) );
  NAND2_X1 U13176 ( .A1(n12094), .A2(n12093), .ZN(n15133) );
  BUF_X1 U13177 ( .A(n11158), .Z(n14540) );
  INV_X1 U13178 ( .A(n17099), .ZN(n13591) );
  NOR2_X2 U13179 ( .A1(n14374), .A2(n14372), .ZN(n14463) );
  INV_X1 U13180 ( .A(n13622), .ZN(n14297) );
  AOI21_X1 U13181 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19777), .A(
        n13302), .ZN(n13304) );
  INV_X1 U13182 ( .A(n15904), .ZN(n15901) );
  NAND2_X1 U13183 ( .A1(n15344), .A2(n15343), .ZN(n15345) );
  AND2_X1 U13184 ( .A1(n13204), .A2(n13203), .ZN(n15153) );
  INV_X1 U13185 ( .A(n14884), .ZN(n13193) );
  INV_X1 U13186 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12959) );
  NAND2_X1 U13187 ( .A1(n15689), .A2(n15690), .ZN(n15688) );
  AND2_X1 U13188 ( .A1(n13210), .A2(n13209), .ZN(n15187) );
  AND2_X1 U13189 ( .A1(n14402), .A2(n11255), .ZN(n13150) );
  NOR2_X1 U13190 ( .A1(n17162), .A2(n16076), .ZN(n17128) );
  INV_X1 U13191 ( .A(n17297), .ZN(n14339) );
  INV_X1 U13192 ( .A(n15549), .ZN(n17585) );
  NAND2_X1 U13193 ( .A1(n18386), .A2(n21152), .ZN(n18389) );
  NOR2_X1 U13194 ( .A1(n18757), .A2(n18756), .ZN(n18755) );
  NAND2_X1 U13195 ( .A1(n18765), .A2(n18766), .ZN(n18764) );
  XNOR2_X1 U13196 ( .A(n18365), .B(n18364), .ZN(n18812) );
  NAND2_X1 U13197 ( .A1(n22095), .A2(n14068), .ZN(n22103) );
  NOR2_X1 U13198 ( .A1(n12193), .A2(n22037), .ZN(n12207) );
  XNOR2_X1 U13199 ( .A(n12061), .B(n12060), .ZN(n12179) );
  AND2_X2 U13200 ( .A1(n15391), .A2(n11177), .ZN(n21857) );
  NAND2_X1 U13201 ( .A1(n12396), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12432) );
  AND2_X1 U13202 ( .A1(n14798), .A2(n12187), .ZN(n14840) );
  AND2_X1 U13203 ( .A1(n20552), .A2(n16758), .ZN(n16836) );
  INV_X1 U13204 ( .A(n22015), .ZN(n16851) );
  XNOR2_X1 U13205 ( .A(n12170), .B(n12169), .ZN(n15132) );
  AND2_X1 U13206 ( .A1(n15286), .A2(n15285), .ZN(n22428) );
  INV_X1 U13207 ( .A(n22428), .ZN(n22442) );
  OR2_X1 U13208 ( .A1(n16178), .A2(n15112), .ZN(n15498) );
  INV_X1 U13209 ( .A(n22427), .ZN(n15470) );
  AOI21_X1 U13210 ( .B1(n22485), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n22411), 
        .ZN(n22447) );
  AND2_X1 U13211 ( .A1(n14397), .A2(n14396), .ZN(n15254) );
  NAND2_X1 U13212 ( .A1(n14361), .A2(n14362), .ZN(n14359) );
  OR2_X1 U13213 ( .A1(n18968), .A2(n13611), .ZN(n19111) );
  INV_X1 U13214 ( .A(n16307), .ZN(n16305) );
  NAND2_X1 U13215 ( .A1(n13337), .A2(n16136), .ZN(n13572) );
  AND2_X1 U13216 ( .A1(n16117), .A2(n16126), .ZN(n16118) );
  OR2_X1 U13217 ( .A1(n14503), .A2(n19182), .ZN(n14441) );
  AND2_X1 U13218 ( .A1(n15932), .A2(n14343), .ZN(n17283) );
  INV_X1 U13219 ( .A(n17570), .ZN(n17571) );
  INV_X1 U13220 ( .A(n19189), .ZN(n17622) );
  INV_X1 U13221 ( .A(n19888), .ZN(n19895) );
  INV_X1 U13222 ( .A(n19824), .ZN(n19836) );
  INV_X1 U13223 ( .A(n20234), .ZN(n19914) );
  INV_X1 U13224 ( .A(n19790), .ZN(n19791) );
  INV_X1 U13225 ( .A(n19823), .ZN(n19884) );
  INV_X1 U13226 ( .A(n19880), .ZN(n19908) );
  NOR2_X1 U13227 ( .A1(n21369), .A2(n21339), .ZN(n16001) );
  NAND2_X1 U13228 ( .A1(n21067), .A2(n11844), .ZN(n21068) );
  INV_X1 U13229 ( .A(n21108), .ZN(n21062) );
  NAND2_X1 U13230 ( .A1(n20682), .A2(n21115), .ZN(n20686) );
  NOR2_X1 U13231 ( .A1(n15982), .A2(n21321), .ZN(n18393) );
  INV_X1 U13232 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18752) );
  INV_X1 U13233 ( .A(n18391), .ZN(n18390) );
  INV_X2 U13234 ( .A(n21606), .ZN(n21775) );
  INV_X1 U13235 ( .A(n21366), .ZN(n21369) );
  INV_X1 U13236 ( .A(n16422), .ZN(n16421) );
  NAND2_X1 U13237 ( .A1(n12283), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12311) );
  NOR2_X1 U13238 ( .A1(n22082), .A2(n22083), .ZN(n22095) );
  INV_X1 U13239 ( .A(n22152), .ZN(n22206) );
  AND2_X1 U13240 ( .A1(n12451), .A2(n12450), .ZN(n16573) );
  INV_X1 U13241 ( .A(n22337), .ZN(n22400) );
  AOI21_X1 U13242 ( .B1(n20520), .B2(n16453), .A(n13654), .ZN(n13655) );
  NAND2_X1 U13243 ( .A1(n12516), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12554) );
  NAND2_X1 U13244 ( .A1(n12414), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12467) );
  INV_X1 U13245 ( .A(n20506), .ZN(n20551) );
  AND2_X1 U13246 ( .A1(n17733), .A2(n15124), .ZN(n20556) );
  INV_X1 U13247 ( .A(n22010), .ZN(n22004) );
  AND2_X1 U13248 ( .A1(n14583), .A2(n15125), .ZN(n22015) );
  AND2_X1 U13249 ( .A1(n22428), .A2(n15463), .ZN(n22743) );
  INV_X1 U13250 ( .A(n22760), .ZN(n15633) );
  INV_X1 U13251 ( .A(n22710), .ZN(n22713) );
  INV_X1 U13252 ( .A(n22795), .ZN(n22781) );
  AND2_X1 U13253 ( .A1(n15436), .A2(n15463), .ZN(n22791) );
  AND2_X1 U13254 ( .A1(n17744), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17718) );
  OR2_X1 U13255 ( .A1(n15257), .A2(n13317), .ZN(n15270) );
  INV_X1 U13256 ( .A(n19111), .ZN(n19155) );
  INV_X1 U13257 ( .A(n14864), .ZN(n17757) );
  AND2_X1 U13258 ( .A1(n19929), .A2(n14747), .ZN(n20223) );
  INV_X1 U13259 ( .A(n14216), .ZN(n18958) );
  NOR2_X1 U13260 ( .A1(n14599), .A2(n11178), .ZN(n14678) );
  INV_X1 U13261 ( .A(n17762), .ZN(n17780) );
  AND2_X1 U13262 ( .A1(n14279), .A2(n18966), .ZN(n14421) );
  NAND2_X1 U13263 ( .A1(n17641), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17659) );
  OAI21_X1 U13264 ( .B1(n20335), .B2(n19915), .A(n19914), .ZN(n20341) );
  NOR2_X1 U13265 ( .A1(n19863), .A2(n19845), .ZN(n19888) );
  OAI21_X1 U13266 ( .B1(n19857), .B2(n19856), .A(n19855), .ZN(n20309) );
  NOR2_X1 U13267 ( .A1(n19745), .A2(n19732), .ZN(n19823) );
  OAI21_X1 U13268 ( .B1(n19806), .B2(n20283), .A(n19914), .ZN(n20286) );
  AND2_X1 U13269 ( .A1(n19745), .A2(n19743), .ZN(n19801) );
  NOR2_X1 U13270 ( .A1(n19791), .A2(n19884), .ZN(n20190) );
  AND2_X1 U13271 ( .A1(n19745), .A2(n19732), .ZN(n19860) );
  NOR2_X1 U13272 ( .A1(n19791), .A2(n19846), .ZN(n20040) );
  NOR2_X1 U13273 ( .A1(n19746), .A2(n19835), .ZN(n20261) );
  NAND2_X1 U13274 ( .A1(n21043), .A2(n21042), .ZN(n21055) );
  INV_X1 U13275 ( .A(n21072), .ZN(n21106) );
  INV_X1 U13276 ( .A(n21107), .ZN(n21087) );
  NOR2_X1 U13277 ( .A1(n21828), .A2(n20686), .ZN(n20980) );
  AND2_X1 U13278 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18219), .ZN(n18145) );
  NOR3_X1 U13279 ( .A1(n21179), .A2(n21271), .A3(n21218), .ZN(n21206) );
  NOR3_X1 U13280 ( .A1(n22290), .A2(n21797), .A3(n21847), .ZN(n21118) );
  INV_X2 U13281 ( .A(n18620), .ZN(n18672) );
  INV_X1 U13282 ( .A(n21720), .ZN(n21673) );
  NOR2_X1 U13283 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18669), .ZN(
        n18668) );
  NOR2_X2 U13284 ( .A1(n21655), .A2(n21476), .ZN(n21779) );
  INV_X1 U13285 ( .A(n21728), .ZN(n21789) );
  INV_X1 U13286 ( .A(n21755), .ZN(n21681) );
  INV_X1 U13287 ( .A(n18834), .ZN(n19584) );
  INV_X1 U13288 ( .A(U212), .ZN(n20608) );
  NAND2_X1 U13289 ( .A1(n14763), .A2(n16421), .ZN(n22813) );
  OR2_X1 U13290 ( .A1(n16434), .A2(n13752), .ZN(n12840) );
  INV_X1 U13291 ( .A(n22165), .ZN(n22208) );
  NAND2_X1 U13292 ( .A1(n14075), .A2(n12729), .ZN(n22209) );
  INV_X1 U13293 ( .A(n22166), .ZN(n22201) );
  NAND2_X1 U13294 ( .A1(n14894), .A2(n14893), .ZN(n16659) );
  INV_X1 U13295 ( .A(n20381), .ZN(n20401) );
  OR2_X1 U13296 ( .A1(n22813), .A2(n14765), .ZN(n22399) );
  NAND2_X2 U13297 ( .A1(n14766), .A2(n15391), .ZN(n22405) );
  INV_X1 U13298 ( .A(n20520), .ZN(n20561) );
  OR2_X1 U13299 ( .A1(n20556), .A2(n12945), .ZN(n20506) );
  INV_X1 U13300 ( .A(n22170), .ZN(n21975) );
  INV_X1 U13301 ( .A(n21993), .ZN(n22009) );
  INV_X1 U13302 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22485) );
  AOI22_X1 U13303 ( .A1(n22409), .A2(n22419), .B1(n22408), .B2(n22481), .ZN(
        n22741) );
  INV_X1 U13304 ( .A(n22743), .ZN(n22693) );
  INV_X1 U13305 ( .A(n22445), .ZN(n22754) );
  OR2_X1 U13306 ( .A1(n15461), .A2(n15471), .ZN(n22760) );
  NAND2_X1 U13307 ( .A1(n15310), .A2(n15435), .ZN(n22772) );
  AOI22_X1 U13308 ( .A1(n22483), .A2(n22491), .B1(n22482), .B2(n22481), .ZN(
        n22779) );
  INV_X1 U13309 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n17744) );
  INV_X1 U13310 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n22225) );
  OR2_X1 U13311 ( .A1(n15257), .A2(n13612), .ZN(n14599) );
  INV_X1 U13312 ( .A(n19156), .ZN(n19144) );
  AND4_X1 U13313 ( .A1(n15968), .A2(n15967), .A3(n15966), .A4(n15965), .ZN(
        n15969) );
  INV_X1 U13314 ( .A(n19845), .ZN(n17805) );
  NAND2_X1 U13315 ( .A1(n14746), .A2(n14745), .ZN(n19929) );
  INV_X1 U13316 ( .A(n19972), .ZN(n20176) );
  INV_X1 U13317 ( .A(n17823), .ZN(n17853) );
  INV_X1 U13318 ( .A(n14678), .ZN(n14732) );
  INV_X1 U13319 ( .A(n17754), .ZN(n17790) );
  INV_X1 U13320 ( .A(n17633), .ZN(n19184) );
  NAND2_X1 U13321 ( .A1(n19888), .A2(n19887), .ZN(n20334) );
  NAND2_X1 U13322 ( .A1(n19888), .A2(n19860), .ZN(n20326) );
  INV_X1 U13323 ( .A(n20315), .ZN(n20313) );
  NAND2_X1 U13324 ( .A1(n19824), .A2(n19823), .ZN(n20306) );
  NAND2_X1 U13325 ( .A1(n19801), .A2(n19824), .ZN(n20294) );
  INV_X1 U13326 ( .A(n20190), .ZN(n20282) );
  INV_X1 U13327 ( .A(n20040), .ZN(n20270) );
  INV_X1 U13328 ( .A(n20109), .ZN(n20119) );
  INV_X1 U13329 ( .A(n20011), .ZN(n20019) );
  OR2_X1 U13330 ( .A1(n19746), .A2(n19846), .ZN(n20344) );
  AND2_X1 U13331 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18183), .ZN(n18177) );
  INV_X1 U13332 ( .A(n18271), .ZN(n18248) );
  NOR3_X1 U13333 ( .A1(n20684), .A2(n19589), .A3(n21114), .ZN(n18273) );
  INV_X1 U13334 ( .A(n21270), .ZN(n21253) );
  INV_X1 U13335 ( .A(n21290), .ZN(n21295) );
  INV_X1 U13336 ( .A(n18400), .ZN(n21655) );
  NOR2_X1 U13337 ( .A1(n18299), .A2(n18298), .ZN(n21156) );
  INV_X1 U13338 ( .A(n21302), .ZN(n21300) );
  INV_X1 U13339 ( .A(n18888), .ZN(n18887) );
  INV_X1 U13340 ( .A(n21779), .ZN(n21741) );
  INV_X1 U13341 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21815) );
  AOI22_X1 U13342 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11865) );
  AND2_X2 U13343 ( .A1(n11867), .A2(n15098), .ZN(n12456) );
  AOI22_X1 U13344 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U13345 ( .A1(n11907), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11863) );
  AND2_X2 U13346 ( .A1(n15076), .A2(n15098), .ZN(n11914) );
  AOI22_X1 U13347 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11914), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11862) );
  NAND4_X1 U13348 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11874) );
  AND2_X2 U13349 ( .A1(n11867), .A2(n15090), .ZN(n11885) );
  AND2_X4 U13350 ( .A1(n11868), .A2(n15076), .ZN(n12525) );
  AOI22_X1 U13351 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11872) );
  AND2_X2 U13352 ( .A1(n15090), .A2(n11866), .ZN(n11908) );
  AND2_X2 U13353 ( .A1(n11867), .A2(n11868), .ZN(n12108) );
  AOI22_X1 U13354 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11871) );
  AND2_X2 U13355 ( .A1(n16896), .A2(n11868), .ZN(n11937) );
  AOI22_X1 U13356 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11937), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11870) );
  AND2_X2 U13357 ( .A1(n16896), .A2(n15098), .ZN(n12037) );
  AOI22_X1 U13358 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11869) );
  NAND4_X1 U13359 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11873) );
  OR2_X2 U13360 ( .A1(n11874), .A2(n11873), .ZN(n11922) );
  AOI22_X1 U13361 ( .A1(n12626), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U13362 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U13363 ( .A1(n11907), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U13364 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11914), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11875) );
  NAND4_X1 U13365 ( .A1(n11878), .A2(n11877), .A3(n11876), .A4(n11875), .ZN(
        n11884) );
  AOI22_X1 U13366 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U13367 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U13368 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11937), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U13369 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11879) );
  NAND4_X1 U13370 ( .A1(n11882), .A2(n11881), .A3(n11880), .A4(n11879), .ZN(
        n11883) );
  AOI22_X1 U13371 ( .A1(n11907), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12626), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U13372 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11888) );
  BUF_X2 U13373 ( .A(n11914), .Z(n12629) );
  AOI22_X1 U13374 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11937), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U13375 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U13376 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U13377 ( .A1(n11913), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U13378 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U13379 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12048), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U13380 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U13381 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11937), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U13382 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11914), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U13383 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U13384 ( .A1(n11913), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11899) );
  NAND2_X1 U13385 ( .A1(n11900), .A2(n11899), .ZN(n11904) );
  AOI22_X1 U13386 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U13387 ( .A1(n11907), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11901) );
  NAND2_X1 U13388 ( .A1(n11902), .A2(n11901), .ZN(n11903) );
  NOR2_X1 U13389 ( .A1(n11904), .A2(n11903), .ZN(n11905) );
  AOI22_X1 U13390 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11907), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U13391 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U13392 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U13393 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11909) );
  NAND4_X1 U13394 ( .A1(n11912), .A2(n11911), .A3(n11910), .A4(n11909), .ZN(
        n11920) );
  AOI22_X1 U13395 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12048), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11918) );
  BUF_X4 U13396 ( .A(n11937), .Z(n12380) );
  AOI22_X1 U13397 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11916) );
  BUF_X4 U13398 ( .A(n11914), .Z(n12582) );
  AOI22_X1 U13399 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11915) );
  NAND4_X1 U13400 ( .A1(n11918), .A2(n11917), .A3(n11916), .A4(n11915), .ZN(
        n11919) );
  OR2_X2 U13401 ( .A1(n11920), .A2(n11919), .ZN(n15309) );
  NAND2_X1 U13402 ( .A1(n14580), .A2(n15309), .ZN(n11979) );
  INV_X2 U13403 ( .A(n11922), .ZN(n15529) );
  NAND2_X2 U13404 ( .A1(n15529), .A2(n16595), .ZN(n14895) );
  AOI22_X1 U13405 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U13406 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U13407 ( .A1(n11907), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U13408 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11923) );
  NAND4_X1 U13409 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11932) );
  AOI22_X1 U13410 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U13411 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U13412 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U13413 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11927) );
  NAND4_X1 U13414 ( .A1(n11930), .A2(n11929), .A3(n11928), .A4(n11927), .ZN(
        n11931) );
  OR2_X2 U13415 ( .A1(n11932), .A2(n11931), .ZN(n12842) );
  NAND2_X1 U13416 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11935) );
  NAND2_X1 U13417 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11934) );
  NAND2_X1 U13418 ( .A1(n12629), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11933) );
  NAND2_X1 U13419 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U13420 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11940) );
  NAND2_X1 U13421 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11939) );
  NAND2_X1 U13422 ( .A1(n12630), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11938) );
  NAND2_X1 U13423 ( .A1(n12626), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11945) );
  NAND2_X1 U13424 ( .A1(n11907), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11944) );
  NAND2_X1 U13425 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11943) );
  NAND2_X1 U13426 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11949) );
  NAND2_X1 U13427 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11948) );
  NAND2_X1 U13428 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11947) );
  NAND2_X1 U13429 ( .A1(n12037), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11946) );
  NAND4_X4 U13430 ( .A1(n11953), .A2(n11952), .A3(n11951), .A4(n11950), .ZN(
        n15127) );
  NOR2_X1 U13431 ( .A1(n14559), .A2(n15127), .ZN(n11954) );
  AOI22_X1 U13432 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U13433 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11937), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U13434 ( .A1(n11907), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U13435 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U13436 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U13437 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U13438 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U13439 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11960) );
  INV_X1 U13440 ( .A(n12662), .ZN(n11971) );
  OR2_X2 U13441 ( .A1(n14783), .A2(n16591), .ZN(n14581) );
  AND2_X1 U13442 ( .A1(n15309), .A2(n15127), .ZN(n11965) );
  AND2_X2 U13443 ( .A1(n11966), .A2(n11965), .ZN(n16423) );
  INV_X1 U13444 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20562) );
  NAND2_X1 U13445 ( .A1(n20562), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22266) );
  INV_X1 U13446 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n11967) );
  NAND2_X1 U13447 ( .A1(n11967), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n11968) );
  NAND2_X1 U13448 ( .A1(n22266), .A2(n11968), .ZN(n12732) );
  NAND2_X1 U13449 ( .A1(n14581), .A2(n11969), .ZN(n11970) );
  NOR2_X1 U13450 ( .A1(n11971), .A2(n11970), .ZN(n11986) );
  NAND2_X1 U13451 ( .A1(n11973), .A2(n14548), .ZN(n14567) );
  NAND2_X1 U13452 ( .A1(n15592), .A2(n11922), .ZN(n11974) );
  NAND2_X1 U13453 ( .A1(n11974), .A2(n15309), .ZN(n12939) );
  OR2_X1 U13454 ( .A1(n12939), .A2(n14580), .ZN(n11977) );
  NAND2_X1 U13455 ( .A1(n12842), .A2(n14764), .ZN(n12745) );
  OR2_X1 U13456 ( .A1(n14559), .A2(n12745), .ZN(n14784) );
  NAND2_X1 U13457 ( .A1(n22414), .A2(n14764), .ZN(n14777) );
  NAND2_X1 U13458 ( .A1(n14784), .A2(n14777), .ZN(n11975) );
  AOI21_X1 U13459 ( .B1(n21857), .B2(n11977), .A(n11975), .ZN(n11976) );
  INV_X1 U13460 ( .A(n11977), .ZN(n11978) );
  NAND2_X1 U13461 ( .A1(n14554), .A2(n11177), .ZN(n14561) );
  INV_X1 U13462 ( .A(n14558), .ZN(n11996) );
  NAND2_X1 U13463 ( .A1(n14561), .A2(n11996), .ZN(n11980) );
  NAND3_X1 U13464 ( .A1(n11986), .A2(n11993), .A3(n11981), .ZN(n11982) );
  NAND2_X1 U13465 ( .A1(n11982), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11989) );
  NAND2_X1 U13466 ( .A1(n22464), .A2(n17744), .ZN(n17669) );
  XNOR2_X1 U13467 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22432) );
  INV_X1 U13468 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15451) );
  OR2_X1 U13469 ( .A1(n17718), .A2(n15451), .ZN(n12002) );
  OAI21_X1 U13470 ( .B1(n12947), .B2(n22432), .A(n12002), .ZN(n11984) );
  INV_X1 U13471 ( .A(n11984), .ZN(n11985) );
  OAI21_X1 U13472 ( .B1(n11989), .B2(n11983), .A(n11985), .ZN(n11988) );
  INV_X1 U13473 ( .A(n11986), .ZN(n11987) );
  INV_X1 U13474 ( .A(n11989), .ZN(n12006) );
  NAND2_X1 U13475 ( .A1(n12006), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11992) );
  INV_X1 U13476 ( .A(n17718), .ZN(n12091) );
  INV_X1 U13477 ( .A(n12947), .ZN(n12092) );
  MUX2_X1 U13478 ( .A(n12091), .B(n12092), .S(n22485), .Z(n11990) );
  INV_X1 U13479 ( .A(n11990), .ZN(n11991) );
  INV_X1 U13480 ( .A(n11993), .ZN(n12001) );
  NAND3_X1 U13481 ( .A1(n14535), .A2(n14764), .A3(n14789), .ZN(n11999) );
  OR2_X1 U13482 ( .A1(n17669), .A2(n22225), .ZN(n11994) );
  AOI21_X1 U13483 ( .B1(n14776), .B2(n15127), .A(n11994), .ZN(n11998) );
  INV_X1 U13484 ( .A(n14548), .ZN(n15406) );
  NAND2_X1 U13485 ( .A1(n14730), .A2(n11995), .ZN(n11997) );
  OR2_X1 U13486 ( .A1(n11996), .A2(n11922), .ZN(n14568) );
  NAND4_X1 U13487 ( .A1(n11999), .A2(n11998), .A3(n11997), .A4(n14568), .ZN(
        n12000) );
  NAND2_X1 U13489 ( .A1(n12061), .A2(n12059), .ZN(n12031) );
  INV_X1 U13490 ( .A(n12002), .ZN(n12004) );
  NAND2_X1 U13491 ( .A1(n12006), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12012) );
  NAND2_X1 U13492 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12007) );
  NAND2_X1 U13493 ( .A1(n12665), .A2(n12007), .ZN(n12009) );
  NAND2_X1 U13494 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22463) );
  INV_X1 U13495 ( .A(n22463), .ZN(n12008) );
  NAND2_X1 U13496 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12008), .ZN(
        n15375) );
  NAND2_X1 U13497 ( .A1(n12009), .A2(n15375), .ZN(n15138) );
  OAI22_X1 U13498 ( .A1(n12947), .A2(n15138), .B1(n17718), .B2(n12665), .ZN(
        n12010) );
  INV_X1 U13499 ( .A(n12010), .ZN(n12011) );
  NAND2_X1 U13500 ( .A1(n12012), .A2(n12011), .ZN(n12013) );
  INV_X1 U13501 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U13502 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12626), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U13503 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U13504 ( .A1(n12637), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U13505 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U13506 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12025) );
  AOI22_X1 U13507 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U13508 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U13509 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U13510 ( .A1(n12062), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12020) );
  NAND4_X1 U13511 ( .A1(n12023), .A2(n12022), .A3(n12021), .A4(n12020), .ZN(
        n12024) );
  NOR2_X1 U13512 ( .A1(n12025), .A2(n12024), .ZN(n12858) );
  OAI22_X1 U13513 ( .A1(n12695), .A2(n12026), .B1(n12705), .B2(n12858), .ZN(
        n12027) );
  NAND2_X1 U13515 ( .A1(n12030), .A2(n12031), .ZN(n15397) );
  OR2_X2 U13516 ( .A1(n15134), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12084) );
  NOR2_X1 U13517 ( .A1(n14580), .A2(n22225), .ZN(n12081) );
  AOI22_X1 U13518 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U13519 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U13520 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U13521 ( .A1(n12062), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12033) );
  NAND4_X1 U13522 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        n12043) );
  AOI22_X1 U13523 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U13524 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11370), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U13525 ( .A1(n12637), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U13527 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12038) );
  NAND4_X1 U13528 ( .A1(n12041), .A2(n12040), .A3(n12039), .A4(n12038), .ZN(
        n12042) );
  NOR2_X1 U13529 ( .A1(n15127), .A2(n22225), .ZN(n12055) );
  AOI22_X1 U13530 ( .A1(n12062), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U13531 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U13532 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12044) );
  NAND4_X1 U13533 ( .A1(n12047), .A2(n12046), .A3(n12045), .A4(n12044), .ZN(
        n12054) );
  CLKBUF_X1 U13534 ( .A(n12048), .Z(n12605) );
  AOI22_X1 U13535 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U13536 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U13537 ( .A1(n12630), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U13538 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12049) );
  NAND4_X1 U13539 ( .A1(n12052), .A2(n12051), .A3(n12050), .A4(n12049), .ZN(
        n12053) );
  AOI22_X1 U13540 ( .A1(n12081), .A2(n12146), .B1(n12055), .B2(n12855), .ZN(
        n12057) );
  NAND2_X1 U13541 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12056) );
  NAND2_X1 U13542 ( .A1(n12081), .A2(n12855), .ZN(n12083) );
  AND2_X1 U13543 ( .A1(n12085), .A2(n12083), .ZN(n12058) );
  NAND2_X1 U13544 ( .A1(n12179), .A2(n22225), .ZN(n12076) );
  AOI22_X1 U13545 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12626), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U13546 ( .A1(n11885), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12065) );
  BUF_X1 U13547 ( .A(n12108), .Z(n12062) );
  AOI22_X1 U13548 ( .A1(n12062), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U13549 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U13550 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12073) );
  AOI22_X1 U13551 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U13552 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U13553 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U13554 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12068) );
  NAND4_X1 U13555 ( .A1(n12071), .A2(n12070), .A3(n12069), .A4(n12068), .ZN(
        n12072) );
  XNOR2_X1 U13556 ( .A(n12146), .B(n12856), .ZN(n12074) );
  NAND2_X1 U13557 ( .A1(n12074), .A2(n12081), .ZN(n12075) );
  NAND2_X1 U13558 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12080) );
  NAND2_X1 U13559 ( .A1(n22414), .A2(n12856), .ZN(n12077) );
  OAI211_X1 U13560 ( .C1(n12146), .C2(n14580), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n12077), .ZN(n12078) );
  INV_X1 U13561 ( .A(n12078), .ZN(n12079) );
  NAND2_X1 U13562 ( .A1(n12080), .A2(n12079), .ZN(n12176) );
  NAND2_X1 U13563 ( .A1(n12177), .A2(n12176), .ZN(n12082) );
  NAND2_X1 U13564 ( .A1(n12081), .A2(n12909), .ZN(n12907) );
  NAND2_X1 U13565 ( .A1(n12170), .A2(n12168), .ZN(n12088) );
  NAND2_X1 U13566 ( .A1(n12084), .A2(n12083), .ZN(n12845) );
  INV_X1 U13567 ( .A(n12085), .ZN(n12086) );
  NAND2_X1 U13568 ( .A1(n12845), .A2(n12086), .ZN(n12087) );
  NAND2_X1 U13569 ( .A1(n12088), .A2(n12087), .ZN(n12162) );
  NAND2_X1 U13570 ( .A1(n12163), .A2(n12162), .ZN(n12191) );
  NAND2_X1 U13571 ( .A1(n12006), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12094) );
  INV_X1 U13572 ( .A(n15375), .ZN(n12089) );
  INV_X1 U13573 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U13574 ( .A1(n12089), .A2(n12668), .ZN(n15467) );
  NAND2_X1 U13575 ( .A1(n15375), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12090) );
  NAND2_X1 U13576 ( .A1(n15467), .A2(n12090), .ZN(n15314) );
  AOI22_X1 U13577 ( .A1(n12092), .A2(n15314), .B1(n12091), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12093) );
  NAND2_X1 U13578 ( .A1(n15080), .A2(n22225), .ZN(n12106) );
  AOI22_X1 U13579 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U13580 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U13581 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U13582 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12104) );
  AOI22_X1 U13583 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U13584 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U13585 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U13586 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U13587 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12103) );
  AOI22_X1 U13588 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12720), .B1(
        n12696), .B2(n12868), .ZN(n12105) );
  NAND2_X1 U13589 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12120) );
  AOI22_X1 U13590 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12610), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U13591 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12635), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U13592 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U13593 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12109) );
  NAND4_X1 U13594 ( .A1(n12112), .A2(n12111), .A3(n12110), .A4(n12109), .ZN(
        n12118) );
  AOI22_X1 U13595 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12587), .B1(
        n12456), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U13596 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U13597 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U13598 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12525), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12113) );
  NAND4_X1 U13599 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12117) );
  NAND2_X1 U13600 ( .A1(n12696), .A2(n12881), .ZN(n12119) );
  NAND2_X1 U13601 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12132) );
  AOI22_X1 U13602 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U13603 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U13604 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U13605 ( .A1(n12637), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12121) );
  NAND4_X1 U13606 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12130) );
  AOI22_X1 U13607 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U13608 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U13609 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U13610 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12125) );
  NAND4_X1 U13611 ( .A1(n12128), .A2(n12127), .A3(n12126), .A4(n12125), .ZN(
        n12129) );
  OR2_X1 U13612 ( .A1(n12130), .A2(n12129), .ZN(n12884) );
  NAND2_X1 U13613 ( .A1(n12696), .A2(n12884), .ZN(n12131) );
  NAND2_X1 U13614 ( .A1(n12132), .A2(n12131), .ZN(n12156) );
  NAND2_X1 U13615 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12145) );
  AOI22_X1 U13616 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U13617 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U13618 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12134) );
  NAND4_X1 U13619 ( .A1(n12137), .A2(n12136), .A3(n12135), .A4(n12134), .ZN(
        n12143) );
  AOI22_X1 U13620 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U13621 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U13622 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U13623 ( .A1(n12062), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12138) );
  NAND4_X1 U13624 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n12138), .ZN(
        n12142) );
  OR2_X1 U13625 ( .A1(n12143), .A2(n12142), .ZN(n12900) );
  NAND2_X1 U13626 ( .A1(n12696), .A2(n12900), .ZN(n12144) );
  INV_X1 U13627 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12147) );
  OAI22_X1 U13628 ( .A1(n12695), .A2(n12147), .B1(n12705), .B2(n12146), .ZN(
        n12148) );
  NOR2_X2 U13629 ( .A1(n11922), .A2(n21855), .ZN(n12338) );
  NOR2_X1 U13630 ( .A1(n15309), .A2(n21855), .ZN(n12180) );
  INV_X1 U13631 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12149) );
  NOR2_X1 U13632 ( .A1(n12264), .A2(n12149), .ZN(n12153) );
  OR2_X1 U13633 ( .A1(n12218), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12150) );
  NAND2_X1 U13634 ( .A1(n12239), .A2(n12150), .ZN(n22091) );
  NOR2_X1 U13635 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17711) );
  AOI22_X1 U13636 ( .A1(n22091), .A2(n12657), .B1(n12660), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12151) );
  INV_X1 U13637 ( .A(n12151), .ZN(n12152) );
  INV_X1 U13638 ( .A(n12156), .ZN(n12157) );
  NAND2_X1 U13639 ( .A1(n12202), .A2(n12157), .ZN(n12158) );
  INV_X1 U13640 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12160) );
  OAI21_X1 U13641 ( .B1(n12209), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n12217), .ZN(n22075) );
  AOI22_X1 U13642 ( .A1(n22075), .A2(n12657), .B1(n12660), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12159) );
  OAI21_X1 U13643 ( .B1(n12264), .B2(n12160), .A(n12159), .ZN(n12161) );
  NAND2_X1 U13644 ( .A1(n12854), .A2(n12338), .ZN(n14870) );
  OR2_X1 U13645 ( .A1(n16591), .A2(n21855), .ZN(n12206) );
  XNOR2_X1 U13646 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n22020) );
  AOI21_X1 U13647 ( .B1(n17711), .B2(n22020), .A(n12660), .ZN(n12166) );
  NAND2_X1 U13648 ( .A1(n12652), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12165) );
  OAI211_X1 U13649 ( .C1(n12206), .C2(n11775), .A(n12166), .B(n12165), .ZN(
        n12167) );
  INV_X1 U13650 ( .A(n12167), .ZN(n14868) );
  INV_X1 U13651 ( .A(n12168), .ZN(n12169) );
  NAND2_X1 U13652 ( .A1(n15132), .A2(n12338), .ZN(n12175) );
  NAND2_X1 U13653 ( .A1(n12180), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n12172) );
  NAND2_X1 U13654 ( .A1(n21855), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12171) );
  OAI211_X1 U13655 ( .C1(n12206), .C2(n11983), .A(n12172), .B(n12171), .ZN(
        n12173) );
  INV_X1 U13656 ( .A(n12173), .ZN(n12174) );
  NAND2_X1 U13657 ( .A1(n12175), .A2(n12174), .ZN(n14839) );
  NAND2_X1 U13658 ( .A1(n15112), .A2(n15529), .ZN(n12178) );
  NAND2_X1 U13659 ( .A1(n12178), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14800) );
  NAND2_X1 U13660 ( .A1(n15412), .A2(n12338), .ZN(n12183) );
  INV_X1 U13661 ( .A(n12206), .ZN(n12181) );
  AOI22_X1 U13662 ( .A1(n12181), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n12180), .B2(P1_EAX_REG_0__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U13663 ( .A1(n12183), .A2(n12182), .ZN(n14799) );
  AND2_X1 U13664 ( .A1(n21855), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12184) );
  NAND2_X1 U13665 ( .A1(n14800), .A2(n12185), .ZN(n14798) );
  INV_X1 U13666 ( .A(n12185), .ZN(n12186) );
  NAND2_X1 U13667 ( .A1(n12186), .A2(n12650), .ZN(n12187) );
  NAND2_X1 U13668 ( .A1(n14839), .A2(n14840), .ZN(n14871) );
  INV_X1 U13669 ( .A(n14871), .ZN(n12188) );
  NOR2_X1 U13670 ( .A1(n11858), .A2(n12188), .ZN(n12189) );
  NOR2_X2 U13671 ( .A1(n12190), .A2(n12189), .ZN(n14890) );
  NAND2_X1 U13672 ( .A1(n12191), .A2(n15171), .ZN(n12192) );
  NAND2_X1 U13673 ( .A1(n12200), .A2(n12192), .ZN(n15285) );
  INV_X1 U13674 ( .A(n12338), .ZN(n12203) );
  INV_X1 U13675 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15088) );
  INV_X1 U13676 ( .A(n12193), .ZN(n12195) );
  INV_X1 U13677 ( .A(n12207), .ZN(n12194) );
  OAI21_X1 U13678 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12195), .A(
        n12194), .ZN(n22043) );
  AOI22_X1 U13679 ( .A1(n17711), .A2(n22043), .B1(n12660), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12197) );
  NAND2_X1 U13680 ( .A1(n12652), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12196) );
  OAI211_X1 U13681 ( .C1(n12206), .C2(n15088), .A(n12197), .B(n12196), .ZN(
        n12198) );
  INV_X1 U13682 ( .A(n12198), .ZN(n12199) );
  AND2_X2 U13683 ( .A1(n14890), .A2(n14889), .ZN(n14888) );
  NAND2_X1 U13684 ( .A1(n12200), .A2(n11285), .ZN(n12201) );
  NAND2_X1 U13685 ( .A1(n12202), .A2(n12201), .ZN(n12873) );
  INV_X1 U13686 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17673) );
  INV_X1 U13687 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21856) );
  OAI21_X1 U13688 ( .B1(n21856), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21855), .ZN(n12205) );
  NAND2_X1 U13689 ( .A1(n12652), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12204) );
  OAI211_X1 U13690 ( .C1(n12206), .C2(n17673), .A(n12205), .B(n12204), .ZN(
        n12211) );
  NOR2_X1 U13691 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12207), .ZN(
        n12208) );
  NOR2_X1 U13692 ( .A1(n12209), .A2(n12208), .ZN(n15162) );
  NAND2_X1 U13693 ( .A1(n15162), .A2(n12657), .ZN(n12210) );
  NAND2_X1 U13694 ( .A1(n12211), .A2(n12210), .ZN(n12212) );
  NAND2_X1 U13695 ( .A1(n12216), .A2(n12215), .ZN(n12891) );
  INV_X1 U13696 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n22351) );
  AND2_X1 U13697 ( .A1(n12217), .A2(n12220), .ZN(n12219) );
  OR2_X1 U13698 ( .A1(n12219), .A2(n12218), .ZN(n22087) );
  INV_X1 U13699 ( .A(n12660), .ZN(n12221) );
  NOR2_X1 U13700 ( .A1(n12221), .A2(n12220), .ZN(n12222) );
  AOI21_X1 U13701 ( .B1(n22087), .B2(n12657), .A(n12222), .ZN(n12223) );
  OAI21_X1 U13702 ( .B1(n12264), .B2(n22351), .A(n12223), .ZN(n12224) );
  AOI22_X1 U13703 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U13704 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U13705 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12225) );
  NAND4_X1 U13706 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12234) );
  AOI22_X1 U13707 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U13708 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U13709 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U13710 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12229) );
  NAND4_X1 U13711 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12233) );
  OAI21_X1 U13712 ( .B1(n12234), .B2(n12233), .A(n12338), .ZN(n12238) );
  NAND2_X1 U13713 ( .A1(n12652), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12237) );
  XNOR2_X1 U13714 ( .A(n12239), .B(n15488), .ZN(n15698) );
  NAND2_X1 U13715 ( .A1(n15698), .A2(n12657), .ZN(n12236) );
  NAND2_X1 U13716 ( .A1(n12660), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12235) );
  NAND4_X1 U13717 ( .A1(n12238), .A2(n12237), .A3(n12236), .A4(n12235), .ZN(
        n15427) );
  XOR2_X1 U13718 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12253), .Z(n15783) );
  AOI22_X1 U13719 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U13720 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U13721 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U13722 ( .A1(n12638), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12240) );
  NAND4_X1 U13723 ( .A1(n12243), .A2(n12242), .A3(n12241), .A4(n12240), .ZN(
        n12249) );
  AOI22_X1 U13724 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12626), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U13725 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U13726 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U13727 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12244) );
  NAND4_X1 U13728 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n12248) );
  OR2_X1 U13729 ( .A1(n12249), .A2(n12248), .ZN(n12250) );
  AOI22_X1 U13730 ( .A1(n12338), .A2(n12250), .B1(n12660), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12252) );
  NAND2_X1 U13731 ( .A1(n12652), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12251) );
  OAI211_X1 U13732 ( .C1(n15783), .C2(n12650), .A(n12252), .B(n12251), .ZN(
        n15562) );
  INV_X1 U13733 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14072) );
  XNOR2_X1 U13734 ( .A(n12282), .B(n14072), .ZN(n20507) );
  AOI22_X1 U13735 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U13736 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U13737 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U13738 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12254) );
  NAND4_X1 U13739 ( .A1(n12257), .A2(n12256), .A3(n12255), .A4(n12254), .ZN(
        n12263) );
  AOI22_X1 U13740 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U13741 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U13742 ( .A1(n12637), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U13743 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U13744 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12262) );
  OAI21_X1 U13745 ( .B1(n12263), .B2(n12262), .A(n12338), .ZN(n12267) );
  NAND2_X1 U13746 ( .A1(n12652), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12266) );
  NAND2_X1 U13747 ( .A1(n12660), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12265) );
  NAND3_X1 U13748 ( .A1(n12267), .A2(n12266), .A3(n12265), .ZN(n12268) );
  AOI21_X1 U13749 ( .B1(n20507), .B2(n12657), .A(n12268), .ZN(n14064) );
  INV_X1 U13750 ( .A(n14064), .ZN(n12269) );
  AOI22_X1 U13751 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U13752 ( .A1(n12637), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U13753 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12271) );
  NAND4_X1 U13754 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(
        n12280) );
  AOI22_X1 U13755 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U13756 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U13757 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U13758 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12275) );
  NAND4_X1 U13759 ( .A1(n12278), .A2(n12277), .A3(n12276), .A4(n12275), .ZN(
        n12279) );
  OR2_X1 U13760 ( .A1(n12280), .A2(n12279), .ZN(n12281) );
  NAND2_X1 U13761 ( .A1(n12338), .A2(n12281), .ZN(n15885) );
  NAND2_X1 U13762 ( .A1(n12652), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n12285) );
  OAI21_X1 U13763 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12283), .A(
        n12311), .ZN(n22108) );
  AOI22_X1 U13764 ( .A1(n12657), .A2(n22108), .B1(n12660), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U13765 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U13766 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U13767 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12588), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U13768 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12286) );
  NAND4_X1 U13769 ( .A1(n12289), .A2(n12288), .A3(n12287), .A4(n12286), .ZN(
        n12295) );
  AOI22_X1 U13770 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12635), .B1(
        n12626), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U13771 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U13772 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U13773 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12290) );
  NAND4_X1 U13774 ( .A1(n12293), .A2(n12292), .A3(n12291), .A4(n12290), .ZN(
        n12294) );
  OAI21_X1 U13775 ( .B1(n12295), .B2(n12294), .A(n12338), .ZN(n12299) );
  NAND2_X1 U13776 ( .A1(n12652), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12298) );
  XNOR2_X1 U13777 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12311), .ZN(
        n22117) );
  INV_X1 U13778 ( .A(n22117), .ZN(n12296) );
  AOI22_X1 U13779 ( .A1(n12296), .A2(n12657), .B1(n12660), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12297) );
  NAND3_X1 U13780 ( .A1(n12299), .A2(n12298), .A3(n12297), .ZN(n15937) );
  AOI22_X1 U13781 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U13782 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U13783 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12300) );
  NAND4_X1 U13784 ( .A1(n12303), .A2(n12302), .A3(n12301), .A4(n12300), .ZN(
        n12309) );
  AOI22_X1 U13785 ( .A1(n12062), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U13786 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U13787 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U13788 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12304) );
  NAND4_X1 U13789 ( .A1(n12307), .A2(n12306), .A3(n12305), .A4(n12304), .ZN(
        n12308) );
  OAI21_X1 U13790 ( .B1(n12309), .B2(n12308), .A(n12338), .ZN(n12314) );
  NAND2_X1 U13791 ( .A1(n12652), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12313) );
  INV_X1 U13792 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12310) );
  XNOR2_X1 U13793 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12315), .ZN(
        n16776) );
  AOI22_X1 U13794 ( .A1(n12657), .A2(n16776), .B1(n12660), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12312) );
  NAND3_X1 U13795 ( .A1(n12314), .A2(n12313), .A3(n12312), .ZN(n15936) );
  INV_X1 U13796 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n22123) );
  XOR2_X1 U13797 ( .A(n22123), .B(n12329), .Z(n22126) );
  AOI22_X1 U13798 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U13799 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U13800 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U13801 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12316) );
  NAND4_X1 U13802 ( .A1(n12319), .A2(n12318), .A3(n12317), .A4(n12316), .ZN(
        n12325) );
  AOI22_X1 U13803 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12626), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U13804 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U13805 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U13806 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12320) );
  NAND4_X1 U13807 ( .A1(n12323), .A2(n12322), .A3(n12321), .A4(n12320), .ZN(
        n12324) );
  OR2_X1 U13808 ( .A1(n12325), .A2(n12324), .ZN(n12326) );
  AOI22_X1 U13809 ( .A1(n12338), .A2(n12326), .B1(n12660), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U13810 ( .A1(n12652), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12327) );
  OAI211_X1 U13811 ( .C1(n22126), .C2(n12650), .A(n12328), .B(n12327), .ZN(
        n15879) );
  XNOR2_X1 U13812 ( .A(n12359), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n22131) );
  AOI22_X1 U13813 ( .A1(n12652), .A2(P1_EAX_REG_15__SCAN_IN), .B1(n12660), 
        .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U13814 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U13815 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U13816 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U13817 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12330) );
  NAND4_X1 U13818 ( .A1(n12333), .A2(n12332), .A3(n12331), .A4(n12330), .ZN(
        n12340) );
  AOI22_X1 U13819 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U13820 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U13821 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12334) );
  NAND4_X1 U13822 ( .A1(n12337), .A2(n12336), .A3(n12335), .A4(n12334), .ZN(
        n12339) );
  OAI21_X1 U13823 ( .B1(n12340), .B2(n12339), .A(n12338), .ZN(n12341) );
  OAI211_X1 U13824 ( .C1(n22131), .C2(n12650), .A(n12342), .B(n12341), .ZN(
        n12343) );
  INV_X1 U13825 ( .A(n12343), .ZN(n15951) );
  NOR2_X2 U13826 ( .A1(n15878), .A2(n15951), .ZN(n15950) );
  INV_X1 U13827 ( .A(n14789), .ZN(n16888) );
  NAND2_X1 U13828 ( .A1(n16888), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U13829 ( .A1(n12456), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U13830 ( .A1(n12062), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U13831 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U13832 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12344) );
  NAND4_X1 U13833 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12354) );
  AOI22_X1 U13834 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U13835 ( .A1(n11908), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U13836 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U13837 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12349) );
  NAND4_X1 U13838 ( .A1(n12352), .A2(n12351), .A3(n12350), .A4(n12349), .ZN(
        n12353) );
  NOR2_X1 U13839 ( .A1(n12354), .A2(n12353), .ZN(n12358) );
  NAND2_X1 U13840 ( .A1(n21855), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12355) );
  NAND2_X1 U13841 ( .A1(n12650), .A2(n12355), .ZN(n12356) );
  AOI21_X1 U13842 ( .B1(n12652), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12356), .ZN(
        n12357) );
  OAI21_X1 U13843 ( .B1(n12654), .B2(n12358), .A(n12357), .ZN(n12363) );
  INV_X1 U13844 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16762) );
  OAI21_X1 U13845 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12360), .A(
        n12395), .ZN(n22143) );
  INV_X1 U13846 ( .A(n22143), .ZN(n12361) );
  NAND2_X1 U13847 ( .A1(n12361), .A2(n12657), .ZN(n12362) );
  NAND2_X1 U13848 ( .A1(n12363), .A2(n12362), .ZN(n16658) );
  AND2_X2 U13849 ( .A1(n15950), .A2(n12364), .ZN(n16585) );
  AOI22_X1 U13850 ( .A1(n12637), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U13851 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U13852 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12365) );
  NAND4_X1 U13853 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12374) );
  AOI22_X1 U13854 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12456), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U13855 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U13856 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U13857 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12369) );
  NAND4_X1 U13858 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12373) );
  OR2_X1 U13859 ( .A1(n12374), .A2(n12373), .ZN(n12375) );
  NAND2_X1 U13860 ( .A1(n12619), .A2(n12375), .ZN(n12379) );
  XNOR2_X1 U13861 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12395), .ZN(
        n22155) );
  NAND2_X1 U13862 ( .A1(n12660), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12376) );
  OAI21_X1 U13863 ( .B1(n12650), .B2(n22155), .A(n12376), .ZN(n12377) );
  AOI21_X1 U13864 ( .B1(n12652), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12377), .ZN(
        n12378) );
  NAND2_X1 U13865 ( .A1(n12379), .A2(n12378), .ZN(n16586) );
  AND2_X2 U13866 ( .A1(n16585), .A2(n16586), .ZN(n16584) );
  AOI22_X1 U13867 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U13868 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U13869 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12380), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12381) );
  NAND4_X1 U13870 ( .A1(n12384), .A2(n12383), .A3(n12382), .A4(n12381), .ZN(
        n12390) );
  AOI22_X1 U13871 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U13872 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U13873 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U13874 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12385) );
  NAND4_X1 U13875 ( .A1(n12388), .A2(n12387), .A3(n12386), .A4(n12385), .ZN(
        n12389) );
  NOR2_X1 U13876 ( .A1(n12390), .A2(n12389), .ZN(n12394) );
  NAND2_X1 U13877 ( .A1(n21855), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12391) );
  NAND2_X1 U13878 ( .A1(n12650), .A2(n12391), .ZN(n12392) );
  AOI21_X1 U13879 ( .B1(n12652), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12392), .ZN(
        n12393) );
  OAI21_X1 U13880 ( .B1(n12654), .B2(n12394), .A(n12393), .ZN(n12399) );
  INV_X1 U13881 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n22153) );
  OAI21_X1 U13882 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12396), .A(
        n12432), .ZN(n22168) );
  INV_X1 U13883 ( .A(n22168), .ZN(n12397) );
  NAND2_X1 U13884 ( .A1(n12397), .A2(n12657), .ZN(n12398) );
  AOI22_X1 U13885 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12587), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U13886 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U13887 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12400) );
  NAND4_X1 U13888 ( .A1(n12403), .A2(n12402), .A3(n12401), .A4(n12400), .ZN(
        n12409) );
  AOI22_X1 U13889 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U13890 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U13891 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12062), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12405) );
  AOI22_X1 U13892 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12404) );
  NAND4_X1 U13893 ( .A1(n12407), .A2(n12406), .A3(n12405), .A4(n12404), .ZN(
        n12408) );
  NOR2_X1 U13894 ( .A1(n12409), .A2(n12408), .ZN(n12413) );
  OAI21_X1 U13895 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21856), .A(
        n21855), .ZN(n12410) );
  INV_X1 U13896 ( .A(n12410), .ZN(n12411) );
  AOI21_X1 U13897 ( .B1(n12652), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12411), .ZN(
        n12412) );
  OAI21_X1 U13898 ( .B1(n12654), .B2(n12413), .A(n12412), .ZN(n12417) );
  INV_X1 U13899 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16737) );
  OAI21_X1 U13900 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12414), .A(
        n12467), .ZN(n20543) );
  INV_X1 U13901 ( .A(n20543), .ZN(n12415) );
  NAND2_X1 U13902 ( .A1(n12415), .A2(n12657), .ZN(n12416) );
  NAND2_X1 U13903 ( .A1(n12417), .A2(n12416), .ZN(n16530) );
  AOI22_X1 U13904 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U13905 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U13906 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12419) );
  AOI22_X1 U13907 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12418) );
  NAND4_X1 U13908 ( .A1(n12421), .A2(n12420), .A3(n12419), .A4(n12418), .ZN(
        n12427) );
  AOI22_X1 U13909 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U13910 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U13911 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12422) );
  NAND4_X1 U13912 ( .A1(n12425), .A2(n12424), .A3(n12423), .A4(n12422), .ZN(
        n12426) );
  NOR2_X1 U13913 ( .A1(n12427), .A2(n12426), .ZN(n12431) );
  NOR2_X1 U13914 ( .A1(n16737), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12428) );
  OR2_X1 U13915 ( .A1(n12657), .A2(n12428), .ZN(n12429) );
  AOI21_X1 U13916 ( .B1(n12652), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12429), .ZN(
        n12430) );
  OAI21_X1 U13917 ( .B1(n12654), .B2(n12431), .A(n12430), .ZN(n12434) );
  XNOR2_X1 U13918 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12432), .ZN(
        n16739) );
  NAND2_X1 U13919 ( .A1(n12657), .A2(n16739), .ZN(n12433) );
  NAND2_X1 U13920 ( .A1(n12434), .A2(n12433), .ZN(n16546) );
  AOI22_X1 U13921 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12626), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U13922 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U13923 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U13924 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12436) );
  NAND4_X1 U13925 ( .A1(n12439), .A2(n12438), .A3(n12437), .A4(n12436), .ZN(
        n12445) );
  AOI22_X1 U13926 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U13927 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U13928 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U13929 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12440) );
  NAND4_X1 U13930 ( .A1(n12443), .A2(n12442), .A3(n12441), .A4(n12440), .ZN(
        n12444) );
  NOR2_X1 U13931 ( .A1(n12445), .A2(n12444), .ZN(n12449) );
  INV_X1 U13932 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16730) );
  NOR2_X1 U13933 ( .A1(n16730), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12446) );
  OR2_X1 U13934 ( .A1(n12657), .A2(n12446), .ZN(n12447) );
  AOI21_X1 U13935 ( .B1(n12652), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12447), .ZN(
        n12448) );
  OAI21_X1 U13936 ( .B1(n12654), .B2(n12449), .A(n12448), .ZN(n12451) );
  XNOR2_X1 U13937 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12467), .ZN(
        n22178) );
  NAND2_X1 U13938 ( .A1(n12657), .A2(n22178), .ZN(n12450) );
  AOI22_X1 U13939 ( .A1(n12637), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U13940 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U13941 ( .A1(n12037), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U13942 ( .A1(n12455), .A2(n12454), .A3(n12453), .A4(n12452), .ZN(
        n12462) );
  AOI22_X1 U13943 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12456), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U13944 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U13945 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U13946 ( .A1(n12062), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12457) );
  NAND4_X1 U13947 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(
        n12461) );
  NOR2_X1 U13948 ( .A1(n12462), .A2(n12461), .ZN(n12466) );
  OAI21_X1 U13949 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21856), .A(
        n21855), .ZN(n12463) );
  INV_X1 U13950 ( .A(n12463), .ZN(n12464) );
  AOI21_X1 U13951 ( .B1(n12652), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12464), .ZN(
        n12465) );
  OAI21_X1 U13952 ( .B1(n12654), .B2(n12466), .A(n12465), .ZN(n12471) );
  OAI21_X1 U13953 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12468), .A(
        n12515), .ZN(n20550) );
  INV_X1 U13954 ( .A(n20550), .ZN(n12469) );
  NAND2_X1 U13955 ( .A1(n12469), .A2(n12657), .ZN(n12470) );
  AOI22_X1 U13956 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U13957 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U13958 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U13959 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12472) );
  NAND4_X1 U13960 ( .A1(n12475), .A2(n12474), .A3(n12473), .A4(n12472), .ZN(
        n12481) );
  AOI22_X1 U13961 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U13962 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U13963 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12476) );
  NAND4_X1 U13964 ( .A1(n12479), .A2(n12478), .A3(n12477), .A4(n12476), .ZN(
        n12480) );
  NOR2_X1 U13965 ( .A1(n12481), .A2(n12480), .ZN(n12499) );
  AOI22_X1 U13966 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U13967 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U13968 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12482) );
  NAND4_X1 U13969 ( .A1(n12485), .A2(n12484), .A3(n12483), .A4(n12482), .ZN(
        n12491) );
  AOI22_X1 U13970 ( .A1(n12637), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U13971 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U13972 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U13973 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12037), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12486) );
  NAND4_X1 U13974 ( .A1(n12489), .A2(n12488), .A3(n12487), .A4(n12486), .ZN(
        n12490) );
  NOR2_X1 U13975 ( .A1(n12491), .A2(n12490), .ZN(n12500) );
  XOR2_X1 U13976 ( .A(n12499), .B(n12500), .Z(n12492) );
  NAND2_X1 U13977 ( .A1(n12492), .A2(n12619), .ZN(n12496) );
  INV_X1 U13978 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16719) );
  NOR2_X1 U13979 ( .A1(n16719), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12493) );
  OR2_X1 U13980 ( .A1(n12657), .A2(n12493), .ZN(n12494) );
  AOI21_X1 U13981 ( .B1(n12652), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12494), .ZN(
        n12495) );
  NAND2_X1 U13982 ( .A1(n12496), .A2(n12495), .ZN(n12498) );
  XNOR2_X1 U13983 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12515), .ZN(
        n22188) );
  NAND2_X1 U13984 ( .A1(n12657), .A2(n22188), .ZN(n12497) );
  NAND2_X1 U13985 ( .A1(n12498), .A2(n12497), .ZN(n16569) );
  NOR2_X2 U13986 ( .A1(n16513), .A2(n16569), .ZN(n16570) );
  NOR2_X1 U13987 ( .A1(n12500), .A2(n12499), .ZN(n12533) );
  AOI22_X1 U13988 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U13989 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U13990 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12501) );
  NAND4_X1 U13991 ( .A1(n12504), .A2(n12503), .A3(n12502), .A4(n12501), .ZN(
        n12510) );
  AOI22_X1 U13992 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U13993 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U13994 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U13995 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12505) );
  NAND4_X1 U13996 ( .A1(n12508), .A2(n12507), .A3(n12506), .A4(n12505), .ZN(
        n12509) );
  OR2_X1 U13997 ( .A1(n12510), .A2(n12509), .ZN(n12532) );
  XNOR2_X1 U13998 ( .A(n12533), .B(n12532), .ZN(n12514) );
  NAND2_X1 U13999 ( .A1(n21855), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12511) );
  NAND2_X1 U14000 ( .A1(n12650), .A2(n12511), .ZN(n12512) );
  AOI21_X1 U14001 ( .B1(n12652), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12512), .ZN(
        n12513) );
  OAI21_X1 U14002 ( .B1(n12514), .B2(n12654), .A(n12513), .ZN(n12519) );
  OAI21_X1 U14003 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12516), .A(
        n12554), .ZN(n22204) );
  INV_X1 U14004 ( .A(n22204), .ZN(n12517) );
  NAND2_X1 U14005 ( .A1(n12517), .A2(n12657), .ZN(n12518) );
  NAND2_X1 U14006 ( .A1(n12519), .A2(n12518), .ZN(n16616) );
  INV_X1 U14007 ( .A(n16616), .ZN(n12520) );
  AND2_X2 U14008 ( .A1(n16570), .A2(n12520), .ZN(n16499) );
  AOI22_X1 U14009 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U14010 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12062), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U14011 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12522) );
  AOI22_X1 U14012 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12521) );
  NAND4_X1 U14013 ( .A1(n12524), .A2(n12523), .A3(n12522), .A4(n12521), .ZN(
        n12531) );
  AOI22_X1 U14014 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U14015 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U14016 ( .A1(n12637), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U14017 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12526) );
  NAND4_X1 U14018 ( .A1(n12529), .A2(n12528), .A3(n12527), .A4(n12526), .ZN(
        n12530) );
  NOR2_X1 U14019 ( .A1(n12531), .A2(n12530), .ZN(n12540) );
  NAND2_X1 U14020 ( .A1(n12533), .A2(n12532), .ZN(n12539) );
  XOR2_X1 U14021 ( .A(n12540), .B(n12539), .Z(n12534) );
  NAND2_X1 U14022 ( .A1(n12534), .A2(n12619), .ZN(n12538) );
  INV_X1 U14023 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16711) );
  AOI21_X1 U14024 ( .B1(n16711), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12535) );
  AOI21_X1 U14025 ( .B1(n12652), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12535), .ZN(
        n12537) );
  XNOR2_X1 U14026 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n12554), .ZN(
        n16715) );
  AOI21_X1 U14027 ( .B1(n12538), .B2(n12537), .A(n12536), .ZN(n16501) );
  AND2_X2 U14028 ( .A1(n16499), .A2(n16501), .ZN(n16485) );
  NOR2_X1 U14029 ( .A1(n12540), .A2(n12539), .ZN(n12572) );
  AOI22_X1 U14030 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U14031 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U14032 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12541) );
  NAND4_X1 U14033 ( .A1(n12544), .A2(n12543), .A3(n12542), .A4(n12541), .ZN(
        n12550) );
  AOI22_X1 U14034 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U14035 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U14036 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U14037 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12545) );
  NAND4_X1 U14038 ( .A1(n12548), .A2(n12547), .A3(n12546), .A4(n12545), .ZN(
        n12549) );
  OR2_X1 U14039 ( .A1(n12550), .A2(n12549), .ZN(n12571) );
  INV_X1 U14040 ( .A(n12571), .ZN(n12551) );
  XNOR2_X1 U14041 ( .A(n12572), .B(n12551), .ZN(n12552) );
  NAND2_X1 U14042 ( .A1(n12552), .A2(n12619), .ZN(n12559) );
  INV_X1 U14043 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16492) );
  AOI21_X1 U14044 ( .B1(n16492), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12553) );
  AOI21_X1 U14045 ( .B1(n12652), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12553), .ZN(
        n12558) );
  INV_X1 U14046 ( .A(n12554), .ZN(n12555) );
  OAI21_X1 U14047 ( .B1(n12556), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n12599), .ZN(n16704) );
  NOR2_X1 U14048 ( .A1(n16704), .A2(n12650), .ZN(n12557) );
  AOI21_X1 U14049 ( .B1(n12559), .B2(n12558), .A(n12557), .ZN(n16487) );
  NAND2_X1 U14050 ( .A1(n16485), .A2(n16487), .ZN(n16473) );
  AOI22_X1 U14051 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12610), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U14052 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12588), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U14053 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12561) );
  NAND4_X1 U14054 ( .A1(n12564), .A2(n12563), .A3(n12562), .A4(n12561), .ZN(
        n12570) );
  AOI22_X1 U14055 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U14056 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U14057 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12627), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U14058 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12565) );
  NAND4_X1 U14059 ( .A1(n12568), .A2(n12567), .A3(n12566), .A4(n12565), .ZN(
        n12569) );
  NOR2_X1 U14060 ( .A1(n12570), .A2(n12569), .ZN(n12580) );
  NAND2_X1 U14061 ( .A1(n12572), .A2(n12571), .ZN(n12579) );
  XOR2_X1 U14062 ( .A(n12580), .B(n12579), .Z(n12575) );
  INV_X1 U14063 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16698) );
  NAND2_X1 U14064 ( .A1(n12180), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12573) );
  OAI211_X1 U14065 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n16698), .A(n12573), 
        .B(n12650), .ZN(n12574) );
  AOI21_X1 U14066 ( .B1(n12575), .B2(n12619), .A(n12574), .ZN(n12576) );
  INV_X1 U14067 ( .A(n12576), .ZN(n12578) );
  XNOR2_X1 U14068 ( .A(n12599), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16696) );
  NAND2_X1 U14069 ( .A1(n16696), .A2(n12657), .ZN(n12577) );
  NAND2_X1 U14070 ( .A1(n12578), .A2(n12577), .ZN(n16474) );
  NOR2_X1 U14071 ( .A1(n12580), .A2(n12579), .ZN(n12618) );
  AOI22_X1 U14072 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U14073 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U14074 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11913), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U14075 ( .A1(n12637), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12583) );
  NAND4_X1 U14076 ( .A1(n12586), .A2(n12585), .A3(n12584), .A4(n12583), .ZN(
        n12594) );
  AOI22_X1 U14077 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U14078 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U14079 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U14080 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12589) );
  NAND4_X1 U14081 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n12593) );
  OR2_X1 U14082 ( .A1(n12594), .A2(n12593), .ZN(n12617) );
  INV_X1 U14083 ( .A(n12617), .ZN(n12595) );
  XNOR2_X1 U14084 ( .A(n12618), .B(n12595), .ZN(n12598) );
  INV_X1 U14085 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16466) );
  NAND2_X1 U14086 ( .A1(n12180), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n12596) );
  OAI211_X1 U14087 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n16466), .A(n12596), 
        .B(n12650), .ZN(n12597) );
  AOI21_X1 U14088 ( .B1(n12598), .B2(n12619), .A(n12597), .ZN(n12603) );
  NOR2_X1 U14089 ( .A1(n12600), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12601) );
  OR2_X1 U14090 ( .A1(n12656), .A2(n12601), .ZN(n16689) );
  NOR2_X1 U14091 ( .A1(n16689), .A2(n12650), .ZN(n12602) );
  INV_X1 U14092 ( .A(n16462), .ZN(n12604) );
  AOI22_X1 U14093 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12637), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U14094 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12588), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U14095 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U14096 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12606) );
  NAND4_X1 U14097 ( .A1(n12609), .A2(n12608), .A3(n12607), .A4(n12606), .ZN(
        n12616) );
  AOI22_X1 U14098 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U14099 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U14100 ( .A1(n12037), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12611) );
  NAND4_X1 U14101 ( .A1(n12614), .A2(n12613), .A3(n12612), .A4(n12611), .ZN(
        n12615) );
  NOR2_X1 U14102 ( .A1(n12616), .A2(n12615), .ZN(n12646) );
  NAND2_X1 U14103 ( .A1(n12618), .A2(n12617), .ZN(n12645) );
  XOR2_X1 U14104 ( .A(n12646), .B(n12645), .Z(n12620) );
  NAND2_X1 U14105 ( .A1(n12620), .A2(n12619), .ZN(n12625) );
  NAND2_X1 U14106 ( .A1(n21855), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12621) );
  NAND2_X1 U14107 ( .A1(n12650), .A2(n12621), .ZN(n12622) );
  AOI21_X1 U14108 ( .B1(n12652), .B2(P1_EAX_REG_29__SCAN_IN), .A(n12622), .ZN(
        n12624) );
  INV_X1 U14109 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13653) );
  XNOR2_X1 U14110 ( .A(n12656), .B(n13653), .ZN(n16453) );
  AND2_X1 U14111 ( .A1(n16453), .A2(n17711), .ZN(n12623) );
  AOI21_X1 U14112 ( .B1(n12625), .B2(n12624), .A(n12623), .ZN(n13650) );
  AOI22_X1 U14113 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12626), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U14114 ( .A1(n12628), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U14115 ( .A1(n12587), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12629), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U14116 ( .A1(n12588), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12630), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12631) );
  NAND4_X1 U14117 ( .A1(n12634), .A2(n12633), .A3(n12632), .A4(n12631), .ZN(
        n12644) );
  AOI22_X1 U14118 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U14119 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12641) );
  AOI22_X1 U14120 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U14121 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12638), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12639) );
  NAND4_X1 U14122 ( .A1(n12642), .A2(n12641), .A3(n12640), .A4(n12639), .ZN(
        n12643) );
  NOR2_X1 U14123 ( .A1(n12644), .A2(n12643), .ZN(n12648) );
  NOR2_X1 U14124 ( .A1(n12646), .A2(n12645), .ZN(n12647) );
  XOR2_X1 U14125 ( .A(n12648), .B(n12647), .Z(n12655) );
  NAND2_X1 U14126 ( .A1(n21855), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12649) );
  NAND2_X1 U14127 ( .A1(n12650), .A2(n12649), .ZN(n12651) );
  AOI21_X1 U14128 ( .B1(n12652), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12651), .ZN(
        n12653) );
  OAI21_X1 U14129 ( .B1(n12655), .B2(n12654), .A(n12653), .ZN(n12659) );
  INV_X1 U14130 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16676) );
  XNOR2_X1 U14131 ( .A(n12727), .B(n16676), .ZN(n16674) );
  NAND2_X1 U14132 ( .A1(n16674), .A2(n12657), .ZN(n12658) );
  NAND2_X1 U14133 ( .A1(n12659), .A2(n12658), .ZN(n16433) );
  AOI22_X1 U14134 ( .A1(n12180), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12660), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12661) );
  INV_X1 U14135 ( .A(n16590), .ZN(n12730) );
  NAND2_X1 U14136 ( .A1(n22485), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12700) );
  XNOR2_X1 U14137 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12677) );
  NAND2_X1 U14138 ( .A1(n12679), .A2(n12677), .ZN(n12664) );
  NAND2_X1 U14139 ( .A1(n15451), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12663) );
  NAND2_X1 U14140 ( .A1(n12664), .A2(n12663), .ZN(n12676) );
  MUX2_X1 U14141 ( .A(n12665), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12674) );
  NAND2_X1 U14142 ( .A1(n12676), .A2(n12674), .ZN(n12667) );
  NAND2_X1 U14143 ( .A1(n12665), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12666) );
  NAND2_X1 U14144 ( .A1(n12667), .A2(n12666), .ZN(n12673) );
  MUX2_X1 U14145 ( .A(n12668), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12671) );
  NAND2_X1 U14146 ( .A1(n12673), .A2(n12671), .ZN(n12670) );
  NAND2_X1 U14147 ( .A1(n12668), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12669) );
  NAND2_X1 U14148 ( .A1(n12670), .A2(n12669), .ZN(n12682) );
  NAND2_X1 U14149 ( .A1(n17673), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12683) );
  OR2_X1 U14150 ( .A1(n12682), .A2(n12683), .ZN(n12687) );
  INV_X1 U14151 ( .A(n12671), .ZN(n12672) );
  XNOR2_X1 U14152 ( .A(n12673), .B(n12672), .ZN(n12718) );
  INV_X1 U14153 ( .A(n12674), .ZN(n12675) );
  XNOR2_X1 U14154 ( .A(n12676), .B(n12675), .ZN(n12693) );
  INV_X1 U14155 ( .A(n12677), .ZN(n12678) );
  XNOR2_X1 U14156 ( .A(n12679), .B(n12678), .ZN(n12703) );
  AND2_X1 U14157 ( .A1(n12693), .A2(n12703), .ZN(n12680) );
  NAND2_X1 U14158 ( .A1(n12721), .A2(n12680), .ZN(n12685) );
  INV_X1 U14159 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17748) );
  AND2_X1 U14160 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17748), .ZN(
        n12681) );
  NAND2_X1 U14161 ( .A1(n12685), .A2(n12686), .ZN(n16419) );
  NAND2_X1 U14162 ( .A1(n16595), .A2(n14764), .ZN(n12906) );
  NAND2_X1 U14163 ( .A1(n12720), .A2(n14533), .ZN(n12704) );
  INV_X1 U14164 ( .A(n12687), .ZN(n12692) );
  NAND2_X1 U14165 ( .A1(n15592), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12694) );
  NAND3_X1 U14166 ( .A1(n12705), .A2(n12694), .A3(n14764), .ZN(n12698) );
  INV_X1 U14167 ( .A(n12698), .ZN(n12691) );
  INV_X1 U14168 ( .A(n12693), .ZN(n12688) );
  AND2_X1 U14169 ( .A1(n15391), .A2(n16595), .ZN(n12689) );
  INV_X1 U14170 ( .A(n12711), .ZN(n12690) );
  AOI22_X1 U14171 ( .A1(n12692), .A2(n12691), .B1(n12715), .B2(n12690), .ZN(
        n12717) );
  OAI21_X1 U14172 ( .B1(n12693), .B2(n12695), .A(n12711), .ZN(n12714) );
  INV_X1 U14173 ( .A(n12703), .ZN(n12699) );
  AOI21_X1 U14174 ( .B1(n12696), .B2(n14764), .A(n12702), .ZN(n12697) );
  AOI21_X1 U14175 ( .B1(n12699), .B2(n12698), .A(n12697), .ZN(n12713) );
  INV_X1 U14176 ( .A(n14559), .ZN(n12701) );
  OAI21_X1 U14177 ( .B1(n22485), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12700), .ZN(n12706) );
  OAI21_X1 U14178 ( .B1(n12701), .B2(n12706), .A(n11177), .ZN(n12710) );
  NOR3_X1 U14179 ( .A1(n14764), .A2(n12703), .A3(n12702), .ZN(n12709) );
  OAI21_X1 U14180 ( .B1(n12706), .B2(n12705), .A(n12704), .ZN(n12707) );
  INV_X1 U14181 ( .A(n12707), .ZN(n12708) );
  AOI211_X1 U14182 ( .C1(n12711), .C2(n12710), .A(n12709), .B(n12708), .ZN(
        n12712) );
  OAI22_X1 U14183 ( .A1(n12715), .A2(n12714), .B1(n12713), .B2(n12712), .ZN(
        n12716) );
  OAI211_X1 U14184 ( .C1(n12718), .C2(n12906), .A(n12717), .B(n12716), .ZN(
        n12719) );
  OAI21_X1 U14185 ( .B1(n12721), .B2(n12720), .A(n12719), .ZN(n12722) );
  OAI22_X1 U14186 ( .A1(n15103), .A2(n16419), .B1(n16422), .B2(n14762), .ZN(
        n14770) );
  NAND2_X1 U14187 ( .A1(n22810), .A2(n14764), .ZN(n16890) );
  NAND2_X1 U14188 ( .A1(n17718), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22234) );
  INV_X1 U14189 ( .A(n22234), .ZN(n22809) );
  NAND2_X1 U14190 ( .A1(n17744), .A2(n21855), .ZN(n21858) );
  INV_X1 U14191 ( .A(n21858), .ZN(n22229) );
  NAND2_X1 U14192 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22229), .ZN(n17743) );
  NAND2_X1 U14193 ( .A1(n21855), .A2(n22225), .ZN(n12725) );
  NAND2_X1 U14194 ( .A1(n21856), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12946) );
  AND3_X1 U14195 ( .A1(n17669), .A2(n12946), .A3(n22225), .ZN(n12724) );
  AOI21_X1 U14196 ( .B1(n17743), .B2(n12725), .A(n12724), .ZN(n12726) );
  NAND2_X1 U14197 ( .A1(n12727), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12728) );
  XNOR2_X1 U14198 ( .A(n12728), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14073) );
  NAND2_X1 U14199 ( .A1(n12730), .A2(n22172), .ZN(n12841) );
  INV_X1 U14200 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n22191) );
  INV_X1 U14201 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n16533) );
  INV_X1 U14202 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n16548) );
  INV_X1 U14203 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n16547) );
  INV_X1 U14204 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21908) );
  INV_X1 U14205 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n22139) );
  NOR4_X1 U14206 ( .A1(n16548), .A2(n16547), .A3(n21908), .A4(n22139), .ZN(
        n12731) );
  NAND3_X1 U14207 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(n12731), .ZN(n16535) );
  NOR2_X1 U14208 ( .A1(n16533), .A2(n16535), .ZN(n16515) );
  NAND3_X1 U14209 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .ZN(n16516) );
  INV_X1 U14210 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n22082) );
  INV_X1 U14211 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n22055) );
  INV_X1 U14212 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n22259) );
  AND2_X1 U14213 ( .A1(n12732), .A2(n22259), .ZN(n22261) );
  INV_X1 U14214 ( .A(n22261), .ZN(n17713) );
  NAND2_X1 U14215 ( .A1(n15391), .A2(n17713), .ZN(n14541) );
  NAND2_X1 U14216 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n22253) );
  NAND2_X1 U14217 ( .A1(n22253), .A2(n21856), .ZN(n17714) );
  INV_X1 U14218 ( .A(n17714), .ZN(n12733) );
  NAND2_X1 U14219 ( .A1(n14541), .A2(n12733), .ZN(n12832) );
  NAND4_X1 U14220 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(n22034), .ZN(n22056) );
  NAND2_X1 U14221 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22072), .ZN(n22083) );
  INV_X1 U14222 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15485) );
  INV_X1 U14223 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15578) );
  INV_X1 U14224 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n16881) );
  INV_X1 U14225 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n22094) );
  NOR4_X1 U14226 ( .A1(n15485), .A2(n15578), .A3(n16881), .A4(n22094), .ZN(
        n14068) );
  NAND2_X1 U14227 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n12734) );
  NAND2_X1 U14228 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n12735) );
  NAND2_X1 U14229 ( .A1(n16455), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n12836) );
  NAND2_X1 U14230 ( .A1(n12836), .A2(n22200), .ZN(n16434) );
  INV_X1 U14231 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n13752) );
  INV_X1 U14232 ( .A(n12842), .ZN(n15383) );
  NAND2_X1 U14233 ( .A1(n12786), .A2(n12820), .ZN(n15301) );
  OR2_X1 U14234 ( .A1(n15301), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12737) );
  INV_X1 U14235 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n16559) );
  NAND2_X1 U14236 ( .A1(n15304), .A2(n16559), .ZN(n12736) );
  NAND2_X1 U14237 ( .A1(n12737), .A2(n12736), .ZN(n16440) );
  NAND2_X1 U14238 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12738) );
  OAI211_X1 U14239 ( .C1(n12752), .C2(P1_EBX_REG_1__SCAN_IN), .A(n12786), .B(
        n12738), .ZN(n12739) );
  MUX2_X1 U14240 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_0__SCAN_IN), .Z(
        n15303) );
  INV_X1 U14241 ( .A(n15303), .ZN(n12740) );
  OR2_X1 U14242 ( .A1(n12819), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U14243 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12742) );
  OAI211_X1 U14244 ( .C1(n12752), .C2(P1_EBX_REG_2__SCAN_IN), .A(n12786), .B(
        n12742), .ZN(n12743) );
  INV_X1 U14245 ( .A(n12745), .ZN(n16435) );
  MUX2_X1 U14246 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12748) );
  NAND2_X1 U14247 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12752), .ZN(
        n12746) );
  AND2_X1 U14248 ( .A1(n12794), .A2(n12746), .ZN(n12747) );
  NAND2_X1 U14249 ( .A1(n12748), .A2(n12747), .ZN(n12749) );
  MUX2_X1 U14250 ( .A(n12819), .B(n12820), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12751) );
  OAI21_X1 U14251 ( .B1(n15301), .B2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n12751), .ZN(n15358) );
  MUX2_X1 U14252 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12755) );
  NAND2_X1 U14253 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12752), .ZN(
        n12753) );
  AND2_X1 U14254 ( .A1(n12794), .A2(n12753), .ZN(n12754) );
  NAND2_X1 U14255 ( .A1(n12755), .A2(n12754), .ZN(n15479) );
  MUX2_X1 U14256 ( .A(n12819), .B(n12820), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12756) );
  OAI21_X1 U14257 ( .B1(n15301), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n12756), .ZN(n15356) );
  MUX2_X1 U14258 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n12759) );
  NAND2_X1 U14259 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n12752), .ZN(
        n12757) );
  AND2_X1 U14260 ( .A1(n12794), .A2(n12757), .ZN(n12758) );
  OR2_X1 U14261 ( .A1(n12819), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n12762) );
  NAND2_X1 U14262 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12760) );
  OAI211_X1 U14263 ( .C1(n12752), .C2(P1_EBX_REG_8__SCAN_IN), .A(n12786), .B(
        n12760), .ZN(n12761) );
  NAND2_X1 U14264 ( .A1(n12762), .A2(n12761), .ZN(n15487) );
  MUX2_X1 U14265 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12765) );
  NAND2_X1 U14266 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n12752), .ZN(
        n12763) );
  AND2_X1 U14267 ( .A1(n12794), .A2(n12763), .ZN(n12764) );
  NAND2_X1 U14268 ( .A1(n12765), .A2(n12764), .ZN(n15579) );
  OR2_X1 U14269 ( .A1(n12819), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n12768) );
  NAND2_X1 U14270 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12766) );
  OAI211_X1 U14271 ( .C1(n12752), .C2(P1_EBX_REG_10__SCAN_IN), .A(n12786), .B(
        n12766), .ZN(n12767) );
  NAND2_X1 U14272 ( .A1(n12768), .A2(n12767), .ZN(n14070) );
  MUX2_X1 U14273 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12771) );
  NAND2_X1 U14274 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n12752), .ZN(
        n12769) );
  AND2_X1 U14275 ( .A1(n12794), .A2(n12769), .ZN(n12770) );
  OR2_X1 U14276 ( .A1(n15301), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12773) );
  MUX2_X1 U14277 ( .A(n12819), .B(n12820), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12772) );
  AND2_X1 U14278 ( .A1(n12773), .A2(n12772), .ZN(n15920) );
  MUX2_X1 U14279 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12776) );
  NAND2_X1 U14280 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12752), .ZN(
        n12774) );
  AND2_X1 U14281 ( .A1(n12794), .A2(n12774), .ZN(n12775) );
  AND2_X1 U14282 ( .A1(n12776), .A2(n12775), .ZN(n15941) );
  OR2_X1 U14283 ( .A1(n12819), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U14284 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12777) );
  OAI211_X1 U14285 ( .C1(n12752), .C2(P1_EBX_REG_14__SCAN_IN), .A(n12786), .B(
        n12777), .ZN(n12778) );
  NAND2_X1 U14286 ( .A1(n12779), .A2(n12778), .ZN(n16848) );
  INV_X1 U14287 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21901) );
  NAND2_X1 U14288 ( .A1(n12786), .A2(n21901), .ZN(n12780) );
  OAI211_X1 U14289 ( .C1(n12752), .C2(P1_EBX_REG_15__SCAN_IN), .A(n12780), .B(
        n12820), .ZN(n12781) );
  OAI21_X1 U14290 ( .B1(n12820), .B2(P1_EBX_REG_15__SCAN_IN), .A(n12781), .ZN(
        n12782) );
  INV_X1 U14291 ( .A(n12782), .ZN(n15970) );
  OR2_X1 U14292 ( .A1(n12819), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n12785) );
  NAND2_X1 U14293 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12783) );
  OAI211_X1 U14294 ( .C1(n12752), .C2(P1_EBX_REG_16__SCAN_IN), .A(n12786), .B(
        n12783), .ZN(n12784) );
  AND2_X1 U14295 ( .A1(n12785), .A2(n12784), .ZN(n20466) );
  MUX2_X1 U14296 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12789) );
  NAND2_X1 U14297 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n12752), .ZN(
        n12787) );
  AND2_X1 U14298 ( .A1(n12794), .A2(n12787), .ZN(n12788) );
  AND2_X1 U14299 ( .A1(n12789), .A2(n12788), .ZN(n16581) );
  OR2_X1 U14300 ( .A1(n12819), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U14301 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12790) );
  OAI211_X1 U14302 ( .C1(n12752), .C2(P1_EBX_REG_18__SCAN_IN), .A(n12786), .B(
        n12790), .ZN(n12791) );
  NAND2_X1 U14303 ( .A1(n12792), .A2(n12791), .ZN(n14578) );
  MUX2_X1 U14304 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12796) );
  NAND2_X1 U14305 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n12752), .ZN(
        n12793) );
  AND2_X1 U14306 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  NAND2_X1 U14307 ( .A1(n12796), .A2(n12795), .ZN(n16549) );
  OR2_X1 U14308 ( .A1(n12819), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U14309 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12797) );
  OAI211_X1 U14310 ( .C1(n12752), .C2(P1_EBX_REG_20__SCAN_IN), .A(n12786), .B(
        n12797), .ZN(n12798) );
  NAND2_X1 U14311 ( .A1(n12799), .A2(n12798), .ZN(n16537) );
  INV_X1 U14312 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12800) );
  NAND2_X1 U14313 ( .A1(n12786), .A2(n12800), .ZN(n12801) );
  OAI211_X1 U14314 ( .C1(n12752), .C2(P1_EBX_REG_21__SCAN_IN), .A(n12801), .B(
        n12820), .ZN(n12802) );
  OAI21_X1 U14315 ( .B1(n12820), .B2(P1_EBX_REG_21__SCAN_IN), .A(n12802), .ZN(
        n12803) );
  INV_X1 U14316 ( .A(n12803), .ZN(n16574) );
  OR2_X1 U14317 ( .A1(n12819), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n12806) );
  NAND2_X1 U14318 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12804) );
  OAI211_X1 U14319 ( .C1(n12752), .C2(P1_EBX_REG_22__SCAN_IN), .A(n12786), .B(
        n12804), .ZN(n12805) );
  AND2_X1 U14320 ( .A1(n12806), .A2(n12805), .ZN(n16518) );
  MUX2_X1 U14321 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12808) );
  NAND2_X1 U14322 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n12752), .ZN(
        n12807) );
  NAND2_X1 U14323 ( .A1(n12808), .A2(n12807), .ZN(n16566) );
  OR2_X1 U14324 ( .A1(n12819), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n12811) );
  NAND2_X1 U14325 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12809) );
  OAI211_X1 U14326 ( .C1(n12752), .C2(P1_EBX_REG_24__SCAN_IN), .A(n12786), .B(
        n12809), .ZN(n12810) );
  NAND2_X1 U14327 ( .A1(n12811), .A2(n12810), .ZN(n20476) );
  MUX2_X1 U14328 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12813) );
  NAND2_X1 U14329 ( .A1(n12752), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12812) );
  AND2_X1 U14330 ( .A1(n12813), .A2(n12812), .ZN(n16503) );
  OR2_X1 U14331 ( .A1(n12819), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n12816) );
  NAND2_X1 U14332 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12814) );
  OAI211_X1 U14333 ( .C1(n12752), .C2(P1_EBX_REG_26__SCAN_IN), .A(n12786), .B(
        n12814), .ZN(n12815) );
  NAND2_X1 U14334 ( .A1(n12816), .A2(n12815), .ZN(n16489) );
  MUX2_X1 U14335 ( .A(n12820), .B(n12786), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12818) );
  NAND2_X1 U14336 ( .A1(n12752), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12817) );
  NAND2_X1 U14337 ( .A1(n12818), .A2(n12817), .ZN(n16476) );
  OR2_X1 U14338 ( .A1(n12819), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n12823) );
  NAND2_X1 U14339 ( .A1(n12820), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12821) );
  OAI211_X1 U14340 ( .C1(n12752), .C2(P1_EBX_REG_28__SCAN_IN), .A(n12786), .B(
        n12821), .ZN(n12822) );
  AND2_X1 U14341 ( .A1(n12823), .A2(n12822), .ZN(n16463) );
  OR2_X1 U14342 ( .A1(n15301), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12825) );
  INV_X1 U14343 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n16561) );
  NAND2_X1 U14344 ( .A1(n15304), .A2(n16561), .ZN(n12824) );
  NAND2_X1 U14345 ( .A1(n12825), .A2(n12824), .ZN(n16436) );
  OAI22_X1 U14346 ( .A1(n16436), .A2(n16435), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12820), .ZN(n16452) );
  NOR2_X1 U14347 ( .A1(n16451), .A2(n16440), .ZN(n12829) );
  OR2_X1 U14348 ( .A1(n15301), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12827) );
  INV_X1 U14349 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16557) );
  NAND2_X1 U14350 ( .A1(n15304), .A2(n16557), .ZN(n12826) );
  NAND2_X1 U14351 ( .A1(n12827), .A2(n12826), .ZN(n12828) );
  NOR2_X1 U14352 ( .A1(n12752), .A2(n16557), .ZN(n12833) );
  NAND2_X1 U14353 ( .A1(n12833), .A2(n17714), .ZN(n12831) );
  NAND2_X1 U14354 ( .A1(n12832), .A2(n15127), .ZN(n12834) );
  OR2_X1 U14355 ( .A1(n12834), .A2(n12833), .ZN(n12835) );
  NOR2_X2 U14356 ( .A1(n15410), .A2(n12835), .ZN(n22166) );
  INV_X1 U14357 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12948) );
  OAI22_X1 U14358 ( .A1(n22201), .A2(n16557), .B1(n22152), .B2(n12948), .ZN(
        n12838) );
  NOR2_X1 U14359 ( .A1(n12836), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n12837) );
  AOI211_X1 U14360 ( .C1(n16804), .C2(n22165), .A(n12838), .B(n12837), .ZN(
        n12839) );
  NAND3_X1 U14361 ( .A1(n12841), .A2(n12840), .A3(n12839), .ZN(P1_U2809) );
  INV_X1 U14362 ( .A(n12856), .ZN(n12843) );
  AND2_X1 U14363 ( .A1(n22414), .A2(n12842), .ZN(n12859) );
  AOI21_X1 U14364 ( .B1(n12843), .B2(n21857), .A(n12859), .ZN(n12844) );
  NAND2_X1 U14365 ( .A1(n14801), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14803) );
  INV_X1 U14366 ( .A(n21857), .ZN(n12850) );
  XNOR2_X1 U14367 ( .A(n12856), .B(n12855), .ZN(n12849) );
  INV_X1 U14368 ( .A(n12845), .ZN(n12846) );
  NAND2_X1 U14369 ( .A1(n12846), .A2(n14764), .ZN(n12848) );
  NOR2_X1 U14370 ( .A1(n14554), .A2(n15592), .ZN(n12847) );
  NAND2_X1 U14371 ( .A1(n14838), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12853) );
  OR2_X1 U14372 ( .A1(n14803), .A2(n12851), .ZN(n12852) );
  NAND2_X1 U14373 ( .A1(n12853), .A2(n12852), .ZN(n12863) );
  INV_X1 U14374 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15361) );
  XNOR2_X1 U14375 ( .A(n12863), .B(n15361), .ZN(n14866) );
  NAND2_X1 U14376 ( .A1(n15172), .A2(n14533), .ZN(n12862) );
  NAND2_X1 U14377 ( .A1(n12856), .A2(n12855), .ZN(n12857) );
  NAND2_X1 U14378 ( .A1(n12857), .A2(n12858), .ZN(n12867) );
  OAI21_X1 U14379 ( .B1(n12858), .B2(n12857), .A(n12867), .ZN(n12860) );
  AOI21_X1 U14380 ( .B1(n12860), .B2(n21857), .A(n12859), .ZN(n12861) );
  NAND2_X1 U14381 ( .A1(n12862), .A2(n12861), .ZN(n14867) );
  NAND2_X1 U14382 ( .A1(n14866), .A2(n14867), .ZN(n12865) );
  NAND2_X1 U14383 ( .A1(n12863), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12864) );
  NAND2_X1 U14384 ( .A1(n12865), .A2(n12864), .ZN(n12870) );
  INV_X1 U14385 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12866) );
  XNOR2_X1 U14386 ( .A(n12870), .B(n12866), .ZN(n14954) );
  NAND2_X1 U14387 ( .A1(n12867), .A2(n12868), .ZN(n12883) );
  OAI211_X1 U14388 ( .C1(n12868), .C2(n12867), .A(n12883), .B(n21857), .ZN(
        n12869) );
  OAI21_X1 U14389 ( .B1(n15285), .B2(n12906), .A(n12869), .ZN(n14955) );
  NAND2_X1 U14390 ( .A1(n14954), .A2(n14955), .ZN(n12872) );
  NAND2_X1 U14391 ( .A1(n12870), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12871) );
  NAND2_X1 U14392 ( .A1(n12872), .A2(n12871), .ZN(n15161) );
  OR2_X1 U14393 ( .A1(n12873), .A2(n12906), .ZN(n12876) );
  XNOR2_X1 U14394 ( .A(n12883), .B(n12881), .ZN(n12874) );
  NAND2_X1 U14395 ( .A1(n12874), .A2(n21857), .ZN(n12875) );
  NAND2_X1 U14396 ( .A1(n12876), .A2(n12875), .ZN(n12878) );
  INV_X1 U14397 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12877) );
  XNOR2_X1 U14398 ( .A(n12878), .B(n12877), .ZN(n15160) );
  NAND2_X1 U14399 ( .A1(n12878), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12879) );
  NAND2_X1 U14400 ( .A1(n12880), .A2(n14533), .ZN(n12887) );
  INV_X1 U14401 ( .A(n12881), .ZN(n12882) );
  NOR2_X1 U14402 ( .A1(n12883), .A2(n12882), .ZN(n12885) );
  NAND2_X1 U14403 ( .A1(n12885), .A2(n12884), .ZN(n12899) );
  OAI211_X1 U14404 ( .C1(n12885), .C2(n12884), .A(n12899), .B(n21857), .ZN(
        n12886) );
  NAND2_X1 U14405 ( .A1(n12887), .A2(n12886), .ZN(n12889) );
  INV_X1 U14406 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12888) );
  XNOR2_X1 U14407 ( .A(n12889), .B(n12888), .ZN(n15515) );
  NAND3_X1 U14408 ( .A1(n12890), .A2(n12891), .A3(n14533), .ZN(n12894) );
  XNOR2_X1 U14409 ( .A(n12899), .B(n12900), .ZN(n12892) );
  NAND2_X1 U14410 ( .A1(n12892), .A2(n21857), .ZN(n12893) );
  NAND2_X1 U14411 ( .A1(n12894), .A2(n12893), .ZN(n12896) );
  INV_X1 U14412 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12895) );
  XNOR2_X1 U14413 ( .A(n12896), .B(n12895), .ZN(n15605) );
  NAND2_X1 U14414 ( .A1(n12896), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12897) );
  NAND2_X1 U14415 ( .A1(n12898), .A2(n14533), .ZN(n12904) );
  INV_X1 U14416 ( .A(n12899), .ZN(n12901) );
  NAND2_X1 U14417 ( .A1(n12901), .A2(n12900), .ZN(n12911) );
  XNOR2_X1 U14418 ( .A(n12911), .B(n12909), .ZN(n12902) );
  NAND2_X1 U14419 ( .A1(n12902), .A2(n21857), .ZN(n12903) );
  NAND2_X1 U14420 ( .A1(n12904), .A2(n12903), .ZN(n12905) );
  XNOR2_X1 U14421 ( .A(n12905), .B(n15719), .ZN(n15716) );
  NOR2_X1 U14422 ( .A1(n12907), .A2(n12906), .ZN(n12908) );
  NAND2_X1 U14423 ( .A1(n21857), .A2(n12909), .ZN(n12910) );
  OR2_X1 U14424 ( .A1(n12911), .A2(n12910), .ZN(n12912) );
  NAND2_X1 U14425 ( .A1(n20552), .A2(n12912), .ZN(n12913) );
  XNOR2_X1 U14426 ( .A(n12913), .B(n15709), .ZN(n15695) );
  NAND2_X1 U14427 ( .A1(n12913), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12914) );
  NAND2_X1 U14428 ( .A1(n11861), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12915) );
  XNOR2_X1 U14429 ( .A(n20552), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16773) );
  INV_X1 U14430 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21889) );
  NAND2_X1 U14431 ( .A1(n20552), .A2(n21889), .ZN(n16772) );
  NAND2_X1 U14432 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12916) );
  NAND2_X1 U14433 ( .A1(n20552), .A2(n12916), .ZN(n16770) );
  AND2_X1 U14434 ( .A1(n16772), .A2(n16770), .ZN(n12917) );
  NAND2_X1 U14435 ( .A1(n16773), .A2(n12917), .ZN(n16837) );
  INV_X1 U14436 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16758) );
  NOR2_X1 U14437 ( .A1(n16837), .A2(n16836), .ZN(n12918) );
  AND2_X1 U14438 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12919) );
  NAND2_X1 U14439 ( .A1(n12919), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14577) );
  INV_X1 U14440 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16879) );
  INV_X1 U14441 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16867) );
  AND2_X1 U14442 ( .A1(n16879), .A2(n16867), .ZN(n12920) );
  NAND2_X1 U14443 ( .A1(n16768), .A2(n16771), .ZN(n16747) );
  INV_X1 U14444 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16757) );
  NAND3_X1 U14445 ( .A1(n21901), .A2(n16758), .A3(n16757), .ZN(n16749) );
  INV_X1 U14446 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21911) );
  INV_X1 U14447 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16752) );
  NAND2_X1 U14448 ( .A1(n21911), .A2(n16752), .ZN(n21902) );
  NOR2_X1 U14449 ( .A1(n16749), .A2(n21902), .ZN(n12921) );
  NOR2_X1 U14450 ( .A1(n20552), .A2(n12921), .ZN(n12922) );
  NAND2_X1 U14451 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21944) );
  INV_X1 U14452 ( .A(n21944), .ZN(n21941) );
  AND2_X1 U14453 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21941), .ZN(
        n21946) );
  NAND3_X1 U14454 ( .A1(n14529), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n21946), .ZN(n12923) );
  NAND2_X1 U14455 ( .A1(n12923), .A2(n20552), .ZN(n20545) );
  NOR2_X1 U14456 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21930) );
  INV_X1 U14457 ( .A(n21930), .ZN(n12924) );
  INV_X1 U14458 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21997) );
  INV_X1 U14459 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21960) );
  NAND2_X1 U14460 ( .A1(n21997), .A2(n21960), .ZN(n16682) );
  NAND2_X1 U14461 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21969) );
  INV_X1 U14462 ( .A(n21969), .ZN(n12926) );
  NAND2_X1 U14463 ( .A1(n12926), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16787) );
  NAND2_X1 U14464 ( .A1(n20552), .A2(n16787), .ZN(n16681) );
  NAND2_X1 U14465 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16808) );
  INV_X1 U14466 ( .A(n16808), .ZN(n12927) );
  NAND2_X1 U14467 ( .A1(n12928), .A2(n20552), .ZN(n16672) );
  NOR2_X1 U14468 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21979) );
  AND2_X1 U14469 ( .A1(n16693), .A2(n21979), .ZN(n12930) );
  INV_X1 U14470 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16823) );
  INV_X1 U14471 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16894) );
  XNOR2_X1 U14472 ( .A(n20552), .B(n16894), .ZN(n12936) );
  INV_X1 U14473 ( .A(n12936), .ZN(n12932) );
  NOR2_X1 U14474 ( .A1(n11861), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12933) );
  INV_X1 U14475 ( .A(n12933), .ZN(n12931) );
  NAND2_X1 U14476 ( .A1(n12932), .A2(n12931), .ZN(n12938) );
  OAI21_X1 U14477 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n11861), .ZN(n12935) );
  INV_X1 U14478 ( .A(n12935), .ZN(n12934) );
  OAI21_X1 U14479 ( .B1(n12934), .B2(n12933), .A(n16894), .ZN(n12937) );
  INV_X1 U14480 ( .A(n12939), .ZN(n12941) );
  OR2_X1 U14481 ( .A1(n14895), .A2(n14580), .ZN(n12940) );
  AND2_X1 U14482 ( .A1(n12941), .A2(n12940), .ZN(n14556) );
  NAND2_X1 U14483 ( .A1(n14789), .A2(n22414), .ZN(n12942) );
  NAND3_X1 U14484 ( .A1(n14556), .A2(n12943), .A3(n12942), .ZN(n14532) );
  NOR2_X1 U14485 ( .A1(n14532), .A2(n14559), .ZN(n17733) );
  NOR2_X1 U14486 ( .A1(n16422), .A2(n22234), .ZN(n15124) );
  NAND3_X1 U14487 ( .A1(n22225), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(
        P1_STATEBS16_REG_SCAN_IN), .ZN(n22220) );
  INV_X1 U14488 ( .A(n22220), .ZN(n12944) );
  NOR2_X2 U14489 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22440) );
  NAND2_X1 U14490 ( .A1(n12944), .A2(n22440), .ZN(n20538) );
  OR2_X1 U14491 ( .A1(n16590), .A2(n20538), .ZN(n12951) );
  INV_X1 U14492 ( .A(n22440), .ZN(n22497) );
  NAND2_X1 U14493 ( .A1(n22497), .A2(n12947), .ZN(n21861) );
  AND2_X1 U14494 ( .A1(n21861), .A2(n22225), .ZN(n12945) );
  NAND2_X1 U14495 ( .A1(n22225), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17712) );
  NAND2_X1 U14496 ( .A1(n12946), .A2(n17712), .ZN(n14804) );
  NOR2_X2 U14497 ( .A1(n12947), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22170) );
  NAND2_X1 U14498 ( .A1(n22170), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n16801) );
  OAI21_X1 U14499 ( .B1(n20506), .B2(n12948), .A(n16801), .ZN(n12949) );
  NAND3_X1 U14500 ( .A1(n12952), .A2(n12951), .A3(n12950), .ZN(P1_U2968) );
  INV_X1 U14501 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16097) );
  INV_X1 U14502 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17288) );
  INV_X1 U14503 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17277) );
  INV_X1 U14504 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17221) );
  INV_X1 U14505 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17200) );
  INV_X1 U14506 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17194) );
  INV_X1 U14507 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17183) );
  INV_X1 U14508 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17158) );
  INV_X1 U14509 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13275) );
  INV_X1 U14510 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12956) );
  AOI21_X1 U14511 ( .B1(n16097), .B2(n12958), .A(n13002), .ZN(n16099) );
  NAND2_X1 U14512 ( .A1(n12955), .A2(n12956), .ZN(n12957) );
  NAND2_X1 U14513 ( .A1(n12958), .A2(n12957), .ZN(n19169) );
  INV_X1 U14514 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16155) );
  INV_X1 U14515 ( .A(n12998), .ZN(n12961) );
  AOI21_X1 U14516 ( .B1(n17158), .B2(n12960), .A(n12961), .ZN(n17161) );
  AND2_X1 U14517 ( .A1(n12965), .A2(n17183), .ZN(n12962) );
  NOR2_X1 U14518 ( .A1(n12996), .A2(n12962), .ZN(n19106) );
  NAND2_X1 U14519 ( .A1(n12967), .A2(n17194), .ZN(n12964) );
  AND2_X1 U14520 ( .A1(n12965), .A2(n12964), .ZN(n19094) );
  AOI21_X1 U14521 ( .B1(n17200), .B2(n12966), .A(n11666), .ZN(n19080) );
  OAI21_X1 U14522 ( .B1(n12968), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n12966), .ZN(n14479) );
  INV_X1 U14523 ( .A(n14479), .ZN(n16941) );
  AOI21_X1 U14524 ( .B1(n17221), .B2(n12969), .A(n12968), .ZN(n19066) );
  OAI21_X1 U14525 ( .B1(n12970), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n12969), .ZN(n16960) );
  INV_X1 U14526 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19038) );
  INV_X1 U14527 ( .A(n12971), .ZN(n12972) );
  AOI21_X1 U14528 ( .B1(n19038), .B2(n12972), .A(n12990), .ZN(n19034) );
  AND2_X1 U14529 ( .A1(n12987), .A2(n17277), .ZN(n12973) );
  OR2_X1 U14530 ( .A1(n12973), .A2(n12988), .ZN(n19026) );
  INV_X1 U14531 ( .A(n19026), .ZN(n17280) );
  NAND2_X1 U14532 ( .A1(n12975), .A2(n11682), .ZN(n12976) );
  NAND2_X1 U14533 ( .A1(n12974), .A2(n12976), .ZN(n17299) );
  AOI21_X1 U14534 ( .B1(n17318), .B2(n12977), .A(n12978), .ZN(n17317) );
  AOI21_X1 U14535 ( .B1(n17338), .B2(n12979), .A(n12980), .ZN(n18995) );
  AOI21_X1 U14536 ( .B1(n15755), .B2(n12981), .A(n11209), .ZN(n18978) );
  AOI21_X1 U14537 ( .B1(n17763), .B2(n12982), .A(n12983), .ZN(n17753) );
  OAI22_X1 U14538 ( .A1(n17752), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n12984) );
  INV_X1 U14539 ( .A(n12984), .ZN(n17642) );
  INV_X1 U14540 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14719) );
  AOI22_X1 U14541 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14719), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17752), .ZN(n16963) );
  NOR2_X1 U14542 ( .A1(n17642), .A2(n16963), .ZN(n16962) );
  OAI21_X1 U14543 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12982), .ZN(n15825) );
  NAND2_X1 U14544 ( .A1(n16962), .A2(n15825), .ZN(n15726) );
  NOR2_X1 U14545 ( .A1(n17753), .A2(n15726), .ZN(n16017) );
  OAI21_X1 U14546 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12983), .A(
        n12981), .ZN(n17769) );
  NAND2_X1 U14547 ( .A1(n16017), .A2(n17769), .ZN(n18976) );
  NOR2_X1 U14548 ( .A1(n18978), .A2(n18976), .ZN(n18987) );
  OAI21_X1 U14549 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11209), .A(
        n12979), .ZN(n18988) );
  NAND2_X1 U14550 ( .A1(n18987), .A2(n18988), .ZN(n18994) );
  NOR2_X1 U14551 ( .A1(n18995), .A2(n18994), .ZN(n15835) );
  OAI21_X1 U14552 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12980), .A(
        n12977), .ZN(n17789) );
  NAND2_X1 U14553 ( .A1(n15835), .A2(n17789), .ZN(n19008) );
  NOR2_X1 U14554 ( .A1(n17317), .A2(n19008), .ZN(n15814) );
  OR2_X1 U14555 ( .A1(n12978), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12985) );
  NAND2_X1 U14556 ( .A1(n12975), .A2(n12985), .ZN(n17312) );
  AND2_X1 U14557 ( .A1(n15814), .A2(n17312), .ZN(n15910) );
  NAND2_X1 U14558 ( .A1(n17299), .A2(n15910), .ZN(n15925) );
  INV_X1 U14559 ( .A(n15925), .ZN(n15909) );
  NAND2_X1 U14560 ( .A1(n12974), .A2(n17288), .ZN(n12986) );
  NAND2_X1 U14561 ( .A1(n12987), .A2(n12986), .ZN(n17289) );
  NAND2_X1 U14562 ( .A1(n15909), .A2(n17289), .ZN(n19016) );
  NOR2_X1 U14563 ( .A1(n17280), .A2(n19016), .ZN(n19017) );
  NOR2_X1 U14564 ( .A1(n12988), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12989) );
  OR2_X1 U14565 ( .A1(n12971), .A2(n12989), .ZN(n17268) );
  NAND2_X1 U14566 ( .A1(n19017), .A2(n17268), .ZN(n19031) );
  NOR2_X1 U14567 ( .A1(n19034), .A2(n19031), .ZN(n15785) );
  OR2_X1 U14568 ( .A1(n12990), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12991) );
  NAND2_X1 U14569 ( .A1(n12991), .A2(n12992), .ZN(n17239) );
  AND2_X1 U14570 ( .A1(n15785), .A2(n17239), .ZN(n19058) );
  INV_X1 U14571 ( .A(n12970), .ZN(n12994) );
  NAND2_X1 U14572 ( .A1(n12953), .A2(n12992), .ZN(n12993) );
  NAND2_X1 U14573 ( .A1(n12994), .A2(n12993), .ZN(n19057) );
  NAND2_X1 U14574 ( .A1(n19058), .A2(n19057), .ZN(n12995) );
  NOR2_X1 U14575 ( .A1(n19066), .A2(n19065), .ZN(n19064) );
  NOR2_X1 U14576 ( .A1(n19134), .A2(n19064), .ZN(n16940) );
  NOR2_X1 U14577 ( .A1(n16941), .A2(n16940), .ZN(n16939) );
  NOR2_X1 U14578 ( .A1(n19134), .A2(n16939), .ZN(n19079) );
  NOR2_X1 U14579 ( .A1(n19080), .A2(n19079), .ZN(n19078) );
  NOR2_X1 U14580 ( .A1(n19134), .A2(n19078), .ZN(n19093) );
  NOR2_X1 U14581 ( .A1(n19094), .A2(n19093), .ZN(n19092) );
  NOR2_X1 U14582 ( .A1(n19134), .A2(n19092), .ZN(n19105) );
  NOR2_X1 U14583 ( .A1(n19106), .A2(n19105), .ZN(n19104) );
  OR2_X1 U14584 ( .A1(n12996), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12997) );
  NAND2_X1 U14585 ( .A1(n12960), .A2(n12997), .ZN(n19121) );
  AOI21_X1 U14586 ( .B1(n19104), .B2(n19121), .A(n19134), .ZN(n16934) );
  NOR2_X1 U14587 ( .A1(n17161), .A2(n16934), .ZN(n19137) );
  AND2_X1 U14588 ( .A1(n12998), .A2(n13275), .ZN(n12999) );
  OR2_X1 U14589 ( .A1(n12999), .A2(n11309), .ZN(n19133) );
  AOI21_X1 U14590 ( .B1(n19137), .B2(n19133), .A(n19134), .ZN(n13000) );
  INV_X1 U14591 ( .A(n13000), .ZN(n19147) );
  OR2_X1 U14592 ( .A1(n11309), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13001) );
  NAND2_X1 U14593 ( .A1(n12955), .A2(n13001), .ZN(n19148) );
  XNOR2_X1 U14594 ( .A(n13002), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16913) );
  INV_X1 U14595 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n17690) );
  INV_X1 U14596 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n22239) );
  NAND4_X1 U14597 ( .A1(n17752), .A2(n17690), .A3(n22239), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19201) );
  INV_X1 U14598 ( .A(n19201), .ZN(n19167) );
  NAND2_X1 U14599 ( .A1(n16914), .A2(n16913), .ZN(n13003) );
  OAI211_X1 U14600 ( .C1(n16914), .C2(n16913), .A(n19167), .B(n13003), .ZN(
        n13648) );
  NAND2_X2 U14601 ( .A1(n13329), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16394) );
  INV_X2 U14602 ( .A(n16394), .ZN(n16386) );
  AOI22_X1 U14603 ( .A1(n16386), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U14604 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13004) );
  AND2_X1 U14605 ( .A1(n13005), .A2(n13004), .ZN(n13008) );
  NOR2_X1 U14606 ( .A1(n15234), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13326) );
  AOI22_X1 U14607 ( .A1(n11162), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13007) );
  AND2_X4 U14608 ( .A1(n15192), .A2(n14219), .ZN(n13021) );
  AOI22_X1 U14609 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11190), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13006) );
  NAND3_X1 U14610 ( .A1(n13008), .A2(n13007), .A3(n13006), .ZN(n13009) );
  NAND2_X1 U14611 ( .A1(n13009), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13017) );
  AOI22_X1 U14612 ( .A1(n16386), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U14613 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13010) );
  AND2_X1 U14614 ( .A1(n13011), .A2(n13010), .ZN(n13014) );
  AOI22_X1 U14615 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U14616 ( .A1(n16399), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11192), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13012) );
  NAND3_X1 U14617 ( .A1(n13014), .A2(n13013), .A3(n13012), .ZN(n13015) );
  NAND2_X1 U14618 ( .A1(n13015), .A2(n15200), .ZN(n13016) );
  INV_X2 U14619 ( .A(n13064), .ZN(n14700) );
  INV_X4 U14620 ( .A(n16394), .ZN(n16376) );
  BUF_X4 U14621 ( .A(n13021), .Z(n16385) );
  AOI22_X1 U14622 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11189), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U14623 ( .A1(n16386), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U14624 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13024) );
  AOI22_X1 U14625 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13023) );
  AOI22_X1 U14626 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11191), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13026) );
  NAND2_X1 U14627 ( .A1(n13064), .A2(n11183), .ZN(n13105) );
  AOI22_X1 U14628 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11190), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U14629 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13029) );
  AOI22_X1 U14630 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13028) );
  NAND4_X1 U14631 ( .A1(n13031), .A2(n13030), .A3(n13029), .A4(n13028), .ZN(
        n13032) );
  NAND2_X1 U14632 ( .A1(n13032), .A2(n15200), .ZN(n13039) );
  AOI22_X1 U14633 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11196), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U14634 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U14635 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13033) );
  NAND4_X1 U14636 ( .A1(n13036), .A2(n13035), .A3(n13034), .A4(n13033), .ZN(
        n13037) );
  NAND2_X1 U14637 ( .A1(n13037), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13038) );
  NAND2_X2 U14638 ( .A1(n13039), .A2(n13038), .ZN(n13111) );
  INV_X2 U14639 ( .A(n13111), .ZN(n20030) );
  NAND2_X1 U14640 ( .A1(n14252), .A2(n20030), .ZN(n13041) );
  NAND2_X1 U14641 ( .A1(n13358), .A2(n13111), .ZN(n13040) );
  NAND2_X1 U14642 ( .A1(n13041), .A2(n13040), .ZN(n13053) );
  AOI22_X1 U14643 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13042), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U14644 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11189), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U14645 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13044) );
  AOI22_X1 U14646 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11185), .B1(
        n16400), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13043) );
  NAND4_X1 U14647 ( .A1(n13046), .A2(n13045), .A3(n13044), .A4(n13043), .ZN(
        n13052) );
  AOI22_X1 U14648 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11192), .B1(
        n16399), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U14649 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U14650 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13047) );
  NAND4_X1 U14651 ( .A1(n13050), .A2(n13049), .A3(n13048), .A4(n13047), .ZN(
        n13051) );
  MUX2_X2 U14652 ( .A(n13052), .B(n13051), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14710) );
  NAND2_X1 U14653 ( .A1(n13053), .A2(n14710), .ZN(n14407) );
  AOI22_X1 U14654 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U14655 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U14656 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16400), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U14657 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13054) );
  NAND4_X1 U14658 ( .A1(n13057), .A2(n13056), .A3(n13055), .A4(n13054), .ZN(
        n13063) );
  AOI22_X1 U14659 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13061) );
  AOI22_X1 U14660 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11189), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U14661 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U14662 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13058) );
  NAND4_X1 U14663 ( .A1(n13061), .A2(n13060), .A3(n13059), .A4(n13058), .ZN(
        n13062) );
  NAND2_X1 U14664 ( .A1(n14407), .A2(n14410), .ZN(n13066) );
  AOI22_X1 U14665 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U14666 ( .A1(n11193), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16400), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U14667 ( .A1(n16399), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13067) );
  NAND2_X1 U14668 ( .A1(n13071), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13077) );
  AOI22_X1 U14669 ( .A1(n11162), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U14670 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13074) );
  NAND2_X1 U14671 ( .A1(n13075), .A2(n11233), .ZN(n13076) );
  NAND2_X2 U14672 ( .A1(n13077), .A2(n13076), .ZN(n13109) );
  AOI22_X1 U14673 ( .A1(n16386), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13079) );
  AOI22_X1 U14674 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13078) );
  NAND4_X1 U14675 ( .A1(n13081), .A2(n13080), .A3(n13079), .A4(n13078), .ZN(
        n13087) );
  AOI22_X1 U14676 ( .A1(n16399), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11194), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U14677 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U14678 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13082) );
  NAND4_X1 U14679 ( .A1(n13085), .A2(n13084), .A3(n13083), .A4(n13082), .ZN(
        n13086) );
  MUX2_X2 U14680 ( .A(n13087), .B(n13086), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13113) );
  NAND2_X2 U14681 ( .A1(n19175), .A2(n13113), .ZN(n13619) );
  NAND2_X1 U14682 ( .A1(n13110), .A2(n14410), .ZN(n13089) );
  NAND2_X1 U14683 ( .A1(n13089), .A2(n13088), .ZN(n13124) );
  NAND3_X1 U14684 ( .A1(n20079), .A2(n20030), .A3(n14878), .ZN(n13090) );
  NAND2_X1 U14685 ( .A1(n13124), .A2(n13090), .ZN(n13118) );
  AOI22_X1 U14686 ( .A1(n11162), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U14687 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11191), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U14688 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U14689 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13091) );
  NAND4_X1 U14690 ( .A1(n13094), .A2(n13093), .A3(n13092), .A4(n13091), .ZN(
        n13095) );
  NAND2_X1 U14691 ( .A1(n13095), .A2(n15200), .ZN(n13103) );
  AOI22_X1 U14692 ( .A1(n16400), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13097) );
  AOI22_X1 U14693 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13096) );
  NAND3_X1 U14694 ( .A1(n13098), .A2(n13097), .A3(n13096), .ZN(n13101) );
  AOI22_X1 U14695 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11190), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13099) );
  NAND2_X1 U14696 ( .A1(n13118), .A2(n13107), .ZN(n13108) );
  NAND2_X1 U14697 ( .A1(n13113), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14216) );
  NOR2_X1 U14698 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13609) );
  INV_X1 U14699 ( .A(n13609), .ZN(n19195) );
  NAND2_X2 U14700 ( .A1(n20079), .A2(n14257), .ZN(n14404) );
  AND2_X1 U14701 ( .A1(n14878), .A2(n14710), .ZN(n14748) );
  NAND4_X1 U14702 ( .A1(n13115), .A2(n14412), .A3(n19982), .A4(n14748), .ZN(
        n13119) );
  NAND2_X1 U14703 ( .A1(n13118), .A2(n13117), .ZN(n13314) );
  OAI211_X1 U14704 ( .C1(n19195), .C2(n19889), .A(n13127), .B(n13126), .ZN(
        n13120) );
  INV_X1 U14705 ( .A(n13120), .ZN(n13121) );
  INV_X1 U14706 ( .A(n14412), .ZN(n13122) );
  AOI21_X1 U14707 ( .B1(n11563), .B2(n20237), .A(n14410), .ZN(n13125) );
  INV_X1 U14708 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n16969) );
  NAND2_X1 U14709 ( .A1(n16146), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n13129) );
  AOI22_X1 U14710 ( .A1(n13164), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13128) );
  NAND2_X1 U14711 ( .A1(n13131), .A2(n13130), .ZN(n13132) );
  AND2_X2 U14712 ( .A1(n13151), .A2(n13132), .ZN(n14088) );
  NAND2_X1 U14713 ( .A1(n13624), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13133) );
  NOR2_X1 U14714 ( .A1(n13133), .A2(n14404), .ZN(n13134) );
  NAND2_X1 U14715 ( .A1(n13609), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13135) );
  AND2_X1 U14716 ( .A1(n13136), .A2(n13135), .ZN(n13137) );
  NAND2_X1 U14717 ( .A1(n13138), .A2(n13137), .ZN(n14090) );
  NAND2_X1 U14718 ( .A1(n13140), .A2(n13139), .ZN(n14402) );
  NAND2_X1 U14719 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13141) );
  NAND3_X1 U14720 ( .A1(n13142), .A2(n19195), .A3(n13141), .ZN(n13145) );
  INV_X1 U14721 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13617) );
  NOR2_X1 U14722 ( .A1(n13143), .A2(n13617), .ZN(n13144) );
  NOR2_X1 U14723 ( .A1(n13145), .A2(n13144), .ZN(n13147) );
  NAND2_X1 U14724 ( .A1(n13163), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13148) );
  NAND2_X2 U14725 ( .A1(n14090), .A2(n14089), .ZN(n14092) );
  NAND2_X1 U14726 ( .A1(n14088), .A2(n14092), .ZN(n13152) );
  NAND2_X1 U14727 ( .A1(n13152), .A2(n13151), .ZN(n14087) );
  NAND2_X1 U14728 ( .A1(n13161), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13154) );
  AOI21_X1 U14729 ( .B1(n17752), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13153) );
  INV_X1 U14730 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13621) );
  NAND2_X1 U14731 ( .A1(n13163), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13156) );
  AOI22_X1 U14732 ( .A1(n13164), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13155) );
  NAND2_X1 U14733 ( .A1(n13158), .A2(n13157), .ZN(n13159) );
  NOR2_X1 U14734 ( .A1(n19195), .A2(n19777), .ZN(n13162) );
  INV_X1 U14735 ( .A(n13163), .ZN(n16149) );
  INV_X1 U14736 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13623) );
  NAND2_X1 U14737 ( .A1(n13164), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13166) );
  NAND2_X1 U14738 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13165) );
  OAI211_X1 U14739 ( .C1(n13143), .C2(n13623), .A(n13166), .B(n13165), .ZN(
        n13167) );
  NAND2_X1 U14740 ( .A1(n13168), .A2(n13169), .ZN(n13173) );
  INV_X1 U14741 ( .A(n13168), .ZN(n13171) );
  INV_X1 U14742 ( .A(n13169), .ZN(n13170) );
  NAND2_X1 U14743 ( .A1(n13171), .A2(n13170), .ZN(n13172) );
  INV_X1 U14744 ( .A(n14085), .ZN(n13175) );
  INV_X1 U14745 ( .A(n13173), .ZN(n13174) );
  INV_X1 U14746 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U14747 ( .A1(n13176), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13178) );
  AOI22_X1 U14748 ( .A1(n13164), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13177) );
  OAI211_X1 U14749 ( .C1(n13289), .C2(n13625), .A(n13178), .B(n13177), .ZN(
        n15654) );
  NAND2_X1 U14750 ( .A1(n15655), .A2(n15654), .ZN(n15739) );
  NAND2_X1 U14751 ( .A1(n13176), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13183) );
  INV_X1 U14752 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18972) );
  INV_X2 U14753 ( .A(n16146), .ZN(n13289) );
  NAND2_X1 U14754 ( .A1(n13164), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n13180) );
  NAND2_X1 U14755 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13179) );
  OAI211_X1 U14756 ( .C1(n18972), .C2(n13289), .A(n13180), .B(n13179), .ZN(
        n13181) );
  INV_X1 U14757 ( .A(n13181), .ZN(n13182) );
  NAND2_X1 U14758 ( .A1(n13176), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13189) );
  INV_X1 U14759 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n13185) );
  INV_X1 U14760 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13184) );
  OAI22_X1 U14761 ( .A1(n13287), .A2(n13185), .B1(n13265), .B2(n13184), .ZN(
        n13187) );
  INV_X1 U14762 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n14942) );
  NOR2_X1 U14763 ( .A1(n13289), .A2(n14942), .ZN(n13186) );
  NOR2_X1 U14764 ( .A1(n13187), .A2(n13186), .ZN(n13188) );
  NAND2_X1 U14765 ( .A1(n13189), .A2(n13188), .ZN(n14939) );
  NAND2_X1 U14766 ( .A1(n14937), .A2(n14939), .ZN(n14938) );
  INV_X1 U14767 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13629) );
  NAND2_X1 U14768 ( .A1(n13164), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n13191) );
  NAND2_X1 U14769 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13190) );
  OAI211_X1 U14770 ( .C1(n13289), .C2(n13629), .A(n13191), .B(n13190), .ZN(
        n13192) );
  AOI21_X1 U14771 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n13176), .A(
        n13192), .ZN(n14884) );
  NAND2_X1 U14772 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13199) );
  INV_X1 U14773 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n15841) );
  INV_X1 U14774 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13195) );
  OAI22_X1 U14775 ( .A1(n13287), .A2(n15841), .B1(n13265), .B2(n13195), .ZN(
        n13197) );
  INV_X1 U14776 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n15842) );
  NOR2_X1 U14777 ( .A1(n13289), .A2(n15842), .ZN(n13196) );
  NOR2_X1 U14778 ( .A1(n13197), .A2(n13196), .ZN(n13198) );
  OR2_X2 U14779 ( .A1(n15118), .A2(n15117), .ZN(n15154) );
  NAND2_X1 U14780 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13204) );
  INV_X1 U14781 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n13200) );
  OAI22_X1 U14782 ( .A1(n13287), .A2(n13200), .B1(n13265), .B2(n17318), .ZN(
        n13202) );
  INV_X1 U14783 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13630) );
  NOR2_X1 U14784 ( .A1(n13289), .A2(n13630), .ZN(n13201) );
  NOR2_X1 U14785 ( .A1(n13202), .A2(n13201), .ZN(n13203) );
  NOR2_X4 U14786 ( .A1(n15154), .A2(n15153), .ZN(n15178) );
  INV_X1 U14787 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n15819) );
  NAND2_X1 U14788 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13206) );
  AOI22_X1 U14789 ( .A1(n13164), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n13205) );
  OAI211_X1 U14790 ( .C1(n13289), .C2(n15819), .A(n13206), .B(n13205), .ZN(
        n15177) );
  NAND2_X1 U14791 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13210) );
  INV_X1 U14792 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n17872) );
  INV_X1 U14793 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13265) );
  OAI22_X1 U14794 ( .A1(n13287), .A2(n17872), .B1(n13265), .B2(n11682), .ZN(
        n13208) );
  INV_X1 U14795 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13632) );
  NOR2_X1 U14796 ( .A1(n13289), .A2(n13632), .ZN(n13207) );
  NOR2_X1 U14797 ( .A1(n13208), .A2(n13207), .ZN(n13209) );
  NAND2_X1 U14798 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13214) );
  INV_X1 U14799 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n13531) );
  OAI22_X1 U14800 ( .A1(n13287), .A2(n13531), .B1(n13265), .B2(n17288), .ZN(
        n13212) );
  INV_X1 U14801 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13633) );
  NOR2_X1 U14802 ( .A1(n13289), .A2(n13633), .ZN(n13211) );
  NOR2_X1 U14803 ( .A1(n13212), .A2(n13211), .ZN(n13213) );
  INV_X1 U14804 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13634) );
  NAND2_X1 U14805 ( .A1(n13176), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13216) );
  AOI22_X1 U14806 ( .A1(n13164), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n13215) );
  OAI211_X1 U14807 ( .C1(n13289), .C2(n13634), .A(n13216), .B(n13215), .ZN(
        n15445) );
  NAND2_X1 U14808 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13223) );
  INV_X1 U14809 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n13218) );
  INV_X1 U14810 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13217) );
  OAI22_X1 U14811 ( .A1(n13287), .A2(n13218), .B1(n13265), .B2(n13217), .ZN(
        n13221) );
  INV_X1 U14812 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13219) );
  NOR2_X1 U14813 ( .A1(n13289), .A2(n13219), .ZN(n13220) );
  NOR2_X1 U14814 ( .A1(n13221), .A2(n13220), .ZN(n13222) );
  NAND2_X1 U14815 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13229) );
  INV_X1 U14816 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n13224) );
  OAI22_X1 U14817 ( .A1(n13287), .A2(n13224), .B1(n13265), .B2(n19038), .ZN(
        n13227) );
  INV_X1 U14818 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13225) );
  NOR2_X1 U14819 ( .A1(n13289), .A2(n13225), .ZN(n13226) );
  NOR2_X1 U14820 ( .A1(n13227), .A2(n13226), .ZN(n13228) );
  INV_X1 U14821 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n13232) );
  NAND2_X1 U14822 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13231) );
  AOI22_X1 U14823 ( .A1(n13164), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n13230) );
  OAI211_X1 U14824 ( .C1(n13289), .C2(n13232), .A(n13231), .B(n13230), .ZN(
        n15690) );
  NAND2_X1 U14825 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13236) );
  INV_X1 U14826 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n17880) );
  OAI22_X1 U14827 ( .A1(n13287), .A2(n17880), .B1(n13265), .B2(n12953), .ZN(
        n13234) );
  INV_X1 U14828 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n19053) );
  NOR2_X1 U14829 ( .A1(n13289), .A2(n19053), .ZN(n13233) );
  NOR2_X1 U14830 ( .A1(n13234), .A2(n13233), .ZN(n13235) );
  NAND2_X1 U14831 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13242) );
  INV_X1 U14832 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n13238) );
  INV_X1 U14833 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13237) );
  OAI22_X1 U14834 ( .A1(n13287), .A2(n13238), .B1(n13265), .B2(n13237), .ZN(
        n13240) );
  INV_X1 U14835 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n13635) );
  NOR2_X1 U14836 ( .A1(n13289), .A2(n13635), .ZN(n13239) );
  NOR2_X1 U14837 ( .A1(n13240), .A2(n13239), .ZN(n13241) );
  NAND2_X1 U14838 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13247) );
  INV_X1 U14839 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19070) );
  OAI22_X1 U14840 ( .A1(n13287), .A2(n19070), .B1(n13265), .B2(n17221), .ZN(
        n13245) );
  INV_X1 U14841 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n13243) );
  NOR2_X1 U14842 ( .A1(n13289), .A2(n13243), .ZN(n13244) );
  NOR2_X1 U14843 ( .A1(n13245), .A2(n13244), .ZN(n13246) );
  INV_X1 U14844 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n13250) );
  NAND2_X1 U14845 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13249) );
  AOI22_X1 U14846 ( .A1(n13164), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n13248) );
  OAI211_X1 U14847 ( .C1(n13289), .C2(n13250), .A(n13249), .B(n13248), .ZN(
        n14473) );
  NAND2_X1 U14848 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13254) );
  INV_X1 U14849 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19083) );
  OAI22_X1 U14850 ( .A1(n13287), .A2(n19083), .B1(n13265), .B2(n17200), .ZN(
        n13252) );
  INV_X1 U14851 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n19082) );
  NOR2_X1 U14852 ( .A1(n13289), .A2(n19082), .ZN(n13251) );
  NOR2_X1 U14853 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  AND2_X1 U14854 ( .A1(n13254), .A2(n13253), .ZN(n17035) );
  NAND2_X1 U14855 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13260) );
  INV_X1 U14856 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n13255) );
  OAI22_X1 U14857 ( .A1(n13287), .A2(n13255), .B1(n13265), .B2(n17194), .ZN(
        n13258) );
  INV_X1 U14858 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n13256) );
  NOR2_X1 U14859 ( .A1(n13289), .A2(n13256), .ZN(n13257) );
  NOR2_X1 U14860 ( .A1(n13258), .A2(n13257), .ZN(n13259) );
  NOR2_X4 U14861 ( .A1(n11223), .A2(n17029), .ZN(n17030) );
  NAND2_X1 U14862 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13264) );
  INV_X1 U14863 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19110) );
  OAI22_X1 U14864 ( .A1(n13287), .A2(n19110), .B1(n13265), .B2(n17183), .ZN(
        n13262) );
  INV_X1 U14865 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n19109) );
  NOR2_X1 U14866 ( .A1(n13289), .A2(n19109), .ZN(n13261) );
  NOR2_X1 U14867 ( .A1(n13262), .A2(n13261), .ZN(n13263) );
  NAND2_X1 U14868 ( .A1(n13264), .A2(n13263), .ZN(n17022) );
  NAND2_X1 U14869 ( .A1(n13176), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13270) );
  INV_X1 U14870 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n17888) );
  OAI22_X1 U14871 ( .A1(n13287), .A2(n17888), .B1(n13265), .B2(n11716), .ZN(
        n13268) );
  INV_X1 U14872 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n13266) );
  NOR2_X1 U14873 ( .A1(n13289), .A2(n13266), .ZN(n13267) );
  NOR2_X1 U14874 ( .A1(n13268), .A2(n13267), .ZN(n13269) );
  NAND2_X1 U14875 ( .A1(n13270), .A2(n13269), .ZN(n17017) );
  NAND2_X1 U14876 ( .A1(n13176), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13274) );
  INV_X1 U14877 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n17891) );
  OAI22_X1 U14878 ( .A1(n13287), .A2(n17891), .B1(n13265), .B2(n17158), .ZN(
        n13272) );
  INV_X1 U14879 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16931) );
  NOR2_X1 U14880 ( .A1(n13289), .A2(n16931), .ZN(n13271) );
  NOR2_X1 U14881 ( .A1(n13272), .A2(n13271), .ZN(n13273) );
  AND2_X1 U14882 ( .A1(n13274), .A2(n13273), .ZN(n16925) );
  NAND2_X1 U14883 ( .A1(n13176), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13279) );
  INV_X1 U14884 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n17892) );
  OAI22_X1 U14885 ( .A1(n13287), .A2(n17892), .B1(n13265), .B2(n13275), .ZN(
        n13277) );
  INV_X1 U14886 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n13637) );
  NOR2_X1 U14887 ( .A1(n13289), .A2(n13637), .ZN(n13276) );
  NOR2_X1 U14888 ( .A1(n13277), .A2(n13276), .ZN(n13278) );
  AND2_X1 U14889 ( .A1(n13279), .A2(n13278), .ZN(n17000) );
  NAND2_X1 U14890 ( .A1(n13163), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13283) );
  INV_X1 U14891 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n17895) );
  OAI22_X1 U14892 ( .A1(n13287), .A2(n17895), .B1(n13265), .B2(n11717), .ZN(
        n13281) );
  INV_X1 U14893 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n13638) );
  NOR2_X1 U14894 ( .A1(n13289), .A2(n13638), .ZN(n13280) );
  NOR2_X1 U14895 ( .A1(n13281), .A2(n13280), .ZN(n13282) );
  NAND2_X1 U14896 ( .A1(n13283), .A2(n13282), .ZN(n16996) );
  INV_X1 U14897 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n13286) );
  NAND2_X1 U14898 ( .A1(n13163), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13285) );
  AOI22_X1 U14899 ( .A1(n13164), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n13284) );
  OAI211_X1 U14900 ( .C1(n13289), .C2(n13286), .A(n13285), .B(n13284), .ZN(
        n16987) );
  NAND2_X1 U14901 ( .A1(n13163), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13293) );
  INV_X1 U14902 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17899) );
  OAI22_X1 U14903 ( .A1(n13287), .A2(n17899), .B1(n13265), .B2(n16097), .ZN(
        n13291) );
  INV_X1 U14904 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n13288) );
  NOR2_X1 U14905 ( .A1(n13289), .A2(n13288), .ZN(n13290) );
  NOR2_X1 U14906 ( .A1(n13291), .A2(n13290), .ZN(n13292) );
  AND2_X1 U14907 ( .A1(n13293), .A2(n13292), .ZN(n14445) );
  INV_X1 U14908 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n13297) );
  NAND2_X1 U14909 ( .A1(n13294), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13296) );
  AOI22_X1 U14910 ( .A1(n13164), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n13295) );
  OAI211_X1 U14911 ( .C1(n13289), .C2(n13297), .A(n13296), .B(n13295), .ZN(
        n16144) );
  XNOR2_X1 U14912 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14266) );
  NAND2_X1 U14913 ( .A1(n14266), .A2(n14218), .ZN(n13299) );
  NAND2_X1 U14914 ( .A1(n19889), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13298) );
  NAND2_X1 U14915 ( .A1(n13299), .A2(n13298), .ZN(n13307) );
  XNOR2_X1 U14916 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13308) );
  NAND2_X1 U14917 ( .A1(n13307), .A2(n13308), .ZN(n13311) );
  NAND2_X1 U14918 ( .A1(n19766), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13300) );
  XNOR2_X1 U14919 ( .A(n15200), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13305) );
  INV_X1 U14920 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19179) );
  INV_X1 U14921 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17695) );
  NOR2_X1 U14922 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17695), .ZN(
        n13303) );
  AOI221_X1 U14923 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n13304), 
        .C1(n19179), .C2(n13304), .A(n13303), .ZN(n14269) );
  NAND3_X1 U14924 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13304), .A3(
        n19179), .ZN(n14212) );
  XNOR2_X1 U14925 ( .A(n13306), .B(n13305), .ZN(n14234) );
  INV_X1 U14926 ( .A(n13307), .ZN(n13310) );
  INV_X1 U14927 ( .A(n13308), .ZN(n13309) );
  NAND2_X1 U14928 ( .A1(n13310), .A2(n13309), .ZN(n13312) );
  AND2_X1 U14929 ( .A1(n13312), .A2(n13311), .ZN(n14223) );
  NAND3_X1 U14930 ( .A1(n14212), .A2(n14234), .A3(n14223), .ZN(n14246) );
  XNOR2_X1 U14931 ( .A(n14266), .B(n14218), .ZN(n14224) );
  NOR2_X1 U14932 ( .A1(n14246), .A2(n14224), .ZN(n13313) );
  OR2_X1 U14933 ( .A1(n14269), .A2(n13313), .ZN(n15257) );
  INV_X1 U14934 ( .A(n13315), .ZN(n13316) );
  OR2_X1 U14935 ( .A1(n14383), .A2(n13316), .ZN(n15256) );
  INV_X1 U14936 ( .A(n15256), .ZN(n13317) );
  AND3_X1 U14937 ( .A1(n13265), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18966) );
  INV_X1 U14938 ( .A(n18966), .ZN(n19219) );
  AND2_X1 U14939 ( .A1(n18968), .A2(n13624), .ZN(n13644) );
  NAND2_X1 U14940 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19213) );
  AND2_X1 U14941 ( .A1(n19213), .A2(n22239), .ZN(n13642) );
  INV_X1 U14942 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n22289) );
  INV_X1 U14943 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n17685) );
  INV_X1 U14944 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n17684) );
  NAND2_X1 U14945 ( .A1(n17685), .A2(n17684), .ZN(n13318) );
  NAND2_X1 U14946 ( .A1(n17684), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n22278) );
  OAI21_X1 U14947 ( .B1(n22289), .B2(n13318), .A(n17904), .ZN(n18957) );
  NAND2_X1 U14948 ( .A1(n19213), .A2(n18957), .ZN(n14239) );
  NOR2_X1 U14949 ( .A1(n14239), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n13613) );
  NAND2_X1 U14950 ( .A1(n20178), .A2(n13113), .ZN(n14271) );
  INV_X1 U14951 ( .A(n14271), .ZN(n13319) );
  AND2_X1 U14952 ( .A1(n13613), .A2(n13319), .ZN(n15281) );
  NAND2_X1 U14953 ( .A1(n18968), .A2(n15281), .ZN(n19161) );
  INV_X1 U14954 ( .A(n19161), .ZN(n19118) );
  INV_X1 U14955 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19876) );
  AND2_X2 U14956 ( .A1(n16398), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13369) );
  AOI22_X1 U14958 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13325) );
  AND2_X2 U14959 ( .A1(n13042), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16210) );
  AOI22_X1 U14961 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13324) );
  AND2_X2 U14962 ( .A1(n11184), .A2(n15200), .ZN(n13344) );
  AND2_X2 U14963 ( .A1(n13321), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13442) );
  AOI22_X1 U14964 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13323) );
  AND2_X2 U14965 ( .A1(n16384), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13447) );
  AOI22_X1 U14966 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13322) );
  NAND4_X1 U14967 ( .A1(n13325), .A2(n13324), .A3(n13323), .A4(n13322), .ZN(
        n13336) );
  AND2_X2 U14968 ( .A1(n16386), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16194) );
  AND2_X2 U14969 ( .A1(n16376), .A2(n15200), .ZN(n16239) );
  AOI22_X1 U14970 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13334) );
  AOI22_X1 U14971 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11159), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13333) );
  AND2_X2 U14972 ( .A1(n13327), .A2(n16249), .ZN(n16241) );
  AOI22_X1 U14973 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U14974 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13331) );
  NAND4_X1 U14975 ( .A1(n13334), .A2(n13333), .A3(n13332), .A4(n13331), .ZN(
        n13335) );
  INV_X1 U14976 ( .A(n14190), .ZN(n13437) );
  INV_X1 U14977 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n13343) );
  INV_X1 U14978 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13340) );
  NAND2_X1 U14979 ( .A1(n13338), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n13339) );
  OAI211_X1 U14980 ( .C1(n20178), .C2(n13340), .A(n13339), .B(n19876), .ZN(
        n13341) );
  INV_X1 U14981 ( .A(n13341), .ZN(n13342) );
  AOI22_X1 U14982 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U14983 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13347) );
  INV_X1 U14984 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14751) );
  AOI22_X1 U14985 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U14986 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13345) );
  NAND4_X1 U14987 ( .A1(n13348), .A2(n13347), .A3(n13346), .A4(n13345), .ZN(
        n13354) );
  AOI22_X1 U14988 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13352) );
  AOI22_X1 U14989 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11159), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13351) );
  AOI22_X1 U14990 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U14991 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13349) );
  NAND4_X1 U14992 ( .A1(n13352), .A2(n13351), .A3(n13350), .A4(n13349), .ZN(
        n13353) );
  INV_X1 U14993 ( .A(n14264), .ZN(n13360) );
  AND2_X1 U14994 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13356) );
  NOR2_X1 U14995 ( .A1(n13355), .A2(n13356), .ZN(n13359) );
  NAND2_X1 U14996 ( .A1(n13357), .A2(n13358), .ZN(n13389) );
  AOI22_X1 U14997 ( .A1(n13357), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13355), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13362) );
  NAND2_X1 U14998 ( .A1(n13362), .A2(n13361), .ZN(n13380) );
  INV_X1 U14999 ( .A(n13380), .ZN(n13363) );
  AOI22_X1 U15000 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16234), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U15001 ( .A1(n16239), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13366) );
  AOI22_X1 U15002 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16194), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U15003 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13364) );
  NAND4_X1 U15004 ( .A1(n13367), .A2(n13366), .A3(n13365), .A4(n13364), .ZN(
        n13375) );
  AOI22_X1 U15005 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16240), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13373) );
  AOI22_X1 U15006 ( .A1(n16242), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13372) );
  AOI22_X1 U15007 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13371) );
  AOI22_X1 U15008 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13370) );
  NAND4_X1 U15009 ( .A1(n13373), .A2(n13372), .A3(n13371), .A4(n13370), .ZN(
        n13374) );
  OR2_X1 U15010 ( .A1(n14133), .A2(n13572), .ZN(n13378) );
  NAND2_X1 U15011 ( .A1(n13110), .A2(n14710), .ZN(n13376) );
  MUX2_X1 U15012 ( .A(n13376), .B(n19889), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13377) );
  NAND2_X1 U15013 ( .A1(n13378), .A2(n13377), .ZN(n14944) );
  INV_X1 U15014 ( .A(n14944), .ZN(n13379) );
  NAND2_X1 U15015 ( .A1(n14943), .A2(n13379), .ZN(n14947) );
  AOI22_X1 U15016 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13383) );
  AOI22_X1 U15017 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13382) );
  AOI22_X1 U15018 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13381) );
  AOI22_X1 U15019 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13387) );
  AOI22_X1 U15020 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16234), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13386) );
  AOI22_X1 U15021 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13385) );
  AOI22_X1 U15022 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13384) );
  NAND4_X1 U15023 ( .A1(n13387), .A2(n13386), .A3(n13385), .A4(n13384), .ZN(
        n13388) );
  INV_X1 U15024 ( .A(n14132), .ZN(n14114) );
  NAND2_X1 U15025 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13390) );
  OAI211_X1 U15026 ( .C1(n13572), .C2(n14114), .A(n13390), .B(n13389), .ZN(
        n13392) );
  INV_X1 U15027 ( .A(n13392), .ZN(n13393) );
  INV_X2 U15028 ( .A(n13469), .ZN(n13595) );
  AOI22_X1 U15029 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13396) );
  NAND2_X1 U15030 ( .A1(n13394), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13395) );
  NAND2_X1 U15031 ( .A1(n13396), .A2(n13395), .ZN(n14826) );
  AOI22_X1 U15032 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13400) );
  AOI22_X1 U15033 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13399) );
  AOI22_X1 U15034 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13398) );
  AOI22_X1 U15035 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13397) );
  NAND4_X1 U15036 ( .A1(n13400), .A2(n13399), .A3(n13398), .A4(n13397), .ZN(
        n13406) );
  AOI22_X1 U15037 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13404) );
  AOI22_X1 U15038 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11159), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U15039 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U15040 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13401) );
  NAND4_X1 U15041 ( .A1(n13404), .A2(n13403), .A3(n13402), .A4(n13401), .ZN(
        n13405) );
  NAND2_X1 U15042 ( .A1(n13534), .A2(n14127), .ZN(n13410) );
  NAND2_X1 U15043 ( .A1(n13394), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13409) );
  AOI22_X1 U15044 ( .A1(n13595), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13408) );
  NAND2_X1 U15045 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13407) );
  NAND4_X1 U15046 ( .A1(n13410), .A2(n13409), .A3(n13408), .A4(n13407), .ZN(
        n15321) );
  AOI22_X1 U15047 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13414) );
  AOI22_X1 U15048 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U15049 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U15050 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13411) );
  NAND4_X1 U15051 ( .A1(n13414), .A2(n13413), .A3(n13412), .A4(n13411), .ZN(
        n13420) );
  AOI22_X1 U15052 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U15053 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11159), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U15054 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U15055 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13415) );
  NAND4_X1 U15056 ( .A1(n13418), .A2(n13417), .A3(n13416), .A4(n13415), .ZN(
        n13419) );
  NAND2_X1 U15057 ( .A1(n13534), .A2(n14140), .ZN(n13423) );
  NAND2_X1 U15058 ( .A1(n13394), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n13422) );
  INV_X2 U15059 ( .A(n13470), .ZN(n13577) );
  AOI22_X1 U15060 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13421) );
  AOI22_X1 U15061 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13427) );
  AOI22_X1 U15062 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13426) );
  AOI22_X1 U15063 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13344), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U15064 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13424) );
  NAND4_X1 U15065 ( .A1(n13427), .A2(n13426), .A3(n13425), .A4(n13424), .ZN(
        n13433) );
  AOI22_X1 U15066 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13431) );
  AOI22_X1 U15067 ( .A1(n11159), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U15068 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16240), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13429) );
  AOI22_X1 U15069 ( .A1(n16242), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13428) );
  NAND4_X1 U15070 ( .A1(n13431), .A2(n13430), .A3(n13429), .A4(n13428), .ZN(
        n13432) );
  INV_X1 U15071 ( .A(n14169), .ZN(n13626) );
  AOI22_X1 U15072 ( .A1(n13534), .A2(n13626), .B1(n13394), .B2(
        P2_REIP_REG_5__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U15073 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U15074 ( .A1(n13435), .A2(n13434), .ZN(n15748) );
  AOI21_X1 U15075 ( .B1(n13534), .B2(n13437), .A(n13436), .ZN(n17621) );
  AOI222_X1 U15076 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n13394), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n13577), .C1(
        P2_EAX_REG_6__SCAN_IN), .C2(n13595), .ZN(n17620) );
  NAND2_X1 U15077 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13441) );
  NAND2_X1 U15078 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13440) );
  NAND2_X1 U15079 ( .A1(n16232), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13439) );
  NAND2_X1 U15080 ( .A1(n16211), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n13438) );
  NAND4_X1 U15081 ( .A1(n13441), .A2(n13440), .A3(n13439), .A4(n13438), .ZN(
        n13455) );
  INV_X1 U15082 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13445) );
  INV_X1 U15083 ( .A(n13442), .ZN(n13444) );
  INV_X1 U15084 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16393) );
  OAI22_X1 U15085 ( .A1(n13445), .A2(n13444), .B1(n13443), .B2(n16393), .ZN(
        n13453) );
  INV_X1 U15086 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13451) );
  INV_X1 U15087 ( .A(n13446), .ZN(n13450) );
  INV_X1 U15088 ( .A(n13447), .ZN(n13449) );
  INV_X1 U15089 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13448) );
  OAI22_X1 U15090 ( .A1(n13451), .A2(n13450), .B1(n13449), .B2(n13448), .ZN(
        n13452) );
  OR2_X1 U15091 ( .A1(n13453), .A2(n13452), .ZN(n13454) );
  AOI22_X1 U15092 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n16241), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13459) );
  AOI22_X1 U15093 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n16240), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13458) );
  NAND2_X1 U15094 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13457) );
  NAND2_X1 U15095 ( .A1(n16239), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13456) );
  NAND4_X1 U15096 ( .A1(n13459), .A2(n13458), .A3(n13457), .A4(n13456), .ZN(
        n13466) );
  INV_X1 U15097 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13464) );
  INV_X1 U15098 ( .A(n13460), .ZN(n13463) );
  INV_X1 U15099 ( .A(n11159), .ZN(n13462) );
  INV_X1 U15100 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13461) );
  OAI22_X1 U15101 ( .A1(n13464), .A2(n13463), .B1(n13462), .B2(n13461), .ZN(
        n13465) );
  NOR2_X1 U15102 ( .A1(n13466), .A2(n13465), .ZN(n13467) );
  INV_X1 U15103 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17605) );
  INV_X1 U15104 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19715) );
  INV_X1 U15105 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n18999) );
  OAI222_X1 U15106 ( .A1(n13470), .A2(n17605), .B1(n13469), .B2(n19715), .C1(
        n13532), .C2(n18999), .ZN(n17601) );
  NAND2_X1 U15107 ( .A1(n13394), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U15108 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13482) );
  AOI22_X1 U15109 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13369), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13474) );
  AOI22_X1 U15110 ( .A1(n16232), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13473) );
  AOI22_X1 U15111 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13472) );
  AOI22_X1 U15112 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13471) );
  NAND4_X1 U15113 ( .A1(n13474), .A2(n13473), .A3(n13472), .A4(n13471), .ZN(
        n13480) );
  AOI22_X1 U15114 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13478) );
  AOI22_X1 U15115 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11159), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13477) );
  AOI22_X1 U15116 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16240), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13476) );
  AOI22_X1 U15117 ( .A1(n16242), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13475) );
  NAND4_X1 U15118 ( .A1(n13478), .A2(n13477), .A3(n13476), .A4(n13475), .ZN(
        n13479) );
  NOR2_X1 U15119 ( .A1(n13480), .A2(n13479), .ZN(n15342) );
  OR2_X1 U15120 ( .A1(n13572), .A2(n15342), .ZN(n13481) );
  AOI22_X1 U15121 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13487) );
  AOI22_X1 U15122 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13486) );
  AOI22_X1 U15123 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13485) );
  AOI22_X1 U15124 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13484) );
  NAND4_X1 U15125 ( .A1(n13487), .A2(n13486), .A3(n13485), .A4(n13484), .ZN(
        n13493) );
  AOI22_X1 U15126 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13491) );
  AOI22_X1 U15127 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16234), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13490) );
  AOI22_X1 U15128 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13489) );
  AOI22_X1 U15129 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13488) );
  NAND4_X1 U15130 ( .A1(n13491), .A2(n13490), .A3(n13489), .A4(n13488), .ZN(
        n13492) );
  OR2_X1 U15131 ( .A1(n13493), .A2(n13492), .ZN(n15181) );
  AOI22_X1 U15132 ( .A1(n13534), .A2(n15181), .B1(n13394), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n13495) );
  AOI22_X1 U15133 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13494) );
  NAND2_X1 U15134 ( .A1(n13495), .A2(n13494), .ZN(n17558) );
  AOI22_X1 U15135 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13499) );
  AOI22_X1 U15136 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13498) );
  AOI22_X1 U15137 ( .A1(n11159), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13344), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13497) );
  AOI22_X1 U15138 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13496) );
  NAND4_X1 U15139 ( .A1(n13499), .A2(n13498), .A3(n13497), .A4(n13496), .ZN(
        n13505) );
  AOI22_X1 U15140 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13503) );
  AOI22_X1 U15141 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13502) );
  AOI22_X1 U15142 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16240), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13501) );
  AOI22_X1 U15143 ( .A1(n16242), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13500) );
  NAND4_X1 U15144 ( .A1(n13503), .A2(n13502), .A3(n13501), .A4(n13500), .ZN(
        n13504) );
  OR2_X1 U15145 ( .A1(n13505), .A2(n13504), .ZN(n15183) );
  INV_X1 U15146 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U15147 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n13506) );
  OAI21_X1 U15148 ( .B1(n13532), .B2(n17308), .A(n13506), .ZN(n13507) );
  AOI21_X1 U15149 ( .B1(n13534), .B2(n15183), .A(n13507), .ZN(n15813) );
  AOI22_X1 U15150 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13511) );
  AOI22_X1 U15151 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13510) );
  AOI22_X1 U15152 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13509) );
  AOI22_X1 U15153 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13508) );
  NAND4_X1 U15154 ( .A1(n13511), .A2(n13510), .A3(n13509), .A4(n13508), .ZN(
        n13517) );
  AOI22_X1 U15155 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13515) );
  AOI22_X1 U15156 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16234), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13514) );
  AOI22_X1 U15157 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13513) );
  AOI22_X1 U15158 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13512) );
  NAND4_X1 U15159 ( .A1(n13515), .A2(n13514), .A3(n13513), .A4(n13512), .ZN(
        n13516) );
  OR2_X1 U15160 ( .A1(n13517), .A2(n13516), .ZN(n15339) );
  AOI22_X1 U15161 ( .A1(n13534), .A2(n15339), .B1(n13394), .B2(
        P2_REIP_REG_11__SCAN_IN), .ZN(n13519) );
  AOI22_X1 U15162 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13518) );
  NAND2_X1 U15163 ( .A1(n13519), .A2(n13518), .ZN(n15908) );
  AOI22_X1 U15164 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13523) );
  AOI22_X1 U15165 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13522) );
  AOI22_X1 U15166 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13521) );
  AOI22_X1 U15167 ( .A1(n11159), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13344), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13520) );
  NAND4_X1 U15168 ( .A1(n13523), .A2(n13522), .A3(n13521), .A4(n13520), .ZN(
        n13529) );
  AOI22_X1 U15169 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U15170 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13526) );
  AOI22_X1 U15171 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16240), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13525) );
  AOI22_X1 U15172 ( .A1(n16242), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13524) );
  NAND4_X1 U15173 ( .A1(n13527), .A2(n13526), .A3(n13525), .A4(n13524), .ZN(
        n13528) );
  OR2_X1 U15174 ( .A1(n13529), .A2(n13528), .ZN(n15348) );
  AOI22_X1 U15175 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n13530) );
  OAI21_X1 U15176 ( .B1(n13532), .B2(n13531), .A(n13530), .ZN(n13533) );
  AOI21_X1 U15177 ( .B1(n13534), .B2(n15348), .A(n13533), .ZN(n15924) );
  AOI22_X1 U15178 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13538) );
  AOI22_X1 U15179 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13537) );
  AOI22_X1 U15180 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13536) );
  AOI22_X1 U15181 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13535) );
  NAND4_X1 U15182 ( .A1(n13538), .A2(n13537), .A3(n13536), .A4(n13535), .ZN(
        n13544) );
  AOI22_X1 U15183 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13542) );
  AOI22_X1 U15184 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16234), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U15185 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13540) );
  AOI22_X1 U15186 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13539) );
  NAND4_X1 U15187 ( .A1(n13542), .A2(n13541), .A3(n13540), .A4(n13539), .ZN(
        n13543) );
  OR2_X1 U15188 ( .A1(n13544), .A2(n13543), .ZN(n15443) );
  INV_X1 U15189 ( .A(n15443), .ZN(n13547) );
  AOI22_X1 U15190 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13546) );
  NAND2_X1 U15191 ( .A1(n13394), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n13545) );
  OAI211_X1 U15192 ( .C1(n13547), .C2(n13572), .A(n13546), .B(n13545), .ZN(
        n17509) );
  AOI22_X1 U15193 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13551) );
  AOI22_X1 U15194 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13550) );
  AOI22_X1 U15195 ( .A1(n13442), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13549) );
  AOI22_X1 U15196 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13344), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13548) );
  NAND4_X1 U15197 ( .A1(n13551), .A2(n13550), .A3(n13549), .A4(n13548), .ZN(
        n13557) );
  AOI22_X1 U15198 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13555) );
  AOI22_X1 U15199 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11159), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13554) );
  AOI22_X1 U15200 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16240), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13553) );
  AOI22_X1 U15201 ( .A1(n16242), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13552) );
  NAND4_X1 U15202 ( .A1(n13555), .A2(n13554), .A3(n13553), .A4(n13552), .ZN(
        n13556) );
  NOR2_X1 U15203 ( .A1(n13557), .A2(n13556), .ZN(n15420) );
  AOI22_X1 U15204 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n13559) );
  NAND2_X1 U15205 ( .A1(n13394), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n13558) );
  OAI211_X1 U15206 ( .C1(n15420), .C2(n13572), .A(n13559), .B(n13558), .ZN(
        n15805) );
  AOI22_X1 U15207 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n16232), .B1(
        n13369), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13563) );
  AOI22_X1 U15208 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13562) );
  AOI22_X1 U15209 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n13344), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13561) );
  AOI22_X1 U15210 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13560) );
  NAND4_X1 U15211 ( .A1(n13563), .A2(n13562), .A3(n13561), .A4(n13560), .ZN(
        n13569) );
  AOI22_X1 U15212 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U15213 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11159), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13566) );
  AOI22_X1 U15214 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n16242), .B1(
        n16241), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13565) );
  AOI22_X1 U15215 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13368), .B1(
        n16240), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13564) );
  NAND4_X1 U15216 ( .A1(n13567), .A2(n13566), .A3(n13565), .A4(n13564), .ZN(
        n13568) );
  NOR2_X1 U15217 ( .A1(n13569), .A2(n13568), .ZN(n15705) );
  AOI22_X1 U15218 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n13571) );
  NAND2_X1 U15219 ( .A1(n13394), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n13570) );
  OAI211_X1 U15220 ( .C1(n15705), .C2(n13572), .A(n13571), .B(n13570), .ZN(
        n17475) );
  NAND2_X1 U15221 ( .A1(n15803), .A2(n17475), .ZN(n15787) );
  NAND2_X1 U15222 ( .A1(n13394), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n13574) );
  AOI22_X1 U15223 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13573) );
  AND2_X1 U15224 ( .A1(n13574), .A2(n13573), .ZN(n15788) );
  NAND2_X1 U15225 ( .A1(n13394), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n13576) );
  AOI22_X1 U15226 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13575) );
  AND2_X1 U15227 ( .A1(n13576), .A2(n13575), .ZN(n15850) );
  AOI22_X1 U15228 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13579) );
  NAND2_X1 U15229 ( .A1(n13394), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n13578) );
  NAND2_X1 U15230 ( .A1(n13579), .A2(n13578), .ZN(n14393) );
  NAND2_X1 U15231 ( .A1(n13394), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n13581) );
  AOI22_X1 U15232 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13580) );
  AND2_X1 U15233 ( .A1(n13581), .A2(n13580), .ZN(n17118) );
  NAND2_X1 U15234 ( .A1(n13394), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n13584) );
  AOI22_X1 U15235 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13583) );
  AND2_X1 U15236 ( .A1(n13584), .A2(n13583), .ZN(n14486) );
  AOI22_X1 U15237 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13586) );
  NAND2_X1 U15238 ( .A1(n13394), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n13585) );
  NAND2_X1 U15239 ( .A1(n13586), .A2(n13585), .ZN(n17111) );
  AOI22_X1 U15240 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13588) );
  NAND2_X1 U15241 ( .A1(n13394), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n13587) );
  NAND2_X1 U15242 ( .A1(n13588), .A2(n13587), .ZN(n17410) );
  NAND2_X1 U15243 ( .A1(n13394), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n13590) );
  AOI22_X1 U15244 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13589) );
  AND2_X1 U15245 ( .A1(n13590), .A2(n13589), .ZN(n17099) );
  NAND2_X1 U15246 ( .A1(n13394), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U15247 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n13593) );
  AND2_X1 U15248 ( .A1(n13594), .A2(n13593), .ZN(n17091) );
  AOI22_X1 U15249 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13597) );
  NAND2_X1 U15250 ( .A1(n13394), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n13596) );
  NAND2_X1 U15251 ( .A1(n13597), .A2(n13596), .ZN(n16928) );
  AOI22_X1 U15252 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n13599) );
  NAND2_X1 U15253 ( .A1(n13394), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n13598) );
  NAND2_X1 U15254 ( .A1(n13599), .A2(n13598), .ZN(n17077) );
  NAND2_X1 U15255 ( .A1(n13394), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n13601) );
  AOI22_X1 U15256 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n13600) );
  AND2_X1 U15257 ( .A1(n13601), .A2(n13600), .ZN(n17065) );
  NAND2_X1 U15258 ( .A1(n13394), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n13603) );
  AOI22_X1 U15259 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n13602) );
  AND2_X1 U15260 ( .A1(n13603), .A2(n13602), .ZN(n17058) );
  NAND2_X1 U15261 ( .A1(n13394), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n13605) );
  AOI22_X1 U15262 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n13604) );
  AND2_X1 U15263 ( .A1(n13605), .A2(n13604), .ZN(n14447) );
  AOI22_X1 U15264 ( .A1(n13577), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n13595), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n13607) );
  NAND2_X1 U15265 ( .A1(n13394), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13606) );
  NAND2_X1 U15266 ( .A1(n13607), .A2(n13606), .ZN(n13608) );
  AOI22_X1 U15267 ( .A1(n16414), .A2(n19131), .B1(n19118), .B2(n16115), .ZN(
        n13647) );
  NAND2_X1 U15268 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17690), .ZN(n19204) );
  NOR3_X1 U15269 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19876), .A3(n19204), 
        .ZN(n19207) );
  NOR2_X2 U15270 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19880) );
  AND2_X1 U15271 ( .A1(n13609), .A2(n19880), .ZN(n19040) );
  OR2_X1 U15272 ( .A1(n19047), .A2(n19167), .ZN(n13610) );
  OR2_X1 U15273 ( .A1(n19207), .A2(n13610), .ZN(n13611) );
  NAND2_X1 U15274 ( .A1(n19111), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19037) );
  INV_X2 U15275 ( .A(n19037), .ZN(n19159) );
  NAND2_X1 U15276 ( .A1(n14383), .A2(n18966), .ZN(n13612) );
  INV_X1 U15277 ( .A(n13613), .ZN(n13614) );
  NAND2_X1 U15278 ( .A1(n14682), .A2(n13614), .ZN(n16915) );
  INV_X1 U15279 ( .A(n14599), .ZN(n14600) );
  NOR2_X1 U15280 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13642), .ZN(n13615) );
  NAND2_X1 U15281 ( .A1(n14600), .A2(n13615), .ZN(n13616) );
  NAND2_X1 U15282 ( .A1(n16915), .A2(n13616), .ZN(n19158) );
  AOI22_X1 U15283 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19159), .B1(
        P2_EBX_REG_30__SCAN_IN), .B2(n19158), .ZN(n13646) );
  NAND2_X1 U15284 ( .A1(n13617), .A2(n16969), .ZN(n13618) );
  MUX2_X1 U15285 ( .A(n13618), .B(n14133), .S(n16136), .Z(n14298) );
  NAND2_X1 U15286 ( .A1(n13619), .A2(n14223), .ZN(n14217) );
  NAND2_X1 U15287 ( .A1(n13620), .A2(n14217), .ZN(n14265) );
  MUX2_X1 U15288 ( .A(n14265), .B(n13621), .S(n19982), .Z(n13622) );
  MUX2_X1 U15289 ( .A(n14127), .B(n14234), .S(n13619), .Z(n14214) );
  MUX2_X1 U15290 ( .A(n14214), .B(n13623), .S(n19982), .Z(n14290) );
  MUX2_X1 U15291 ( .A(n14212), .B(n14140), .S(n13624), .Z(n14215) );
  MUX2_X1 U15292 ( .A(n13625), .B(n14215), .S(n16136), .Z(n14300) );
  MUX2_X1 U15293 ( .A(n18972), .B(n13626), .S(n16136), .Z(n14282) );
  MUX2_X1 U15294 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n14190), .S(n16136), .Z(
        n14313) );
  INV_X1 U15295 ( .A(n14313), .ZN(n13627) );
  MUX2_X1 U15296 ( .A(n13629), .B(n14287), .S(n16136), .Z(n14322) );
  NAND2_X1 U15297 ( .A1(n19982), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14318) );
  NOR2_X1 U15298 ( .A1(n16136), .A2(n13630), .ZN(n14325) );
  NAND2_X1 U15299 ( .A1(n19982), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14329) );
  NOR2_X1 U15300 ( .A1(n16136), .A2(n13632), .ZN(n14336) );
  NOR2_X1 U15301 ( .A1(n16136), .A2(n13634), .ZN(n14348) );
  NAND2_X1 U15302 ( .A1(n19982), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14345) );
  NAND2_X1 U15303 ( .A1(n19982), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14353) );
  NAND2_X1 U15304 ( .A1(n19982), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n14362) );
  NOR2_X1 U15305 ( .A1(n16136), .A2(n19053), .ZN(n14357) );
  NOR2_X1 U15306 ( .A1(n16136), .A2(n13635), .ZN(n14372) );
  NAND2_X1 U15307 ( .A1(n19982), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14464) );
  AND2_X2 U15308 ( .A1(n14463), .A2(n14464), .ZN(n14468) );
  NAND2_X1 U15309 ( .A1(n19982), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14469) );
  NOR2_X1 U15310 ( .A1(n16136), .A2(n19082), .ZN(n16032) );
  NAND2_X1 U15311 ( .A1(n19982), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16048) );
  NOR2_X1 U15312 ( .A1(n16136), .A2(n19109), .ZN(n16050) );
  NAND2_X1 U15313 ( .A1(n19982), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16055) );
  NOR2_X1 U15314 ( .A1(n16136), .A2(n16931), .ZN(n16064) );
  NOR2_X1 U15315 ( .A1(n16136), .A2(n13637), .ZN(n16058) );
  NOR2_X1 U15316 ( .A1(n16136), .A2(n13638), .ZN(n16068) );
  INV_X1 U15317 ( .A(n16072), .ZN(n13639) );
  NAND2_X1 U15318 ( .A1(n19982), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16071) );
  INV_X1 U15319 ( .A(n14453), .ZN(n13640) );
  NAND2_X1 U15320 ( .A1(n19982), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14452) );
  NAND2_X1 U15321 ( .A1(n13640), .A2(n14452), .ZN(n16135) );
  NAND2_X1 U15322 ( .A1(n19982), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13641) );
  XNOR2_X1 U15323 ( .A(n16135), .B(n13641), .ZN(n16108) );
  INV_X1 U15324 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16975) );
  NOR2_X1 U15325 ( .A1(n16975), .A2(n13642), .ZN(n13643) );
  AOI22_X1 U15326 ( .A1(n16108), .A2(n19156), .B1(n19155), .B2(
        P2_REIP_REG_30__SCAN_IN), .ZN(n13645) );
  NAND2_X1 U15327 ( .A1(n13648), .A2(n11830), .ZN(P2_U2825) );
  NOR2_X1 U15328 ( .A1(n16450), .A2(n20538), .ZN(n13656) );
  XNOR2_X1 U15329 ( .A(n20552), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16670) );
  NAND2_X1 U15330 ( .A1(n22170), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n16822) );
  OAI21_X1 U15331 ( .B1(n20506), .B2(n13653), .A(n16822), .ZN(n13654) );
  INV_X1 U15332 ( .A(keyinput_117), .ZN(n13855) );
  INV_X1 U15333 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n22402) );
  INV_X1 U15334 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n13854) );
  INV_X1 U15335 ( .A(keyinput_116), .ZN(n13853) );
  INV_X1 U15336 ( .A(keyinput_77), .ZN(n13799) );
  AOI22_X1 U15337 ( .A1(n16729), .A2(keyinput_62), .B1(n16533), .B2(
        keyinput_63), .ZN(n13657) );
  OAI221_X1 U15338 ( .B1(n16729), .B2(keyinput_62), .C1(n16533), .C2(
        keyinput_63), .A(n13657), .ZN(n13768) );
  INV_X1 U15339 ( .A(keyinput_61), .ZN(n13766) );
  INV_X1 U15340 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n16526) );
  INV_X1 U15341 ( .A(keyinput_60), .ZN(n13765) );
  INV_X1 U15342 ( .A(keyinput_52), .ZN(n13751) );
  INV_X1 U15343 ( .A(keyinput_48), .ZN(n13748) );
  INV_X1 U15344 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20459) );
  OAI22_X1 U15345 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_43), .B1(
        P1_D_C_N_REG_SCAN_IN), .B2(keyinput_42), .ZN(n13658) );
  AOI221_X1 U15346 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_43), 
        .C1(keyinput_42), .C2(P1_D_C_N_REG_SCAN_IN), .A(n13658), .ZN(n13746)
         );
  INV_X1 U15347 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17749) );
  XNOR2_X1 U15348 ( .A(n17749), .B(keyinput_39), .ZN(n13740) );
  INV_X1 U15349 ( .A(DATAI_3_), .ZN(n13917) );
  INV_X1 U15350 ( .A(keyinput_29), .ZN(n13718) );
  INV_X1 U15351 ( .A(keyinput_18), .ZN(n13659) );
  INV_X1 U15352 ( .A(DATAI_14_), .ZN(n13897) );
  INV_X1 U15353 ( .A(DATAI_19_), .ZN(n16641) );
  INV_X1 U15354 ( .A(keyinput_13), .ZN(n13687) );
  AOI22_X1 U15355 ( .A1(DATAI_25_), .A2(keyinput_7), .B1(DATAI_26_), .B2(
        keyinput_6), .ZN(n13660) );
  OAI221_X1 U15356 ( .B1(DATAI_25_), .B2(keyinput_7), .C1(DATAI_26_), .C2(
        keyinput_6), .A(n13660), .ZN(n13676) );
  NAND2_X1 U15357 ( .A1(n13664), .A2(n13663), .ZN(n13667) );
  INV_X1 U15358 ( .A(keyinput_2), .ZN(n13665) );
  MUX2_X1 U15359 ( .A(n13665), .B(keyinput_2), .S(DATAI_30_), .Z(n13666) );
  NAND2_X1 U15360 ( .A1(n13667), .A2(n13666), .ZN(n13675) );
  XNOR2_X1 U15361 ( .A(n13668), .B(DATAI_28_), .ZN(n13673) );
  XNOR2_X1 U15362 ( .A(DATAI_27_), .B(keyinput_5), .ZN(n13672) );
  INV_X1 U15363 ( .A(DATAI_22_), .ZN(n16629) );
  INV_X1 U15364 ( .A(keyinput_10), .ZN(n13679) );
  XNOR2_X1 U15365 ( .A(DATAI_23_), .B(keyinput_9), .ZN(n13678) );
  XNOR2_X1 U15366 ( .A(DATAI_21_), .B(keyinput_11), .ZN(n13677) );
  OAI211_X1 U15367 ( .C1(n16629), .C2(n13679), .A(n13678), .B(n13677), .ZN(
        n13680) );
  INV_X1 U15368 ( .A(DATAI_20_), .ZN(n22633) );
  INV_X1 U15369 ( .A(keyinput_12), .ZN(n13682) );
  OAI221_X1 U15370 ( .B1(DATAI_19_), .B2(keyinput_13), .C1(n16641), .C2(n13687), .A(n13686), .ZN(n13691) );
  INV_X1 U15371 ( .A(DATAI_18_), .ZN(n22558) );
  INV_X1 U15372 ( .A(keyinput_14), .ZN(n13688) );
  NAND2_X1 U15373 ( .A1(n13691), .A2(n13690), .ZN(n13695) );
  INV_X1 U15374 ( .A(DATAI_16_), .ZN(n22422) );
  OAI22_X1 U15375 ( .A1(n22422), .A2(keyinput_16), .B1(DATAI_17_), .B2(
        keyinput_15), .ZN(n13692) );
  AOI221_X1 U15376 ( .B1(n22422), .B2(keyinput_16), .C1(keyinput_15), .C2(
        DATAI_17_), .A(n13692), .ZN(n13694) );
  AOI21_X1 U15377 ( .B1(n13695), .B2(n13694), .A(n13693), .ZN(n13696) );
  INV_X1 U15378 ( .A(keyinput_19), .ZN(n13697) );
  OR2_X1 U15379 ( .A1(DATAI_13_), .A2(n13697), .ZN(n13699) );
  INV_X1 U15380 ( .A(DATAI_13_), .ZN(n13901) );
  OR2_X1 U15381 ( .A1(n13901), .A2(keyinput_19), .ZN(n13698) );
  NAND3_X1 U15382 ( .A1(n13700), .A2(n13699), .A3(n13698), .ZN(n13704) );
  INV_X1 U15383 ( .A(DATAI_12_), .ZN(n13902) );
  INV_X1 U15384 ( .A(keyinput_20), .ZN(n13701) );
  INV_X1 U15385 ( .A(n13702), .ZN(n13703) );
  NAND2_X1 U15386 ( .A1(n13704), .A2(n13703), .ZN(n13716) );
  OAI22_X1 U15387 ( .A1(DATAI_9_), .A2(keyinput_23), .B1(keyinput_21), .B2(
        DATAI_11_), .ZN(n13705) );
  AOI221_X1 U15388 ( .B1(DATAI_9_), .B2(keyinput_23), .C1(DATAI_11_), .C2(
        keyinput_21), .A(n13705), .ZN(n13709) );
  INV_X1 U15389 ( .A(DATAI_7_), .ZN(n13707) );
  OAI22_X1 U15390 ( .A1(n13707), .A2(keyinput_25), .B1(DATAI_10_), .B2(
        keyinput_22), .ZN(n13706) );
  AOI221_X1 U15391 ( .B1(n13707), .B2(keyinput_25), .C1(keyinput_22), .C2(
        DATAI_10_), .A(n13706), .ZN(n13708) );
  OAI211_X1 U15392 ( .C1(DATAI_8_), .C2(keyinput_24), .A(n13709), .B(n13708), 
        .ZN(n13710) );
  AOI21_X1 U15393 ( .B1(DATAI_8_), .B2(keyinput_24), .A(n13710), .ZN(n13715)
         );
  INV_X1 U15394 ( .A(DATAI_6_), .ZN(n13712) );
  AOI22_X1 U15395 ( .A1(DATAI_4_), .A2(keyinput_28), .B1(n13712), .B2(
        keyinput_26), .ZN(n13711) );
  OAI221_X1 U15396 ( .B1(DATAI_4_), .B2(keyinput_28), .C1(n13712), .C2(
        keyinput_26), .A(n13711), .ZN(n13714) );
  XOR2_X1 U15397 ( .A(DATAI_5_), .B(keyinput_27), .Z(n13713) );
  AOI21_X1 U15398 ( .B1(n13716), .B2(n13715), .A(n11838), .ZN(n13717) );
  AOI221_X1 U15399 ( .B1(DATAI_3_), .B2(keyinput_29), .C1(n13917), .C2(n13718), 
        .A(n13717), .ZN(n13723) );
  INV_X1 U15400 ( .A(DATAI_1_), .ZN(n15147) );
  AOI22_X1 U15401 ( .A1(DATAI_2_), .A2(keyinput_30), .B1(n15147), .B2(
        keyinput_31), .ZN(n13719) );
  OAI221_X1 U15402 ( .B1(DATAI_2_), .B2(keyinput_30), .C1(n15147), .C2(
        keyinput_31), .A(n13719), .ZN(n13722) );
  OAI22_X1 U15403 ( .A1(HOLD), .A2(keyinput_33), .B1(keyinput_32), .B2(
        DATAI_0_), .ZN(n13720) );
  AOI221_X1 U15404 ( .B1(HOLD), .B2(keyinput_33), .C1(DATAI_0_), .C2(
        keyinput_32), .A(n13720), .ZN(n13721) );
  INV_X1 U15405 ( .A(NA), .ZN(n22302) );
  INV_X1 U15406 ( .A(keyinput_34), .ZN(n13724) );
  OR2_X1 U15407 ( .A1(n22302), .A2(n13724), .ZN(n13726) );
  OR2_X1 U15408 ( .A1(NA), .A2(keyinput_34), .ZN(n13725) );
  NAND3_X1 U15409 ( .A1(n13727), .A2(n13726), .A3(n13725), .ZN(n13731) );
  INV_X1 U15410 ( .A(BS16), .ZN(n17708) );
  INV_X1 U15411 ( .A(keyinput_35), .ZN(n13728) );
  INV_X1 U15412 ( .A(n13729), .ZN(n13730) );
  OAI22_X1 U15413 ( .A1(READY1), .A2(keyinput_36), .B1(keyinput_37), .B2(
        READY2), .ZN(n13732) );
  AOI221_X1 U15414 ( .B1(READY1), .B2(keyinput_36), .C1(READY2), .C2(
        keyinput_37), .A(n13732), .ZN(n13735) );
  INV_X1 U15415 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n14596) );
  OAI22_X1 U15416 ( .A1(n14596), .A2(keyinput_40), .B1(P1_M_IO_N_REG_SCAN_IN), 
        .B2(keyinput_41), .ZN(n13737) );
  AOI221_X1 U15417 ( .B1(n14596), .B2(keyinput_40), .C1(keyinput_41), .C2(
        P1_M_IO_N_REG_SCAN_IN), .A(n13737), .ZN(n13738) );
  OAI21_X1 U15418 ( .B1(n13740), .B2(n13739), .A(n13738), .ZN(n13745) );
  INV_X1 U15419 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n22217) );
  INV_X1 U15420 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20628) );
  AOI22_X1 U15421 ( .A1(n22217), .A2(keyinput_46), .B1(n20628), .B2(
        keyinput_47), .ZN(n13741) );
  OAI221_X1 U15422 ( .B1(n22217), .B2(keyinput_46), .C1(n20628), .C2(
        keyinput_47), .A(n13741), .ZN(n13744) );
  AOI22_X1 U15423 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_45), .B1(n21856), 
        .B2(keyinput_44), .ZN(n13742) );
  OAI221_X1 U15424 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_45), .C1(n21856), 
        .C2(keyinput_44), .A(n13742), .ZN(n13743) );
  INV_X1 U15425 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20452) );
  AOI22_X1 U15426 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_49), .B1(
        n20452), .B2(keyinput_50), .ZN(n13749) );
  OAI221_X1 U15427 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_49), .C1(
        n20452), .C2(keyinput_50), .A(n13749), .ZN(n13750) );
  INV_X1 U15428 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n13755) );
  INV_X1 U15429 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n13754) );
  AOI22_X1 U15430 ( .A1(n13755), .A2(keyinput_54), .B1(n13754), .B2(
        keyinput_53), .ZN(n13753) );
  OAI221_X1 U15431 ( .B1(n13755), .B2(keyinput_54), .C1(n13754), .C2(
        keyinput_53), .A(n13753), .ZN(n13758) );
  OAI22_X1 U15432 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput_55), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_56), .ZN(n13756) );
  AOI221_X1 U15433 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_55), .C1(
        keyinput_56), .C2(P1_REIP_REG_27__SCAN_IN), .A(n13756), .ZN(n13757) );
  OAI21_X1 U15434 ( .B1(n13759), .B2(n13758), .A(n13757), .ZN(n13763) );
  INV_X1 U15435 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21976) );
  OAI22_X1 U15436 ( .A1(n21976), .A2(keyinput_57), .B1(keyinput_58), .B2(
        P1_REIP_REG_25__SCAN_IN), .ZN(n13760) );
  AOI221_X1 U15437 ( .B1(n21976), .B2(keyinput_57), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_58), .A(n13760), .ZN(n13762) );
  NOR2_X1 U15438 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_59), .ZN(n13761)
         );
  AOI221_X1 U15439 ( .B1(n13763), .B2(n13762), .C1(keyinput_59), .C2(
        P1_REIP_REG_24__SCAN_IN), .A(n13761), .ZN(n13764) );
  NAND2_X1 U15440 ( .A1(n16548), .A2(keyinput_64), .ZN(n13767) );
  INV_X1 U15441 ( .A(keyinput_65), .ZN(n13769) );
  INV_X1 U15442 ( .A(n13770), .ZN(n13775) );
  INV_X1 U15443 ( .A(keyinput_66), .ZN(n13771) );
  OR2_X1 U15444 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n13771), .ZN(n13773) );
  INV_X1 U15445 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n22158) );
  OR2_X1 U15446 ( .A1(n22158), .A2(keyinput_66), .ZN(n13772) );
  INV_X1 U15447 ( .A(keyinput_67), .ZN(n13776) );
  OR3_X1 U15448 ( .A1(n13777), .A2(n11855), .A3(n11839), .ZN(n13782) );
  OR2_X1 U15449 ( .A1(n22139), .A2(keyinput_68), .ZN(n13780) );
  INV_X1 U15450 ( .A(keyinput_68), .ZN(n13778) );
  OR2_X1 U15451 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n13778), .ZN(n13779) );
  AND2_X1 U15452 ( .A1(n13780), .A2(n13779), .ZN(n13781) );
  INV_X1 U15453 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n16849) );
  INV_X1 U15454 ( .A(keyinput_69), .ZN(n13783) );
  INV_X1 U15455 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n15940) );
  INV_X1 U15456 ( .A(keyinput_70), .ZN(n13785) );
  INV_X1 U15457 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n22113) );
  INV_X1 U15458 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n22114) );
  AOI22_X1 U15459 ( .A1(n16881), .A2(keyinput_73), .B1(n22114), .B2(
        keyinput_72), .ZN(n13788) );
  OAI221_X1 U15460 ( .B1(n16881), .B2(keyinput_73), .C1(n22114), .C2(
        keyinput_72), .A(n13788), .ZN(n13791) );
  AOI22_X1 U15461 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(keyinput_74), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(keyinput_75), .ZN(n13789) );
  OAI221_X1 U15462 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(keyinput_74), .C1(
        P1_REIP_REG_8__SCAN_IN), .C2(keyinput_75), .A(n13789), .ZN(n13790) );
  NOR2_X1 U15463 ( .A1(n13791), .A2(n13790), .ZN(n13796) );
  NAND2_X1 U15464 ( .A1(n22094), .A2(keyinput_76), .ZN(n13794) );
  INV_X1 U15465 ( .A(keyinput_76), .ZN(n13792) );
  AOI21_X1 U15466 ( .B1(n13797), .B2(n13796), .A(n13795), .ZN(n13798) );
  INV_X1 U15467 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n22031) );
  AOI22_X1 U15468 ( .A1(n22031), .A2(keyinput_82), .B1(n16557), .B2(
        keyinput_84), .ZN(n13800) );
  OAI221_X1 U15469 ( .B1(n22031), .B2(keyinput_82), .C1(n16557), .C2(
        keyinput_84), .A(n13800), .ZN(n13805) );
  INV_X1 U15470 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13802) );
  OAI22_X1 U15471 ( .A1(n13802), .A2(keyinput_83), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(keyinput_81), .ZN(n13801) );
  AOI221_X1 U15472 ( .B1(n13802), .B2(keyinput_83), .C1(keyinput_81), .C2(
        P1_REIP_REG_2__SCAN_IN), .A(n13801), .ZN(n13803) );
  OAI21_X1 U15473 ( .B1(keyinput_80), .B2(P1_REIP_REG_3__SCAN_IN), .A(n13803), 
        .ZN(n13804) );
  AOI211_X1 U15474 ( .C1(keyinput_80), .C2(P1_REIP_REG_3__SCAN_IN), .A(n13805), 
        .B(n13804), .ZN(n13810) );
  INV_X1 U15475 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n22071) );
  AOI22_X1 U15476 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(keyinput_79), .B1(n22071), 
        .B2(keyinput_78), .ZN(n13806) );
  OAI221_X1 U15477 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(keyinput_79), .C1(n22071), .C2(keyinput_78), .A(n13806), .ZN(n13809) );
  INV_X1 U15478 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n16564) );
  AOI22_X1 U15479 ( .A1(P1_EBX_REG_28__SCAN_IN), .A2(keyinput_87), .B1(n16564), 
        .B2(keyinput_89), .ZN(n13807) );
  OAI221_X1 U15480 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(keyinput_87), .C1(n16564), .C2(keyinput_89), .A(n13807), .ZN(n13808) );
  AOI22_X1 U15481 ( .A1(n16561), .A2(keyinput_86), .B1(keyinput_85), .B2(
        n16559), .ZN(n13811) );
  OAI221_X1 U15482 ( .B1(n16561), .B2(keyinput_86), .C1(n16559), .C2(
        keyinput_85), .A(n13811), .ZN(n13812) );
  AOI21_X1 U15483 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput_88), .A(n13812), 
        .ZN(n13813) );
  INV_X1 U15484 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n22151) );
  AOI22_X1 U15485 ( .A1(P1_EBX_REG_23__SCAN_IN), .A2(keyinput_92), .B1(n22151), 
        .B2(keyinput_98), .ZN(n13814) );
  OAI221_X1 U15486 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(keyinput_92), .C1(n22151), .C2(keyinput_98), .A(n13814), .ZN(n13821) );
  AOI22_X1 U15487 ( .A1(P1_EBX_REG_18__SCAN_IN), .A2(keyinput_97), .B1(
        P1_EBX_REG_25__SCAN_IN), .B2(keyinput_90), .ZN(n13815) );
  OAI221_X1 U15488 ( .B1(P1_EBX_REG_18__SCAN_IN), .B2(keyinput_97), .C1(
        P1_EBX_REG_25__SCAN_IN), .C2(keyinput_90), .A(n13815), .ZN(n13820) );
  INV_X1 U15489 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15973) );
  INV_X1 U15490 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n20486) );
  AOI22_X1 U15491 ( .A1(n15973), .A2(keyinput_100), .B1(n20486), .B2(
        keyinput_95), .ZN(n13816) );
  OAI221_X1 U15492 ( .B1(n15973), .B2(keyinput_100), .C1(n20486), .C2(
        keyinput_95), .A(n13816), .ZN(n13819) );
  INV_X1 U15493 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n22142) );
  INV_X1 U15494 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n16579) );
  AOI22_X1 U15495 ( .A1(n22142), .A2(keyinput_99), .B1(n16579), .B2(
        keyinput_96), .ZN(n13817) );
  OAI221_X1 U15496 ( .B1(n22142), .B2(keyinput_99), .C1(n16579), .C2(
        keyinput_96), .A(n13817), .ZN(n13818) );
  NOR4_X1 U15497 ( .A1(n13821), .A2(n13820), .A3(n13819), .A4(n13818), .ZN(
        n13824) );
  INV_X1 U15498 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n20475) );
  INV_X1 U15499 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n22180) );
  OAI22_X1 U15500 ( .A1(n20475), .A2(keyinput_93), .B1(n22180), .B2(
        keyinput_94), .ZN(n13822) );
  AOI221_X1 U15501 ( .B1(n20475), .B2(keyinput_93), .C1(keyinput_94), .C2(
        n22180), .A(n13822), .ZN(n13823) );
  OAI211_X1 U15502 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(keyinput_91), .A(n13824), 
        .B(n13823), .ZN(n13825) );
  AOI21_X1 U15503 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(keyinput_91), .A(n13825), 
        .ZN(n13826) );
  AOI22_X1 U15504 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(keyinput_103), .B1(
        P1_EBX_REG_13__SCAN_IN), .B2(keyinput_102), .ZN(n13827) );
  OAI221_X1 U15505 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(keyinput_103), .C1(
        P1_EBX_REG_13__SCAN_IN), .C2(keyinput_102), .A(n13827), .ZN(n13829) );
  INV_X1 U15506 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n22122) );
  NAND2_X1 U15507 ( .A1(n13831), .A2(n13830), .ZN(n13837) );
  INV_X1 U15508 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15884) );
  INV_X1 U15509 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n20492) );
  OAI22_X1 U15510 ( .A1(n15884), .A2(keyinput_104), .B1(n20492), .B2(
        keyinput_107), .ZN(n13832) );
  AOI221_X1 U15511 ( .B1(n15884), .B2(keyinput_104), .C1(keyinput_107), .C2(
        n20492), .A(n13832), .ZN(n13835) );
  INV_X1 U15512 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15674) );
  OAI22_X1 U15513 ( .A1(n15674), .A2(keyinput_106), .B1(keyinput_108), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n13833) );
  AOI221_X1 U15514 ( .B1(n15674), .B2(keyinput_106), .C1(P1_EBX_REG_7__SCAN_IN), .C2(keyinput_108), .A(n13833), .ZN(n13834) );
  AND2_X1 U15515 ( .A1(n13835), .A2(n13834), .ZN(n13836) );
  NAND2_X1 U15516 ( .A1(n13837), .A2(n13836), .ZN(n13842) );
  INV_X1 U15517 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n22079) );
  INV_X1 U15518 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15725) );
  AOI22_X1 U15519 ( .A1(n22079), .A2(keyinput_109), .B1(n15725), .B2(
        keyinput_105), .ZN(n13838) );
  OAI221_X1 U15520 ( .B1(n22079), .B2(keyinput_109), .C1(n15725), .C2(
        keyinput_105), .A(n13838), .ZN(n13841) );
  OAI21_X1 U15521 ( .B1(n13842), .B2(n13841), .A(n13840), .ZN(n13848) );
  INV_X1 U15522 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n22064) );
  AOI22_X1 U15523 ( .A1(n22064), .A2(keyinput_111), .B1(keyinput_114), .B2(
        n11742), .ZN(n13843) );
  OAI221_X1 U15524 ( .B1(n22064), .B2(keyinput_111), .C1(n11742), .C2(
        keyinput_114), .A(n13843), .ZN(n13844) );
  INV_X1 U15525 ( .A(n13844), .ZN(n13847) );
  INV_X1 U15526 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n22038) );
  INV_X1 U15527 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n20465) );
  OAI22_X1 U15528 ( .A1(n22038), .A2(keyinput_112), .B1(n20465), .B2(
        keyinput_113), .ZN(n13845) );
  AOI221_X1 U15529 ( .B1(n22038), .B2(keyinput_112), .C1(keyinput_113), .C2(
        n20465), .A(n13845), .ZN(n13846) );
  NAND3_X1 U15530 ( .A1(n13848), .A2(n13847), .A3(n13846), .ZN(n13852) );
  INV_X1 U15531 ( .A(keyinput_115), .ZN(n13850) );
  INV_X1 U15532 ( .A(n13856), .ZN(n13860) );
  INV_X1 U15533 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n22385) );
  INV_X1 U15534 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n22393) );
  AOI22_X1 U15535 ( .A1(n22385), .A2(keyinput_119), .B1(n22393), .B2(
        keyinput_118), .ZN(n13857) );
  OAI221_X1 U15536 ( .B1(n22385), .B2(keyinput_119), .C1(n22393), .C2(
        keyinput_118), .A(n13857), .ZN(n13858) );
  INV_X1 U15537 ( .A(n13858), .ZN(n13859) );
  NAND2_X1 U15538 ( .A1(n13860), .A2(n13859), .ZN(n13865) );
  OAI22_X1 U15539 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(keyinput_120), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(keyinput_121), .ZN(n13861) );
  AOI221_X1 U15540 ( .B1(P1_EAX_REG_27__SCAN_IN), .B2(keyinput_120), .C1(
        keyinput_121), .C2(P1_EAX_REG_26__SCAN_IN), .A(n13861), .ZN(n13864) );
  AOI22_X1 U15541 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_123), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(keyinput_122), .ZN(n13862) );
  OAI221_X1 U15542 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_123), .C1(
        P1_EAX_REG_25__SCAN_IN), .C2(keyinput_122), .A(n13862), .ZN(n13863) );
  AOI21_X1 U15543 ( .B1(n13865), .B2(n13864), .A(n13863), .ZN(n13873) );
  INV_X1 U15544 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n22354) );
  AOI22_X1 U15545 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(keyinput_125), .B1(n22354), .B2(keyinput_124), .ZN(n13867) );
  OR2_X1 U15546 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(keyinput_125), .ZN(n13866)
         );
  OAI211_X1 U15547 ( .C1(n22354), .C2(keyinput_124), .A(n13867), .B(n13866), 
        .ZN(n13872) );
  INV_X1 U15548 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n22336) );
  OAI22_X1 U15549 ( .A1(n22336), .A2(keyinput_127), .B1(keyinput_126), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n13870) );
  INV_X1 U15550 ( .A(keyinput_127), .ZN(n13868) );
  NOR2_X1 U15551 ( .A1(n13868), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n13869) );
  AOI211_X1 U15552 ( .C1(P1_EAX_REG_21__SCAN_IN), .C2(keyinput_126), .A(n13870), .B(n13869), .ZN(n13871) );
  OAI21_X1 U15553 ( .B1(n13873), .B2(n13872), .A(n13871), .ZN(n14060) );
  XNOR2_X1 U15554 ( .A(keyinput_128), .B(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(
        n13876) );
  XNOR2_X1 U15555 ( .A(DATAI_31_), .B(keyinput_129), .ZN(n13875) );
  XNOR2_X1 U15556 ( .A(DATAI_30_), .B(keyinput_130), .ZN(n13874) );
  OAI21_X1 U15557 ( .B1(n13876), .B2(n13875), .A(n13874), .ZN(n13880) );
  XOR2_X1 U15558 ( .A(DATAI_28_), .B(keyinput_132), .Z(n13879) );
  XNOR2_X1 U15559 ( .A(DATAI_27_), .B(keyinput_133), .ZN(n13878) );
  XNOR2_X1 U15560 ( .A(DATAI_29_), .B(keyinput_131), .ZN(n13877) );
  NAND4_X1 U15561 ( .A1(n13880), .A2(n13879), .A3(n13878), .A4(n13877), .ZN(
        n13883) );
  XOR2_X1 U15562 ( .A(DATAI_26_), .B(keyinput_134), .Z(n13882) );
  XNOR2_X1 U15563 ( .A(DATAI_25_), .B(keyinput_135), .ZN(n13881) );
  NAND3_X1 U15564 ( .A1(n13883), .A2(n13882), .A3(n13881), .ZN(n13889) );
  XOR2_X1 U15565 ( .A(DATAI_24_), .B(keyinput_136), .Z(n13888) );
  XNOR2_X1 U15566 ( .A(keyinput_138), .B(DATAI_22_), .ZN(n13886) );
  XNOR2_X1 U15567 ( .A(keyinput_139), .B(DATAI_21_), .ZN(n13885) );
  XNOR2_X1 U15568 ( .A(keyinput_137), .B(DATAI_23_), .ZN(n13884) );
  NAND3_X1 U15569 ( .A1(n13886), .A2(n13885), .A3(n13884), .ZN(n13887) );
  AOI21_X1 U15570 ( .B1(n13889), .B2(n13888), .A(n13887), .ZN(n13892) );
  XNOR2_X1 U15571 ( .A(keyinput_140), .B(DATAI_20_), .ZN(n13891) );
  XNOR2_X1 U15572 ( .A(keyinput_141), .B(DATAI_19_), .ZN(n13890) );
  OAI21_X1 U15573 ( .B1(n13892), .B2(n13891), .A(n13890), .ZN(n13896) );
  XOR2_X1 U15574 ( .A(keyinput_142), .B(DATAI_18_), .Z(n13895) );
  XNOR2_X1 U15575 ( .A(DATAI_17_), .B(keyinput_143), .ZN(n13894) );
  XNOR2_X1 U15576 ( .A(DATAI_16_), .B(keyinput_144), .ZN(n13893) );
  AOI211_X1 U15577 ( .C1(n13896), .C2(n13895), .A(n13894), .B(n13893), .ZN(
        n13900) );
  XOR2_X1 U15578 ( .A(DATAI_15_), .B(keyinput_145), .Z(n13899) );
  XNOR2_X1 U15579 ( .A(n13897), .B(keyinput_146), .ZN(n13898) );
  OAI21_X1 U15580 ( .B1(n13900), .B2(n13899), .A(n13898), .ZN(n13905) );
  XNOR2_X1 U15581 ( .A(n13901), .B(keyinput_147), .ZN(n13904) );
  XNOR2_X1 U15582 ( .A(n13902), .B(keyinput_148), .ZN(n13903) );
  AOI21_X1 U15583 ( .B1(n13905), .B2(n13904), .A(n13903), .ZN(n13912) );
  INV_X1 U15584 ( .A(DATAI_10_), .ZN(n13907) );
  AOI22_X1 U15585 ( .A1(DATAI_7_), .A2(keyinput_153), .B1(n13907), .B2(
        keyinput_150), .ZN(n13906) );
  OAI221_X1 U15586 ( .B1(DATAI_7_), .B2(keyinput_153), .C1(n13907), .C2(
        keyinput_150), .A(n13906), .ZN(n13911) );
  AOI22_X1 U15587 ( .A1(DATAI_11_), .A2(keyinput_149), .B1(DATAI_8_), .B2(
        keyinput_152), .ZN(n13908) );
  OAI221_X1 U15588 ( .B1(DATAI_11_), .B2(keyinput_149), .C1(DATAI_8_), .C2(
        keyinput_152), .A(n13908), .ZN(n13910) );
  XNOR2_X1 U15589 ( .A(DATAI_9_), .B(keyinput_151), .ZN(n13909) );
  NOR4_X1 U15590 ( .A1(n13912), .A2(n13911), .A3(n13910), .A4(n13909), .ZN(
        n13916) );
  XOR2_X1 U15591 ( .A(keyinput_154), .B(DATAI_6_), .Z(n13915) );
  XNOR2_X1 U15592 ( .A(DATAI_4_), .B(keyinput_156), .ZN(n13914) );
  XNOR2_X1 U15593 ( .A(DATAI_5_), .B(keyinput_155), .ZN(n13913) );
  NOR4_X1 U15594 ( .A1(n13916), .A2(n13915), .A3(n13914), .A4(n13913), .ZN(
        n13921) );
  XNOR2_X1 U15595 ( .A(n13917), .B(keyinput_157), .ZN(n13920) );
  XOR2_X1 U15596 ( .A(DATAI_1_), .B(keyinput_159), .Z(n13919) );
  XNOR2_X1 U15597 ( .A(keyinput_158), .B(DATAI_2_), .ZN(n13918) );
  OAI211_X1 U15598 ( .C1(n13921), .C2(n13920), .A(n13919), .B(n13918), .ZN(
        n13924) );
  XOR2_X1 U15599 ( .A(DATAI_0_), .B(keyinput_160), .Z(n13923) );
  XOR2_X1 U15600 ( .A(HOLD), .B(keyinput_161), .Z(n13922) );
  NAND3_X1 U15601 ( .A1(n13924), .A2(n13923), .A3(n13922), .ZN(n13927) );
  XNOR2_X1 U15602 ( .A(keyinput_162), .B(NA), .ZN(n13926) );
  XNOR2_X1 U15603 ( .A(keyinput_163), .B(BS16), .ZN(n13925) );
  AOI21_X1 U15604 ( .B1(n13927), .B2(n13926), .A(n13925), .ZN(n13931) );
  XOR2_X1 U15605 ( .A(READY2), .B(keyinput_165), .Z(n13930) );
  XOR2_X1 U15606 ( .A(keyinput_166), .B(P1_READREQUEST_REG_SCAN_IN), .Z(n13929) );
  XNOR2_X1 U15607 ( .A(READY1), .B(keyinput_164), .ZN(n13928) );
  NOR4_X1 U15608 ( .A1(n13931), .A2(n13930), .A3(n13929), .A4(n13928), .ZN(
        n13935) );
  XOR2_X1 U15609 ( .A(keyinput_167), .B(P1_ADS_N_REG_SCAN_IN), .Z(n13934) );
  XOR2_X1 U15610 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_169), .Z(n13933) );
  XNOR2_X1 U15611 ( .A(keyinput_168), .B(P1_CODEFETCH_REG_SCAN_IN), .ZN(n13932) );
  OAI211_X1 U15612 ( .C1(n13935), .C2(n13934), .A(n13933), .B(n13932), .ZN(
        n13945) );
  INV_X1 U15613 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20564) );
  XNOR2_X1 U15614 ( .A(n20564), .B(keyinput_170), .ZN(n13937) );
  INV_X1 U15615 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22255) );
  XNOR2_X1 U15616 ( .A(n22255), .B(keyinput_171), .ZN(n13936) );
  NOR2_X1 U15617 ( .A1(n13937), .A2(n13936), .ZN(n13944) );
  INV_X1 U15618 ( .A(keyinput_172), .ZN(n13938) );
  XNOR2_X1 U15619 ( .A(n13938), .B(P1_STATEBS16_REG_SCAN_IN), .ZN(n13942) );
  XNOR2_X1 U15620 ( .A(keyinput_174), .B(P1_FLUSH_REG_SCAN_IN), .ZN(n13941) );
  XNOR2_X1 U15621 ( .A(keyinput_173), .B(P1_MORE_REG_SCAN_IN), .ZN(n13940) );
  XNOR2_X1 U15622 ( .A(keyinput_175), .B(P1_W_R_N_REG_SCAN_IN), .ZN(n13939) );
  NAND4_X1 U15623 ( .A1(n13942), .A2(n13941), .A3(n13940), .A4(n13939), .ZN(
        n13943) );
  AOI21_X1 U15624 ( .B1(n13945), .B2(n13944), .A(n13943), .ZN(n13949) );
  XOR2_X1 U15625 ( .A(keyinput_176), .B(P1_BYTEENABLE_REG_0__SCAN_IN), .Z(
        n13948) );
  XOR2_X1 U15626 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_177), .Z(
        n13947) );
  XNOR2_X1 U15627 ( .A(keyinput_178), .B(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(
        n13946) );
  OAI211_X1 U15628 ( .C1(n13949), .C2(n13948), .A(n13947), .B(n13946), .ZN(
        n13952) );
  XNOR2_X1 U15629 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_179), .ZN(
        n13951) );
  XNOR2_X1 U15630 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_180), .ZN(n13950)
         );
  AOI21_X1 U15631 ( .B1(n13952), .B2(n13951), .A(n13950), .ZN(n13955) );
  XOR2_X1 U15632 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_182), .Z(n13954)
         );
  XNOR2_X1 U15633 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_181), .ZN(n13953)
         );
  NOR3_X1 U15634 ( .A1(n13955), .A2(n13954), .A3(n13953), .ZN(n13958) );
  XOR2_X1 U15635 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_183), .Z(n13957)
         );
  XNOR2_X1 U15636 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_184), .ZN(n13956)
         );
  NOR3_X1 U15637 ( .A1(n13958), .A2(n13957), .A3(n13956), .ZN(n13961) );
  XOR2_X1 U15638 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_185), .Z(n13960)
         );
  XNOR2_X1 U15639 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_186), .ZN(n13959)
         );
  NOR3_X1 U15640 ( .A1(n13961), .A2(n13960), .A3(n13959), .ZN(n13964) );
  XNOR2_X1 U15641 ( .A(P1_REIP_REG_24__SCAN_IN), .B(keyinput_187), .ZN(n13963)
         );
  XNOR2_X1 U15642 ( .A(keyinput_188), .B(P1_REIP_REG_23__SCAN_IN), .ZN(n13962)
         );
  OAI21_X1 U15643 ( .B1(n13964), .B2(n13963), .A(n13962), .ZN(n13968) );
  XNOR2_X1 U15644 ( .A(keyinput_189), .B(P1_REIP_REG_22__SCAN_IN), .ZN(n13967)
         );
  XNOR2_X1 U15645 ( .A(keyinput_190), .B(P1_REIP_REG_21__SCAN_IN), .ZN(n13966)
         );
  XNOR2_X1 U15646 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_191), .ZN(n13965)
         );
  AOI211_X1 U15647 ( .C1(n13968), .C2(n13967), .A(n13966), .B(n13965), .ZN(
        n13971) );
  XNOR2_X1 U15648 ( .A(P1_REIP_REG_19__SCAN_IN), .B(keyinput_192), .ZN(n13970)
         );
  XNOR2_X1 U15649 ( .A(keyinput_193), .B(P1_REIP_REG_18__SCAN_IN), .ZN(n13969)
         );
  OAI21_X1 U15650 ( .B1(n13971), .B2(n13970), .A(n13969), .ZN(n13974) );
  XNOR2_X1 U15651 ( .A(keyinput_194), .B(P1_REIP_REG_17__SCAN_IN), .ZN(n13973)
         );
  XNOR2_X1 U15652 ( .A(keyinput_195), .B(P1_REIP_REG_16__SCAN_IN), .ZN(n13972)
         );
  AOI21_X1 U15653 ( .B1(n13974), .B2(n13973), .A(n13972), .ZN(n13977) );
  XOR2_X1 U15654 ( .A(keyinput_196), .B(P1_REIP_REG_15__SCAN_IN), .Z(n13976)
         );
  XNOR2_X1 U15655 ( .A(keyinput_197), .B(P1_REIP_REG_14__SCAN_IN), .ZN(n13975)
         );
  OAI21_X1 U15656 ( .B1(n13977), .B2(n13976), .A(n13975), .ZN(n13980) );
  XNOR2_X1 U15657 ( .A(keyinput_198), .B(P1_REIP_REG_13__SCAN_IN), .ZN(n13979)
         );
  XOR2_X1 U15658 ( .A(keyinput_199), .B(P1_REIP_REG_12__SCAN_IN), .Z(n13978)
         );
  AOI21_X1 U15659 ( .B1(n13980), .B2(n13979), .A(n13978), .ZN(n13987) );
  XOR2_X1 U15660 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_203), .Z(n13984) );
  XOR2_X1 U15661 ( .A(P1_REIP_REG_11__SCAN_IN), .B(keyinput_200), .Z(n13983)
         );
  XOR2_X1 U15662 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_202), .Z(n13982) );
  XNOR2_X1 U15663 ( .A(keyinput_201), .B(P1_REIP_REG_10__SCAN_IN), .ZN(n13981)
         );
  NAND4_X1 U15664 ( .A1(n13984), .A2(n13983), .A3(n13982), .A4(n13981), .ZN(
        n13986) );
  XNOR2_X1 U15665 ( .A(keyinput_204), .B(P1_REIP_REG_7__SCAN_IN), .ZN(n13985)
         );
  OAI21_X1 U15666 ( .B1(n13987), .B2(n13986), .A(n13985), .ZN(n13991) );
  XOR2_X1 U15667 ( .A(keyinput_205), .B(P1_REIP_REG_6__SCAN_IN), .Z(n13990) );
  XOR2_X1 U15668 ( .A(keyinput_206), .B(P1_REIP_REG_5__SCAN_IN), .Z(n13989) );
  XNOR2_X1 U15669 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_207), .ZN(n13988)
         );
  AOI211_X1 U15670 ( .C1(n13991), .C2(n13990), .A(n13989), .B(n13988), .ZN(
        n13999) );
  XNOR2_X1 U15671 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_210), .ZN(n13998)
         );
  XNOR2_X1 U15672 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_212), .ZN(n13997)
         );
  INV_X1 U15673 ( .A(keyinput_208), .ZN(n13992) );
  XNOR2_X1 U15674 ( .A(n13992), .B(P1_REIP_REG_3__SCAN_IN), .ZN(n13995) );
  XNOR2_X1 U15675 ( .A(keyinput_211), .B(P1_REIP_REG_0__SCAN_IN), .ZN(n13994)
         );
  XNOR2_X1 U15676 ( .A(keyinput_209), .B(P1_REIP_REG_2__SCAN_IN), .ZN(n13993)
         );
  NAND3_X1 U15677 ( .A1(n13995), .A2(n13994), .A3(n13993), .ZN(n13996) );
  NOR4_X1 U15678 ( .A1(n13999), .A2(n13998), .A3(n13997), .A4(n13996), .ZN(
        n14005) );
  AOI22_X1 U15679 ( .A1(n16559), .A2(keyinput_213), .B1(n16564), .B2(
        keyinput_217), .ZN(n14000) );
  OAI221_X1 U15680 ( .B1(n16559), .B2(keyinput_213), .C1(n16564), .C2(
        keyinput_217), .A(n14000), .ZN(n14004) );
  INV_X1 U15681 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n16562) );
  AOI22_X1 U15682 ( .A1(P1_EBX_REG_29__SCAN_IN), .A2(keyinput_214), .B1(n16562), .B2(keyinput_215), .ZN(n14001) );
  OAI221_X1 U15683 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(keyinput_214), .C1(
        n16562), .C2(keyinput_215), .A(n14001), .ZN(n14003) );
  XNOR2_X1 U15684 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_216), .ZN(n14002)
         );
  NOR4_X1 U15685 ( .A1(n14005), .A2(n14004), .A3(n14003), .A4(n14002), .ZN(
        n14018) );
  INV_X1 U15686 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n22198) );
  AOI22_X1 U15687 ( .A1(n22198), .A2(keyinput_220), .B1(keyinput_221), .B2(
        n20475), .ZN(n14006) );
  OAI221_X1 U15688 ( .B1(n22198), .B2(keyinput_220), .C1(n20475), .C2(
        keyinput_221), .A(n14006), .ZN(n14017) );
  INV_X1 U15689 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n16565) );
  AOI22_X1 U15690 ( .A1(n16565), .A2(keyinput_218), .B1(keyinput_223), .B2(
        n20486), .ZN(n14007) );
  OAI221_X1 U15691 ( .B1(n16565), .B2(keyinput_218), .C1(n20486), .C2(
        keyinput_223), .A(n14007), .ZN(n14016) );
  AOI22_X1 U15692 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(keyinput_222), .B1(n22142), .B2(keyinput_227), .ZN(n14008) );
  OAI221_X1 U15693 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(keyinput_222), .C1(
        n22142), .C2(keyinput_227), .A(n14008), .ZN(n14014) );
  AOI22_X1 U15694 ( .A1(P1_EBX_REG_17__SCAN_IN), .A2(keyinput_226), .B1(n15973), .B2(keyinput_228), .ZN(n14009) );
  OAI221_X1 U15695 ( .B1(P1_EBX_REG_17__SCAN_IN), .B2(keyinput_226), .C1(
        n15973), .C2(keyinput_228), .A(n14009), .ZN(n14013) );
  INV_X1 U15696 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n20471) );
  AOI22_X1 U15697 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(keyinput_224), .B1(n20471), .B2(keyinput_225), .ZN(n14010) );
  OAI221_X1 U15698 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(keyinput_224), .C1(
        n20471), .C2(keyinput_225), .A(n14010), .ZN(n14012) );
  XOR2_X1 U15699 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_219), .Z(n14011) );
  OR4_X1 U15700 ( .A1(n14014), .A2(n14013), .A3(n14012), .A4(n14011), .ZN(
        n14015) );
  NOR4_X1 U15701 ( .A1(n14018), .A2(n14017), .A3(n14016), .A4(n14015), .ZN(
        n14022) );
  XOR2_X1 U15702 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_229), .Z(n14021) );
  XOR2_X1 U15703 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_230), .Z(n14020) );
  XNOR2_X1 U15704 ( .A(P1_EBX_REG_12__SCAN_IN), .B(keyinput_231), .ZN(n14019)
         );
  NOR4_X1 U15705 ( .A1(n14022), .A2(n14021), .A3(n14020), .A4(n14019), .ZN(
        n14034) );
  XNOR2_X1 U15706 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_232), .ZN(n14024)
         );
  XNOR2_X1 U15707 ( .A(P1_EBX_REG_10__SCAN_IN), .B(keyinput_233), .ZN(n14023)
         );
  NOR2_X1 U15708 ( .A1(n14024), .A2(n14023), .ZN(n14031) );
  XNOR2_X1 U15709 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_234), .ZN(n14026)
         );
  XNOR2_X1 U15710 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_235), .ZN(n14025)
         );
  NOR2_X1 U15711 ( .A1(n14026), .A2(n14025), .ZN(n14030) );
  INV_X1 U15712 ( .A(keyinput_236), .ZN(n14027) );
  XNOR2_X1 U15713 ( .A(n14027), .B(P1_EBX_REG_7__SCAN_IN), .ZN(n14029) );
  XNOR2_X1 U15714 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_237), .ZN(n14028)
         );
  NAND4_X1 U15715 ( .A1(n14031), .A2(n14030), .A3(n14029), .A4(n14028), .ZN(
        n14033) );
  XOR2_X1 U15716 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_238), .Z(n14032) );
  OAI21_X1 U15717 ( .B1(n14034), .B2(n14033), .A(n14032), .ZN(n14041) );
  XOR2_X1 U15718 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_242), .Z(n14038) );
  XOR2_X1 U15719 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_239), .Z(n14037) );
  XNOR2_X1 U15720 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_240), .ZN(n14036)
         );
  XNOR2_X1 U15721 ( .A(P1_EBX_REG_2__SCAN_IN), .B(keyinput_241), .ZN(n14035)
         );
  NOR4_X1 U15722 ( .A1(n14038), .A2(n14037), .A3(n14036), .A4(n14035), .ZN(
        n14040) );
  XNOR2_X1 U15723 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_243), .ZN(n14039)
         );
  AOI21_X1 U15724 ( .B1(n14041), .B2(n14040), .A(n14039), .ZN(n14044) );
  XNOR2_X1 U15725 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_244), .ZN(n14043)
         );
  XOR2_X1 U15726 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_245), .Z(n14042) );
  OAI21_X1 U15727 ( .B1(n14044), .B2(n14043), .A(n14042), .ZN(n14047) );
  XOR2_X1 U15728 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_247), .Z(n14046) );
  XNOR2_X1 U15729 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_246), .ZN(n14045)
         );
  NAND3_X1 U15730 ( .A1(n14047), .A2(n14046), .A3(n14045), .ZN(n14050) );
  XOR2_X1 U15731 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_248), .Z(n14049) );
  XNOR2_X1 U15732 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_249), .ZN(n14048)
         );
  NAND3_X1 U15733 ( .A1(n14050), .A2(n14049), .A3(n14048), .ZN(n14053) );
  XOR2_X1 U15734 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_250), .Z(n14052) );
  XOR2_X1 U15735 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_251), .Z(n14051) );
  NAND3_X1 U15736 ( .A1(n14053), .A2(n14052), .A3(n14051), .ZN(n14056) );
  XOR2_X1 U15737 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_252), .Z(n14055) );
  XOR2_X1 U15738 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_253), .Z(n14054) );
  NAND3_X1 U15739 ( .A1(n14056), .A2(n14055), .A3(n14054), .ZN(n14059) );
  XOR2_X1 U15740 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_254), .Z(n14058) );
  XNOR2_X1 U15741 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_255), .ZN(n14057)
         );
  NAND2_X1 U15742 ( .A1(n14060), .A2(n11845), .ZN(n14084) );
  NAND2_X1 U15743 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n22095), .ZN(n15484) );
  NOR2_X1 U15744 ( .A1(n15485), .A2(n15484), .ZN(n15483) );
  NAND2_X1 U15745 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15483), .ZN(n15585) );
  NAND2_X1 U15746 ( .A1(n14063), .A2(n14064), .ZN(n14065) );
  AND2_X1 U15747 ( .A1(n14061), .A2(n14065), .ZN(n20509) );
  NAND2_X1 U15748 ( .A1(n20509), .A2(n22172), .ZN(n14082) );
  NAND3_X1 U15749 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .ZN(n14066) );
  NOR3_X1 U15750 ( .A1(n22030), .A2(n22055), .A3(n14066), .ZN(n22054) );
  NAND3_X1 U15751 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n22054), .ZN(n22077) );
  INV_X1 U15752 ( .A(n22077), .ZN(n14067) );
  NAND2_X1 U15753 ( .A1(n14068), .A2(n14067), .ZN(n22112) );
  AND2_X1 U15754 ( .A1(n22200), .A2(n22112), .ZN(n22099) );
  NAND2_X1 U15755 ( .A1(n14069), .A2(n14070), .ZN(n14071) );
  NAND2_X1 U15756 ( .A1(n15882), .A2(n14071), .ZN(n16882) );
  OAI21_X1 U15757 ( .B1(n22152), .B2(n14072), .A(n21975), .ZN(n14077) );
  NOR2_X1 U15758 ( .A1(n14073), .A2(n17744), .ZN(n14074) );
  NOR2_X1 U15759 ( .A1(n22203), .A2(n20507), .ZN(n14076) );
  NOR2_X1 U15760 ( .A1(n14077), .A2(n14076), .ZN(n14079) );
  NAND2_X1 U15761 ( .A1(n22166), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n14078) );
  OAI211_X1 U15762 ( .C1(n16882), .C2(n22208), .A(n14079), .B(n14078), .ZN(
        n14080) );
  AOI21_X1 U15763 ( .B1(n22099), .B2(P1_REIP_REG_10__SCAN_IN), .A(n14080), 
        .ZN(n14081) );
  OAI211_X1 U15764 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n15585), .A(n14082), 
        .B(n14081), .ZN(n14083) );
  XNOR2_X1 U15765 ( .A(n14084), .B(n14083), .ZN(P1_U2830) );
  INV_X1 U15766 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14422) );
  XNOR2_X2 U15767 ( .A(n14087), .B(n14086), .ZN(n14808) );
  OR2_X1 U15768 ( .A1(n14090), .A2(n14089), .ZN(n14091) );
  NAND2_X2 U15769 ( .A1(n14092), .A2(n14091), .ZN(n19183) );
  AND2_X2 U15770 ( .A1(n14104), .A2(n14108), .ZN(n14148) );
  NOR2_X2 U15771 ( .A1(n14844), .A2(n14686), .ZN(n14109) );
  AOI22_X1 U15772 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14148), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14097) );
  AOI22_X1 U15773 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14146), .B1(
        n14149), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14096) );
  AOI22_X1 U15774 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14150), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14095) );
  AND2_X2 U15775 ( .A1(n14099), .A2(n14108), .ZN(n14153) );
  AND2_X2 U15776 ( .A1(n14107), .A2(n14105), .ZN(n14159) );
  AOI22_X1 U15777 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14153), .B1(
        n14159), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14094) );
  INV_X1 U15778 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14098) );
  NAND2_X1 U15779 ( .A1(n14099), .A2(n14103), .ZN(n14116) );
  INV_X1 U15780 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14100) );
  NOR2_X1 U15781 ( .A1(n14102), .A2(n14101), .ZN(n14113) );
  AOI22_X1 U15782 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n14158), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14112) );
  AND2_X2 U15783 ( .A1(n14104), .A2(n14105), .ZN(n14162) );
  AOI22_X1 U15784 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n14162), .B1(
        n14160), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14111) );
  NAND2_X1 U15785 ( .A1(n20178), .A2(n14264), .ZN(n14623) );
  OR2_X1 U15786 ( .A1(n14133), .A2(n14623), .ZN(n14130) );
  NAND2_X1 U15787 ( .A1(n14130), .A2(n14114), .ZN(n14115) );
  AOI22_X1 U15788 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14163), .B1(
        n14164), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14120) );
  AOI22_X1 U15789 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19796), .B1(
        n14162), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14119) );
  AOI22_X1 U15790 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n14158), .B1(
        n14159), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14118) );
  AOI22_X1 U15791 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n14160), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14117) );
  NOR2_X1 U15792 ( .A1(n14147), .A2(n14121), .ZN(n14122) );
  AOI21_X1 U15793 ( .B1(n14146), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n14122), .ZN(n14126) );
  AOI22_X1 U15794 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n14148), .B1(
        n14149), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U15795 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n14151), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14124) );
  AOI22_X1 U15796 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14152), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14123) );
  INV_X1 U15797 ( .A(n14127), .ZN(n14128) );
  NAND2_X1 U15798 ( .A1(n14128), .A2(n20178), .ZN(n14129) );
  INV_X1 U15799 ( .A(n14130), .ZN(n14131) );
  XOR2_X1 U15800 ( .A(n14132), .B(n14131), .Z(n14692) );
  XOR2_X1 U15801 ( .A(n14264), .B(n14133), .Z(n14134) );
  NAND2_X1 U15802 ( .A1(n14623), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14622) );
  NOR2_X1 U15803 ( .A1(n14134), .A2(n14622), .ZN(n14135) );
  XNOR2_X1 U15804 ( .A(n14134), .B(n14622), .ZN(n14718) );
  NOR2_X1 U15805 ( .A1(n14719), .A2(n14718), .ZN(n14717) );
  NOR2_X1 U15806 ( .A1(n14135), .A2(n14717), .ZN(n14136) );
  XOR2_X1 U15807 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n14136), .Z(
        n14691) );
  NOR2_X1 U15808 ( .A1(n14692), .A2(n14691), .ZN(n14690) );
  INV_X1 U15809 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14424) );
  NOR2_X1 U15810 ( .A1(n14136), .A2(n14424), .ZN(n14137) );
  OR2_X1 U15811 ( .A1(n14690), .A2(n14137), .ZN(n14138) );
  XNOR2_X1 U15812 ( .A(n14138), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15557) );
  NAND2_X1 U15813 ( .A1(n14138), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14139) );
  INV_X1 U15814 ( .A(n14140), .ZN(n14141) );
  NAND2_X1 U15815 ( .A1(n14173), .A2(n14142), .ZN(n14143) );
  INV_X1 U15816 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15743) );
  INV_X1 U15817 ( .A(n14143), .ZN(n14144) );
  AOI21_X2 U15818 ( .B1(n15649), .B2(n15743), .A(n14145), .ZN(n14193) );
  INV_X1 U15819 ( .A(n14173), .ZN(n14172) );
  INV_X1 U15820 ( .A(n14147), .ZN(n14179) );
  AOI22_X1 U15821 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n14146), .B1(
        n14179), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14157) );
  AOI22_X1 U15822 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n14148), .B1(
        n14149), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14156) );
  AOI22_X1 U15823 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14150), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14155) );
  AOI22_X1 U15824 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n14152), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14154) );
  AOI22_X1 U15825 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n14158), .B1(
        n14159), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14168) );
  AOI22_X1 U15826 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n14160), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14167) );
  AOI22_X1 U15827 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n14162), .B1(
        n19796), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14166) );
  AOI22_X1 U15828 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n14163), .B1(
        n14164), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14165) );
  NAND2_X1 U15829 ( .A1(n11841), .A2(n11847), .ZN(n14171) );
  NAND2_X1 U15830 ( .A1(n14169), .A2(n20178), .ZN(n14170) );
  NAND2_X1 U15831 ( .A1(n14172), .A2(n14174), .ZN(n14178) );
  INV_X1 U15832 ( .A(n14174), .ZN(n14175) );
  NAND2_X1 U15833 ( .A1(n14173), .A2(n14175), .ZN(n14176) );
  INV_X1 U15834 ( .A(n14280), .ZN(n14177) );
  NAND2_X1 U15835 ( .A1(n14193), .A2(n14177), .ZN(n14200) );
  INV_X1 U15836 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15742) );
  AOI22_X1 U15837 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14148), .B1(
        n14179), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14183) );
  AOI22_X1 U15838 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14150), .B1(
        n14158), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14182) );
  AOI22_X1 U15839 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n14160), .B1(
        n14159), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14181) );
  AOI22_X1 U15840 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14163), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14180) );
  NAND4_X1 U15841 ( .A1(n14183), .A2(n14182), .A3(n14181), .A4(n14180), .ZN(
        n14189) );
  AOI22_X1 U15842 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14146), .B1(
        n14149), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14187) );
  AOI22_X1 U15843 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n14151), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14186) );
  AOI22_X1 U15844 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19796), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14185) );
  AOI22_X1 U15845 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n14164), .B1(
        n14162), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14184) );
  NAND4_X1 U15846 ( .A1(n14187), .A2(n14186), .A3(n14185), .A4(n14184), .ZN(
        n14188) );
  NAND2_X1 U15847 ( .A1(n14190), .A2(n20178), .ZN(n14191) );
  NOR2_X1 U15848 ( .A1(n11206), .A2(n14201), .ZN(n14195) );
  AOI21_X1 U15849 ( .B1(n14280), .B2(n15742), .A(n14312), .ZN(n14194) );
  MUX2_X1 U15850 ( .A(n14195), .B(n14194), .S(n14193), .Z(n14199) );
  MUX2_X1 U15851 ( .A(n14204), .B(n15742), .S(n14280), .Z(n14197) );
  NAND2_X1 U15852 ( .A1(n14201), .A2(n15742), .ZN(n14196) );
  INV_X1 U15853 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17616) );
  INV_X1 U15854 ( .A(n11206), .ZN(n15754) );
  INV_X1 U15855 ( .A(n14206), .ZN(n14207) );
  XNOR2_X1 U15856 ( .A(n14209), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17572) );
  INV_X1 U15857 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17532) );
  INV_X1 U15858 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17533) );
  INV_X1 U15859 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17504) );
  NOR2_X1 U15860 ( .A1(n17516), .A2(n17504), .ZN(n17276) );
  NAND2_X1 U15861 ( .A1(n17276), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17263) );
  INV_X1 U15862 ( .A(n17263), .ZN(n17250) );
  NAND3_X1 U15863 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14438) );
  INV_X1 U15864 ( .A(n14438), .ZN(n14427) );
  NAND2_X1 U15865 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14211) );
  INV_X1 U15866 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17461) );
  NOR2_X1 U15867 ( .A1(n14212), .A2(n13619), .ZN(n14213) );
  OR2_X1 U15868 ( .A1(n14269), .A2(n14213), .ZN(n14236) );
  NAND2_X1 U15869 ( .A1(n14215), .A2(n14214), .ZN(n14268) );
  AOI21_X1 U15870 ( .B1(n11178), .B2(n14216), .A(n14223), .ZN(n14232) );
  INV_X1 U15871 ( .A(n14217), .ZN(n14231) );
  INV_X1 U15872 ( .A(n14266), .ZN(n14222) );
  INV_X1 U15873 ( .A(n14218), .ZN(n14221) );
  NAND2_X1 U15874 ( .A1(n14219), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n14220) );
  NAND2_X1 U15875 ( .A1(n14221), .A2(n14220), .ZN(n14262) );
  NOR2_X1 U15876 ( .A1(n14222), .A2(n14262), .ZN(n14229) );
  NAND2_X1 U15877 ( .A1(n14412), .A2(n14223), .ZN(n14228) );
  NAND2_X1 U15878 ( .A1(n20178), .A2(n14262), .ZN(n14226) );
  INV_X1 U15879 ( .A(n14224), .ZN(n14225) );
  NAND3_X1 U15880 ( .A1(n14226), .A2(n20237), .A3(n14225), .ZN(n14227) );
  OAI211_X1 U15881 ( .C1(n14229), .C2(n13619), .A(n14228), .B(n14227), .ZN(
        n14230) );
  OAI21_X1 U15882 ( .B1(n14232), .B2(n14231), .A(n14230), .ZN(n14233) );
  AOI22_X1 U15883 ( .A1(n14268), .A2(n13619), .B1(n14234), .B2(n14233), .ZN(
        n14235) );
  NOR2_X1 U15884 ( .A1(n14236), .A2(n14235), .ZN(n14237) );
  MUX2_X1 U15885 ( .A(n19179), .B(n14237), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n14240) );
  AND2_X1 U15886 ( .A1(n14269), .A2(n18958), .ZN(n14238) );
  NAND2_X1 U15887 ( .A1(n17641), .A2(n11178), .ZN(n14731) );
  INV_X1 U15888 ( .A(n14239), .ZN(n15268) );
  NAND2_X1 U15889 ( .A1(n15268), .A2(n14405), .ZN(n14278) );
  OAI21_X1 U15890 ( .B1(n14240), .B2(n13113), .A(n13111), .ZN(n14241) );
  INV_X1 U15891 ( .A(n14241), .ZN(n14242) );
  NAND2_X1 U15892 ( .A1(n14242), .A2(n14731), .ZN(n14277) );
  NOR2_X1 U15893 ( .A1(n14378), .A2(n20178), .ZN(n14275) );
  NAND2_X1 U15894 ( .A1(n14243), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14244) );
  NAND2_X1 U15895 ( .A1(n14244), .A2(n19179), .ZN(n19174) );
  INV_X1 U15896 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n14245) );
  OAI21_X1 U15897 ( .B1(n16210), .B2(n19174), .A(n14245), .ZN(n17791) );
  NOR2_X1 U15898 ( .A1(n14246), .A2(n14262), .ZN(n14247) );
  NOR2_X1 U15899 ( .A1(n15257), .A2(n14247), .ZN(n14248) );
  MUX2_X1 U15900 ( .A(n17791), .B(n14248), .S(n13265), .Z(n19203) );
  MUX2_X1 U15901 ( .A(n14249), .B(n14257), .S(n20178), .Z(n14250) );
  INV_X1 U15902 ( .A(n19213), .ZN(n22274) );
  OR2_X1 U15903 ( .A1(n14250), .A2(n22274), .ZN(n14273) );
  NAND2_X1 U15904 ( .A1(n15280), .A2(n15268), .ZN(n14251) );
  OR2_X1 U15905 ( .A1(n15257), .A2(n14251), .ZN(n14261) );
  AOI21_X1 U15906 ( .B1(n14252), .B2(n14710), .A(n14271), .ZN(n14408) );
  NAND2_X1 U15907 ( .A1(n20178), .A2(n13111), .ZN(n14395) );
  NAND2_X1 U15908 ( .A1(n14395), .A2(n20237), .ZN(n14253) );
  NAND2_X1 U15909 ( .A1(n14253), .A2(n14710), .ZN(n14254) );
  NAND2_X1 U15910 ( .A1(n14254), .A2(n14257), .ZN(n14255) );
  OAI211_X1 U15911 ( .C1(n14252), .C2(n13111), .A(n14255), .B(n14404), .ZN(
        n14256) );
  NOR2_X1 U15912 ( .A1(n14408), .A2(n14256), .ZN(n14260) );
  OAI21_X1 U15913 ( .B1(n13358), .B2(n20030), .A(n14257), .ZN(n14258) );
  NAND2_X1 U15914 ( .A1(n13315), .A2(n14258), .ZN(n14259) );
  AND2_X1 U15915 ( .A1(n14260), .A2(n14259), .ZN(n14397) );
  AND2_X1 U15916 ( .A1(n14261), .A2(n14397), .ZN(n15209) );
  INV_X1 U15917 ( .A(n14262), .ZN(n14263) );
  MUX2_X1 U15918 ( .A(n14264), .B(n14263), .S(n13619), .Z(n14294) );
  AOI21_X1 U15919 ( .B1(n14294), .B2(n14266), .A(n14265), .ZN(n14267) );
  NOR2_X1 U15920 ( .A1(n14268), .A2(n14267), .ZN(n14270) );
  OR2_X1 U15921 ( .A1(n14270), .A2(n14269), .ZN(n15258) );
  INV_X1 U15922 ( .A(n15258), .ZN(n14272) );
  NOR2_X1 U15923 ( .A1(n14378), .A2(n14271), .ZN(n15259) );
  NAND2_X1 U15924 ( .A1(n14272), .A2(n15259), .ZN(n14461) );
  OAI211_X1 U15925 ( .C1(n15257), .C2(n14273), .A(n15209), .B(n14461), .ZN(
        n14274) );
  AOI21_X1 U15926 ( .B1(n14275), .B2(n19203), .A(n14274), .ZN(n14276) );
  OAI211_X1 U15927 ( .C1(n14731), .C2(n14278), .A(n14277), .B(n14276), .ZN(
        n14279) );
  NAND2_X1 U15928 ( .A1(n14421), .A2(n15259), .ZN(n19193) );
  INV_X1 U15929 ( .A(n14281), .ZN(n14284) );
  INV_X1 U15930 ( .A(n14282), .ZN(n14283) );
  NAND2_X1 U15931 ( .A1(n14284), .A2(n14283), .ZN(n14285) );
  NAND2_X1 U15932 ( .A1(n14314), .A2(n14285), .ZN(n18973) );
  INV_X1 U15933 ( .A(n14288), .ZN(n14302) );
  INV_X1 U15934 ( .A(n14289), .ZN(n14292) );
  INV_X1 U15935 ( .A(n14290), .ZN(n14291) );
  NAND2_X1 U15936 ( .A1(n14292), .A2(n14291), .ZN(n14293) );
  NAND2_X1 U15937 ( .A1(n14302), .A2(n14293), .ZN(n15729) );
  MUX2_X1 U15938 ( .A(n14294), .B(P2_EBX_REG_0__SCAN_IN), .S(n19982), .Z(
        n15957) );
  NAND2_X1 U15939 ( .A1(n15957), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14621) );
  NAND3_X1 U15940 ( .A1(n19982), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n14295) );
  NAND2_X1 U15941 ( .A1(n14298), .A2(n14295), .ZN(n16965) );
  AND2_X1 U15942 ( .A1(n14621), .A2(n16965), .ZN(n14720) );
  NOR2_X1 U15943 ( .A1(n14621), .A2(n16965), .ZN(n14721) );
  NOR2_X1 U15944 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14721), .ZN(
        n14296) );
  NOR2_X1 U15945 ( .A1(n14720), .A2(n14296), .ZN(n14687) );
  XNOR2_X1 U15946 ( .A(n14298), .B(n14297), .ZN(n15831) );
  XNOR2_X1 U15947 ( .A(n15831), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14688) );
  NOR2_X1 U15948 ( .A1(n15831), .A2(n14424), .ZN(n14299) );
  AOI21_X1 U15949 ( .B1(n14687), .B2(n14688), .A(n14299), .ZN(n15547) );
  INV_X1 U15950 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15546) );
  INV_X1 U15951 ( .A(n14300), .ZN(n14301) );
  XNOR2_X1 U15952 ( .A(n14302), .B(n14301), .ZN(n16025) );
  AND2_X1 U15953 ( .A1(n16025), .A2(n15743), .ZN(n14303) );
  AOI21_X1 U15954 ( .B1(n15547), .B2(n15546), .A(n14303), .ZN(n14308) );
  INV_X1 U15955 ( .A(n15547), .ZN(n15645) );
  INV_X1 U15956 ( .A(n14303), .ZN(n14304) );
  NAND3_X1 U15957 ( .A1(n15645), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n14304), .ZN(n14307) );
  INV_X1 U15958 ( .A(n16025), .ZN(n14305) );
  NAND2_X1 U15959 ( .A1(n14305), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14306) );
  NAND3_X1 U15960 ( .A1(n14309), .A2(n15742), .A3(n18973), .ZN(n14310) );
  NAND2_X1 U15961 ( .A1(n14312), .A2(n16060), .ZN(n14315) );
  XNOR2_X1 U15962 ( .A(n14314), .B(n14313), .ZN(n18984) );
  XNOR2_X1 U15963 ( .A(n14316), .B(n17616), .ZN(n17610) );
  NAND2_X1 U15964 ( .A1(n14316), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14317) );
  INV_X1 U15965 ( .A(n14318), .ZN(n14319) );
  NAND2_X1 U15966 ( .A1(n11250), .A2(n14319), .ZN(n14320) );
  NAND2_X1 U15967 ( .A1(n14326), .A2(n14320), .ZN(n15848) );
  INV_X1 U15968 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17591) );
  OR3_X1 U15969 ( .A1(n15848), .A2(n16060), .A3(n17591), .ZN(n17575) );
  INV_X1 U15970 ( .A(n14321), .ZN(n16137) );
  XNOR2_X1 U15971 ( .A(n16137), .B(n14322), .ZN(n18997) );
  NAND2_X1 U15972 ( .A1(n18997), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17573) );
  OR2_X1 U15973 ( .A1(n15848), .A2(n16060), .ZN(n14323) );
  NAND2_X1 U15974 ( .A1(n14323), .A2(n17591), .ZN(n17576) );
  INV_X1 U15975 ( .A(n18997), .ZN(n14324) );
  NAND2_X1 U15976 ( .A1(n14324), .A2(n17605), .ZN(n17333) );
  AND2_X1 U15977 ( .A1(n17576), .A2(n17333), .ZN(n17320) );
  NAND2_X1 U15978 ( .A1(n14326), .A2(n14325), .ZN(n14327) );
  NAND2_X1 U15979 ( .A1(n14331), .A2(n14327), .ZN(n19005) );
  OAI21_X1 U15980 ( .B1(n19005), .B2(n16060), .A(n17532), .ZN(n17323) );
  AND2_X1 U15981 ( .A1(n17320), .A2(n17323), .ZN(n14328) );
  INV_X1 U15982 ( .A(n14329), .ZN(n14330) );
  NAND2_X1 U15983 ( .A1(n14331), .A2(n14330), .ZN(n14332) );
  NAND2_X1 U15984 ( .A1(n14337), .A2(n14332), .ZN(n15820) );
  OR2_X1 U15985 ( .A1(n15820), .A2(n16060), .ZN(n14333) );
  INV_X1 U15986 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17547) );
  NAND2_X1 U15987 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14334) );
  OR2_X1 U15988 ( .A1(n15820), .A2(n14334), .ZN(n17305) );
  NAND2_X1 U15989 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14335) );
  INV_X1 U15990 ( .A(n17294), .ZN(n14340) );
  NAND2_X1 U15991 ( .A1(n14337), .A2(n14336), .ZN(n14338) );
  NAND2_X1 U15992 ( .A1(n14342), .A2(n14338), .ZN(n15911) );
  NOR2_X1 U15993 ( .A1(n14341), .A2(n17533), .ZN(n17297) );
  NAND2_X1 U15994 ( .A1(n14341), .A2(n17533), .ZN(n17295) );
  XNOR2_X1 U15995 ( .A(n14342), .B(n11306), .ZN(n15932) );
  AND2_X1 U15996 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14343) );
  NAND2_X1 U15997 ( .A1(n15932), .A2(n14287), .ZN(n16035) );
  INV_X1 U15998 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17523) );
  NAND2_X1 U15999 ( .A1(n16035), .A2(n17523), .ZN(n17284) );
  INV_X1 U16000 ( .A(n14344), .ZN(n14346) );
  XNOR2_X1 U16001 ( .A(n14346), .B(n14345), .ZN(n15799) );
  INV_X1 U16002 ( .A(n15799), .ZN(n14347) );
  INV_X1 U16003 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17496) );
  OR3_X1 U16004 ( .A1(n14347), .A2(n16060), .A3(n17496), .ZN(n17255) );
  INV_X1 U16005 ( .A(n14348), .ZN(n14349) );
  XNOR2_X1 U16006 ( .A(n14350), .B(n14349), .ZN(n19025) );
  AND2_X1 U16007 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14351) );
  NAND2_X1 U16008 ( .A1(n19025), .A2(n14351), .ZN(n17272) );
  AND2_X1 U16009 ( .A1(n17255), .A2(n17272), .ZN(n14356) );
  INV_X1 U16010 ( .A(n14352), .ZN(n14354) );
  XNOR2_X1 U16011 ( .A(n14354), .B(n14353), .ZN(n19035) );
  AND2_X1 U16012 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14355) );
  NAND2_X1 U16013 ( .A1(n19035), .A2(n14355), .ZN(n17251) );
  AND2_X1 U16014 ( .A1(n14356), .A2(n17251), .ZN(n16044) );
  NAND2_X1 U16015 ( .A1(n17275), .A2(n16044), .ZN(n17227) );
  INV_X1 U16016 ( .A(n14357), .ZN(n14358) );
  XNOR2_X1 U16017 ( .A(n14359), .B(n14358), .ZN(n19055) );
  NAND2_X1 U16018 ( .A1(n19055), .A2(n14287), .ZN(n14360) );
  NAND2_X1 U16019 ( .A1(n14360), .A2(n17461), .ZN(n17230) );
  INV_X1 U16020 ( .A(n14361), .ZN(n14363) );
  XNOR2_X1 U16021 ( .A(n14363), .B(n14362), .ZN(n15790) );
  NAND2_X1 U16022 ( .A1(n15790), .A2(n14287), .ZN(n14364) );
  XNOR2_X1 U16023 ( .A(n14364), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17243) );
  NAND2_X1 U16024 ( .A1(n15799), .A2(n14287), .ZN(n14365) );
  NAND2_X1 U16025 ( .A1(n14365), .A2(n17496), .ZN(n17256) );
  NAND2_X1 U16026 ( .A1(n19025), .A2(n14287), .ZN(n14366) );
  NAND2_X1 U16027 ( .A1(n14366), .A2(n17504), .ZN(n17273) );
  AND2_X1 U16028 ( .A1(n17256), .A2(n17273), .ZN(n14368) );
  NAND2_X1 U16029 ( .A1(n19035), .A2(n14287), .ZN(n14367) );
  INV_X1 U16030 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17478) );
  NAND2_X1 U16031 ( .A1(n14367), .A2(n17478), .ZN(n17252) );
  AND2_X1 U16032 ( .A1(n14368), .A2(n17252), .ZN(n17226) );
  AND2_X1 U16033 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14369) );
  NAND2_X1 U16034 ( .A1(n19055), .A2(n14369), .ZN(n17229) );
  AND2_X1 U16035 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14370) );
  NAND2_X1 U16036 ( .A1(n15790), .A2(n14370), .ZN(n17228) );
  AND2_X1 U16037 ( .A1(n17229), .A2(n17228), .ZN(n16045) );
  INV_X1 U16038 ( .A(n16045), .ZN(n14371) );
  INV_X1 U16039 ( .A(n14372), .ZN(n14373) );
  XNOR2_X1 U16040 ( .A(n14374), .B(n14373), .ZN(n16950) );
  NAND2_X1 U16041 ( .A1(n16950), .A2(n14287), .ZN(n14375) );
  NAND2_X1 U16042 ( .A1(n14375), .A2(n14422), .ZN(n17213) );
  AND2_X1 U16043 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14376) );
  NAND2_X1 U16044 ( .A1(n16950), .A2(n14376), .ZN(n17215) );
  NAND2_X1 U16045 ( .A1(n17213), .A2(n17215), .ZN(n14377) );
  XNOR2_X1 U16046 ( .A(n17216), .B(n14377), .ZN(n14503) );
  NOR2_X1 U16047 ( .A1(n14378), .A2(n13619), .ZN(n15255) );
  NAND2_X1 U16048 ( .A1(n14421), .A2(n15255), .ZN(n19182) );
  INV_X1 U16049 ( .A(n15889), .ZN(n14379) );
  AOI21_X1 U16050 ( .B1(n14381), .B2(n14380), .A(n14379), .ZN(n16954) );
  OR2_X1 U16051 ( .A1(n14383), .A2(n14382), .ZN(n15235) );
  NAND2_X1 U16052 ( .A1(n15235), .A2(n20178), .ZN(n14385) );
  NAND2_X1 U16053 ( .A1(n14385), .A2(n14384), .ZN(n14386) );
  NAND2_X1 U16054 ( .A1(n15256), .A2(n11178), .ZN(n14390) );
  INV_X1 U16055 ( .A(n14387), .ZN(n14389) );
  NAND2_X1 U16056 ( .A1(n14389), .A2(n14388), .ZN(n14707) );
  NAND2_X1 U16057 ( .A1(n14390), .A2(n14707), .ZN(n14391) );
  OR2_X1 U16058 ( .A1(n15852), .A2(n14393), .ZN(n14394) );
  NAND2_X1 U16059 ( .A1(n14392), .A2(n14394), .ZN(n20121) );
  INV_X1 U16060 ( .A(n14395), .ZN(n14396) );
  NAND2_X1 U16061 ( .A1(n14421), .A2(n15254), .ZN(n15549) );
  NAND3_X1 U16062 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17613) );
  NOR2_X1 U16063 ( .A1(n17616), .A2(n17613), .ZN(n14435) );
  AND2_X1 U16064 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17587) );
  NAND2_X1 U16065 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17637) );
  NAND2_X1 U16066 ( .A1(n14424), .A2(n17637), .ZN(n15548) );
  NAND3_X1 U16067 ( .A1(n14435), .A2(n17587), .A3(n15548), .ZN(n14425) );
  INV_X1 U16068 ( .A(n14425), .ZN(n14399) );
  INV_X1 U16069 ( .A(n14421), .ZN(n14398) );
  INV_X2 U16070 ( .A(n19040), .ZN(n19068) );
  NAND2_X1 U16071 ( .A1(n14398), .A2(n19068), .ZN(n17631) );
  OAI21_X1 U16072 ( .B1(n15549), .B2(n14399), .A(n17631), .ZN(n16085) );
  NAND3_X1 U16073 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17489) );
  INV_X1 U16074 ( .A(n17489), .ZN(n14400) );
  AND4_X1 U16075 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n14400), .ZN(n17449) );
  NOR2_X1 U16076 ( .A1(n15549), .A2(n17449), .ZN(n14401) );
  OR2_X1 U16077 ( .A1(n16085), .A2(n14401), .ZN(n17452) );
  INV_X1 U16078 ( .A(n17452), .ZN(n14430) );
  INV_X1 U16079 ( .A(n14402), .ZN(n14418) );
  INV_X1 U16080 ( .A(n14403), .ZN(n14594) );
  NAND2_X1 U16081 ( .A1(n14404), .A2(n20030), .ZN(n14406) );
  AOI22_X1 U16082 ( .A1(n14594), .A2(n14406), .B1(n13113), .B2(n14405), .ZN(
        n14415) );
  NAND2_X1 U16083 ( .A1(n14407), .A2(n11178), .ZN(n15229) );
  INV_X1 U16084 ( .A(n14408), .ZN(n14409) );
  NAND2_X1 U16085 ( .A1(n15229), .A2(n14409), .ZN(n14411) );
  NAND2_X1 U16086 ( .A1(n14411), .A2(n14410), .ZN(n14414) );
  NAND2_X1 U16087 ( .A1(n14413), .A2(n14412), .ZN(n14743) );
  NAND4_X1 U16088 ( .A1(n14416), .A2(n14415), .A3(n14414), .A4(n14743), .ZN(
        n14417) );
  AOI21_X1 U16089 ( .B1(n14418), .B2(n13115), .A(n14417), .ZN(n15238) );
  NAND2_X1 U16090 ( .A1(n15238), .A2(n14419), .ZN(n14420) );
  NAND2_X1 U16091 ( .A1(n14421), .A2(n14420), .ZN(n17579) );
  AND2_X1 U16092 ( .A1(n15549), .A2(n17579), .ZN(n17581) );
  INV_X1 U16093 ( .A(n17581), .ZN(n19186) );
  NOR2_X1 U16094 ( .A1(n14438), .A2(n14422), .ZN(n14423) );
  NAND2_X1 U16095 ( .A1(n14423), .A2(n17449), .ZN(n14493) );
  INV_X1 U16096 ( .A(n14493), .ZN(n14426) );
  NOR2_X1 U16097 ( .A1(n14424), .A2(n17637), .ZN(n14432) );
  INV_X1 U16098 ( .A(n14432), .ZN(n15551) );
  NOR2_X1 U16099 ( .A1(n14425), .A2(n15551), .ZN(n16084) );
  AOI22_X1 U16100 ( .A1(n17579), .A2(n14427), .B1(n14426), .B2(n16084), .ZN(
        n14428) );
  NAND2_X1 U16101 ( .A1(n19186), .A2(n14428), .ZN(n14429) );
  NAND2_X1 U16102 ( .A1(n14430), .A2(n14429), .ZN(n14491) );
  NAND2_X1 U16103 ( .A1(n14491), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14431) );
  NAND2_X1 U16104 ( .A1(n19047), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n14500) );
  OAI211_X1 U16105 ( .C1(n17622), .C2(n20121), .A(n14431), .B(n14500), .ZN(
        n14439) );
  NAND2_X1 U16106 ( .A1(n17585), .A2(n15548), .ZN(n14434) );
  INV_X1 U16107 ( .A(n17579), .ZN(n15552) );
  NAND2_X1 U16108 ( .A1(n15552), .A2(n14432), .ZN(n14433) );
  INV_X1 U16109 ( .A(n14435), .ZN(n14436) );
  NOR2_X1 U16110 ( .A1(n17614), .A2(n14436), .ZN(n17606) );
  NAND2_X1 U16111 ( .A1(n17606), .A2(n17587), .ZN(n17563) );
  INV_X1 U16112 ( .A(n17449), .ZN(n14437) );
  OR2_X1 U16113 ( .A1(n17563), .A2(n14437), .ZN(n17484) );
  NOR3_X1 U16114 ( .A1(n17484), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n14438), .ZN(n14492) );
  AOI211_X1 U16115 ( .C1(n16954), .C2(n17633), .A(n14439), .B(n14492), .ZN(
        n14440) );
  INV_X1 U16116 ( .A(n16099), .ZN(n14442) );
  NAND2_X1 U16117 ( .A1(n19166), .A2(n19032), .ZN(n14443) );
  AOI21_X1 U16118 ( .B1(n14442), .B2(n14443), .A(n19201), .ZN(n14444) );
  NAND2_X1 U16119 ( .A1(n14444), .A2(n11243), .ZN(n14458) );
  AND2_X1 U16120 ( .A1(n16989), .A2(n14445), .ZN(n14446) );
  OR2_X2 U16121 ( .A1(n16145), .A2(n14446), .ZN(n16980) );
  AND2_X1 U16122 ( .A1(n17060), .A2(n14447), .ZN(n14448) );
  NOR2_X1 U16123 ( .A1(n14449), .A2(n14448), .ZN(n17053) );
  INV_X1 U16124 ( .A(n17053), .ZN(n14450) );
  OAI22_X1 U16125 ( .A1(n16980), .A2(n19163), .B1(n14450), .B2(n19161), .ZN(
        n14451) );
  INV_X1 U16126 ( .A(n14451), .ZN(n14457) );
  XNOR2_X1 U16127 ( .A(n14453), .B(n14452), .ZN(n16029) );
  AOI22_X1 U16128 ( .A1(n16029), .A2(n19156), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n19158), .ZN(n14455) );
  AOI22_X1 U16129 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19159), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19155), .ZN(n14454) );
  AND2_X1 U16130 ( .A1(n14455), .A2(n14454), .ZN(n14456) );
  NAND2_X1 U16131 ( .A1(n14458), .A2(n11829), .ZN(P2_U2826) );
  NAND2_X1 U16132 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14459) );
  OR2_X1 U16133 ( .A1(n14493), .A2(n14459), .ZN(n17422) );
  NAND2_X1 U16134 ( .A1(n19203), .A2(n15255), .ZN(n14462) );
  NAND2_X1 U16135 ( .A1(n14462), .A2(n14461), .ZN(n15267) );
  NAND2_X1 U16136 ( .A1(n15267), .A2(n18966), .ZN(n19222) );
  OR2_X1 U16137 ( .A1(n19222), .A2(n11178), .ZN(n17770) );
  NAND2_X1 U16138 ( .A1(n14484), .A2(n17782), .ZN(n14483) );
  INV_X1 U16139 ( .A(n14463), .ZN(n14465) );
  XNOR2_X1 U16140 ( .A(n14465), .B(n14464), .ZN(n19067) );
  NAND2_X1 U16141 ( .A1(n19067), .A2(n14287), .ZN(n14466) );
  INV_X1 U16142 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17442) );
  OR2_X1 U16143 ( .A1(n14466), .A2(n17442), .ZN(n17218) );
  AND2_X1 U16144 ( .A1(n17218), .A2(n17215), .ZN(n16046) );
  NAND2_X1 U16145 ( .A1(n14466), .A2(n17442), .ZN(n17217) );
  AND2_X1 U16146 ( .A1(n17217), .A2(n17213), .ZN(n16038) );
  INV_X1 U16147 ( .A(n16038), .ZN(n14467) );
  INV_X1 U16148 ( .A(n14468), .ZN(n14470) );
  NAND2_X1 U16149 ( .A1(n14470), .A2(n11663), .ZN(n14471) );
  NAND2_X1 U16150 ( .A1(n16033), .A2(n14471), .ZN(n16948) );
  XNOR2_X1 U16151 ( .A(n17206), .B(n17205), .ZN(n17207) );
  XNOR2_X1 U16152 ( .A(n17207), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14485) );
  OR2_X1 U16153 ( .A1(n19222), .A2(n13109), .ZN(n17774) );
  OR2_X1 U16154 ( .A1(n14485), .A2(n17774), .ZN(n14482) );
  OR2_X1 U16155 ( .A1(n14472), .A2(n14473), .ZN(n14474) );
  AND2_X1 U16156 ( .A1(n14474), .A2(n17036), .ZN(n17045) );
  NAND2_X1 U16157 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17693) );
  NAND2_X1 U16158 ( .A1(n19876), .A2(n17693), .ZN(n18965) );
  OR2_X1 U16159 ( .A1(n18965), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14475) );
  AND2_X1 U16160 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n14476) );
  NAND2_X1 U16161 ( .A1(n17752), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17692) );
  NAND2_X1 U16162 ( .A1(n22239), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14477) );
  NAND2_X1 U16163 ( .A1(n17692), .A2(n14477), .ZN(n14626) );
  NAND2_X1 U16164 ( .A1(n19047), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n14489) );
  NAND2_X1 U16165 ( .A1(n17780), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14478) );
  OAI211_X1 U16166 ( .C1(n17790), .C2(n14479), .A(n14489), .B(n14478), .ZN(
        n14480) );
  AOI21_X1 U16167 ( .B1(n17045), .B2(n17784), .A(n14480), .ZN(n14481) );
  NAND2_X1 U16168 ( .A1(n14483), .A2(n11833), .ZN(P2_U2994) );
  NAND2_X1 U16169 ( .A1(n14484), .A2(n17628), .ZN(n14498) );
  OR2_X1 U16170 ( .A1(n14485), .A2(n19182), .ZN(n14497) );
  AND2_X1 U16171 ( .A1(n17120), .A2(n14486), .ZN(n14487) );
  OR2_X1 U16172 ( .A1(n14487), .A2(n11267), .ZN(n20022) );
  INV_X1 U16173 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16047) );
  NAND2_X1 U16174 ( .A1(n16047), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14488) );
  OR3_X1 U16175 ( .A1(n17563), .A2(n14493), .A3(n14488), .ZN(n14490) );
  OAI211_X1 U16176 ( .C1(n17622), .C2(n20022), .A(n14490), .B(n14489), .ZN(
        n14495) );
  NOR2_X1 U16177 ( .A1(n14492), .A2(n14491), .ZN(n17443) );
  OR3_X1 U16178 ( .A1(n17563), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14493), .ZN(n17438) );
  AOI21_X1 U16179 ( .B1(n17443), .B2(n17438), .A(n16047), .ZN(n14494) );
  AOI211_X1 U16180 ( .C1(n17045), .C2(n17633), .A(n14495), .B(n14494), .ZN(
        n14496) );
  NAND2_X1 U16181 ( .A1(n14498), .A2(n11834), .ZN(P2_U3026) );
  NAND2_X1 U16182 ( .A1(n17780), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14499) );
  OAI211_X1 U16183 ( .C1(n17790), .C2(n16960), .A(n14500), .B(n14499), .ZN(
        n14501) );
  AOI21_X1 U16184 ( .B1(n16954), .B2(n17784), .A(n14501), .ZN(n14502) );
  OAI21_X1 U16185 ( .B1(n14503), .B2(n17774), .A(n14502), .ZN(n14504) );
  INV_X1 U16186 ( .A(n14504), .ZN(n14505) );
  NOR4_X1 U16187 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n14509) );
  NOR4_X1 U16188 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n14508) );
  NOR4_X1 U16189 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n14507) );
  NOR4_X1 U16190 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n14506) );
  NAND4_X1 U16191 ( .A1(n14509), .A2(n14508), .A3(n14507), .A4(n14506), .ZN(
        n14514) );
  NOR4_X1 U16192 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n14512) );
  NOR4_X1 U16193 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n14511) );
  NOR4_X1 U16194 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n14510) );
  INV_X1 U16195 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20403) );
  NAND4_X1 U16196 ( .A1(n14512), .A2(n14511), .A3(n14510), .A4(n20403), .ZN(
        n14513) );
  OAI21_X2 U16197 ( .B1(n14514), .B2(n14513), .A(P1_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n16592) );
  NOR3_X1 U16198 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20628), .ZN(n14516) );
  NOR4_X1 U16199 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14515) );
  NAND4_X1 U16200 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(n16588), .A3(n14516), .A4(
        n14515), .ZN(U214) );
  NOR4_X1 U16201 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n14520) );
  NOR4_X1 U16202 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n14519) );
  NOR4_X1 U16203 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n14518) );
  NOR4_X1 U16204 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n14517) );
  NAND4_X1 U16205 ( .A1(n14520), .A2(n14519), .A3(n14518), .A4(n14517), .ZN(
        n14525) );
  NOR4_X1 U16206 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n14523) );
  NOR4_X1 U16207 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n14522) );
  NOR4_X1 U16208 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n14521) );
  INV_X1 U16209 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n17858) );
  NAND4_X1 U16210 ( .A1(n14523), .A2(n14522), .A3(n14521), .A4(n17858), .ZN(
        n14524) );
  OAI21_X1 U16211 ( .B1(n14525), .B2(n14524), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14712) );
  NOR2_X1 U16212 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14527) );
  NOR4_X1 U16213 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14526) );
  NAND4_X1 U16214 ( .A1(n14527), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14526), .ZN(n14528) );
  OR2_X1 U16215 ( .A1(n19718), .A2(n14528), .ZN(n20565) );
  OR2_X1 U16216 ( .A1(n20565), .A2(n20615), .ZN(U212) );
  NOR2_X1 U16217 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14528), .ZN(n19247)
         );
  INV_X1 U16218 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14530) );
  MUX2_X1 U16219 ( .A(n14530), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .S(
        n20552), .Z(n14531) );
  NAND2_X1 U16220 ( .A1(n16734), .A2(n14531), .ZN(n16723) );
  OAI21_X1 U16221 ( .B1(n16734), .B2(n14531), .A(n16723), .ZN(n16746) );
  INV_X1 U16222 ( .A(n22810), .ZN(n14538) );
  INV_X1 U16223 ( .A(n14532), .ZN(n14536) );
  AOI21_X1 U16224 ( .B1(n14533), .B2(n15529), .A(n22414), .ZN(n14534) );
  NAND2_X1 U16225 ( .A1(n14535), .A2(n14534), .ZN(n14565) );
  NAND2_X1 U16226 ( .A1(n14536), .A2(n14565), .ZN(n14537) );
  NAND2_X1 U16227 ( .A1(n14538), .A2(n14537), .ZN(n14775) );
  INV_X1 U16228 ( .A(n16419), .ZN(n22808) );
  NAND2_X1 U16229 ( .A1(n14764), .A2(n17713), .ZN(n14539) );
  NAND4_X1 U16230 ( .A1(n22808), .A2(n14776), .A3(n22253), .A4(n14539), .ZN(
        n14546) );
  NAND2_X1 U16231 ( .A1(n14541), .A2(n22253), .ZN(n14542) );
  OAI211_X1 U16232 ( .C1(n14785), .C2(n14542), .A(n15127), .B(n16591), .ZN(
        n14543) );
  NAND3_X1 U16233 ( .A1(n16421), .A2(n14540), .A3(n14543), .ZN(n14545) );
  NAND3_X1 U16234 ( .A1(n16422), .A2(n16888), .A3(n14764), .ZN(n14544) );
  NAND4_X1 U16235 ( .A1(n14775), .A2(n14546), .A3(n14545), .A4(n14544), .ZN(
        n14547) );
  NOR2_X1 U16236 ( .A1(n14789), .A2(n14554), .ZN(n15075) );
  NAND2_X1 U16237 ( .A1(n15075), .A2(n14548), .ZN(n14771) );
  INV_X1 U16238 ( .A(n14771), .ZN(n14549) );
  NOR2_X1 U16239 ( .A1(n17733), .A2(n14549), .ZN(n16418) );
  OAI22_X1 U16240 ( .A1(n14581), .A2(n14550), .B1(n15391), .B2(n14762), .ZN(
        n14551) );
  INV_X1 U16241 ( .A(n14551), .ZN(n14552) );
  NAND3_X1 U16242 ( .A1(n16418), .A2(n14552), .A3(n15103), .ZN(n14553) );
  NOR2_X1 U16243 ( .A1(n16746), .A2(n22010), .ZN(n14588) );
  OR2_X1 U16244 ( .A1(n14554), .A2(n12752), .ZN(n14555) );
  NOR2_X1 U16245 ( .A1(n14789), .A2(n14555), .ZN(n16420) );
  NAND2_X1 U16246 ( .A1(n16420), .A2(n14583), .ZN(n16788) );
  INV_X1 U16247 ( .A(n16890), .ZN(n15125) );
  INV_X1 U16248 ( .A(n14556), .ZN(n14564) );
  OAI21_X1 U16249 ( .B1(n14540), .B2(n11922), .A(n15309), .ZN(n14557) );
  OAI21_X1 U16250 ( .B1(n14558), .B2(n14557), .A(n14764), .ZN(n14562) );
  INV_X1 U16251 ( .A(n14777), .ZN(n15411) );
  NAND2_X1 U16252 ( .A1(n15411), .A2(n14559), .ZN(n14560) );
  NAND3_X1 U16253 ( .A1(n14562), .A2(n14561), .A3(n14560), .ZN(n14563) );
  AOI21_X1 U16254 ( .B1(n14564), .B2(n16435), .A(n14563), .ZN(n14566) );
  NAND3_X1 U16255 ( .A1(n14567), .A2(n14566), .A3(n14565), .ZN(n14787) );
  OAI21_X1 U16256 ( .B1(n14784), .B2(n11177), .A(n14568), .ZN(n14569) );
  OR2_X1 U16257 ( .A1(n14787), .A2(n14569), .ZN(n14570) );
  NAND2_X1 U16258 ( .A1(n16788), .A2(n21922), .ZN(n16798) );
  INV_X1 U16259 ( .A(n16798), .ZN(n16878) );
  INV_X1 U16260 ( .A(n14577), .ZN(n16781) );
  INV_X1 U16261 ( .A(n21922), .ZN(n16793) );
  NOR2_X1 U16262 ( .A1(n16758), .A2(n16757), .ZN(n14576) );
  INV_X1 U16263 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15709) );
  INV_X1 U16264 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15719) );
  NOR3_X1 U16265 ( .A1(n15709), .A2(n15719), .A3(n12895), .ZN(n16877) );
  AND3_X1 U16266 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n16877), .ZN(n16868) );
  AND2_X1 U16267 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16868), .ZN(
        n21890) );
  NAND2_X1 U16268 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21890), .ZN(
        n16844) );
  INV_X1 U16269 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16893) );
  NAND2_X1 U16270 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14571) );
  NOR3_X1 U16271 ( .A1(n15361), .A2(n16893), .A3(n14571), .ZN(n15520) );
  NAND2_X1 U16272 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15520), .ZN(
        n15610) );
  NOR2_X1 U16273 ( .A1(n16844), .A2(n15610), .ZN(n16852) );
  NAND2_X1 U16274 ( .A1(n14576), .A2(n16852), .ZN(n16785) );
  INV_X1 U16275 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16895) );
  OAI21_X1 U16276 ( .B1(n16895), .B2(n16893), .A(n15361), .ZN(n15363) );
  NAND3_X1 U16277 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n15363), .ZN(n15517) );
  OR2_X1 U16278 ( .A1(n12888), .A2(n15517), .ZN(n15611) );
  NOR2_X1 U16279 ( .A1(n16844), .A2(n15611), .ZN(n16850) );
  AND2_X1 U16280 ( .A1(n14576), .A2(n16850), .ZN(n16782) );
  NAND2_X1 U16281 ( .A1(n14900), .A2(n16895), .ZN(n14573) );
  INV_X2 U16282 ( .A(n21975), .ZN(n21999) );
  NOR2_X1 U16283 ( .A1(n21999), .A2(n14583), .ZN(n16854) );
  INV_X1 U16284 ( .A(n16854), .ZN(n14572) );
  OAI21_X1 U16285 ( .B1(n16782), .B2(n16788), .A(n21920), .ZN(n14574) );
  AOI21_X1 U16286 ( .B1(n16793), .B2(n16785), .A(n14574), .ZN(n21907) );
  OAI21_X1 U16287 ( .B1(n16878), .B2(n16781), .A(n21907), .ZN(n21903) );
  AND2_X1 U16288 ( .A1(n21903), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14587) );
  INV_X1 U16289 ( .A(n16852), .ZN(n14575) );
  NOR2_X1 U16290 ( .A1(n16895), .A2(n14575), .ZN(n16858) );
  AOI22_X1 U16291 ( .A1(n21918), .A2(n16850), .B1(n14900), .B2(n16858), .ZN(
        n16859) );
  OAI21_X1 U16292 ( .B1(n14575), .B2(n16851), .A(n16859), .ZN(n21866) );
  NAND2_X1 U16293 ( .A1(n14576), .A2(n21866), .ZN(n21915) );
  NOR3_X1 U16294 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14577), .A3(
        n21915), .ZN(n14586) );
  AND2_X1 U16295 ( .A1(n16583), .A2(n14578), .ZN(n14579) );
  NOR2_X1 U16296 ( .A1(n16550), .A2(n14579), .ZN(n22164) );
  NAND2_X1 U16297 ( .A1(n16423), .A2(n15391), .ZN(n17715) );
  OAI21_X1 U16298 ( .B1(n14581), .B2(n14580), .A(n17715), .ZN(n14582) );
  NAND2_X1 U16299 ( .A1(n22164), .A2(n21993), .ZN(n14584) );
  NAND2_X1 U16300 ( .A1(n21999), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16743) );
  NAND2_X1 U16301 ( .A1(n14584), .A2(n16743), .ZN(n14585) );
  OR4_X1 U16302 ( .A1(n14588), .A2(n14587), .A3(n14586), .A4(n14585), .ZN(
        P1_U3013) );
  OR2_X1 U16303 ( .A1(n13315), .A2(n19219), .ZN(n14589) );
  OR2_X1 U16304 ( .A1(n15257), .A2(n14589), .ZN(n16973) );
  INV_X1 U16305 ( .A(n16973), .ZN(n14592) );
  INV_X1 U16306 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n14590) );
  NAND2_X1 U16307 ( .A1(n19880), .A2(n13265), .ZN(n17751) );
  OAI211_X1 U16308 ( .C1(n14592), .C2(n14590), .A(n14599), .B(n17751), .ZN(
        P2_U2814) );
  INV_X1 U16309 ( .A(n17751), .ZN(n14591) );
  NOR4_X1 U16310 ( .A1(n14600), .A2(n14592), .A3(P2_READREQUEST_REG_SCAN_IN), 
        .A4(n14591), .ZN(n14593) );
  AOI21_X1 U16311 ( .B1(n18968), .B2(n14594), .A(n14593), .ZN(P2_U3612) );
  NAND2_X1 U16312 ( .A1(n22810), .A2(n22808), .ZN(n14768) );
  AND2_X1 U16313 ( .A1(n16422), .A2(n15406), .ZN(n14595) );
  AOI21_X1 U16314 ( .B1(n14768), .B2(n14762), .A(n14595), .ZN(n16430) );
  AOI21_X1 U16315 ( .B1(n16430), .B2(n22809), .A(n14596), .ZN(n14598) );
  NOR3_X1 U16316 ( .A1(n17669), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n22225), 
        .ZN(n14597) );
  OR2_X1 U16317 ( .A1(n14598), .A2(n14597), .ZN(P1_U2803) );
  INV_X1 U16318 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14923) );
  OAI21_X1 U16319 ( .B1(n22274), .B2(n14599), .A(n14732), .ZN(n14649) );
  INV_X1 U16320 ( .A(n14649), .ZN(n14618) );
  NAND2_X1 U16321 ( .A1(n14618), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14603) );
  NAND3_X1 U16322 ( .A1(n14600), .A2(n11178), .A3(n19213), .ZN(n14713) );
  INV_X1 U16323 ( .A(n14713), .ZN(n14614) );
  NAND2_X1 U16324 ( .A1(n19718), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14602) );
  INV_X1 U16325 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20586) );
  OR2_X1 U16326 ( .A1(n14712), .A2(n20586), .ZN(n14601) );
  NAND2_X1 U16327 ( .A1(n14602), .A2(n14601), .ZN(n19705) );
  NAND2_X1 U16328 ( .A1(n14614), .A2(n19705), .ZN(n14616) );
  OAI211_X1 U16329 ( .C1(n14923), .C2(n14732), .A(n14603), .B(n14616), .ZN(
        P2_U2962) );
  INV_X1 U16330 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14934) );
  NAND2_X1 U16331 ( .A1(n14618), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14604) );
  MUX2_X1 U16332 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n19718), .Z(n19693) );
  NAND2_X1 U16333 ( .A1(n14614), .A2(n19693), .ZN(n14608) );
  OAI211_X1 U16334 ( .C1(n14934), .C2(n14732), .A(n14604), .B(n14608), .ZN(
        P2_U2966) );
  INV_X1 U16335 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14920) );
  NAND2_X1 U16336 ( .A1(n14618), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14605) );
  INV_X1 U16337 ( .A(n14712), .ZN(n19717) );
  AOI22_X1 U16338 ( .A1(n19717), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19718), .ZN(n19702) );
  INV_X1 U16339 ( .A(n19702), .ZN(n17068) );
  NAND2_X1 U16340 ( .A1(n14614), .A2(n17068), .ZN(n14684) );
  OAI211_X1 U16341 ( .C1(n14732), .C2(n14920), .A(n14605), .B(n14684), .ZN(
        P2_U2963) );
  INV_X1 U16342 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n17048) );
  NAND2_X1 U16343 ( .A1(n14618), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14607) );
  AOI22_X1 U16344 ( .A1(n19717), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19718), .ZN(n19696) );
  INV_X1 U16345 ( .A(n19696), .ZN(n14606) );
  NAND2_X1 U16346 ( .A1(n14614), .A2(n14606), .ZN(n14676) );
  OAI211_X1 U16347 ( .C1(n14732), .C2(n17048), .A(n14607), .B(n14676), .ZN(
        P2_U2965) );
  INV_X1 U16348 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17849) );
  NAND2_X1 U16349 ( .A1(n14618), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n14609) );
  OAI211_X1 U16350 ( .C1(n17849), .C2(n14732), .A(n14609), .B(n14608), .ZN(
        P2_U2981) );
  INV_X1 U16351 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14741) );
  NAND2_X1 U16352 ( .A1(n14618), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14613) );
  INV_X1 U16353 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14610) );
  OR2_X1 U16354 ( .A1(n14712), .A2(n14610), .ZN(n14612) );
  NAND2_X1 U16355 ( .A1(n14712), .A2(BUF2_REG_9__SCAN_IN), .ZN(n14611) );
  AND2_X1 U16356 ( .A1(n14612), .A2(n14611), .ZN(n19708) );
  INV_X1 U16357 ( .A(n19708), .ZN(n17083) );
  NAND2_X1 U16358 ( .A1(n14614), .A2(n17083), .ZN(n14680) );
  OAI211_X1 U16359 ( .C1(n14732), .C2(n14741), .A(n14613), .B(n14680), .ZN(
        P2_U2961) );
  INV_X1 U16360 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17846) );
  NAND2_X1 U16361 ( .A1(n14618), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n14615) );
  MUX2_X1 U16362 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n14712), .Z(n19699) );
  NAND2_X1 U16363 ( .A1(n14614), .A2(n19699), .ZN(n14619) );
  OAI211_X1 U16364 ( .C1(n17846), .C2(n14732), .A(n14615), .B(n14619), .ZN(
        P2_U2979) );
  INV_X1 U16365 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17843) );
  NAND2_X1 U16366 ( .A1(n14618), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14617) );
  OAI211_X1 U16367 ( .C1(n17843), .C2(n14732), .A(n14617), .B(n14616), .ZN(
        P2_U2977) );
  INV_X1 U16368 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14925) );
  NAND2_X1 U16369 ( .A1(n14618), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14620) );
  OAI211_X1 U16370 ( .C1(n14925), .C2(n14732), .A(n14620), .B(n14619), .ZN(
        P2_U2964) );
  OAI21_X1 U16371 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15957), .A(
        n14621), .ZN(n19181) );
  INV_X1 U16372 ( .A(n19181), .ZN(n14625) );
  OAI21_X1 U16373 ( .B1(n14623), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14622), .ZN(n19194) );
  NAND2_X1 U16374 ( .A1(n19047), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19191) );
  OAI21_X1 U16375 ( .B1(n17770), .B2(n19194), .A(n19191), .ZN(n14624) );
  AOI21_X1 U16376 ( .B1(n17785), .B2(n14625), .A(n14624), .ZN(n14628) );
  OAI21_X1 U16377 ( .B1(n17780), .B2(n14626), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14627) );
  OAI211_X1 U16378 ( .C1(n17773), .C2(n19183), .A(n14628), .B(n14627), .ZN(
        P2_U3014) );
  INV_X1 U16379 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n14630) );
  AOI22_X1 U16380 ( .A1(n19717), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19718), .ZN(n20077) );
  NOR2_X1 U16381 ( .A1(n14713), .A2(n20077), .ZN(n14635) );
  AOI21_X1 U16382 ( .B1(n14682), .B2(P2_EAX_REG_19__SCAN_IN), .A(n14635), .ZN(
        n14629) );
  OAI21_X1 U16383 ( .B1(n14649), .B2(n14630), .A(n14629), .ZN(P2_U2955) );
  INV_X1 U16384 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n14632) );
  OAI22_X1 U16385 ( .A1(n19718), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19717), .ZN(n20028) );
  NOR2_X1 U16386 ( .A1(n14713), .A2(n20028), .ZN(n14662) );
  AOI21_X1 U16387 ( .B1(n14682), .B2(P2_EAX_REG_20__SCAN_IN), .A(n14662), .ZN(
        n14631) );
  OAI21_X1 U16388 ( .B1(n14649), .B2(n14632), .A(n14631), .ZN(P2_U2956) );
  INV_X1 U16389 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n14634) );
  AOI22_X1 U16390 ( .A1(n19717), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19718), .ZN(n19980) );
  NOR2_X1 U16391 ( .A1(n14713), .A2(n19980), .ZN(n14653) );
  AOI21_X1 U16392 ( .B1(n14682), .B2(P2_EAX_REG_5__SCAN_IN), .A(n14653), .ZN(
        n14633) );
  OAI21_X1 U16393 ( .B1(n14649), .B2(n14634), .A(n14633), .ZN(P2_U2972) );
  INV_X1 U16394 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n14637) );
  AOI21_X1 U16395 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n14678), .A(n14635), .ZN(
        n14636) );
  OAI21_X1 U16396 ( .B1(n14649), .B2(n14637), .A(n14636), .ZN(P2_U2970) );
  INV_X1 U16397 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n14639) );
  AOI22_X1 U16398 ( .A1(n19717), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19718), .ZN(n19712) );
  NOR2_X1 U16399 ( .A1(n14713), .A2(n19712), .ZN(n14659) );
  AOI21_X1 U16400 ( .B1(n14682), .B2(P2_EAX_REG_24__SCAN_IN), .A(n14659), .ZN(
        n14638) );
  OAI21_X1 U16401 ( .B1(n14649), .B2(n14639), .A(n14638), .ZN(P2_U2960) );
  INV_X1 U16402 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n14641) );
  OAI22_X1 U16403 ( .A1(n19718), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19717), .ZN(n20235) );
  NOR2_X1 U16404 ( .A1(n14713), .A2(n20235), .ZN(n14644) );
  AOI21_X1 U16405 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n14682), .A(n14644), .ZN(
        n14640) );
  OAI21_X1 U16406 ( .B1(n14649), .B2(n14641), .A(n14640), .ZN(P2_U2967) );
  INV_X1 U16407 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n14643) );
  AOI22_X1 U16408 ( .A1(n19717), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19718), .ZN(n20177) );
  NOR2_X1 U16409 ( .A1(n14713), .A2(n20177), .ZN(n14656) );
  AOI21_X1 U16410 ( .B1(n14678), .B2(P2_EAX_REG_17__SCAN_IN), .A(n14656), .ZN(
        n14642) );
  OAI21_X1 U16411 ( .B1(n14649), .B2(n14643), .A(n14642), .ZN(P2_U2953) );
  INV_X1 U16412 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n14646) );
  AOI21_X1 U16413 ( .B1(n14682), .B2(P2_EAX_REG_16__SCAN_IN), .A(n14644), .ZN(
        n14645) );
  OAI21_X1 U16414 ( .B1(n14649), .B2(n14646), .A(n14645), .ZN(P2_U2952) );
  INV_X1 U16415 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n14648) );
  OAI22_X1 U16416 ( .A1(n19718), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19717), .ZN(n20128) );
  NOR2_X1 U16417 ( .A1(n14713), .A2(n20128), .ZN(n14650) );
  AOI21_X1 U16418 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n14682), .A(n14650), .ZN(
        n14647) );
  OAI21_X1 U16419 ( .B1(n14715), .B2(n14648), .A(n14647), .ZN(P2_U2969) );
  CLKBUF_X1 U16420 ( .A(n14649), .Z(n14715) );
  INV_X1 U16421 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14652) );
  AOI21_X1 U16422 ( .B1(n14682), .B2(P2_EAX_REG_18__SCAN_IN), .A(n14650), .ZN(
        n14651) );
  OAI21_X1 U16423 ( .B1(n14715), .B2(n14652), .A(n14651), .ZN(P2_U2954) );
  INV_X1 U16424 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n14655) );
  AOI21_X1 U16425 ( .B1(n14682), .B2(P2_EAX_REG_21__SCAN_IN), .A(n14653), .ZN(
        n14654) );
  OAI21_X1 U16426 ( .B1(n14715), .B2(n14655), .A(n14654), .ZN(P2_U2957) );
  INV_X1 U16427 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n14658) );
  AOI21_X1 U16428 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n14682), .A(n14656), .ZN(
        n14657) );
  OAI21_X1 U16429 ( .B1(n14715), .B2(n14658), .A(n14657), .ZN(P2_U2968) );
  INV_X1 U16430 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n14661) );
  AOI21_X1 U16431 ( .B1(P2_EAX_REG_8__SCAN_IN), .B2(n14678), .A(n14659), .ZN(
        n14660) );
  OAI21_X1 U16432 ( .B1(n14715), .B2(n14661), .A(n14660), .ZN(P2_U2975) );
  INV_X1 U16433 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n14664) );
  AOI21_X1 U16434 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n14682), .A(n14662), .ZN(
        n14663) );
  OAI21_X1 U16435 ( .B1(n14715), .B2(n14664), .A(n14663), .ZN(P2_U2971) );
  INV_X1 U16436 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n14666) );
  AOI22_X1 U16437 ( .A1(n19717), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19718), .ZN(n19721) );
  NOR2_X1 U16438 ( .A1(n14713), .A2(n19721), .ZN(n14669) );
  AOI21_X1 U16439 ( .B1(n14682), .B2(P2_EAX_REG_7__SCAN_IN), .A(n14669), .ZN(
        n14665) );
  OAI21_X1 U16440 ( .B1(n14715), .B2(n14666), .A(n14665), .ZN(P2_U2974) );
  INV_X1 U16441 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n14668) );
  INV_X1 U16442 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20579) );
  INV_X1 U16443 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21199) );
  AOI22_X1 U16444 ( .A1(n19717), .A2(n20579), .B1(n21199), .B2(n19718), .ZN(
        n19922) );
  INV_X1 U16445 ( .A(n19922), .ZN(n19932) );
  NOR2_X1 U16446 ( .A1(n14713), .A2(n19932), .ZN(n14672) );
  AOI21_X1 U16447 ( .B1(n14682), .B2(P2_EAX_REG_22__SCAN_IN), .A(n14672), .ZN(
        n14667) );
  OAI21_X1 U16448 ( .B1(n14715), .B2(n14668), .A(n14667), .ZN(P2_U2958) );
  INV_X1 U16449 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n14671) );
  AOI21_X1 U16450 ( .B1(n14678), .B2(P2_EAX_REG_23__SCAN_IN), .A(n14669), .ZN(
        n14670) );
  OAI21_X1 U16451 ( .B1(n14715), .B2(n14671), .A(n14670), .ZN(P2_U2959) );
  INV_X1 U16452 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n14674) );
  AOI21_X1 U16453 ( .B1(n14682), .B2(P2_EAX_REG_6__SCAN_IN), .A(n14672), .ZN(
        n14673) );
  OAI21_X1 U16454 ( .B1(n14715), .B2(n14674), .A(n14673), .ZN(P2_U2973) );
  INV_X1 U16455 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n14677) );
  NAND2_X1 U16456 ( .A1(n14678), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n14675) );
  OAI211_X1 U16457 ( .C1(n14649), .C2(n14677), .A(n14676), .B(n14675), .ZN(
        P2_U2980) );
  INV_X1 U16458 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n14681) );
  NAND2_X1 U16459 ( .A1(n14678), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n14679) );
  OAI211_X1 U16460 ( .C1(n14649), .C2(n14681), .A(n14680), .B(n14679), .ZN(
        P2_U2976) );
  INV_X1 U16461 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n14685) );
  NAND2_X1 U16462 ( .A1(n14682), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n14683) );
  OAI211_X1 U16463 ( .C1(n14715), .C2(n14685), .A(n14684), .B(n14683), .ZN(
        P2_U2978) );
  XOR2_X1 U16464 ( .A(n14688), .B(n14687), .Z(n14836) );
  INV_X1 U16465 ( .A(n15825), .ZN(n14689) );
  AND2_X1 U16466 ( .A1(n17754), .A2(n14689), .ZN(n14696) );
  INV_X1 U16467 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14694) );
  AOI21_X1 U16468 ( .B1(n14692), .B2(n14691), .A(n14690), .ZN(n14828) );
  NAND2_X1 U16469 ( .A1(n17782), .A2(n14828), .ZN(n14693) );
  NAND2_X1 U16470 ( .A1(n19047), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14831) );
  OAI211_X1 U16471 ( .C1(n17762), .C2(n14694), .A(n14693), .B(n14831), .ZN(
        n14695) );
  AOI211_X1 U16472 ( .C1(n14836), .C2(n17785), .A(n14696), .B(n14695), .ZN(
        n14697) );
  OAI21_X1 U16473 ( .B1(n14686), .B2(n17773), .A(n14697), .ZN(P2_U3012) );
  NAND2_X1 U16474 ( .A1(n14878), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14698) );
  NAND2_X1 U16475 ( .A1(n14698), .A2(n19876), .ZN(n14849) );
  AOI22_X1 U16476 ( .A1(n14849), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19880), .B2(n19891), .ZN(n14699) );
  INV_X1 U16477 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14702) );
  NOR2_X1 U16478 ( .A1(n16324), .A2(n14702), .ZN(n14818) );
  AND2_X1 U16479 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n14846) );
  INV_X1 U16480 ( .A(n14846), .ZN(n19861) );
  NAND2_X1 U16481 ( .A1(n19891), .A2(n19889), .ZN(n19905) );
  AND2_X1 U16482 ( .A1(n19861), .A2(n19905), .ZN(n19754) );
  AND2_X1 U16483 ( .A1(n19754), .A2(n19880), .ZN(n19873) );
  AOI21_X1 U16484 ( .B1(n14849), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19873), .ZN(n14703) );
  NAND2_X1 U16485 ( .A1(n14705), .A2(n14704), .ZN(n14706) );
  INV_X1 U16486 ( .A(n19745), .ZN(n17799) );
  INV_X1 U16487 ( .A(n17641), .ZN(n14708) );
  INV_X1 U16488 ( .A(n14707), .ZN(n15263) );
  NAND2_X1 U16489 ( .A1(n14708), .A2(n15263), .ZN(n15210) );
  NAND2_X1 U16490 ( .A1(n15210), .A2(n14419), .ZN(n14709) );
  NAND2_X1 U16491 ( .A1(n17044), .A2(n14710), .ZN(n17034) );
  MUX2_X1 U16492 ( .A(n16969), .B(n15239), .S(n17044), .Z(n14711) );
  OAI21_X1 U16493 ( .B1(n17799), .B2(n17034), .A(n14711), .ZN(P2_U2886) );
  INV_X1 U16494 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14714) );
  AOI22_X1 U16495 ( .A1(n19717), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14712), .ZN(n19690) );
  INV_X1 U16496 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19691) );
  OAI222_X1 U16497 ( .A1(n14715), .A2(n14714), .B1(n14713), .B2(n19690), .C1(
        n14732), .C2(n19691), .ZN(P2_U2982) );
  INV_X1 U16498 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14716) );
  MUX2_X1 U16499 ( .A(n17780), .B(n17754), .S(n14716), .Z(n14726) );
  AOI21_X1 U16500 ( .B1(n14719), .B2(n14718), .A(n14717), .ZN(n17627) );
  INV_X1 U16501 ( .A(n17627), .ZN(n14724) );
  NOR2_X1 U16502 ( .A1(n14721), .A2(n14720), .ZN(n14722) );
  XOR2_X1 U16503 ( .A(n14722), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17635) );
  NAND2_X1 U16504 ( .A1(n17635), .A2(n17785), .ZN(n14723) );
  NAND2_X1 U16505 ( .A1(n19047), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n17629) );
  OAI211_X1 U16506 ( .C1(n14724), .C2(n17770), .A(n14723), .B(n17629), .ZN(
        n14725) );
  AOI211_X1 U16507 ( .C1(n17784), .C2(n17634), .A(n14726), .B(n14725), .ZN(
        n14727) );
  INV_X1 U16508 ( .A(n14727), .ZN(P2_U3013) );
  NAND2_X1 U16509 ( .A1(n17744), .A2(n22440), .ZN(n22814) );
  INV_X1 U16510 ( .A(n22814), .ZN(n14728) );
  OAI21_X1 U16511 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(n14728), .A(n15410), 
        .ZN(n14729) );
  OAI21_X1 U16512 ( .B1(n14730), .B2(n15410), .A(n14729), .ZN(P1_U3487) );
  INV_X1 U16513 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14736) );
  NOR2_X1 U16514 ( .A1(n14731), .A2(n13315), .ZN(n15205) );
  NAND2_X1 U16515 ( .A1(n15205), .A2(n18966), .ZN(n14733) );
  NAND2_X1 U16516 ( .A1(n14733), .A2(n14732), .ZN(n14734) );
  NAND2_X1 U16517 ( .A1(n17823), .A2(n18958), .ZN(n14933) );
  NOR2_X1 U16518 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17693), .ZN(n17841) );
  AOI22_X1 U16519 ( .A1(n17851), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17836), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14735) );
  OAI21_X1 U16520 ( .B1(n14736), .B2(n14933), .A(n14735), .ZN(P2_U2929) );
  INV_X1 U16521 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14738) );
  AOI22_X1 U16522 ( .A1(n17851), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17836), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14737) );
  OAI21_X1 U16523 ( .B1(n14738), .B2(n14933), .A(n14737), .ZN(P2_U2930) );
  INV_X1 U16524 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U16525 ( .A1(n17851), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17836), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14739) );
  OAI21_X1 U16526 ( .B1(n17092), .B2(n14933), .A(n14739), .ZN(P2_U2927) );
  AOI22_X1 U16527 ( .A1(n17851), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17836), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14740) );
  OAI21_X1 U16528 ( .B1(n14741), .B2(n14933), .A(n14740), .ZN(P2_U2926) );
  INV_X1 U16529 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U16530 ( .A1(n17851), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17836), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14742) );
  OAI21_X1 U16531 ( .B1(n17102), .B2(n14933), .A(n14742), .ZN(P2_U2928) );
  NAND2_X1 U16532 ( .A1(n17641), .A2(n15254), .ZN(n15208) );
  NAND2_X1 U16533 ( .A1(n15208), .A2(n14743), .ZN(n14744) );
  NAND2_X1 U16534 ( .A1(n14744), .A2(n18966), .ZN(n14746) );
  AND2_X1 U16535 ( .A1(n14403), .A2(n19213), .ZN(n15269) );
  NAND2_X1 U16536 ( .A1(n18968), .A2(n15269), .ZN(n14745) );
  AND2_X1 U16537 ( .A1(n19929), .A2(n14748), .ZN(n15849) );
  INV_X1 U16538 ( .A(n15849), .ZN(n14749) );
  NAND2_X1 U16539 ( .A1(n17123), .A2(n14749), .ZN(n19972) );
  AND2_X1 U16540 ( .A1(n19876), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14750) );
  OAI211_X1 U16541 ( .C1(n20178), .C2(n14751), .A(n14700), .B(n14750), .ZN(
        n14752) );
  INV_X1 U16542 ( .A(n14752), .ZN(n14753) );
  NOR2_X1 U16543 ( .A1(n14755), .A2(n14754), .ZN(n14756) );
  OR2_X1 U16544 ( .A1(n14757), .A2(n14756), .ZN(n15964) );
  INV_X1 U16545 ( .A(n15964), .ZN(n19190) );
  NOR2_X1 U16546 ( .A1(n19732), .A2(n15964), .ZN(n20172) );
  INV_X1 U16547 ( .A(n20172), .ZN(n14758) );
  NAND2_X1 U16548 ( .A1(n19929), .A2(n13358), .ZN(n20228) );
  OAI211_X1 U16549 ( .C1(n19743), .C2(n19190), .A(n14758), .B(n20123), .ZN(
        n14760) );
  AOI22_X1 U16550 ( .A1(n20169), .A2(n19190), .B1(n20221), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n14759) );
  OAI211_X1 U16551 ( .C1(n20176), .C2(n20235), .A(n14760), .B(n14759), .ZN(
        P2_U2919) );
  MUX2_X1 U16552 ( .A(n13617), .B(n19183), .S(n17044), .Z(n14761) );
  OAI21_X1 U16553 ( .B1(n17034), .B2(n19732), .A(n14761), .ZN(P2_U2887) );
  NOR2_X1 U16554 ( .A1(n14762), .A2(n22234), .ZN(n14763) );
  INV_X1 U16555 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20402) );
  NAND2_X1 U16556 ( .A1(n14764), .A2(n22253), .ZN(n14765) );
  AOI22_X1 U16557 ( .A1(n16588), .A2(BUF1_REG_15__SCAN_IN), .B1(DATAI_15_), 
        .B2(n16592), .ZN(n15953) );
  INV_X1 U16558 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14767) );
  OAI21_X1 U16559 ( .B1(n21857), .B2(n22253), .A(n14766), .ZN(n22387) );
  INV_X1 U16560 ( .A(n22387), .ZN(n22337) );
  OAI222_X1 U16561 ( .A1(n22405), .A2(n20402), .B1(n22399), .B2(n15953), .C1(
        n14767), .C2(n22337), .ZN(P1_U2967) );
  INV_X1 U16562 ( .A(n22253), .ZN(n22254) );
  AOI21_X1 U16563 ( .B1(n14768), .B2(n15391), .A(n22254), .ZN(n14769) );
  NAND2_X1 U16564 ( .A1(n14770), .A2(n14769), .ZN(n14773) );
  OR2_X1 U16565 ( .A1(n14771), .A2(n16422), .ZN(n14772) );
  NAND2_X1 U16566 ( .A1(n14773), .A2(n14772), .ZN(n14892) );
  NAND2_X1 U16567 ( .A1(n16420), .A2(n16422), .ZN(n14774) );
  OAI211_X1 U16568 ( .C1(n14777), .C2(n14776), .A(n14775), .B(n14774), .ZN(
        n14780) );
  NAND3_X1 U16569 ( .A1(n16421), .A2(n22261), .A3(n22253), .ZN(n14778) );
  AOI21_X1 U16570 ( .B1(n16890), .B2(n14785), .A(n14778), .ZN(n14779) );
  NAND2_X1 U16571 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n22224) );
  NOR2_X1 U16572 ( .A1(n22225), .A2(n22224), .ZN(n15109) );
  AND2_X1 U16573 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15109), .ZN(n14781) );
  AOI21_X1 U16574 ( .B1(n15104), .B2(n22809), .A(n14781), .ZN(n17670) );
  NAND2_X1 U16575 ( .A1(n22225), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U16576 ( .A1(n17670), .A2(n14782), .ZN(n17674) );
  INV_X1 U16577 ( .A(n15412), .ZN(n15114) );
  NAND3_X1 U16578 ( .A1(n14783), .A2(n14785), .A3(n14784), .ZN(n14786) );
  NOR2_X1 U16579 ( .A1(n14787), .A2(n14786), .ZN(n14788) );
  NAND2_X1 U16580 ( .A1(n14788), .A2(n15103), .ZN(n16892) );
  INV_X1 U16581 ( .A(n16892), .ZN(n14790) );
  OAI22_X1 U16582 ( .A1(n15114), .A2(n14790), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14789), .ZN(n17720) );
  INV_X1 U16583 ( .A(n17720), .ZN(n14792) );
  INV_X1 U16584 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n22464) );
  AOI22_X1 U16585 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n16895), .B1(n14797), 
        .B2(n22228), .ZN(n14791) );
  OAI21_X1 U16586 ( .B1(n14792), .B2(n17669), .A(n14791), .ZN(n14793) );
  NAND2_X1 U16587 ( .A1(n14793), .A2(n17674), .ZN(n14796) );
  NOR2_X1 U16588 ( .A1(n16890), .A2(n14797), .ZN(n17719) );
  INV_X1 U16589 ( .A(n17669), .ZN(n14794) );
  NAND2_X1 U16590 ( .A1(n17719), .A2(n14794), .ZN(n14795) );
  OAI211_X1 U16591 ( .C1(n17674), .C2(n14797), .A(n14796), .B(n14795), .ZN(
        P1_U3474) );
  OAI21_X1 U16592 ( .B1(n14800), .B2(n14799), .A(n14798), .ZN(n15167) );
  OR2_X1 U16593 ( .A1(n14801), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14802) );
  NAND2_X1 U16594 ( .A1(n14803), .A2(n14802), .ZN(n22011) );
  NAND2_X1 U16595 ( .A1(n21999), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n22017) );
  OAI21_X1 U16596 ( .B1(n20551), .B2(n14804), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14805) );
  OAI211_X1 U16597 ( .C1(n22011), .C2(n22216), .A(n22017), .B(n14805), .ZN(
        n14806) );
  AOI21_X1 U16598 ( .B1(n20557), .B2(n15167), .A(n14806), .ZN(n14807) );
  INV_X1 U16599 ( .A(n14807), .ZN(P1_U2999) );
  INV_X1 U16600 ( .A(n17692), .ZN(n14812) );
  NAND2_X1 U16601 ( .A1(n14846), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19719) );
  NAND2_X1 U16602 ( .A1(n19861), .A2(n19766), .ZN(n14809) );
  NAND2_X1 U16603 ( .A1(n19719), .A2(n14809), .ZN(n19753) );
  NAND2_X1 U16604 ( .A1(n14849), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14810) );
  OAI21_X1 U16605 ( .B1(n19753), .B2(n19908), .A(n14810), .ZN(n14811) );
  NAND2_X1 U16606 ( .A1(n16347), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14814) );
  NAND2_X1 U16607 ( .A1(n14813), .A2(n14814), .ZN(n14817) );
  INV_X1 U16608 ( .A(n14813), .ZN(n14816) );
  INV_X1 U16609 ( .A(n14814), .ZN(n14815) );
  NAND2_X1 U16610 ( .A1(n14817), .A2(n14857), .ZN(n14823) );
  OR2_X1 U16611 ( .A1(n14819), .A2(n14818), .ZN(n14820) );
  NAND2_X1 U16612 ( .A1(n14821), .A2(n14820), .ZN(n14822) );
  NAND2_X1 U16613 ( .A1(n14823), .A2(n14822), .ZN(n14824) );
  MUX2_X1 U16614 ( .A(n13621), .B(n14686), .S(n17044), .Z(n14825) );
  OAI21_X1 U16615 ( .B1(n17805), .B2(n17034), .A(n14825), .ZN(P2_U2885) );
  XNOR2_X1 U16616 ( .A(n14827), .B(n14826), .ZN(n17795) );
  INV_X1 U16617 ( .A(n17795), .ZN(n14830) );
  INV_X1 U16618 ( .A(n14828), .ZN(n14829) );
  OAI22_X1 U16619 ( .A1(n17622), .A2(n14830), .B1(n19193), .B2(n14829), .ZN(
        n14835) );
  NAND2_X1 U16620 ( .A1(n15548), .A2(n15551), .ZN(n14833) );
  INV_X1 U16621 ( .A(n17631), .ZN(n19185) );
  AOI22_X1 U16622 ( .A1(n19185), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n17585), .B2(n14833), .ZN(n14832) );
  OAI211_X1 U16623 ( .C1(n14833), .C2(n17579), .A(n14832), .B(n14831), .ZN(
        n14834) );
  AOI211_X1 U16624 ( .C1(n17636), .C2(n14836), .A(n14835), .B(n14834), .ZN(
        n14837) );
  OAI21_X1 U16625 ( .B1(n14686), .B2(n19184), .A(n14837), .ZN(P2_U3044) );
  XNOR2_X1 U16626 ( .A(n14838), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14905) );
  XOR2_X1 U16627 ( .A(n14840), .B(n14839), .Z(n20462) );
  NOR2_X1 U16628 ( .A1(n21975), .A2(n22031), .ZN(n14902) );
  AOI21_X1 U16629 ( .B1(n20551), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14902), .ZN(n14841) );
  OAI21_X1 U16630 ( .B1(n20561), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14841), .ZN(n14842) );
  AOI21_X1 U16631 ( .B1(n20462), .B2(n20557), .A(n14842), .ZN(n14843) );
  OAI21_X1 U16632 ( .B1(n14905), .B2(n22216), .A(n14843), .ZN(P1_U2998) );
  INV_X1 U16633 ( .A(n14844), .ZN(n14864) );
  NAND2_X1 U16634 ( .A1(n19719), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14847) );
  NAND2_X1 U16635 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19777), .ZN(
        n19847) );
  INV_X1 U16636 ( .A(n19847), .ZN(n14845) );
  NAND2_X1 U16637 ( .A1(n14846), .A2(n14845), .ZN(n19815) );
  NAND2_X1 U16638 ( .A1(n14847), .A2(n19815), .ZN(n14848) );
  AND2_X1 U16639 ( .A1(n14848), .A2(n19880), .ZN(n19756) );
  AOI21_X1 U16640 ( .B1(n14849), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19756), .ZN(n14850) );
  NAND2_X1 U16641 ( .A1(n16347), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14854) );
  INV_X1 U16642 ( .A(n14854), .ZN(n14852) );
  NAND2_X1 U16643 ( .A1(n14855), .A2(n14854), .ZN(n14856) );
  INV_X1 U16644 ( .A(n14862), .ZN(n14860) );
  INV_X1 U16645 ( .A(n14861), .ZN(n14859) );
  NAND2_X1 U16646 ( .A1(n14860), .A2(n14859), .ZN(n14863) );
  INV_X1 U16647 ( .A(n19863), .ZN(n19768) );
  MUX2_X1 U16648 ( .A(n17757), .B(n13623), .S(n15444), .Z(n14865) );
  OAI21_X1 U16649 ( .B1(n19768), .B2(n17034), .A(n14865), .ZN(P2_U2884) );
  XNOR2_X1 U16650 ( .A(n14866), .B(n14867), .ZN(n14916) );
  OR2_X1 U16651 ( .A1(n11858), .A2(n14868), .ZN(n14869) );
  AND2_X1 U16652 ( .A1(n14870), .A2(n14869), .ZN(n14872) );
  OR2_X1 U16653 ( .A1(n14872), .A2(n14871), .ZN(n14874) );
  NAND2_X1 U16654 ( .A1(n14872), .A2(n14871), .ZN(n14873) );
  AND2_X1 U16655 ( .A1(n14874), .A2(n14873), .ZN(n22026) );
  AOI22_X1 U16656 ( .A1(n20551), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21999), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14875) );
  OAI21_X1 U16657 ( .B1(n20561), .B2(n22020), .A(n14875), .ZN(n14876) );
  AOI21_X1 U16658 ( .B1(n22026), .B2(n20557), .A(n14876), .ZN(n14877) );
  OAI21_X1 U16659 ( .B1(n14916), .B2(n22216), .A(n14877), .ZN(P1_U2997) );
  NAND2_X1 U16660 ( .A1(n14878), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14879) );
  INV_X1 U16661 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14883) );
  NOR2_X1 U16662 ( .A1(n16324), .A2(n14883), .ZN(n15329) );
  XNOR2_X1 U16663 ( .A(n15120), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14887) );
  NAND2_X1 U16664 ( .A1(n14938), .A2(n14884), .ZN(n14885) );
  NAND2_X1 U16665 ( .A1(n15118), .A2(n14885), .ZN(n19000) );
  MUX2_X1 U16666 ( .A(n13629), .B(n19000), .S(n17044), .Z(n14886) );
  OAI21_X1 U16667 ( .B1(n14887), .B2(n17034), .A(n14886), .ZN(P2_U2880) );
  NOR2_X1 U16668 ( .A1(n14890), .A2(n14889), .ZN(n14891) );
  OR2_X1 U16669 ( .A1(n14888), .A2(n14891), .ZN(n15355) );
  NAND2_X1 U16670 ( .A1(n14892), .A2(n22809), .ZN(n14894) );
  INV_X1 U16671 ( .A(n15309), .ZN(n16596) );
  NAND4_X1 U16672 ( .A1(n14550), .A2(n16596), .A3(n22809), .A4(n11922), .ZN(
        n15306) );
  OR2_X1 U16673 ( .A1(n14783), .A2(n15306), .ZN(n14893) );
  NAND2_X1 U16674 ( .A1(n14895), .A2(n15309), .ZN(n14896) );
  INV_X1 U16675 ( .A(n14896), .ZN(n14897) );
  OAI22_X1 U16676 ( .A1(n16592), .A2(BUF1_REG_3__SCAN_IN), .B1(DATAI_3_), .B2(
        n16588), .ZN(n22328) );
  INV_X1 U16677 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n22333) );
  OAI222_X1 U16678 ( .A1(n15355), .A2(n16667), .B1(n15954), .B2(n22328), .C1(
        n16659), .C2(n22333), .ZN(P1_U2901) );
  INV_X1 U16679 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14899) );
  AOI22_X1 U16680 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17850), .B1(n17851), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14898) );
  OAI21_X1 U16681 ( .B1(n14899), .B2(n14933), .A(n14898), .ZN(P2_U2935) );
  NAND2_X1 U16682 ( .A1(n16895), .A2(n16851), .ZN(n14912) );
  INV_X1 U16683 ( .A(n14900), .ZN(n16857) );
  NAND2_X1 U16684 ( .A1(n16788), .A2(n16857), .ZN(n22013) );
  AOI21_X1 U16685 ( .B1(n16895), .B2(n22013), .A(n16854), .ZN(n14901) );
  INV_X1 U16686 ( .A(n14901), .ZN(n22014) );
  OAI222_X1 U16687 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16798), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14912), .C1(n16893), .C2(
        n22014), .ZN(n14904) );
  XNOR2_X1 U16688 ( .A(n16184), .B(n15304), .ZN(n20461) );
  AOI21_X1 U16689 ( .B1(n21993), .B2(n20461), .A(n14902), .ZN(n14903) );
  OAI211_X1 U16690 ( .C1(n14905), .C2(n22010), .A(n14904), .B(n14903), .ZN(
        P1_U3030) );
  OR2_X1 U16691 ( .A1(n14907), .A2(n14906), .ZN(n14908) );
  AND2_X1 U16692 ( .A1(n15353), .A2(n14908), .ZN(n22019) );
  INV_X1 U16693 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n22032) );
  NOR2_X1 U16694 ( .A1(n21975), .A2(n22032), .ZN(n14911) );
  NAND2_X1 U16695 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14909) );
  AOI221_X1 U16696 ( .B1(n15361), .B2(n15363), .C1(n14909), .C2(n15363), .A(
        n16788), .ZN(n14910) );
  AOI211_X1 U16697 ( .C1(n21993), .C2(n22019), .A(n14911), .B(n14910), .ZN(
        n14915) );
  OAI21_X1 U16698 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21922), .A(
        n21920), .ZN(n15365) );
  NAND2_X1 U16699 ( .A1(n16793), .A2(n14912), .ZN(n16786) );
  OAI21_X1 U16700 ( .B1(n16893), .B2(n16786), .A(n15361), .ZN(n14913) );
  OAI21_X1 U16701 ( .B1(n15361), .B2(n15365), .A(n14913), .ZN(n14914) );
  OAI211_X1 U16702 ( .C1(n22010), .C2(n14916), .A(n14915), .B(n14914), .ZN(
        P1_U3029) );
  INV_X1 U16703 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14918) );
  AOI22_X1 U16704 ( .A1(n17851), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14917) );
  OAI21_X1 U16705 ( .B1(n14918), .B2(n14933), .A(n14917), .ZN(P2_U2931) );
  AOI22_X1 U16706 ( .A1(n17851), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14919) );
  OAI21_X1 U16707 ( .B1(n14920), .B2(n14933), .A(n14919), .ZN(P2_U2924) );
  AOI22_X1 U16708 ( .A1(n17851), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14921) );
  OAI21_X1 U16709 ( .B1(n17048), .B2(n14933), .A(n14921), .ZN(P2_U2922) );
  AOI22_X1 U16710 ( .A1(n17851), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14922) );
  OAI21_X1 U16711 ( .B1(n14923), .B2(n14933), .A(n14922), .ZN(P2_U2925) );
  AOI22_X1 U16712 ( .A1(n17851), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14924) );
  OAI21_X1 U16713 ( .B1(n14925), .B2(n14933), .A(n14924), .ZN(P2_U2923) );
  INV_X1 U16714 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14927) );
  AOI22_X1 U16715 ( .A1(n17841), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14926) );
  OAI21_X1 U16716 ( .B1(n14927), .B2(n14933), .A(n14926), .ZN(P2_U2933) );
  INV_X1 U16717 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14929) );
  AOI22_X1 U16718 ( .A1(n17841), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14928) );
  OAI21_X1 U16719 ( .B1(n14929), .B2(n14933), .A(n14928), .ZN(P2_U2934) );
  INV_X1 U16720 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14931) );
  AOI22_X1 U16721 ( .A1(n17841), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14930) );
  OAI21_X1 U16722 ( .B1(n14931), .B2(n14933), .A(n14930), .ZN(P2_U2932) );
  AOI22_X1 U16723 ( .A1(n17841), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14932) );
  OAI21_X1 U16724 ( .B1(n14934), .B2(n14933), .A(n14932), .ZN(P2_U2921) );
  NOR2_X1 U16725 ( .A1(n16011), .A2(n16214), .ZN(n14936) );
  INV_X1 U16726 ( .A(n15120), .ZN(n14935) );
  INV_X1 U16727 ( .A(n17034), .ZN(n17039) );
  OAI211_X1 U16728 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14936), .A(
        n14935), .B(n17039), .ZN(n14941) );
  OAI21_X1 U16729 ( .B1(n14939), .B2(n14937), .A(n14938), .ZN(n17772) );
  INV_X1 U16730 ( .A(n17772), .ZN(n18990) );
  NAND2_X1 U16731 ( .A1(n17044), .A2(n18990), .ZN(n14940) );
  OAI211_X1 U16732 ( .C1(n17044), .C2(n14942), .A(n14941), .B(n14940), .ZN(
        P2_U2881) );
  INV_X1 U16733 ( .A(n14943), .ZN(n14945) );
  NAND2_X1 U16734 ( .A1(n14945), .A2(n14944), .ZN(n14946) );
  NAND2_X1 U16735 ( .A1(n14947), .A2(n14946), .ZN(n20168) );
  INV_X1 U16736 ( .A(n20168), .ZN(n14948) );
  XNOR2_X1 U16737 ( .A(n19745), .B(n20168), .ZN(n20171) );
  NOR2_X1 U16738 ( .A1(n20171), .A2(n20172), .ZN(n20170) );
  AOI21_X1 U16739 ( .B1(n14948), .B2(n17799), .A(n20170), .ZN(n15323) );
  XNOR2_X1 U16740 ( .A(n15323), .B(n17795), .ZN(n15325) );
  XNOR2_X1 U16741 ( .A(n15325), .B(n17805), .ZN(n14951) );
  AOI22_X1 U16742 ( .A1(n20169), .A2(n17795), .B1(n20221), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n14950) );
  INV_X1 U16743 ( .A(n20128), .ZN(n20120) );
  NAND2_X1 U16744 ( .A1(n19972), .A2(n20120), .ZN(n14949) );
  OAI211_X1 U16745 ( .C1(n14951), .C2(n20228), .A(n14950), .B(n14949), .ZN(
        P2_U2917) );
  OAI21_X1 U16746 ( .B1(n14888), .B2(n14953), .A(n14952), .ZN(n22059) );
  OAI22_X1 U16747 ( .A1(n16592), .A2(BUF1_REG_4__SCAN_IN), .B1(DATAI_4_), .B2(
        n16588), .ZN(n22334) );
  INV_X1 U16748 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n22340) );
  OAI222_X1 U16749 ( .A1(n22059), .A2(n16667), .B1(n15954), .B2(n22334), .C1(
        n22340), .C2(n16659), .ZN(P1_U2900) );
  XNOR2_X1 U16750 ( .A(n14954), .B(n14955), .ZN(n21872) );
  INV_X1 U16751 ( .A(n15355), .ZN(n22045) );
  AOI22_X1 U16752 ( .A1(n20551), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n22170), .ZN(n14956) );
  OAI21_X1 U16753 ( .B1(n20561), .B2(n22043), .A(n14956), .ZN(n14957) );
  AOI21_X1 U16754 ( .B1(n22045), .B2(n20557), .A(n14957), .ZN(n14958) );
  OAI21_X1 U16755 ( .B1(n21872), .B2(n22216), .A(n14958), .ZN(P1_U2996) );
  INV_X2 U16756 ( .A(n18010), .ZN(n18255) );
  AOI22_X1 U16757 ( .A1(n18323), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14963) );
  NOR2_X2 U16758 ( .A1(n14965), .A2(n14967), .ZN(n15006) );
  AOI22_X1 U16759 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14962) );
  AOI22_X1 U16760 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14961) );
  AND2_X2 U16761 ( .A1(n21361), .A2(n20710), .ZN(n18321) );
  AOI22_X1 U16762 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14960) );
  NAND4_X1 U16763 ( .A1(n14963), .A2(n14962), .A3(n14961), .A4(n14960), .ZN(
        n14973) );
  NOR2_X2 U16764 ( .A1(n21344), .A2(n14965), .ZN(n14985) );
  NOR2_X2 U16765 ( .A1(n14965), .A2(n14964), .ZN(n18026) );
  AOI22_X1 U16766 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11160), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14971) );
  AOI22_X1 U16767 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14970) );
  AOI22_X1 U16768 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14969) );
  AOI22_X1 U16769 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14968) );
  NAND4_X1 U16770 ( .A1(n14971), .A2(n14970), .A3(n14969), .A4(n14968), .ZN(
        n14972) );
  AOI22_X1 U16771 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14977) );
  AOI22_X1 U16772 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14976) );
  AOI22_X1 U16773 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14975) );
  AOI22_X1 U16774 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14974) );
  NAND4_X1 U16775 ( .A1(n14977), .A2(n14976), .A3(n14975), .A4(n14974), .ZN(
        n14983) );
  AOI22_X1 U16776 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18335), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14981) );
  AOI22_X1 U16777 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14980) );
  AOI22_X1 U16778 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14979) );
  AOI22_X1 U16779 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18323), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14978) );
  NAND4_X1 U16780 ( .A1(n14981), .A2(n14980), .A3(n14979), .A4(n14978), .ZN(
        n14982) );
  AOI22_X1 U16781 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14995) );
  AOI22_X1 U16782 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14994) );
  INV_X1 U16783 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19686) );
  AOI22_X1 U16784 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14987) );
  OAI21_X1 U16785 ( .B1(n18099), .B2(n19686), .A(n14987), .ZN(n14993) );
  AOI22_X1 U16786 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U16787 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14991) );
  AOI22_X1 U16788 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14990) );
  AOI22_X1 U16789 ( .A1(n20722), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14989) );
  AOI22_X1 U16790 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18335), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15005) );
  AOI22_X1 U16791 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15004) );
  INV_X1 U16792 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19452) );
  AOI22_X1 U16793 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14996) );
  OAI21_X1 U16794 ( .B1(n18099), .B2(n19452), .A(n14996), .ZN(n15002) );
  AOI22_X1 U16795 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11161), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15000) );
  AOI22_X1 U16796 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14999) );
  AOI22_X1 U16797 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14998) );
  AOI22_X1 U16798 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14997) );
  NAND4_X1 U16799 ( .A1(n15000), .A2(n14999), .A3(n14998), .A4(n14997), .ZN(
        n15001) );
  AOI211_X1 U16800 ( .C1(n18347), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n15002), .B(n15001), .ZN(n15003) );
  NAND3_X1 U16801 ( .A1(n15005), .A2(n15004), .A3(n15003), .ZN(n15988) );
  AOI22_X1 U16802 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15010) );
  AOI22_X1 U16803 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15009) );
  AOI22_X1 U16804 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U16805 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15007) );
  NAND4_X1 U16806 ( .A1(n15010), .A2(n15009), .A3(n15008), .A4(n15007), .ZN(
        n15016) );
  AOI22_X1 U16807 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15014) );
  AOI22_X1 U16808 ( .A1(n18323), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15013) );
  AOI22_X1 U16809 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15012) );
  AOI22_X1 U16810 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15011) );
  NAND4_X1 U16811 ( .A1(n15014), .A2(n15013), .A3(n15012), .A4(n15011), .ZN(
        n15015) );
  AOI22_X1 U16812 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15025) );
  AOI22_X1 U16813 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15024) );
  INV_X1 U16814 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19411) );
  AOI22_X1 U16815 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15017) );
  OAI21_X1 U16816 ( .B1(n18099), .B2(n19411), .A(n15017), .ZN(n15023) );
  AOI22_X1 U16817 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U16818 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U16819 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15019) );
  AOI22_X1 U16820 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15018) );
  NAND4_X1 U16821 ( .A1(n15021), .A2(n15020), .A3(n15019), .A4(n15018), .ZN(
        n15022) );
  AOI22_X1 U16822 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15033) );
  AOI22_X1 U16823 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15032) );
  AOI22_X1 U16824 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15026) );
  OAI21_X1 U16825 ( .B1(n18099), .B2(n19534), .A(n15026), .ZN(n15031) );
  AOI22_X1 U16826 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15030) );
  AOI22_X1 U16827 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15029) );
  AOI22_X1 U16828 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15028) );
  AOI22_X1 U16829 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15027) );
  AOI22_X1 U16830 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15037) );
  AOI22_X1 U16831 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15036) );
  AOI22_X1 U16832 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15035) );
  AOI22_X1 U16833 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15034) );
  NAND4_X1 U16834 ( .A1(n15037), .A2(n15036), .A3(n15035), .A4(n15034), .ZN(
        n15043) );
  AOI22_X1 U16835 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15041) );
  AOI22_X1 U16836 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15040) );
  AOI22_X1 U16837 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15039) );
  AOI22_X1 U16838 ( .A1(n18323), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15038) );
  NAND4_X1 U16839 ( .A1(n15041), .A2(n15040), .A3(n15039), .A4(n15038), .ZN(
        n15042) );
  NAND2_X1 U16840 ( .A1(n21369), .A2(n19455), .ZN(n21320) );
  NOR3_X1 U16841 ( .A1(n21179), .A2(n15988), .A3(n15978), .ZN(n15057) );
  NOR2_X1 U16842 ( .A1(n21366), .A2(n15988), .ZN(n16006) );
  NOR2_X1 U16843 ( .A1(n15979), .A2(n21366), .ZN(n21373) );
  AOI21_X1 U16844 ( .B1(n16006), .B2(n15999), .A(n21373), .ZN(n15044) );
  INV_X1 U16845 ( .A(n15044), .ZN(n15990) );
  NAND2_X1 U16846 ( .A1(n21180), .A2(n15988), .ZN(n21321) );
  INV_X1 U16847 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21819) );
  OAI22_X1 U16848 ( .A1(n21342), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n21815), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15050) );
  NAND2_X1 U16849 ( .A1(n21806), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15993) );
  OAI22_X1 U16850 ( .A1(n21324), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n21809), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15994) );
  NOR2_X1 U16851 ( .A1(n15993), .A2(n15994), .ZN(n15045) );
  AOI21_X1 U16852 ( .B1(n21809), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n15045), .ZN(n15051) );
  OAI21_X1 U16853 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21342), .A(
        n15046), .ZN(n15047) );
  OAI22_X1 U16854 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21819), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n15047), .ZN(n15053) );
  NOR2_X1 U16855 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21819), .ZN(
        n15048) );
  NAND2_X1 U16856 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n15047), .ZN(
        n15052) );
  AOI22_X1 U16857 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15053), .B1(
        n15048), .B2(n15052), .ZN(n15056) );
  OAI21_X1 U16858 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21806), .A(
        n15993), .ZN(n18397) );
  NOR2_X1 U16859 ( .A1(n15994), .A2(n18397), .ZN(n15055) );
  OAI21_X1 U16860 ( .B1(n15051), .B2(n15050), .A(n15056), .ZN(n15049) );
  AOI21_X1 U16861 ( .B1(n15051), .B2(n15050), .A(n15049), .ZN(n18399) );
  INV_X1 U16862 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21802) );
  AND2_X1 U16863 ( .A1(n15052), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15054) );
  OAI22_X1 U16864 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21802), .B1(
        n15054), .B2(n15053), .ZN(n15995) );
  INV_X1 U16865 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20629) );
  NAND2_X1 U16866 ( .A1(n21314), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n21830) );
  NOR2_X1 U16867 ( .A1(n20629), .A2(n21830), .ZN(n21826) );
  OAI221_X1 U16868 ( .B1(n15057), .B2(n18393), .C1(n15057), .C2(n21790), .A(
        n21826), .ZN(n21114) );
  INV_X1 U16869 ( .A(n18273), .ZN(n18265) );
  NOR2_X1 U16870 ( .A1(n21179), .A2(n18265), .ZN(n18270) );
  INV_X1 U16871 ( .A(n18270), .ZN(n18269) );
  NOR2_X2 U16872 ( .A1(n18265), .A2(n21219), .ZN(n18271) );
  INV_X1 U16873 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20802) );
  INV_X1 U16874 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20768) );
  INV_X1 U16875 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20704) );
  NAND2_X1 U16876 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18267) );
  NOR2_X1 U16877 ( .A1(n20704), .A2(n18267), .ZN(n17910) );
  NAND3_X1 U16878 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17910), .ZN(n17909) );
  INV_X1 U16879 ( .A(n17909), .ZN(n17935) );
  AND3_X1 U16880 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17935), .ZN(n18040) );
  NAND2_X1 U16881 ( .A1(n18273), .A2(n18040), .ZN(n17929) );
  NOR2_X1 U16882 ( .A1(n20768), .A2(n17929), .ZN(n17932) );
  NAND2_X1 U16883 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17932), .ZN(n18033) );
  NOR2_X1 U16884 ( .A1(n20802), .A2(n18033), .ZN(n18008) );
  AND2_X1 U16885 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18008), .ZN(n18006) );
  NAND2_X1 U16886 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n18006), .ZN(n17991) );
  INV_X1 U16887 ( .A(n17991), .ZN(n17990) );
  NAND2_X1 U16888 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17990), .ZN(n17939) );
  NAND2_X1 U16889 ( .A1(n18268), .A2(n17939), .ZN(n17977) );
  OAI21_X1 U16890 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n18269), .A(n17977), .ZN(
        n15069) );
  AOI22_X1 U16891 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15068) );
  AOI22_X1 U16892 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15067) );
  INV_X1 U16893 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19371) );
  AOI22_X1 U16894 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15059) );
  OAI21_X1 U16895 ( .B1(n18010), .B2(n19371), .A(n15059), .ZN(n15065) );
  AOI22_X1 U16896 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15063) );
  AOI22_X1 U16897 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15062) );
  AOI22_X1 U16898 ( .A1(n11160), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15061) );
  AOI22_X1 U16899 ( .A1(n18321), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15060) );
  NAND4_X1 U16900 ( .A1(n15063), .A2(n15062), .A3(n15061), .A4(n15060), .ZN(
        n15064) );
  AOI211_X1 U16901 ( .C1(n11164), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n15065), .B(n15064), .ZN(n15066) );
  NAND3_X1 U16902 ( .A1(n15068), .A2(n15067), .A3(n15066), .ZN(n21277) );
  AOI22_X1 U16903 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n15069), .B1(n18271), 
        .B2(n21277), .ZN(n15073) );
  INV_X1 U16904 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n15071) );
  NAND3_X1 U16905 ( .A1(n21219), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17990), 
        .ZN(n17978) );
  INV_X1 U16906 ( .A(n17978), .ZN(n15070) );
  NAND3_X1 U16907 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n15071), .A3(n15070), 
        .ZN(n15072) );
  NAND2_X1 U16908 ( .A1(n15073), .A2(n15072), .ZN(P3_U2689) );
  XNOR2_X1 U16909 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15078) );
  NOR2_X1 U16910 ( .A1(n15411), .A2(n21857), .ZN(n16428) );
  NAND2_X1 U16911 ( .A1(n15075), .A2(n16428), .ZN(n15081) );
  XNOR2_X1 U16912 ( .A(n15076), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16901) );
  MUX2_X1 U16913 ( .A(n15092), .B(n15081), .S(n16901), .Z(n15077) );
  OAI21_X1 U16914 ( .B1(n16890), .B2(n15078), .A(n15077), .ZN(n15079) );
  AOI21_X1 U16915 ( .B1(n15074), .B2(n16892), .A(n15079), .ZN(n16906) );
  MUX2_X1 U16916 ( .A(n11775), .B(n16906), .S(n15104), .Z(n17727) );
  INV_X1 U16917 ( .A(n17727), .ZN(n15097) );
  NAND2_X1 U16918 ( .A1(n22041), .A2(n16892), .ZN(n15096) );
  AND2_X1 U16919 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15084) );
  INV_X1 U16920 ( .A(n15084), .ZN(n15083) );
  NOR2_X1 U16921 ( .A1(n15076), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15082) );
  OAI22_X1 U16922 ( .A1(n16890), .A2(n15083), .B1(n15082), .B2(n15081), .ZN(
        n15086) );
  NOR2_X1 U16923 ( .A1(n16890), .A2(n15084), .ZN(n15085) );
  MUX2_X1 U16924 ( .A(n15086), .B(n15085), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15094) );
  INV_X1 U16925 ( .A(n15090), .ZN(n15087) );
  OAI21_X1 U16926 ( .B1(n15076), .B2(n15088), .A(n15087), .ZN(n15089) );
  NOR2_X1 U16927 ( .A1(n15089), .A2(n11370), .ZN(n16910) );
  INV_X1 U16928 ( .A(n15076), .ZN(n16887) );
  NAND2_X1 U16929 ( .A1(n16887), .A2(n15090), .ZN(n15091) );
  OAI21_X1 U16930 ( .B1(n15092), .B2(n16910), .A(n15091), .ZN(n15093) );
  NOR2_X1 U16931 ( .A1(n15094), .A2(n15093), .ZN(n15095) );
  NAND2_X1 U16932 ( .A1(n15096), .A2(n15095), .ZN(n16908) );
  MUX2_X1 U16933 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16908), .S(
        n15104), .Z(n17728) );
  NAND3_X1 U16934 ( .A1(n15097), .A2(n17728), .A3(n17744), .ZN(n15100) );
  NOR2_X1 U16935 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n17744), .ZN(n15105) );
  NAND2_X1 U16936 ( .A1(n15098), .A2(n15105), .ZN(n15099) );
  INV_X1 U16937 ( .A(n15133), .ZN(n15288) );
  OR2_X1 U16938 ( .A1(n15101), .A2(n15288), .ZN(n15102) );
  XNOR2_X1 U16939 ( .A(n15102), .B(n17673), .ZN(n22051) );
  OR2_X1 U16940 ( .A1(n22051), .A2(n15103), .ZN(n17671) );
  NAND2_X1 U16941 ( .A1(n17671), .A2(n15104), .ZN(n15108) );
  INV_X1 U16942 ( .A(n15104), .ZN(n17722) );
  AOI21_X1 U16943 ( .B1(n17722), .B2(n17673), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n15107) );
  AND2_X1 U16944 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15105), .ZN(
        n15106) );
  AOI21_X1 U16945 ( .B1(n15108), .B2(n15107), .A(n15106), .ZN(n17738) );
  OAI21_X1 U16946 ( .B1(n17739), .B2(n16896), .A(n17738), .ZN(n15111) );
  OAI21_X1 U16947 ( .B1(n15111), .B2(P1_FLUSH_REG_SCAN_IN), .A(n15109), .ZN(
        n15110) );
  NAND2_X1 U16948 ( .A1(n15110), .A2(n22411), .ZN(n17747) );
  NOR2_X1 U16949 ( .A1(n15111), .A2(n22224), .ZN(n22232) );
  NAND2_X1 U16950 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22464), .ZN(n15158) );
  INV_X1 U16951 ( .A(n15158), .ZN(n15113) );
  OAI22_X1 U16952 ( .A1(n15112), .A2(n22497), .B1(n15114), .B2(n15113), .ZN(
        n15115) );
  OAI21_X1 U16953 ( .B1(n22232), .B2(n15115), .A(n17747), .ZN(n15116) );
  OAI21_X1 U16954 ( .B1(n17747), .B2(n22485), .A(n15116), .ZN(P1_U3478) );
  NAND2_X1 U16955 ( .A1(n15118), .A2(n15117), .ZN(n15119) );
  AND2_X1 U16956 ( .A1(n15154), .A2(n15119), .ZN(n17783) );
  INV_X1 U16957 ( .A(n17783), .ZN(n15843) );
  INV_X1 U16958 ( .A(n15346), .ZN(n15121) );
  OR2_X1 U16959 ( .A1(n15346), .A2(n15342), .ZN(n15182) );
  OAI211_X1 U16960 ( .C1(n15121), .C2(n15343), .A(n17039), .B(n15182), .ZN(
        n15123) );
  NAND2_X1 U16961 ( .A1(n15444), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n15122) );
  OAI211_X1 U16962 ( .C1(n15843), .C2(n15444), .A(n15123), .B(n15122), .ZN(
        P2_U2879) );
  INV_X1 U16963 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n22318) );
  NAND2_X1 U16964 ( .A1(n15125), .A2(n15124), .ZN(n15126) );
  NAND2_X1 U16965 ( .A1(n20381), .A2(n15127), .ZN(n15576) );
  NOR2_X1 U16966 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22224), .ZN(n20390) );
  AOI22_X1 U16967 ( .A1(n20390), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20393), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n15128) );
  OAI21_X1 U16968 ( .B1(n22318), .B2(n15576), .A(n15128), .ZN(P1_U2919) );
  INV_X1 U16969 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n22324) );
  AOI22_X1 U16970 ( .A1(n21862), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20393), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n15129) );
  OAI21_X1 U16971 ( .B1(n22324), .B2(n15576), .A(n15129), .ZN(P1_U2918) );
  NAND2_X1 U16972 ( .A1(n14952), .A2(n15130), .ZN(n15131) );
  AND2_X1 U16973 ( .A1(n15298), .A2(n15131), .ZN(n22070) );
  INV_X1 U16974 ( .A(n22070), .ZN(n15482) );
  OAI22_X1 U16975 ( .A1(n16592), .A2(BUF1_REG_5__SCAN_IN), .B1(DATAI_5_), .B2(
        n16588), .ZN(n22341) );
  OAI222_X1 U16976 ( .A1(n15482), .A2(n16667), .B1(n15954), .B2(n22341), .C1(
        n16659), .C2(n12160), .ZN(P1_U2899) );
  NAND2_X1 U16977 ( .A1(n15436), .A2(n22427), .ZN(n22804) );
  INV_X1 U16978 ( .A(n15498), .ZN(n15463) );
  OAI21_X1 U16979 ( .B1(n15639), .B2(n22791), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15135) );
  NAND2_X1 U16980 ( .A1(n15074), .A2(n15133), .ZN(n22501) );
  INV_X1 U16981 ( .A(n22501), .ZN(n15430) );
  INV_X1 U16982 ( .A(n22430), .ZN(n22500) );
  NAND2_X1 U16983 ( .A1(n15430), .A2(n22500), .ZN(n15139) );
  AOI21_X1 U16984 ( .B1(n15135), .B2(n15139), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15137) );
  INV_X1 U16985 ( .A(n15138), .ZN(n15136) );
  NOR2_X1 U16986 ( .A1(n15136), .A2(n21855), .ZN(n22481) );
  NOR2_X1 U16987 ( .A1(n22481), .A2(n22411), .ZN(n22509) );
  INV_X1 U16988 ( .A(n22432), .ZN(n15291) );
  NAND2_X1 U16989 ( .A1(n15291), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22480) );
  NAND2_X1 U16990 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22480), .ZN(n22486) );
  OAI211_X1 U16991 ( .C1(n15137), .C2(n22729), .A(n22509), .B(n22486), .ZN(
        n22733) );
  INV_X1 U16992 ( .A(n22733), .ZN(n15643) );
  INV_X1 U16993 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15146) );
  OAI22_X1 U16994 ( .A1(n16592), .A2(BUF1_REG_7__SCAN_IN), .B1(DATAI_7_), .B2(
        n16588), .ZN(n22352) );
  INV_X1 U16995 ( .A(n22352), .ZN(n16626) );
  NAND2_X1 U16996 ( .A1(n22626), .A2(n16626), .ZN(n22787) );
  NOR2_X1 U16997 ( .A1(n15138), .A2(n21855), .ZN(n22503) );
  INV_X1 U16998 ( .A(n22503), .ZN(n15292) );
  OAI22_X1 U16999 ( .A1(n15139), .A2(n22497), .B1(n15292), .B2(n22480), .ZN(
        n22731) );
  INV_X1 U17000 ( .A(DATAI_31_), .ZN(n15140) );
  NAND2_X1 U17001 ( .A1(n16592), .A2(n20557), .ZN(n22632) );
  INV_X1 U17002 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20625) );
  OAI22_X1 U17003 ( .A1(n15140), .A2(n22632), .B1(n20625), .B2(n22630), .ZN(
        n22782) );
  AOI22_X1 U17004 ( .A1(n22799), .A2(n22731), .B1(n22791), .B2(n11345), .ZN(
        n15145) );
  INV_X1 U17005 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20610) );
  INV_X1 U17006 ( .A(DATAI_23_), .ZN(n16624) );
  OR2_X1 U17007 ( .A1(n22632), .A2(n16624), .ZN(n15141) );
  NOR2_X2 U17008 ( .A1(n22629), .A2(n16596), .ZN(n22797) );
  AOI22_X1 U17009 ( .A1(n15639), .A2(n15142), .B1(n22729), .B2(n22797), .ZN(
        n15144) );
  OAI211_X1 U17010 ( .C1(n15643), .C2(n15146), .A(n15145), .B(n15144), .ZN(
        P1_U3152) );
  INV_X1 U17011 ( .A(n20462), .ZN(n15149) );
  INV_X1 U17012 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20569) );
  AOI22_X1 U17013 ( .A1(n16588), .A2(n20569), .B1(n15147), .B2(n16592), .ZN(
        n22315) );
  AOI22_X1 U17014 ( .A1(n15948), .A2(n22315), .B1(n16653), .B2(
        P1_EAX_REG_1__SCAN_IN), .ZN(n15148) );
  OAI21_X1 U17015 ( .B1(n15149), .B2(n16667), .A(n15148), .ZN(P1_U2903) );
  INV_X1 U17016 ( .A(n22026), .ZN(n15152) );
  INV_X1 U17017 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20571) );
  INV_X1 U17018 ( .A(DATAI_2_), .ZN(n15150) );
  AOI22_X1 U17019 ( .A1(n16588), .A2(n20571), .B1(n15150), .B2(n16592), .ZN(
        n22555) );
  AOI22_X1 U17020 ( .A1(n15948), .A2(n22555), .B1(n16653), .B2(
        P1_EAX_REG_2__SCAN_IN), .ZN(n15151) );
  OAI21_X1 U17021 ( .B1(n15152), .B2(n16667), .A(n15151), .ZN(P1_U2902) );
  XOR2_X1 U17022 ( .A(n15181), .B(n15182), .Z(n15157) );
  AND2_X1 U17023 ( .A1(n15154), .A2(n15153), .ZN(n15155) );
  OR2_X1 U17024 ( .A1(n15155), .A2(n15178), .ZN(n17559) );
  MUX2_X1 U17025 ( .A(n13630), .B(n17559), .S(n17044), .Z(n15156) );
  OAI21_X1 U17026 ( .B1(n15157), .B2(n17034), .A(n15156), .ZN(P2_U2878) );
  NAND2_X1 U17027 ( .A1(n17747), .A2(n15158), .ZN(n16182) );
  INV_X1 U17028 ( .A(n15074), .ZN(n22024) );
  NAND2_X1 U17029 ( .A1(n17747), .A2(n22440), .ZN(n15168) );
  INV_X1 U17030 ( .A(n15172), .ZN(n15286) );
  NAND2_X1 U17031 ( .A1(n16178), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22441) );
  XNOR2_X1 U17032 ( .A(n15286), .B(n22441), .ZN(n15159) );
  OAI222_X1 U17033 ( .A1(n16182), .A2(n22024), .B1(n17747), .B2(n12665), .C1(
        n15168), .C2(n15159), .ZN(P1_U3476) );
  XNOR2_X1 U17034 ( .A(n15161), .B(n15160), .ZN(n15371) );
  INV_X1 U17035 ( .A(n22059), .ZN(n15165) );
  INV_X1 U17036 ( .A(n15162), .ZN(n22057) );
  NOR2_X1 U17037 ( .A1(n21975), .A2(n22055), .ZN(n15368) );
  AOI21_X1 U17038 ( .B1(n20551), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n15368), .ZN(n15163) );
  OAI21_X1 U17039 ( .B1(n20561), .B2(n22057), .A(n15163), .ZN(n15164) );
  AOI21_X1 U17040 ( .B1(n15165), .B2(n20557), .A(n15164), .ZN(n15166) );
  OAI21_X1 U17041 ( .B1(n15371), .B2(n22216), .A(n15166), .ZN(P1_U2995) );
  INV_X1 U17042 ( .A(n15167), .ZN(n15415) );
  OAI22_X1 U17043 ( .A1(n16592), .A2(BUF1_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        n16588), .ZN(n22410) );
  INV_X1 U17044 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n22314) );
  OAI222_X1 U17045 ( .A1(n16667), .A2(n15415), .B1(n15954), .B2(n22410), .C1(
        n16659), .C2(n22314), .ZN(P1_U2904) );
  INV_X1 U17046 ( .A(n22041), .ZN(n15176) );
  INV_X1 U17047 ( .A(n15168), .ZN(n16177) );
  INV_X1 U17048 ( .A(n15285), .ZN(n15169) );
  NAND2_X1 U17049 ( .A1(n15169), .A2(n21856), .ZN(n15173) );
  OR2_X1 U17050 ( .A1(n16178), .A2(n21856), .ZN(n15495) );
  INV_X1 U17051 ( .A(n15495), .ZN(n15170) );
  NAND2_X1 U17052 ( .A1(n15436), .A2(n15170), .ZN(n15431) );
  NAND2_X1 U17053 ( .A1(n15172), .A2(n15171), .ZN(n15471) );
  OR2_X1 U17054 ( .A1(n15471), .A2(n22441), .ZN(n15468) );
  NAND4_X1 U17055 ( .A1(n15499), .A2(n15173), .A3(n15431), .A4(n15468), .ZN(
        n15174) );
  INV_X1 U17056 ( .A(n17747), .ZN(n16179) );
  AOI22_X1 U17057 ( .A1(n16177), .A2(n15174), .B1(n16179), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15175) );
  OAI21_X1 U17058 ( .B1(n15176), .B2(n16182), .A(n15175), .ZN(P1_U3475) );
  OR2_X1 U17059 ( .A1(n15178), .A2(n15177), .ZN(n15179) );
  AND2_X1 U17060 ( .A1(n15179), .A2(n15188), .ZN(n17310) );
  INV_X1 U17061 ( .A(n17310), .ZN(n17544) );
  INV_X1 U17062 ( .A(n15181), .ZN(n15180) );
  NOR2_X1 U17063 ( .A1(n15182), .A2(n15180), .ZN(n15184) );
  NAND2_X1 U17064 ( .A1(n15181), .A2(n15183), .ZN(n15340) );
  OR2_X1 U17065 ( .A1(n15182), .A2(n15340), .ZN(n15338) );
  OAI211_X1 U17066 ( .C1(n15184), .C2(n15183), .A(n17039), .B(n15338), .ZN(
        n15186) );
  NAND2_X1 U17067 ( .A1(n15444), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15185) );
  OAI211_X1 U17068 ( .C1(n17544), .C2(n15444), .A(n15186), .B(n15185), .ZN(
        P2_U2877) );
  INV_X1 U17069 ( .A(n15339), .ZN(n15337) );
  XNOR2_X1 U17070 ( .A(n15338), .B(n15337), .ZN(n15191) );
  NAND2_X1 U17071 ( .A1(n15188), .A2(n15187), .ZN(n15189) );
  AND2_X1 U17072 ( .A1(n15335), .A2(n15189), .ZN(n17534) );
  INV_X1 U17073 ( .A(n17534), .ZN(n15912) );
  MUX2_X1 U17074 ( .A(n15912), .B(n13632), .S(n15444), .Z(n15190) );
  OAI21_X1 U17075 ( .B1(n15191), .B2(n17034), .A(n15190), .ZN(P2_U2876) );
  OR2_X1 U17076 ( .A1(n17757), .A2(n15238), .ZN(n15204) );
  NAND2_X1 U17077 ( .A1(n14384), .A2(n14419), .ZN(n15218) );
  NOR2_X1 U17078 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15193) );
  OR2_X1 U17079 ( .A1(n15192), .A2(n15193), .ZN(n15215) );
  OAI21_X1 U17080 ( .B1(n15218), .B2(n15215), .A(n15214), .ZN(n15196) );
  INV_X1 U17081 ( .A(n14243), .ZN(n15194) );
  NAND2_X1 U17082 ( .A1(n15235), .A2(n15194), .ZN(n15195) );
  AND2_X1 U17083 ( .A1(n15196), .A2(n15195), .ZN(n15202) );
  OR2_X1 U17084 ( .A1(n15254), .A2(n15263), .ZN(n15223) );
  INV_X1 U17085 ( .A(n15215), .ZN(n15199) );
  NAND2_X1 U17086 ( .A1(n15235), .A2(n14243), .ZN(n15197) );
  NAND2_X1 U17087 ( .A1(n15197), .A2(n15214), .ZN(n15198) );
  AOI21_X1 U17088 ( .B1(n15223), .B2(n15199), .A(n15198), .ZN(n15201) );
  MUX2_X1 U17089 ( .A(n15202), .B(n15201), .S(n15200), .Z(n15203) );
  AND2_X1 U17090 ( .A1(n15204), .A2(n15203), .ZN(n17658) );
  NAND2_X1 U17091 ( .A1(n15205), .A2(n15268), .ZN(n15212) );
  INV_X1 U17092 ( .A(n15270), .ZN(n15206) );
  NAND2_X1 U17093 ( .A1(n15206), .A2(n15269), .ZN(n15207) );
  AND4_X1 U17094 ( .A1(n15210), .A2(n15209), .A3(n15208), .A4(n15207), .ZN(
        n15211) );
  MUX2_X1 U17095 ( .A(n17658), .B(n15200), .S(n17645), .Z(n15251) );
  INV_X1 U17096 ( .A(n15238), .ZN(n15213) );
  NAND2_X1 U17097 ( .A1(n14808), .A2(n15213), .ZN(n15225) );
  NOR2_X1 U17098 ( .A1(n15215), .A2(n13321), .ZN(n15217) );
  INV_X1 U17099 ( .A(n15217), .ZN(n15222) );
  NOR2_X1 U17100 ( .A1(n15192), .A2(n14243), .ZN(n15216) );
  NAND2_X1 U17101 ( .A1(n15235), .A2(n15216), .ZN(n15220) );
  NAND2_X1 U17102 ( .A1(n15218), .A2(n15217), .ZN(n15219) );
  NAND2_X1 U17103 ( .A1(n15220), .A2(n15219), .ZN(n15221) );
  AOI21_X1 U17104 ( .B1(n15223), .B2(n15222), .A(n15221), .ZN(n15224) );
  NAND2_X1 U17105 ( .A1(n15225), .A2(n15224), .ZN(n15244) );
  OR2_X1 U17106 ( .A1(n15244), .A2(n17645), .ZN(n15228) );
  NAND2_X1 U17107 ( .A1(n17645), .A2(n15226), .ZN(n15227) );
  NAND2_X1 U17108 ( .A1(n15228), .A2(n15227), .ZN(n15249) );
  AND2_X1 U17109 ( .A1(n14387), .A2(n15229), .ZN(n15232) );
  INV_X1 U17110 ( .A(n15235), .ZN(n15230) );
  MUX2_X1 U17111 ( .A(n15232), .B(n15230), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15231) );
  OAI21_X1 U17112 ( .B1(n19183), .B2(n15238), .A(n15231), .ZN(n17643) );
  NOR2_X1 U17113 ( .A1(n17643), .A2(n19891), .ZN(n15240) );
  NAND2_X1 U17114 ( .A1(n15240), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15242) );
  INV_X1 U17115 ( .A(n15232), .ZN(n15233) );
  OAI21_X1 U17116 ( .B1(n13327), .B2(n13328), .A(n15233), .ZN(n15237) );
  NAND2_X1 U17117 ( .A1(n15235), .A2(n15234), .ZN(n15236) );
  OAI211_X1 U17118 ( .C1(n15239), .C2(n15238), .A(n15237), .B(n15236), .ZN(
        n17650) );
  INV_X1 U17119 ( .A(n15240), .ZN(n15241) );
  AOI22_X1 U17120 ( .A1(n15242), .A2(n17650), .B1(n19889), .B2(n15241), .ZN(
        n15243) );
  OAI22_X1 U17121 ( .A1(n15249), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n15243), .B2(n17645), .ZN(n15246) );
  INV_X1 U17122 ( .A(n15244), .ZN(n17654) );
  NAND2_X1 U17123 ( .A1(n17654), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15245) );
  NAND2_X1 U17124 ( .A1(n15246), .A2(n15245), .ZN(n15250) );
  OR2_X1 U17125 ( .A1(n15250), .A2(n15251), .ZN(n15247) );
  AND2_X1 U17126 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15247), .ZN(
        n15248) );
  OAI22_X1 U17127 ( .A1(n15251), .A2(n15249), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n15248), .ZN(n15253) );
  NAND2_X1 U17128 ( .A1(n15251), .A2(n15250), .ZN(n15252) );
  NAND2_X1 U17129 ( .A1(n15253), .A2(n15252), .ZN(n15278) );
  INV_X1 U17130 ( .A(n15254), .ZN(n15266) );
  INV_X1 U17131 ( .A(n15255), .ZN(n15261) );
  AOI22_X1 U17132 ( .A1(n15259), .A2(n15258), .B1(n15257), .B2(n15256), .ZN(
        n15260) );
  OAI21_X1 U17133 ( .B1(n19203), .B2(n15261), .A(n15260), .ZN(n15262) );
  INV_X1 U17134 ( .A(n15262), .ZN(n15265) );
  NAND2_X1 U17135 ( .A1(n17641), .A2(n15263), .ZN(n15264) );
  OAI211_X1 U17136 ( .C1(n15266), .C2(n17641), .A(n15265), .B(n15264), .ZN(
        n19221) );
  INV_X1 U17137 ( .A(n19221), .ZN(n15275) );
  INV_X1 U17138 ( .A(n15267), .ZN(n15274) );
  NOR3_X1 U17139 ( .A1(n15270), .A2(n15269), .A3(n15268), .ZN(n19220) );
  OAI21_X1 U17140 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19220), .ZN(n15273) );
  NAND2_X1 U17141 ( .A1(n13109), .A2(n19174), .ZN(n15271) );
  OR2_X1 U17142 ( .A1(n13315), .A2(n15271), .ZN(n15272) );
  NAND4_X1 U17143 ( .A1(n15275), .A2(n15274), .A3(n15273), .A4(n15272), .ZN(
        n15276) );
  AOI21_X1 U17144 ( .B1(n17645), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n15276), .ZN(n15277) );
  AND2_X1 U17145 ( .A1(n13265), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15279) );
  NAND2_X1 U17146 ( .A1(n19218), .A2(n15279), .ZN(n15283) );
  AND2_X1 U17147 ( .A1(n15281), .A2(n15280), .ZN(n15282) );
  AOI21_X1 U17148 ( .B1(n15283), .B2(n17692), .A(n15282), .ZN(n19210) );
  OAI21_X1 U17149 ( .B1(n19210), .B2(n17752), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n15284) );
  NOR2_X1 U17150 ( .A1(n17752), .A2(n17693), .ZN(n17689) );
  INV_X1 U17151 ( .A(n17689), .ZN(n19205) );
  NAND2_X1 U17152 ( .A1(n15284), .A2(n19205), .ZN(P2_U3593) );
  INV_X1 U17153 ( .A(n15112), .ZN(n15287) );
  NAND2_X1 U17154 ( .A1(n16178), .A2(n15287), .ZN(n15455) );
  NOR2_X2 U17155 ( .A1(n22442), .A2(n15455), .ZN(n22750) );
  OAI21_X1 U17156 ( .B1(n22750), .B2(n15633), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15289) );
  AND2_X1 U17157 ( .A1(n15074), .A2(n15288), .ZN(n22460) );
  NAND2_X1 U17158 ( .A1(n22460), .A2(n22430), .ZN(n15293) );
  AOI21_X1 U17159 ( .B1(n15289), .B2(n15293), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15290) );
  NOR3_X1 U17160 ( .A1(n12665), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15396) );
  INV_X1 U17161 ( .A(n15396), .ZN(n15398) );
  NOR2_X1 U17162 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15398), .ZN(
        n22698) );
  INV_X1 U17163 ( .A(n22700), .ZN(n15600) );
  INV_X1 U17164 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15296) );
  OR2_X1 U17165 ( .A1(n15314), .A2(n15291), .ZN(n22417) );
  OAI22_X1 U17166 ( .A1(n15293), .A2(n22497), .B1(n15292), .B2(n22417), .ZN(
        n22699) );
  AOI22_X1 U17167 ( .A1(n15633), .A2(n15142), .B1(n22799), .B2(n22699), .ZN(
        n15295) );
  AOI22_X1 U17168 ( .A1(n22750), .A2(n11345), .B1(n22698), .B2(n22797), .ZN(
        n15294) );
  OAI211_X1 U17169 ( .C1(n15600), .C2(n15296), .A(n15295), .B(n15294), .ZN(
        P1_U3072) );
  AND2_X1 U17170 ( .A1(n15298), .A2(n15297), .ZN(n15300) );
  OR2_X1 U17171 ( .A1(n15300), .A2(n15299), .ZN(n22076) );
  OAI22_X1 U17172 ( .A1(n16592), .A2(BUF1_REG_6__SCAN_IN), .B1(DATAI_6_), .B2(
        n16588), .ZN(n22346) );
  OAI222_X1 U17173 ( .A1(n22076), .A2(n16667), .B1(n15954), .B2(n22346), .C1(
        n22351), .C2(n16659), .ZN(P1_U2898) );
  OR2_X1 U17174 ( .A1(n15301), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15302) );
  NAND2_X1 U17175 ( .A1(n15303), .A2(n15302), .ZN(n22008) );
  NAND3_X1 U17176 ( .A1(n16420), .A2(n22809), .A3(n16422), .ZN(n15308) );
  NAND4_X1 U17177 ( .A1(n15304), .A2(n15383), .A3(n14540), .A4(n15592), .ZN(
        n15305) );
  OR2_X1 U17178 ( .A1(n15306), .A2(n15305), .ZN(n15307) );
  NAND2_X2 U17179 ( .A1(n15308), .A2(n15307), .ZN(n20493) );
  NAND2_X2 U17180 ( .A1(n20493), .A2(n16596), .ZN(n20480) );
  OAI222_X1 U17181 ( .A1(n22008), .A2(n20480), .B1(n20483), .B2(n15415), .C1(
        n20493), .C2(n13849), .ZN(P1_U2872) );
  NOR3_X1 U17182 ( .A1(n12668), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15497) );
  INV_X1 U17183 ( .A(n15497), .ZN(n15500) );
  NOR2_X1 U17184 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15500), .ZN(
        n22711) );
  INV_X1 U17185 ( .A(n15499), .ZN(n15310) );
  INV_X1 U17186 ( .A(n15461), .ZN(n15435) );
  INV_X1 U17187 ( .A(n22772), .ZN(n15624) );
  OR2_X1 U17188 ( .A1(n15471), .A2(n15455), .ZN(n22710) );
  OAI21_X1 U17189 ( .B1(n15624), .B2(n22713), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15311) );
  AND2_X1 U17190 ( .A1(n22024), .A2(n22041), .ZN(n22479) );
  AOI21_X1 U17191 ( .B1(n22479), .B2(n22430), .A(n22711), .ZN(n15313) );
  NAND2_X1 U17192 ( .A1(n15311), .A2(n15313), .ZN(n15312) );
  NOR2_X1 U17193 ( .A1(n22503), .A2(n22411), .ZN(n22490) );
  OAI211_X1 U17194 ( .C1(n22464), .C2(n22711), .A(n15312), .B(n22490), .ZN(
        n22714) );
  INV_X1 U17195 ( .A(n15313), .ZN(n15315) );
  NAND2_X1 U17196 ( .A1(n15314), .A2(n22432), .ZN(n22507) );
  INV_X1 U17197 ( .A(n22507), .ZN(n22502) );
  AOI22_X1 U17198 ( .A1(n15315), .A2(n22440), .B1(n22502), .B2(n22481), .ZN(
        n22473) );
  OAI22_X1 U17199 ( .A1(n22787), .A2(n22473), .B1(n11344), .B2(n22710), .ZN(
        n15319) );
  INV_X1 U17200 ( .A(n15142), .ZN(n15317) );
  INV_X1 U17201 ( .A(n22797), .ZN(n15316) );
  INV_X1 U17202 ( .A(n22711), .ZN(n15668) );
  OAI22_X1 U17203 ( .A1(n22772), .A2(n15317), .B1(n15316), .B2(n15668), .ZN(
        n15318) );
  AOI211_X1 U17204 ( .C1(n22714), .C2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n15319), .B(n15318), .ZN(n15320) );
  INV_X1 U17205 ( .A(n15320), .ZN(P1_U3104) );
  OR2_X1 U17206 ( .A1(n11202), .A2(n15321), .ZN(n15322) );
  NAND2_X1 U17207 ( .A1(n15322), .A2(n15327), .ZN(n17806) );
  NAND2_X1 U17208 ( .A1(n15323), .A2(n17795), .ZN(n15324) );
  OAI21_X1 U17209 ( .B1(n15325), .B2(n17805), .A(n15324), .ZN(n20072) );
  XNOR2_X1 U17210 ( .A(n19768), .B(n17806), .ZN(n20073) );
  NOR2_X1 U17211 ( .A1(n20072), .A2(n20073), .ZN(n20071) );
  AOI21_X1 U17212 ( .B1(n17806), .B2(n19768), .A(n20071), .ZN(n15328) );
  XNOR2_X1 U17213 ( .A(n15327), .B(n15326), .ZN(n15651) );
  INV_X1 U17214 ( .A(n15651), .ZN(n16023) );
  NOR2_X1 U17215 ( .A1(n15328), .A2(n16023), .ZN(n19975) );
  OAI21_X1 U17216 ( .B1(n15330), .B2(n15329), .A(n16011), .ZN(n19974) );
  XNOR2_X1 U17217 ( .A(n19975), .B(n19974), .ZN(n15333) );
  AOI22_X1 U17218 ( .A1(n20169), .A2(n16023), .B1(n20221), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n15332) );
  INV_X1 U17219 ( .A(n20028), .ZN(n20020) );
  NAND2_X1 U17220 ( .A1(n19972), .A2(n20020), .ZN(n15331) );
  OAI211_X1 U17221 ( .C1(n15333), .C2(n20228), .A(n15332), .B(n15331), .ZN(
        P2_U2915) );
  AND2_X1 U17222 ( .A1(n15335), .A2(n15334), .ZN(n15336) );
  NOR2_X1 U17223 ( .A1(n15446), .A2(n15336), .ZN(n17520) );
  INV_X1 U17224 ( .A(n17520), .ZN(n15930) );
  NOR2_X1 U17225 ( .A1(n15338), .A2(n15337), .ZN(n15349) );
  NAND2_X1 U17226 ( .A1(n15339), .A2(n15348), .ZN(n15341) );
  NOR2_X1 U17227 ( .A1(n15341), .A2(n15340), .ZN(n15344) );
  INV_X1 U17228 ( .A(n15419), .ZN(n15347) );
  OAI211_X1 U17229 ( .C1(n15349), .C2(n15348), .A(n15347), .B(n17039), .ZN(
        n15351) );
  NAND2_X1 U17230 ( .A1(n15444), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15350) );
  OAI211_X1 U17231 ( .C1(n15930), .C2(n15444), .A(n15351), .B(n15350), .ZN(
        P2_U2875) );
  NAND2_X1 U17232 ( .A1(n15353), .A2(n15352), .ZN(n15354) );
  NAND2_X1 U17233 ( .A1(n15359), .A2(n15354), .ZN(n22036) );
  OAI222_X1 U17234 ( .A1(n22036), .A2(n20480), .B1(n20493), .B2(n22038), .C1(
        n20483), .C2(n15355), .ZN(P1_U2869) );
  NAND2_X1 U17235 ( .A1(n15478), .A2(n15356), .ZN(n15357) );
  NAND2_X1 U17236 ( .A1(n15523), .A2(n15357), .ZN(n22078) );
  OAI222_X1 U17237 ( .A1(n22078), .A2(n20480), .B1(n22079), .B2(n20493), .C1(
        n22076), .C2(n20483), .ZN(P1_U2866) );
  AND2_X1 U17238 ( .A1(n15359), .A2(n15358), .ZN(n15360) );
  OR2_X1 U17239 ( .A1(n15360), .A2(n15480), .ZN(n22052) );
  OAI222_X1 U17240 ( .A1(n22052), .A2(n20480), .B1(n22064), .B2(n20493), .C1(
        n22059), .C2(n20483), .ZN(P1_U2868) );
  INV_X1 U17241 ( .A(n22052), .ZN(n15369) );
  NOR2_X1 U17242 ( .A1(n15361), .A2(n16893), .ZN(n15362) );
  INV_X1 U17243 ( .A(n16786), .ZN(n15519) );
  AOI22_X1 U17244 ( .A1(n21918), .A2(n15363), .B1(n15362), .B2(n15519), .ZN(
        n21873) );
  XNOR2_X1 U17245 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15366) );
  OAI22_X1 U17246 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21922), .B1(
        n15363), .B2(n16788), .ZN(n15364) );
  NOR2_X1 U17247 ( .A1(n15365), .A2(n15364), .ZN(n21871) );
  OAI22_X1 U17248 ( .A1(n21873), .A2(n15366), .B1(n21871), .B2(n12877), .ZN(
        n15367) );
  AOI211_X1 U17249 ( .C1(n21993), .C2(n15369), .A(n15368), .B(n15367), .ZN(
        n15370) );
  OAI21_X1 U17250 ( .B1(n22010), .B2(n15371), .A(n15370), .ZN(P1_U3027) );
  NOR2_X1 U17251 ( .A1(n12668), .A2(n22463), .ZN(n15376) );
  INV_X1 U17252 ( .A(n15436), .ZN(n15372) );
  NOR3_X1 U17253 ( .A1(n15372), .A2(n22497), .A3(n22441), .ZN(n15373) );
  OAI21_X1 U17254 ( .B1(n15376), .B2(n15373), .A(n22447), .ZN(n22801) );
  INV_X1 U17255 ( .A(n22801), .ZN(n15596) );
  INV_X1 U17256 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15386) );
  INV_X1 U17257 ( .A(n22328), .ZN(n16643) );
  NAND2_X1 U17258 ( .A1(n22626), .A2(n16643), .ZN(n22620) );
  INV_X1 U17259 ( .A(n12030), .ZN(n15374) );
  AND2_X1 U17260 ( .A1(n15374), .A2(n15412), .ZN(n22443) );
  NOR2_X1 U17261 ( .A1(n15375), .A2(n12668), .ZN(n22796) );
  AOI21_X1 U17262 ( .B1(n15430), .B2(n22443), .A(n22796), .ZN(n15378) );
  INV_X1 U17263 ( .A(n15376), .ZN(n15377) );
  OAI22_X1 U17264 ( .A1(n15378), .A2(n22497), .B1(n15377), .B2(n21855), .ZN(
        n22798) );
  INV_X1 U17265 ( .A(n15455), .ZN(n15379) );
  INV_X1 U17266 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20602) );
  OAI22_X1 U17267 ( .A1(n16641), .A2(n22632), .B1(n20602), .B2(n22630), .ZN(
        n22617) );
  AOI22_X1 U17268 ( .A1(n22622), .A2(n22798), .B1(n22800), .B2(n11340), .ZN(
        n15385) );
  INV_X1 U17269 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20617) );
  INV_X1 U17270 ( .A(DATAI_27_), .ZN(n15380) );
  OR2_X1 U17271 ( .A1(n22632), .A2(n15380), .ZN(n15381) );
  NOR2_X2 U17272 ( .A1(n22629), .A2(n15383), .ZN(n22621) );
  AOI22_X1 U17273 ( .A1(n15639), .A2(n15382), .B1(n22796), .B2(n22621), .ZN(
        n15384) );
  OAI211_X1 U17274 ( .C1(n15596), .C2(n15386), .A(n15385), .B(n15384), .ZN(
        P1_U3156) );
  INV_X1 U17275 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15394) );
  NAND2_X1 U17276 ( .A1(n22626), .A2(n22315), .ZN(n22550) );
  INV_X1 U17277 ( .A(DATAI_17_), .ZN(n15387) );
  INV_X1 U17278 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20599) );
  OAI22_X1 U17279 ( .A1(n15387), .A2(n22632), .B1(n20599), .B2(n22630), .ZN(
        n22547) );
  AOI22_X1 U17280 ( .A1(n22552), .A2(n22798), .B1(n22800), .B2(n11342), .ZN(
        n15393) );
  INV_X1 U17281 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20613) );
  INV_X1 U17282 ( .A(DATAI_25_), .ZN(n15388) );
  OR2_X1 U17283 ( .A1(n22632), .A2(n15388), .ZN(n15389) );
  NOR2_X2 U17284 ( .A1(n22629), .A2(n15391), .ZN(n22551) );
  AOI22_X1 U17285 ( .A1(n15639), .A2(n15390), .B1(n22796), .B2(n22551), .ZN(
        n15392) );
  OAI211_X1 U17286 ( .C1(n15596), .C2(n15394), .A(n15393), .B(n15392), .ZN(
        P1_U3154) );
  NOR3_X1 U17287 ( .A1(n15471), .A2(n22497), .A3(n15495), .ZN(n15395) );
  OAI21_X1 U17288 ( .B1(n15396), .B2(n15395), .A(n22447), .ZN(n22757) );
  INV_X1 U17289 ( .A(n22757), .ZN(n15637) );
  INV_X1 U17290 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15402) );
  NOR2_X2 U17291 ( .A1(n15498), .A2(n15471), .ZN(n22762) );
  INV_X1 U17292 ( .A(n15397), .ZN(n15494) );
  NOR2_X1 U17293 ( .A1(n22485), .A2(n15398), .ZN(n22755) );
  AOI21_X1 U17294 ( .B1(n22460), .B2(n15494), .A(n22755), .ZN(n15399) );
  OAI22_X1 U17295 ( .A1(n15399), .A2(n22497), .B1(n15398), .B2(n21855), .ZN(
        n22756) );
  AOI22_X1 U17296 ( .A1(n22762), .A2(n11340), .B1(n22622), .B2(n22756), .ZN(
        n15401) );
  AOI22_X1 U17297 ( .A1(n15633), .A2(n15382), .B1(n22755), .B2(n22621), .ZN(
        n15400) );
  OAI211_X1 U17298 ( .C1(n15637), .C2(n15402), .A(n15401), .B(n15400), .ZN(
        P1_U3076) );
  INV_X1 U17299 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15405) );
  AOI22_X1 U17300 ( .A1(n22762), .A2(n11342), .B1(n22552), .B2(n22756), .ZN(
        n15404) );
  AOI22_X1 U17301 ( .A1(n15633), .A2(n15390), .B1(n22755), .B2(n22551), .ZN(
        n15403) );
  OAI211_X1 U17302 ( .C1(n15637), .C2(n15405), .A(n15404), .B(n15403), .ZN(
        P1_U3074) );
  OAI21_X1 U17303 ( .B1(n15410), .B2(n15406), .A(n22209), .ZN(n22069) );
  INV_X1 U17304 ( .A(n22069), .ZN(n22058) );
  INV_X1 U17305 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15407) );
  AOI21_X1 U17306 ( .B1(n22203), .B2(n22152), .A(n15407), .ZN(n15409) );
  NOR2_X1 U17307 ( .A1(n22208), .A2(n22008), .ZN(n15408) );
  AOI211_X1 U17308 ( .C1(P1_EBX_REG_0__SCAN_IN), .C2(n22166), .A(n15409), .B(
        n15408), .ZN(n15414) );
  NAND2_X1 U17309 ( .A1(n21860), .A2(n15411), .ZN(n22050) );
  INV_X1 U17310 ( .A(n22050), .ZN(n22042) );
  AOI22_X1 U17311 ( .A1(n22200), .A2(P1_REIP_REG_0__SCAN_IN), .B1(n22042), 
        .B2(n15412), .ZN(n15413) );
  OAI211_X1 U17312 ( .C1(n15415), .C2(n22058), .A(n15414), .B(n15413), .ZN(
        P1_U2840) );
  NAND2_X1 U17313 ( .A1(n15416), .A2(n15417), .ZN(n15418) );
  NAND2_X1 U17314 ( .A1(n15702), .A2(n15418), .ZN(n17493) );
  INV_X1 U17315 ( .A(n15420), .ZN(n15421) );
  OAI211_X1 U17316 ( .C1(n11835), .C2(n15421), .A(n17039), .B(n15704), .ZN(
        n15423) );
  NAND2_X1 U17317 ( .A1(n15444), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15422) );
  OAI211_X1 U17318 ( .C1(n17493), .C2(n15444), .A(n15423), .B(n15422), .ZN(
        P2_U2873) );
  INV_X1 U17319 ( .A(n15424), .ZN(n15426) );
  INV_X1 U17320 ( .A(n15299), .ZN(n15425) );
  AOI21_X1 U17321 ( .B1(n15426), .B2(n15425), .A(n11274), .ZN(n20500) );
  INV_X1 U17322 ( .A(n20500), .ZN(n22092) );
  OAI222_X1 U17323 ( .A1(n22092), .A2(n16667), .B1(n15954), .B2(n22352), .C1(
        n16659), .C2(n12149), .ZN(P1_U2897) );
  NOR2_X1 U17324 ( .A1(n11274), .A2(n15427), .ZN(n15428) );
  OR2_X1 U17325 ( .A1(n11275), .A2(n15428), .ZN(n15696) );
  OAI22_X1 U17326 ( .A1(n16592), .A2(BUF1_REG_8__SCAN_IN), .B1(DATAI_8_), .B2(
        n16588), .ZN(n22357) );
  INV_X1 U17327 ( .A(n22357), .ZN(n16621) );
  AOI22_X1 U17328 ( .A1(n15948), .A2(n16621), .B1(n16653), .B2(
        P1_EAX_REG_8__SCAN_IN), .ZN(n15429) );
  OAI21_X1 U17329 ( .B1(n15696), .B2(n16667), .A(n15429), .ZN(P1_U2896) );
  NOR3_X1 U17330 ( .A1(n12665), .A2(n12668), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15433) );
  INV_X1 U17331 ( .A(n15433), .ZN(n22505) );
  NOR2_X1 U17332 ( .A1(n22485), .A2(n22505), .ZN(n22789) );
  AOI21_X1 U17333 ( .B1(n15430), .B2(n15494), .A(n22789), .ZN(n15434) );
  NAND3_X1 U17334 ( .A1(n15431), .A2(n22440), .A3(n15434), .ZN(n15432) );
  OAI211_X1 U17335 ( .C1(n22440), .C2(n15433), .A(n22447), .B(n15432), .ZN(
        n22792) );
  INV_X1 U17336 ( .A(n22792), .ZN(n15604) );
  INV_X1 U17337 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15439) );
  OAI22_X1 U17338 ( .A1(n15434), .A2(n22497), .B1(n22505), .B2(n21855), .ZN(
        n22790) );
  AOI22_X1 U17339 ( .A1(n22552), .A2(n22790), .B1(n22791), .B2(n11342), .ZN(
        n15438) );
  NAND2_X1 U17340 ( .A1(n15436), .A2(n15435), .ZN(n22795) );
  AOI22_X1 U17341 ( .A1(n22781), .A2(n15390), .B1(n22789), .B2(n22551), .ZN(
        n15437) );
  OAI211_X1 U17342 ( .C1(n15604), .C2(n15439), .A(n15438), .B(n15437), .ZN(
        P1_U3138) );
  INV_X1 U17343 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15442) );
  AOI22_X1 U17344 ( .A1(n22622), .A2(n22790), .B1(n22791), .B2(n11340), .ZN(
        n15441) );
  AOI22_X1 U17345 ( .A1(n22781), .A2(n15382), .B1(n22789), .B2(n22621), .ZN(
        n15440) );
  OAI211_X1 U17346 ( .C1(n15604), .C2(n15442), .A(n15441), .B(n15440), .ZN(
        P1_U3140) );
  XNOR2_X1 U17347 ( .A(n15419), .B(n15443), .ZN(n15450) );
  OR2_X1 U17348 ( .A1(n15446), .A2(n15445), .ZN(n15447) );
  NAND2_X1 U17349 ( .A1(n15416), .A2(n15447), .ZN(n19027) );
  NOR2_X1 U17350 ( .A1(n19027), .A2(n15444), .ZN(n15448) );
  AOI21_X1 U17351 ( .B1(P2_EBX_REG_13__SCAN_IN), .B2(n15444), .A(n15448), .ZN(
        n15449) );
  OAI21_X1 U17352 ( .B1(n15450), .B2(n17034), .A(n15449), .ZN(P2_U2874) );
  NOR3_X1 U17353 ( .A1(n12668), .A2(n15451), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22484) );
  INV_X1 U17354 ( .A(n22484), .ZN(n15453) );
  NOR2_X1 U17355 ( .A1(n22485), .A2(n15453), .ZN(n22719) );
  AOI21_X1 U17356 ( .B1(n22479), .B2(n22443), .A(n22719), .ZN(n15454) );
  OAI211_X1 U17357 ( .C1(n15499), .C2(n22441), .A(n22440), .B(n15454), .ZN(
        n15452) );
  OAI211_X1 U17358 ( .C1(n22440), .C2(n22484), .A(n22447), .B(n15452), .ZN(
        n22721) );
  INV_X1 U17359 ( .A(n22721), .ZN(n15632) );
  INV_X1 U17360 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15458) );
  NOR2_X2 U17361 ( .A1(n15499), .A2(n15470), .ZN(n22775) );
  OAI22_X1 U17362 ( .A1(n15454), .A2(n22497), .B1(n15453), .B2(n21855), .ZN(
        n22720) );
  AOI22_X1 U17363 ( .A1(n22775), .A2(n11345), .B1(n22799), .B2(n22720), .ZN(
        n15457) );
  AOI22_X1 U17364 ( .A1(n22783), .A2(n15142), .B1(n22719), .B2(n22797), .ZN(
        n15456) );
  OAI211_X1 U17365 ( .C1(n15632), .C2(n15458), .A(n15457), .B(n15456), .ZN(
        P1_U3128) );
  NOR3_X1 U17366 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15460) );
  OR2_X1 U17367 ( .A1(n15074), .A2(n22041), .ZN(n22431) );
  INV_X1 U17368 ( .A(n22431), .ZN(n22444) );
  INV_X1 U17369 ( .A(n15460), .ZN(n22415) );
  NOR2_X1 U17370 ( .A1(n22485), .A2(n22415), .ZN(n22688) );
  AOI21_X1 U17371 ( .B1(n22444), .B2(n15494), .A(n22688), .ZN(n15462) );
  OAI211_X1 U17372 ( .C1(n22442), .C2(n15495), .A(n22440), .B(n15462), .ZN(
        n15459) );
  OAI211_X1 U17373 ( .C1(n22440), .C2(n15460), .A(n22447), .B(n15459), .ZN(
        n22690) );
  INV_X1 U17374 ( .A(n22690), .ZN(n15619) );
  INV_X1 U17375 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15466) );
  NOR2_X2 U17376 ( .A1(n22442), .A2(n15461), .ZN(n22737) );
  OAI22_X1 U17377 ( .A1(n15462), .A2(n22497), .B1(n22415), .B2(n21855), .ZN(
        n22689) );
  AOI22_X1 U17378 ( .A1(n22737), .A2(n11345), .B1(n22799), .B2(n22689), .ZN(
        n15465) );
  AOI22_X1 U17379 ( .A1(n22743), .A2(n15142), .B1(n22688), .B2(n22797), .ZN(
        n15464) );
  OAI211_X1 U17380 ( .C1(n15619), .C2(n15466), .A(n15465), .B(n15464), .ZN(
        P1_U3048) );
  NOR2_X1 U17381 ( .A1(n22463), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15472) );
  INV_X1 U17382 ( .A(n15467), .ZN(n22705) );
  AOI21_X1 U17383 ( .B1(n22460), .B2(n22443), .A(n22705), .ZN(n15474) );
  NAND3_X1 U17384 ( .A1(n15468), .A2(n22440), .A3(n15474), .ZN(n15469) );
  OAI211_X1 U17385 ( .C1(n22440), .C2(n15472), .A(n22447), .B(n15469), .ZN(
        n22707) );
  INV_X1 U17386 ( .A(n22707), .ZN(n15623) );
  INV_X1 U17387 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15477) );
  NOR2_X2 U17388 ( .A1(n15471), .A2(n15470), .ZN(n22761) );
  INV_X1 U17389 ( .A(n15472), .ZN(n15473) );
  OAI22_X1 U17390 ( .A1(n15474), .A2(n22497), .B1(n15473), .B2(n21855), .ZN(
        n22706) );
  AOI22_X1 U17391 ( .A1(n11345), .A2(n22761), .B1(n22799), .B2(n22706), .ZN(
        n15476) );
  AOI22_X1 U17392 ( .A1(n22713), .A2(n15142), .B1(n22705), .B2(n22797), .ZN(
        n15475) );
  OAI211_X1 U17393 ( .C1(n15623), .C2(n15477), .A(n15476), .B(n15475), .ZN(
        P1_U3096) );
  INV_X1 U17394 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n15481) );
  OAI21_X1 U17395 ( .B1(n15480), .B2(n15479), .A(n15478), .ZN(n22067) );
  OAI222_X1 U17396 ( .A1(n15482), .A2(n20483), .B1(n20493), .B2(n15481), .C1(
        n20480), .C2(n22067), .ZN(P1_U2867) );
  INV_X1 U17397 ( .A(n15483), .ZN(n15577) );
  OAI21_X1 U17398 ( .B1(n22189), .B2(n15485), .A(n15484), .ZN(n15486) );
  NAND2_X1 U17399 ( .A1(n15577), .A2(n15486), .ZN(n15493) );
  AOI21_X1 U17400 ( .B1(n15487), .B2(n15525), .A(n15580), .ZN(n20487) );
  OAI22_X1 U17401 ( .A1(n15488), .A2(n22152), .B1(n20492), .B2(n22201), .ZN(
        n15489) );
  NOR2_X1 U17402 ( .A1(n22170), .A2(n15489), .ZN(n15490) );
  OAI21_X1 U17403 ( .B1(n22203), .B2(n15698), .A(n15490), .ZN(n15491) );
  AOI21_X1 U17404 ( .B1(n20487), .B2(n22165), .A(n15491), .ZN(n15492) );
  OAI211_X1 U17405 ( .C1(n15696), .C2(n22209), .A(n15493), .B(n15492), .ZN(
        P1_U2832) );
  NOR2_X1 U17406 ( .A1(n22485), .A2(n15500), .ZN(n22767) );
  AOI21_X1 U17407 ( .B1(n22479), .B2(n15494), .A(n22767), .ZN(n15501) );
  OAI211_X1 U17408 ( .C1(n15499), .C2(n15495), .A(n22440), .B(n15501), .ZN(
        n15496) );
  OAI211_X1 U17409 ( .C1(n22440), .C2(n15497), .A(n22447), .B(n15496), .ZN(
        n22769) );
  INV_X1 U17410 ( .A(n22769), .ZN(n15628) );
  INV_X1 U17411 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15507) );
  NOR2_X2 U17412 ( .A1(n15499), .A2(n15498), .ZN(n22774) );
  OAI22_X1 U17413 ( .A1(n15501), .A2(n22497), .B1(n15500), .B2(n21855), .ZN(
        n22768) );
  AOI22_X1 U17414 ( .A1(n22774), .A2(n11342), .B1(n22552), .B2(n22768), .ZN(
        n15506) );
  INV_X1 U17415 ( .A(n15390), .ZN(n15503) );
  INV_X1 U17416 ( .A(n22551), .ZN(n15502) );
  INV_X1 U17417 ( .A(n22767), .ZN(n15539) );
  OAI22_X1 U17418 ( .A1(n22772), .A2(n15503), .B1(n15502), .B2(n15539), .ZN(
        n15504) );
  INV_X1 U17419 ( .A(n15504), .ZN(n15505) );
  OAI211_X1 U17420 ( .C1(n15628), .C2(n15507), .A(n15506), .B(n15505), .ZN(
        P1_U3106) );
  INV_X1 U17421 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15513) );
  AOI22_X1 U17422 ( .A1(n22774), .A2(n11340), .B1(n22622), .B2(n22768), .ZN(
        n15512) );
  INV_X1 U17423 ( .A(n15382), .ZN(n15509) );
  INV_X1 U17424 ( .A(n22621), .ZN(n15508) );
  OAI22_X1 U17425 ( .A1(n22772), .A2(n15509), .B1(n15508), .B2(n15539), .ZN(
        n15510) );
  INV_X1 U17426 ( .A(n15510), .ZN(n15511) );
  OAI211_X1 U17427 ( .C1(n15628), .C2(n15513), .A(n15512), .B(n15511), .ZN(
        P1_U3108) );
  XOR2_X1 U17428 ( .A(n15514), .B(n15515), .Z(n20495) );
  INV_X1 U17429 ( .A(n20495), .ZN(n15522) );
  NAND2_X1 U17430 ( .A1(n21918), .A2(n15611), .ZN(n15516) );
  OAI211_X1 U17431 ( .C1(n21922), .C2(n15520), .A(n21920), .B(n15516), .ZN(
        n15608) );
  NOR2_X1 U17432 ( .A1(n21975), .A2(n22071), .ZN(n20496) );
  OAI22_X1 U17433 ( .A1(n15517), .A2(n15516), .B1(n22009), .B2(n22067), .ZN(
        n15518) );
  AOI211_X1 U17434 ( .C1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n15608), .A(
        n20496), .B(n15518), .ZN(n15521) );
  NAND3_X1 U17435 ( .A1(n12888), .A2(n15520), .A3(n15519), .ZN(n15607) );
  OAI211_X1 U17436 ( .C1(n15522), .C2(n22010), .A(n15521), .B(n15607), .ZN(
        P1_U3026) );
  NAND2_X1 U17437 ( .A1(n15523), .A2(n11850), .ZN(n15524) );
  NAND2_X1 U17438 ( .A1(n15525), .A2(n15524), .ZN(n22088) );
  INV_X1 U17439 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n22098) );
  OAI222_X1 U17440 ( .A1(n22088), .A2(n20480), .B1(n20493), .B2(n22098), .C1(
        n20483), .C2(n22092), .ZN(P1_U2865) );
  INV_X1 U17441 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15532) );
  INV_X1 U17442 ( .A(n22346), .ZN(n16631) );
  NAND2_X1 U17443 ( .A1(n22626), .A2(n16631), .ZN(n22728) );
  INV_X1 U17444 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20607) );
  OAI22_X1 U17445 ( .A1(n16629), .A2(n22632), .B1(n20607), .B2(n22630), .ZN(
        n22725) );
  AOI22_X1 U17446 ( .A1(n22732), .A2(n22798), .B1(n22800), .B2(n11338), .ZN(
        n15531) );
  INV_X1 U17447 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20623) );
  INV_X1 U17448 ( .A(DATAI_30_), .ZN(n15526) );
  OR2_X1 U17449 ( .A1(n22632), .A2(n15526), .ZN(n15527) );
  NOR2_X2 U17450 ( .A1(n22629), .A2(n15529), .ZN(n22730) );
  AOI22_X1 U17451 ( .A1(n15639), .A2(n15528), .B1(n22796), .B2(n22730), .ZN(
        n15530) );
  OAI211_X1 U17452 ( .C1(n15596), .C2(n15532), .A(n15531), .B(n15530), .ZN(
        P1_U3159) );
  INV_X1 U17453 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15535) );
  AOI22_X1 U17454 ( .A1(n22732), .A2(n22790), .B1(n22791), .B2(n11338), .ZN(
        n15534) );
  AOI22_X1 U17455 ( .A1(n22781), .A2(n15528), .B1(n22789), .B2(n22730), .ZN(
        n15533) );
  OAI211_X1 U17456 ( .C1(n15604), .C2(n15535), .A(n15534), .B(n15533), .ZN(
        P1_U3143) );
  INV_X1 U17457 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15538) );
  AOI22_X1 U17458 ( .A1(n22762), .A2(n11338), .B1(n22732), .B2(n22756), .ZN(
        n15537) );
  AOI22_X1 U17459 ( .A1(n15633), .A2(n15528), .B1(n22755), .B2(n22730), .ZN(
        n15536) );
  OAI211_X1 U17460 ( .C1(n15637), .C2(n15538), .A(n15537), .B(n15536), .ZN(
        P1_U3079) );
  INV_X1 U17461 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15545) );
  AOI22_X1 U17462 ( .A1(n22774), .A2(n11338), .B1(n22732), .B2(n22768), .ZN(
        n15544) );
  INV_X1 U17463 ( .A(n15528), .ZN(n15541) );
  INV_X1 U17464 ( .A(n22730), .ZN(n15540) );
  OAI22_X1 U17465 ( .A1(n22772), .A2(n15541), .B1(n15540), .B2(n15539), .ZN(
        n15542) );
  INV_X1 U17466 ( .A(n15542), .ZN(n15543) );
  OAI211_X1 U17467 ( .C1(n15628), .C2(n15545), .A(n15544), .B(n15543), .ZN(
        P1_U3111) );
  XNOR2_X1 U17468 ( .A(n15644), .B(n15546), .ZN(n15646) );
  XNOR2_X1 U17469 ( .A(n15646), .B(n15547), .ZN(n17759) );
  INV_X1 U17470 ( .A(n17759), .ZN(n15560) );
  INV_X1 U17471 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n17861) );
  OAI22_X1 U17472 ( .A1(n17806), .A2(n17622), .B1(n17861), .B2(n19068), .ZN(
        n15555) );
  INV_X1 U17473 ( .A(n17614), .ZN(n15650) );
  NOR2_X1 U17474 ( .A1(n15549), .A2(n15548), .ZN(n15550) );
  AOI211_X1 U17475 ( .C1(n15552), .C2(n15551), .A(n15550), .B(n19185), .ZN(
        n17584) );
  INV_X1 U17476 ( .A(n17584), .ZN(n15553) );
  MUX2_X1 U17477 ( .A(n15650), .B(n15553), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n15554) );
  AOI211_X1 U17478 ( .C1(n17633), .C2(n14864), .A(n15555), .B(n15554), .ZN(
        n15559) );
  NAND2_X1 U17479 ( .A1(n14286), .A2(n15557), .ZN(n17755) );
  NAND3_X1 U17480 ( .A1(n15556), .A2(n17755), .A3(n17628), .ZN(n15558) );
  OAI211_X1 U17481 ( .C1(n15560), .C2(n19182), .A(n15559), .B(n15558), .ZN(
        P2_U3043) );
  INV_X1 U17482 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n22311) );
  AOI22_X1 U17483 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20399), .B1(n20390), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n15561) );
  OAI21_X1 U17484 ( .B1(n22311), .B2(n15576), .A(n15561), .ZN(P1_U2920) );
  OAI21_X1 U17485 ( .B1(n11275), .B2(n15562), .A(n14063), .ZN(n15780) );
  OAI22_X1 U17486 ( .A1(n16592), .A2(BUF1_REG_9__SCAN_IN), .B1(DATAI_9_), .B2(
        n16588), .ZN(n22362) );
  INV_X1 U17487 ( .A(n22362), .ZN(n16613) );
  AOI22_X1 U17488 ( .A1(n15948), .A2(n16613), .B1(n16653), .B2(
        P1_EAX_REG_9__SCAN_IN), .ZN(n15563) );
  OAI21_X1 U17489 ( .B1(n15780), .B2(n16667), .A(n15563), .ZN(P1_U2895) );
  AOI22_X1 U17490 ( .A1(n20390), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n15564) );
  OAI21_X1 U17491 ( .B1(n22354), .B2(n15576), .A(n15564), .ZN(P1_U2913) );
  AOI22_X1 U17492 ( .A1(n21862), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n15565) );
  OAI21_X1 U17493 ( .B1(n22385), .B2(n15576), .A(n15565), .ZN(P1_U2908) );
  AOI22_X1 U17494 ( .A1(n21862), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n15566) );
  OAI21_X1 U17495 ( .B1(n22393), .B2(n15576), .A(n15566), .ZN(P1_U2907) );
  AOI22_X1 U17496 ( .A1(n21862), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n15567) );
  OAI21_X1 U17497 ( .B1(n22402), .B2(n15576), .A(n15567), .ZN(P1_U2906) );
  INV_X1 U17498 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n22343) );
  AOI22_X1 U17499 ( .A1(n21862), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n15568) );
  OAI21_X1 U17500 ( .B1(n22343), .B2(n15576), .A(n15568), .ZN(P1_U2915) );
  AOI22_X1 U17501 ( .A1(n21862), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n15569) );
  OAI21_X1 U17502 ( .B1(n16619), .B2(n15576), .A(n15569), .ZN(P1_U2912) );
  INV_X1 U17503 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n22364) );
  AOI22_X1 U17504 ( .A1(n21862), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n15570) );
  OAI21_X1 U17505 ( .B1(n22364), .B2(n15576), .A(n15570), .ZN(P1_U2911) );
  AOI22_X1 U17506 ( .A1(n21862), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n15571) );
  OAI21_X1 U17507 ( .B1(n22336), .B2(n15576), .A(n15571), .ZN(P1_U2916) );
  INV_X1 U17508 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n22378) );
  AOI22_X1 U17509 ( .A1(n21862), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n15572) );
  OAI21_X1 U17510 ( .B1(n22378), .B2(n15576), .A(n15572), .ZN(P1_U2909) );
  INV_X1 U17511 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n22348) );
  AOI22_X1 U17512 ( .A1(n21862), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n15573) );
  OAI21_X1 U17513 ( .B1(n22348), .B2(n15576), .A(n15573), .ZN(P1_U2914) );
  INV_X1 U17514 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n22330) );
  AOI22_X1 U17515 ( .A1(n21862), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n15574) );
  OAI21_X1 U17516 ( .B1(n22330), .B2(n15576), .A(n15574), .ZN(P1_U2917) );
  INV_X1 U17517 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n22371) );
  AOI22_X1 U17518 ( .A1(n21862), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n15575) );
  OAI21_X1 U17519 ( .B1(n22371), .B2(n15576), .A(n15575), .ZN(P1_U2910) );
  OAI21_X1 U17520 ( .B1(n22189), .B2(n15578), .A(n15577), .ZN(n15586) );
  INV_X1 U17521 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15779) );
  OR2_X1 U17522 ( .A1(n15580), .A2(n15579), .ZN(n15581) );
  NAND2_X1 U17523 ( .A1(n14069), .A2(n15581), .ZN(n21884) );
  OAI22_X1 U17524 ( .A1(n15674), .A2(n22201), .B1(n22208), .B2(n21884), .ZN(
        n15582) );
  AOI211_X1 U17525 ( .C1(n22187), .C2(n15783), .A(n22170), .B(n15582), .ZN(
        n15583) );
  OAI21_X1 U17526 ( .B1(n15779), .B2(n22152), .A(n15583), .ZN(n15584) );
  AOI21_X1 U17527 ( .B1(n15586), .B2(n15585), .A(n15584), .ZN(n15587) );
  OAI21_X1 U17528 ( .B1(n22209), .B2(n15780), .A(n15587), .ZN(P1_U2831) );
  INV_X1 U17529 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15595) );
  INV_X1 U17530 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20620) );
  OAI22_X1 U17531 ( .A1(n13670), .A2(n22632), .B1(n22630), .B2(n20620), .ZN(
        n15588) );
  CLKBUF_X1 U17532 ( .A(n15588), .Z(n22682) );
  INV_X1 U17533 ( .A(n22341), .ZN(n16635) );
  NAND2_X1 U17534 ( .A1(n22626), .A2(n16635), .ZN(n22685) );
  AOI22_X1 U17535 ( .A1(n15639), .A2(n22682), .B1(n15638), .B2(n22798), .ZN(
        n15594) );
  INV_X1 U17536 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20605) );
  INV_X1 U17537 ( .A(DATAI_21_), .ZN(n15589) );
  OR2_X1 U17538 ( .A1(n22632), .A2(n15589), .ZN(n15590) );
  NOR2_X2 U17539 ( .A1(n22629), .A2(n15592), .ZN(n22681) );
  AOI22_X1 U17540 ( .A1(n22800), .A2(n15591), .B1(n22681), .B2(n22796), .ZN(
        n15593) );
  OAI211_X1 U17541 ( .C1(n15596), .C2(n15595), .A(n15594), .B(n15593), .ZN(
        P1_U3158) );
  INV_X1 U17542 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15599) );
  AOI22_X1 U17543 ( .A1(n15633), .A2(n15591), .B1(n15638), .B2(n22699), .ZN(
        n15598) );
  AOI22_X1 U17544 ( .A1(n22750), .A2(n22682), .B1(n22681), .B2(n22698), .ZN(
        n15597) );
  OAI211_X1 U17545 ( .C1(n15600), .C2(n15599), .A(n15598), .B(n15597), .ZN(
        P1_U3070) );
  INV_X1 U17546 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15603) );
  AOI22_X1 U17547 ( .A1(n22781), .A2(n22682), .B1(n15638), .B2(n22790), .ZN(
        n15602) );
  AOI22_X1 U17548 ( .A1(n22791), .A2(n15591), .B1(n22681), .B2(n22789), .ZN(
        n15601) );
  OAI211_X1 U17549 ( .C1(n15604), .C2(n15603), .A(n15602), .B(n15601), .ZN(
        P1_U3142) );
  XOR2_X1 U17550 ( .A(n15606), .B(n15605), .Z(n15662) );
  INV_X1 U17551 ( .A(n15662), .ZN(n15615) );
  INV_X1 U17552 ( .A(n22078), .ZN(n15613) );
  NOR2_X1 U17553 ( .A1(n21975), .A2(n22082), .ZN(n15664) );
  INV_X1 U17554 ( .A(n15607), .ZN(n15609) );
  NOR2_X1 U17555 ( .A1(n15609), .A2(n15608), .ZN(n16876) );
  OAI22_X1 U17556 ( .A1(n16788), .A2(n15611), .B1(n15610), .B2(n16786), .ZN(
        n21888) );
  INV_X1 U17557 ( .A(n21888), .ZN(n16843) );
  AOI22_X1 U17558 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16876), .B1(
        n16843), .B2(n12895), .ZN(n15612) );
  AOI211_X1 U17559 ( .C1(n21993), .C2(n15613), .A(n15664), .B(n15612), .ZN(
        n15614) );
  OAI21_X1 U17560 ( .B1(n15615), .B2(n22010), .A(n15614), .ZN(P1_U3025) );
  INV_X1 U17561 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15618) );
  AOI22_X1 U17562 ( .A1(n22737), .A2(n22682), .B1(n15638), .B2(n22689), .ZN(
        n15617) );
  AOI22_X1 U17563 ( .A1(n22743), .A2(n15591), .B1(n22688), .B2(n22681), .ZN(
        n15616) );
  OAI211_X1 U17564 ( .C1(n15619), .C2(n15618), .A(n15617), .B(n15616), .ZN(
        P1_U3046) );
  INV_X1 U17565 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15622) );
  AOI22_X1 U17566 ( .A1(n22761), .A2(n22682), .B1(n15638), .B2(n22706), .ZN(
        n15621) );
  AOI22_X1 U17567 ( .A1(n22713), .A2(n15591), .B1(n22705), .B2(n22681), .ZN(
        n15620) );
  OAI211_X1 U17568 ( .C1(n15623), .C2(n15622), .A(n15621), .B(n15620), .ZN(
        P1_U3094) );
  INV_X1 U17569 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15627) );
  AOI22_X1 U17570 ( .A1(n15624), .A2(n22682), .B1(n15638), .B2(n22768), .ZN(
        n15626) );
  AOI22_X1 U17571 ( .A1(n22774), .A2(n15591), .B1(n22767), .B2(n22681), .ZN(
        n15625) );
  OAI211_X1 U17572 ( .C1(n15628), .C2(n15627), .A(n15626), .B(n15625), .ZN(
        P1_U3110) );
  INV_X1 U17573 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15631) );
  AOI22_X1 U17574 ( .A1(n22775), .A2(n22682), .B1(n15638), .B2(n22720), .ZN(
        n15630) );
  AOI22_X1 U17575 ( .A1(n22783), .A2(n15591), .B1(n22719), .B2(n22681), .ZN(
        n15629) );
  OAI211_X1 U17576 ( .C1(n15632), .C2(n15631), .A(n15630), .B(n15629), .ZN(
        P1_U3126) );
  INV_X1 U17577 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15636) );
  AOI22_X1 U17578 ( .A1(n15633), .A2(n22682), .B1(n15638), .B2(n22756), .ZN(
        n15635) );
  AOI22_X1 U17579 ( .A1(n22762), .A2(n15591), .B1(n22755), .B2(n22681), .ZN(
        n15634) );
  OAI211_X1 U17580 ( .C1(n15637), .C2(n15636), .A(n15635), .B(n15634), .ZN(
        P1_U3078) );
  INV_X1 U17581 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15642) );
  AOI22_X1 U17582 ( .A1(n15638), .A2(n22731), .B1(n22791), .B2(n22682), .ZN(
        n15641) );
  AOI22_X1 U17583 ( .A1(n15639), .A2(n15591), .B1(n22729), .B2(n22681), .ZN(
        n15640) );
  OAI211_X1 U17584 ( .C1(n15643), .C2(n15642), .A(n15641), .B(n15640), .ZN(
        P1_U3150) );
  AOI22_X1 U17585 ( .A1(n15646), .A2(n15645), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15644), .ZN(n15648) );
  XNOR2_X1 U17586 ( .A(n16025), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15647) );
  XNOR2_X1 U17587 ( .A(n15648), .B(n15647), .ZN(n17766) );
  INV_X1 U17588 ( .A(n17766), .ZN(n15661) );
  XNOR2_X1 U17589 ( .A(n15649), .B(n15743), .ZN(n17764) );
  NAND2_X1 U17590 ( .A1(n15650), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15741) );
  OAI21_X1 U17591 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17581), .A(
        n17584), .ZN(n15745) );
  INV_X1 U17592 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n17863) );
  NOR2_X1 U17593 ( .A1(n17863), .A2(n19068), .ZN(n15653) );
  NOR2_X1 U17594 ( .A1(n17622), .A2(n15651), .ZN(n15652) );
  AOI211_X1 U17595 ( .C1(n15745), .C2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n15653), .B(n15652), .ZN(n15658) );
  OR2_X1 U17596 ( .A1(n15655), .A2(n15654), .ZN(n15656) );
  AND2_X1 U17597 ( .A1(n15656), .A2(n15739), .ZN(n17765) );
  NAND2_X1 U17598 ( .A1(n17765), .A2(n17633), .ZN(n15657) );
  OAI211_X1 U17599 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n15741), .A(
        n15658), .B(n15657), .ZN(n15659) );
  AOI21_X1 U17600 ( .B1(n17764), .B2(n17628), .A(n15659), .ZN(n15660) );
  OAI21_X1 U17601 ( .B1(n15661), .B2(n19182), .A(n15660), .ZN(P2_U3042) );
  NAND2_X1 U17602 ( .A1(n15662), .A2(n20556), .ZN(n15666) );
  NOR2_X1 U17603 ( .A1(n20561), .A2(n22087), .ZN(n15663) );
  AOI211_X1 U17604 ( .C1(n20551), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n15664), .B(n15663), .ZN(n15665) );
  OAI211_X1 U17605 ( .C1(n20538), .C2(n22076), .A(n15666), .B(n15665), .ZN(
        P1_U2993) );
  INV_X1 U17606 ( .A(n22682), .ZN(n15667) );
  OAI22_X1 U17607 ( .A1(n22685), .A2(n22473), .B1(n15667), .B2(n22710), .ZN(
        n15672) );
  INV_X1 U17608 ( .A(n15591), .ZN(n15670) );
  INV_X1 U17609 ( .A(n22681), .ZN(n15669) );
  OAI22_X1 U17610 ( .A1(n22772), .A2(n15670), .B1(n15669), .B2(n15668), .ZN(
        n15671) );
  AOI211_X1 U17611 ( .C1(n22714), .C2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n15672), .B(n15671), .ZN(n15673) );
  INV_X1 U17612 ( .A(n15673), .ZN(P1_U3102) );
  OAI222_X1 U17613 ( .A1(n21884), .A2(n20480), .B1(n20493), .B2(n15674), .C1(
        n20483), .C2(n15780), .ZN(P1_U2863) );
  AOI22_X1 U17614 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15678) );
  AOI22_X1 U17615 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15677) );
  AOI22_X1 U17616 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15676) );
  AOI22_X1 U17617 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15675) );
  NAND4_X1 U17618 ( .A1(n15678), .A2(n15677), .A3(n15676), .A4(n15675), .ZN(
        n15684) );
  AOI22_X1 U17619 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15682) );
  AOI22_X1 U17620 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11159), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15681) );
  AOI22_X1 U17621 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U17622 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15679) );
  NAND4_X1 U17623 ( .A1(n15682), .A2(n15681), .A3(n15680), .A4(n15679), .ZN(
        n15683) );
  OR2_X1 U17624 ( .A1(n15684), .A2(n15683), .ZN(n15686) );
  NOR2_X1 U17625 ( .A1(n15685), .A2(n15686), .ZN(n15687) );
  OR2_X1 U17626 ( .A1(n15772), .A2(n15687), .ZN(n20229) );
  NAND2_X1 U17627 ( .A1(n15444), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15693) );
  OR2_X1 U17628 ( .A1(n15689), .A2(n15690), .ZN(n15691) );
  AND2_X1 U17629 ( .A1(n15688), .A2(n15691), .ZN(n17466) );
  NAND2_X1 U17630 ( .A1(n17466), .A2(n17044), .ZN(n15692) );
  OAI211_X1 U17631 ( .C1(n20229), .C2(n17034), .A(n15693), .B(n15692), .ZN(
        P2_U2871) );
  XNOR2_X1 U17632 ( .A(n15694), .B(n15695), .ZN(n15714) );
  INV_X1 U17633 ( .A(n15696), .ZN(n20490) );
  AND2_X1 U17634 ( .A1(n21999), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n15711) );
  AOI21_X1 U17635 ( .B1(n20551), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n15711), .ZN(n15697) );
  OAI21_X1 U17636 ( .B1(n20561), .B2(n15698), .A(n15697), .ZN(n15699) );
  AOI21_X1 U17637 ( .B1(n20490), .B2(n20557), .A(n15699), .ZN(n15700) );
  OAI21_X1 U17638 ( .B1(n15714), .B2(n22216), .A(n15700), .ZN(P1_U2991) );
  AND2_X1 U17639 ( .A1(n15702), .A2(n15701), .ZN(n15703) );
  OR2_X1 U17640 ( .A1(n15703), .A2(n15689), .ZN(n19041) );
  INV_X1 U17641 ( .A(n19041), .ZN(n17482) );
  NOR2_X1 U17642 ( .A1(n17044), .A2(n13225), .ZN(n15707) );
  AOI211_X1 U17643 ( .C1(n15705), .C2(n15704), .A(n17034), .B(n15685), .ZN(
        n15706) );
  AOI211_X1 U17644 ( .C1(n17482), .C2(n17044), .A(n15707), .B(n15706), .ZN(
        n15708) );
  INV_X1 U17645 ( .A(n15708), .ZN(P2_U2872) );
  INV_X1 U17646 ( .A(n21920), .ZN(n16791) );
  NOR2_X1 U17647 ( .A1(n16798), .A2(n16791), .ZN(n21940) );
  AOI21_X1 U17648 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16876), .A(
        n21940), .ZN(n15721) );
  NOR2_X1 U17649 ( .A1(n16843), .A2(n12895), .ZN(n15720) );
  XOR2_X1 U17650 ( .A(n15709), .B(n15719), .Z(n15710) );
  AOI22_X1 U17651 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15721), .B1(
        n15720), .B2(n15710), .ZN(n15713) );
  AOI21_X1 U17652 ( .B1(n20487), .B2(n21993), .A(n15711), .ZN(n15712) );
  OAI211_X1 U17653 ( .C1(n15714), .C2(n22010), .A(n15713), .B(n15712), .ZN(
        P1_U3023) );
  INV_X1 U17654 ( .A(n20509), .ZN(n15724) );
  MUX2_X1 U17655 ( .A(BUF1_REG_10__SCAN_IN), .B(DATAI_10_), .S(n16592), .Z(
        n22368) );
  AOI22_X1 U17656 ( .A1(n15948), .A2(n22368), .B1(n16653), .B2(
        P1_EAX_REG_10__SCAN_IN), .ZN(n15715) );
  OAI21_X1 U17657 ( .B1(n15724), .B2(n16667), .A(n15715), .ZN(P1_U2894) );
  XOR2_X1 U17658 ( .A(n15717), .B(n15716), .Z(n20502) );
  INV_X1 U17659 ( .A(n20502), .ZN(n15723) );
  NAND2_X1 U17660 ( .A1(n21999), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n20503) );
  OAI21_X1 U17661 ( .B1(n22009), .B2(n22088), .A(n20503), .ZN(n15718) );
  AOI221_X1 U17662 ( .B1(n15721), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n15720), .C2(n15719), .A(n15718), .ZN(n15722) );
  OAI21_X1 U17663 ( .B1(n15723), .B2(n22010), .A(n15722), .ZN(P1_U3024) );
  OAI222_X1 U17664 ( .A1(n20493), .A2(n15725), .B1(n20483), .B2(n15724), .C1(
        n16882), .C2(n20480), .ZN(P1_U2862) );
  NAND2_X1 U17665 ( .A1(n19032), .A2(n15726), .ZN(n15727) );
  XNOR2_X1 U17666 ( .A(n17753), .B(n15727), .ZN(n15728) );
  NAND2_X1 U17667 ( .A1(n15728), .A2(n19167), .ZN(n15735) );
  OAI22_X1 U17668 ( .A1(n19108), .A2(n13623), .B1(n17861), .B2(n19111), .ZN(
        n15731) );
  NOR2_X1 U17669 ( .A1(n19144), .A2(n15729), .ZN(n15730) );
  AOI211_X1 U17670 ( .C1(n19159), .C2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15731), .B(n15730), .ZN(n15732) );
  OAI21_X1 U17671 ( .B1(n17806), .B2(n19161), .A(n15732), .ZN(n15733) );
  AOI21_X1 U17672 ( .B1(n14864), .B2(n19131), .A(n15733), .ZN(n15734) );
  OAI211_X1 U17673 ( .C1(n16973), .C2(n19768), .A(n15735), .B(n15734), .ZN(
        P2_U2852) );
  XNOR2_X1 U17674 ( .A(n15736), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15737) );
  XNOR2_X1 U17675 ( .A(n15738), .B(n15737), .ZN(n15760) );
  NAND3_X1 U17676 ( .A1(n15754), .A2(n17628), .A3(n15753), .ZN(n15752) );
  AOI21_X1 U17677 ( .B1(n15740), .B2(n15739), .A(n14937), .ZN(n18979) );
  INV_X1 U17678 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n18971) );
  AOI221_X1 U17679 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n15743), .C2(n15742), .A(
        n15741), .ZN(n15744) );
  AOI21_X1 U17680 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n15745), .A(
        n15744), .ZN(n15746) );
  OAI21_X1 U17681 ( .B1(n19068), .B2(n18971), .A(n15746), .ZN(n15750) );
  OAI21_X1 U17682 ( .B1(n11313), .B2(n15748), .A(n15747), .ZN(n19978) );
  NOR2_X1 U17683 ( .A1(n19978), .A2(n17622), .ZN(n15749) );
  AOI211_X1 U17684 ( .C1(n18979), .C2(n17633), .A(n15750), .B(n15749), .ZN(
        n15751) );
  OAI211_X1 U17685 ( .C1(n15760), .C2(n19182), .A(n15752), .B(n15751), .ZN(
        P2_U3041) );
  NAND3_X1 U17686 ( .A1(n15754), .A2(n17782), .A3(n15753), .ZN(n15759) );
  INV_X1 U17687 ( .A(n18979), .ZN(n16012) );
  NOR2_X1 U17688 ( .A1(n17773), .A2(n16012), .ZN(n15757) );
  OAI22_X1 U17689 ( .A1(n15755), .A2(n17762), .B1(n18971), .B2(n19068), .ZN(
        n15756) );
  AOI211_X1 U17690 ( .C1(n18978), .C2(n17754), .A(n15757), .B(n15756), .ZN(
        n15758) );
  OAI211_X1 U17691 ( .C1(n17774), .C2(n15760), .A(n15759), .B(n15758), .ZN(
        P2_U3009) );
  AOI22_X1 U17692 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15764) );
  AOI22_X1 U17693 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15763) );
  AOI22_X1 U17694 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15762) );
  AOI22_X1 U17695 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15761) );
  NAND4_X1 U17696 ( .A1(n15764), .A2(n15763), .A3(n15762), .A4(n15761), .ZN(
        n15770) );
  AOI22_X1 U17697 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15768) );
  AOI22_X1 U17698 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11159), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15767) );
  AOI22_X1 U17699 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15766) );
  AOI22_X1 U17700 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15765) );
  NAND4_X1 U17701 ( .A1(n15768), .A2(n15767), .A3(n15766), .A4(n15765), .ZN(
        n15769) );
  OR2_X1 U17702 ( .A1(n15770), .A2(n15769), .ZN(n15771) );
  OAI21_X1 U17703 ( .B1(n15772), .B2(n15771), .A(n15870), .ZN(n15859) );
  NAND2_X1 U17704 ( .A1(n15444), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15775) );
  XOR2_X1 U17705 ( .A(n15773), .B(n15688), .Z(n19046) );
  NAND2_X1 U17706 ( .A1(n19046), .A2(n17044), .ZN(n15774) );
  OAI211_X1 U17707 ( .C1(n15859), .C2(n17034), .A(n15775), .B(n15774), .ZN(
        P2_U2870) );
  OAI22_X1 U17708 ( .A1(n20506), .A2(n15779), .B1(n15578), .B2(n21975), .ZN(
        n15782) );
  NOR2_X1 U17709 ( .A1(n15780), .A2(n20538), .ZN(n15781) );
  AOI211_X1 U17710 ( .C1(n20520), .C2(n15783), .A(n15782), .B(n15781), .ZN(
        n15784) );
  OAI21_X1 U17711 ( .B1(n22216), .B2(n21879), .A(n15784), .ZN(P1_U2990) );
  NOR2_X1 U17712 ( .A1(n19134), .A2(n15785), .ZN(n15786) );
  XNOR2_X1 U17713 ( .A(n15786), .B(n17239), .ZN(n15796) );
  NAND2_X1 U17714 ( .A1(n15787), .A2(n15788), .ZN(n15789) );
  NAND2_X1 U17715 ( .A1(n15851), .A2(n15789), .ZN(n20226) );
  INV_X1 U17716 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n17878) );
  AOI22_X1 U17717 ( .A1(n15790), .A2(n19156), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19158), .ZN(n15791) );
  OAI211_X1 U17718 ( .C1(n17878), .C2(n19111), .A(n15791), .B(n19068), .ZN(
        n15792) );
  AOI21_X1 U17719 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19159), .A(
        n15792), .ZN(n15794) );
  NAND2_X1 U17720 ( .A1(n17466), .A2(n19131), .ZN(n15793) );
  OAI211_X1 U17721 ( .C1(n19161), .C2(n20226), .A(n15794), .B(n15793), .ZN(
        n15795) );
  AOI21_X1 U17722 ( .B1(n15796), .B2(n19167), .A(n15795), .ZN(n15797) );
  INV_X1 U17723 ( .A(n15797), .ZN(P2_U2839) );
  NOR2_X1 U17724 ( .A1(n19134), .A2(n19017), .ZN(n15798) );
  XNOR2_X1 U17725 ( .A(n15798), .B(n17268), .ZN(n15809) );
  AOI22_X1 U17726 ( .A1(n15799), .A2(n19156), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19158), .ZN(n15800) );
  OAI211_X1 U17727 ( .C1(n13218), .C2(n19111), .A(n15800), .B(n19068), .ZN(
        n15801) );
  AOI21_X1 U17728 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19159), .A(
        n15801), .ZN(n15802) );
  INV_X1 U17729 ( .A(n15802), .ZN(n15808) );
  NOR2_X1 U17730 ( .A1(n15805), .A2(n15804), .ZN(n15806) );
  OR2_X1 U17731 ( .A1(n15803), .A2(n15806), .ZN(n19695) );
  OAI22_X1 U17732 ( .A1(n17493), .A2(n19163), .B1(n19695), .B2(n19161), .ZN(
        n15807) );
  AOI211_X1 U17733 ( .C1(n15809), .C2(n19167), .A(n15808), .B(n15807), .ZN(
        n15810) );
  INV_X1 U17734 ( .A(n15810), .ZN(P2_U2841) );
  AOI21_X1 U17735 ( .B1(n15811), .B2(n15813), .A(n15812), .ZN(n17551) );
  INV_X1 U17736 ( .A(n17551), .ZN(n19707) );
  NOR2_X1 U17737 ( .A1(n19134), .A2(n15814), .ZN(n15815) );
  XNOR2_X1 U17738 ( .A(n15815), .B(n17312), .ZN(n15816) );
  NAND2_X1 U17739 ( .A1(n15816), .A2(n19167), .ZN(n15824) );
  OAI21_X1 U17740 ( .B1(n19037), .B2(n11681), .A(n19068), .ZN(n15817) );
  AOI21_X1 U17741 ( .B1(n19155), .B2(P2_REIP_REG_10__SCAN_IN), .A(n15817), 
        .ZN(n15818) );
  OAI21_X1 U17742 ( .B1(n19108), .B2(n15819), .A(n15818), .ZN(n15822) );
  NOR2_X1 U17743 ( .A1(n15820), .A2(n19144), .ZN(n15821) );
  AOI211_X1 U17744 ( .C1(n19131), .C2(n17310), .A(n15822), .B(n15821), .ZN(
        n15823) );
  OAI211_X1 U17745 ( .C1(n19161), .C2(n19707), .A(n15824), .B(n15823), .ZN(
        P2_U2845) );
  NOR2_X1 U17746 ( .A1(n19134), .A2(n16962), .ZN(n15826) );
  XNOR2_X1 U17747 ( .A(n15826), .B(n15825), .ZN(n15827) );
  NAND2_X1 U17748 ( .A1(n15827), .A2(n19167), .ZN(n15834) );
  INV_X1 U17749 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n17859) );
  OAI22_X1 U17750 ( .A1(n19108), .A2(n13621), .B1(n17859), .B2(n19111), .ZN(
        n15828) );
  AOI21_X1 U17751 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19159), .A(
        n15828), .ZN(n15830) );
  NAND2_X1 U17752 ( .A1(n17795), .A2(n19118), .ZN(n15829) );
  OAI211_X1 U17753 ( .C1(n19144), .C2(n15831), .A(n15830), .B(n15829), .ZN(
        n15832) );
  AOI21_X1 U17754 ( .B1(n14808), .B2(n19131), .A(n15832), .ZN(n15833) );
  OAI211_X1 U17755 ( .C1(n16973), .C2(n17805), .A(n15834), .B(n15833), .ZN(
        P2_U2853) );
  NOR2_X1 U17756 ( .A1(n19134), .A2(n15835), .ZN(n15836) );
  XNOR2_X1 U17757 ( .A(n15836), .B(n17789), .ZN(n15837) );
  NAND2_X1 U17758 ( .A1(n15837), .A2(n19167), .ZN(n15847) );
  AOI21_X1 U17759 ( .B1(n15839), .B2(n17600), .A(n15838), .ZN(n19711) );
  NAND2_X1 U17760 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19159), .ZN(
        n15840) );
  OAI211_X1 U17761 ( .C1(n19111), .C2(n15841), .A(n19068), .B(n15840), .ZN(
        n15845) );
  OAI22_X1 U17762 ( .A1(n19163), .A2(n15843), .B1(n19108), .B2(n15842), .ZN(
        n15844) );
  AOI211_X1 U17763 ( .C1(n19118), .C2(n19711), .A(n15845), .B(n15844), .ZN(
        n15846) );
  OAI211_X1 U17764 ( .C1(n19144), .C2(n15848), .A(n15847), .B(n15846), .ZN(
        P2_U2847) );
  AOI22_X1 U17765 ( .A1(n20225), .A2(BUF2_REG_17__SCAN_IN), .B1(n20224), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n15856) );
  AND2_X1 U17766 ( .A1(n15851), .A2(n15850), .ZN(n15853) );
  OR2_X1 U17767 ( .A1(n15853), .A2(n15852), .ZN(n19061) );
  INV_X1 U17768 ( .A(n19061), .ZN(n15854) );
  AOI22_X1 U17769 ( .A1(n20169), .A2(n15854), .B1(n20221), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15855) );
  OAI211_X1 U17770 ( .C1(n20177), .C2(n17123), .A(n15856), .B(n15855), .ZN(
        n15857) );
  INV_X1 U17771 ( .A(n15857), .ZN(n15858) );
  OAI21_X1 U17772 ( .B1(n15859), .B2(n20228), .A(n15858), .ZN(P2_U2902) );
  INV_X1 U17773 ( .A(n16954), .ZN(n15874) );
  AOI22_X1 U17774 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15863) );
  AOI22_X1 U17775 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15862) );
  AOI22_X1 U17776 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15861) );
  AOI22_X1 U17777 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15860) );
  NAND4_X1 U17778 ( .A1(n15863), .A2(n15862), .A3(n15861), .A4(n15860), .ZN(
        n15869) );
  AOI22_X1 U17779 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15867) );
  AOI22_X1 U17780 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16234), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15866) );
  AOI22_X1 U17781 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15865) );
  AOI22_X1 U17782 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15864) );
  NAND4_X1 U17783 ( .A1(n15867), .A2(n15866), .A3(n15865), .A4(n15864), .ZN(
        n15868) );
  NOR2_X1 U17784 ( .A1(n15869), .A2(n15868), .ZN(n15871) );
  NOR2_X4 U17785 ( .A1(n15870), .A2(n15871), .ZN(n15902) );
  INV_X1 U17786 ( .A(n15902), .ZN(n15903) );
  AOI21_X1 U17787 ( .B1(n15871), .B2(n15870), .A(n15902), .ZN(n20124) );
  NAND2_X1 U17788 ( .A1(n20124), .A2(n17039), .ZN(n15873) );
  NAND2_X1 U17789 ( .A1(n15444), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15872) );
  OAI211_X1 U17790 ( .C1(n15874), .C2(n15444), .A(n15873), .B(n15872), .ZN(
        P2_U2869) );
  OAI21_X1 U17791 ( .B1(n11819), .B2(n11324), .A(n15875), .ZN(n15886) );
  XNOR2_X1 U17792 ( .A(n15886), .B(n15885), .ZN(n22104) );
  MUX2_X1 U17793 ( .A(BUF1_REG_11__SCAN_IN), .B(DATAI_11_), .S(n16592), .Z(
        n22375) );
  AOI22_X1 U17794 ( .A1(n15948), .A2(n22375), .B1(n16653), .B2(
        P1_EAX_REG_11__SCAN_IN), .ZN(n15876) );
  OAI21_X1 U17795 ( .B1(n22104), .B2(n16667), .A(n15876), .ZN(P1_U2893) );
  OAI21_X1 U17796 ( .B1(n15877), .B2(n15879), .A(n15878), .ZN(n20472) );
  MUX2_X1 U17797 ( .A(BUF1_REG_14__SCAN_IN), .B(DATAI_14_), .S(n16592), .Z(
        n22397) );
  AOI22_X1 U17798 ( .A1(n15948), .A2(n22397), .B1(n16653), .B2(
        P1_EAX_REG_14__SCAN_IN), .ZN(n15880) );
  OAI21_X1 U17799 ( .B1(n20472), .B2(n16667), .A(n15880), .ZN(P1_U2890) );
  AND2_X1 U17800 ( .A1(n15882), .A2(n15881), .ZN(n15883) );
  OR2_X1 U17801 ( .A1(n15883), .A2(n15921), .ZN(n22101) );
  OAI222_X1 U17802 ( .A1(n22101), .A2(n20480), .B1(n20493), .B2(n15884), .C1(
        n20483), .C2(n22104), .ZN(P1_U2861) );
  OAI21_X1 U17803 ( .B1(n15886), .B2(n15885), .A(n15875), .ZN(n15938) );
  XNOR2_X1 U17804 ( .A(n15938), .B(n15937), .ZN(n22120) );
  MUX2_X1 U17805 ( .A(BUF1_REG_12__SCAN_IN), .B(DATAI_12_), .S(n16592), .Z(
        n22382) );
  AOI22_X1 U17806 ( .A1(n15948), .A2(n22382), .B1(n16653), .B2(
        P1_EAX_REG_12__SCAN_IN), .ZN(n15887) );
  OAI21_X1 U17807 ( .B1(n22120), .B2(n16667), .A(n15887), .ZN(P1_U2892) );
  AND2_X1 U17808 ( .A1(n15889), .A2(n15888), .ZN(n15890) );
  OR2_X1 U17809 ( .A1(n15890), .A2(n14472), .ZN(n17436) );
  AOI22_X1 U17810 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15894) );
  AOI22_X1 U17811 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15893) );
  AOI22_X1 U17812 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15892) );
  AOI22_X1 U17813 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15891) );
  NAND4_X1 U17814 ( .A1(n15894), .A2(n15893), .A3(n15892), .A4(n15891), .ZN(
        n15900) );
  AOI22_X1 U17815 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15898) );
  AOI22_X1 U17816 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16234), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15897) );
  AOI22_X1 U17817 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15896) );
  AOI22_X1 U17818 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15895) );
  NAND4_X1 U17819 ( .A1(n15898), .A2(n15897), .A3(n15896), .A4(n15895), .ZN(
        n15899) );
  NOR2_X1 U17820 ( .A1(n15900), .A2(n15899), .ZN(n15904) );
  AOI21_X1 U17821 ( .B1(n15904), .B2(n15903), .A(n16201), .ZN(n17125) );
  NAND2_X1 U17822 ( .A1(n17125), .A2(n17039), .ZN(n15906) );
  NAND2_X1 U17823 ( .A1(n15444), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15905) );
  OAI211_X1 U17824 ( .C1(n15444), .C2(n17436), .A(n15906), .B(n15905), .ZN(
        P2_U2868) );
  OAI21_X1 U17825 ( .B1(n15812), .B2(n15908), .A(n15907), .ZN(n19704) );
  NAND2_X1 U17826 ( .A1(n19032), .A2(n19167), .ZN(n15959) );
  NOR2_X1 U17827 ( .A1(n15909), .A2(n15959), .ZN(n15933) );
  OAI21_X1 U17828 ( .B1(n15910), .B2(n17299), .A(n15933), .ZN(n15918) );
  INV_X1 U17829 ( .A(n15911), .ZN(n15916) );
  NAND2_X1 U17830 ( .A1(n19167), .A2(n19134), .ZN(n19049) );
  OAI22_X1 U17831 ( .A1(n15912), .A2(n19163), .B1(n19049), .B2(n17299), .ZN(
        n15915) );
  AOI22_X1 U17832 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19159), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n19158), .ZN(n15913) );
  OAI211_X1 U17833 ( .C1(n17872), .C2(n19111), .A(n15913), .B(n19068), .ZN(
        n15914) );
  AOI211_X1 U17834 ( .C1(n19156), .C2(n15916), .A(n15915), .B(n15914), .ZN(
        n15917) );
  OAI211_X1 U17835 ( .C1(n19704), .C2(n19161), .A(n15918), .B(n15917), .ZN(
        P2_U2844) );
  INV_X1 U17836 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15922) );
  OAI21_X1 U17837 ( .B1(n15921), .B2(n15920), .A(n15919), .ZN(n21885) );
  OAI222_X1 U17838 ( .A1(n22120), .A2(n20483), .B1(n20493), .B2(n15922), .C1(
        n20480), .C2(n21885), .ZN(P1_U2860) );
  AOI21_X1 U17839 ( .B1(n15924), .B2(n15907), .A(n15923), .ZN(n17526) );
  INV_X1 U17840 ( .A(n17526), .ZN(n19701) );
  AOI211_X1 U17841 ( .C1(n19032), .C2(n15925), .A(n19201), .B(n17289), .ZN(
        n15928) );
  AOI22_X1 U17842 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19159), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n19158), .ZN(n15926) );
  NAND2_X1 U17843 ( .A1(n19068), .A2(n15926), .ZN(n15927) );
  AOI211_X1 U17844 ( .C1(n19155), .C2(P2_REIP_REG_12__SCAN_IN), .A(n15928), 
        .B(n15927), .ZN(n15929) );
  OAI21_X1 U17845 ( .B1(n15930), .B2(n19163), .A(n15929), .ZN(n15931) );
  AOI21_X1 U17846 ( .B1(n19156), .B2(n15932), .A(n15931), .ZN(n15935) );
  NAND2_X1 U17847 ( .A1(n15933), .A2(n17289), .ZN(n15934) );
  OAI211_X1 U17848 ( .C1(n19701), .C2(n19161), .A(n15935), .B(n15934), .ZN(
        P2_U2843) );
  AOI21_X1 U17849 ( .B1(n15938), .B2(n15937), .A(n15936), .ZN(n15939) );
  NOR2_X1 U17850 ( .A1(n15939), .A2(n15877), .ZN(n16778) );
  INV_X1 U17851 ( .A(n16778), .ZN(n15955) );
  OR3_X1 U17852 ( .A1(n22114), .A2(n22113), .A3(n22103), .ZN(n22115) );
  OAI21_X1 U17853 ( .B1(n22189), .B2(n15940), .A(n22115), .ZN(n15946) );
  INV_X1 U17854 ( .A(n22121), .ZN(n16534) );
  INV_X1 U17855 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15956) );
  NAND2_X1 U17856 ( .A1(n15919), .A2(n15941), .ZN(n15942) );
  NAND2_X1 U17857 ( .A1(n16847), .A2(n15942), .ZN(n21870) );
  OAI22_X1 U17858 ( .A1(n15956), .A2(n22201), .B1(n22208), .B2(n21870), .ZN(
        n15943) );
  AOI211_X1 U17859 ( .C1(n22206), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n22170), .B(n15943), .ZN(n15944) );
  OAI21_X1 U17860 ( .B1(n22203), .B2(n16776), .A(n15944), .ZN(n15945) );
  AOI21_X1 U17861 ( .B1(n15946), .B2(n16534), .A(n15945), .ZN(n15947) );
  OAI21_X1 U17862 ( .B1(n15955), .B2(n22209), .A(n15947), .ZN(P1_U2827) );
  MUX2_X1 U17863 ( .A(BUF1_REG_13__SCAN_IN), .B(DATAI_13_), .S(n16592), .Z(
        n22390) );
  AOI22_X1 U17864 ( .A1(n15948), .A2(n22390), .B1(n16653), .B2(
        P1_EAX_REG_13__SCAN_IN), .ZN(n15949) );
  OAI21_X1 U17865 ( .B1(n15955), .B2(n16667), .A(n15949), .ZN(P1_U2891) );
  INV_X1 U17866 ( .A(n15950), .ZN(n16657) );
  NAND2_X1 U17867 ( .A1(n15878), .A2(n15951), .ZN(n15952) );
  NAND2_X1 U17868 ( .A1(n16657), .A2(n15952), .ZN(n16766) );
  OAI222_X1 U17869 ( .A1(n16766), .A2(n16667), .B1(n15954), .B2(n15953), .C1(
        n16659), .C2(n20402), .ZN(P1_U2889) );
  OAI222_X1 U17870 ( .A1(n21870), .A2(n20480), .B1(n15956), .B2(n20493), .C1(
        n20483), .C2(n15955), .ZN(P1_U2859) );
  AOI22_X1 U17871 ( .A1(n19156), .A2(n15957), .B1(n19158), .B2(
        P2_EBX_REG_0__SCAN_IN), .ZN(n15968) );
  INV_X1 U17872 ( .A(n19049), .ZN(n15958) );
  OAI21_X1 U17873 ( .B1(n19159), .B2(n15958), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15961) );
  INV_X1 U17874 ( .A(n15959), .ZN(n19019) );
  NAND2_X1 U17875 ( .A1(n17642), .A2(n19019), .ZN(n15960) );
  OAI211_X1 U17876 ( .C1(n19111), .C2(n13343), .A(n15961), .B(n15960), .ZN(
        n15962) );
  INV_X1 U17877 ( .A(n15962), .ZN(n15967) );
  NAND2_X1 U17878 ( .A1(n15963), .A2(n19131), .ZN(n15966) );
  OR2_X1 U17879 ( .A1(n19161), .A2(n15964), .ZN(n15965) );
  OAI21_X1 U17880 ( .B1(n19732), .B2(n16973), .A(n15969), .ZN(P2_U2855) );
  INV_X1 U17881 ( .A(n16766), .ZN(n22136) );
  INV_X1 U17882 ( .A(n20467), .ZN(n15972) );
  NAND2_X1 U17883 ( .A1(n16845), .A2(n15970), .ZN(n15971) );
  NAND2_X1 U17884 ( .A1(n15972), .A2(n15971), .ZN(n22134) );
  OAI22_X1 U17885 ( .A1(n22134), .A2(n20480), .B1(n15973), .B2(n20493), .ZN(
        n15974) );
  AOI21_X1 U17886 ( .B1(n22136), .B2(n20489), .A(n15974), .ZN(n15975) );
  INV_X1 U17887 ( .A(n15975), .ZN(P1_U2857) );
  INV_X1 U17888 ( .A(n15988), .ZN(n21364) );
  INV_X1 U17889 ( .A(n19455), .ZN(n15976) );
  NOR2_X1 U17890 ( .A1(n15976), .A2(n15992), .ZN(n15977) );
  NAND3_X1 U17891 ( .A1(n21364), .A2(n15977), .A3(n21363), .ZN(n21339) );
  NOR2_X1 U17892 ( .A1(n21366), .A2(n20684), .ZN(n21367) );
  INV_X1 U17893 ( .A(n15986), .ZN(n15980) );
  NOR2_X1 U17894 ( .A1(n21115), .A2(n20684), .ZN(n17681) );
  INV_X1 U17895 ( .A(n17681), .ZN(n15984) );
  NAND2_X1 U17896 ( .A1(n20684), .A2(n15983), .ZN(n21827) );
  NOR2_X2 U17897 ( .A1(n16001), .A2(n15983), .ZN(n21798) );
  AOI21_X1 U17898 ( .B1(n15984), .B2(n21827), .A(n21798), .ZN(n17680) );
  NOR2_X1 U17899 ( .A1(n21366), .A2(n17681), .ZN(n15998) );
  NAND2_X1 U17900 ( .A1(n21179), .A2(n21122), .ZN(n21120) );
  NOR2_X1 U17901 ( .A1(n21370), .A2(n19589), .ZN(n17682) );
  NAND2_X1 U17902 ( .A1(n21120), .A2(n17682), .ZN(n15997) );
  OAI211_X1 U17903 ( .C1(n21363), .C2(n15998), .A(n15997), .B(n15986), .ZN(
        n15987) );
  AOI221_X1 U17904 ( .B1(n21219), .B2(n15988), .C1(n21363), .C2(n15988), .A(
        n15987), .ZN(n15989) );
  OAI21_X1 U17905 ( .B1(n15990), .B2(n19455), .A(n15989), .ZN(n15991) );
  OAI21_X1 U17906 ( .B1(n21341), .B2(n21361), .A(n21802), .ZN(n17662) );
  NAND2_X1 U17907 ( .A1(n21327), .A2(n17662), .ZN(n21801) );
  INV_X1 U17908 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21836) );
  NAND2_X1 U17909 ( .A1(n21314), .A2(n21836), .ZN(n21308) );
  NOR2_X1 U17910 ( .A1(n21801), .A2(n21308), .ZN(n16010) );
  INV_X1 U17911 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n22250) );
  NOR2_X1 U17912 ( .A1(n22250), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n22252) );
  INV_X2 U17913 ( .A(n22252), .ZN(n22298) );
  INV_X1 U17914 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n22249) );
  NAND2_X1 U17915 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22249), .ZN(n22295) );
  NAND2_X1 U17916 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22252), .ZN(n18948) );
  INV_X1 U17917 ( .A(n18948), .ZN(n18949) );
  AOI21_X1 U17918 ( .B1(n22298), .B2(n22295), .A(n18949), .ZN(n21371) );
  AOI21_X1 U17919 ( .B1(n21371), .B2(n17680), .A(n21117), .ZN(n16009) );
  XOR2_X1 U17920 ( .A(n15994), .B(n15993), .Z(n15996) );
  NAND2_X1 U17921 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n22297) );
  NAND2_X1 U17922 ( .A1(n21793), .A2(n22297), .ZN(n16008) );
  INV_X1 U17923 ( .A(n15997), .ZN(n16004) );
  OAI211_X1 U17924 ( .C1(n21307), .C2(n21364), .A(n15999), .B(n15998), .ZN(
        n16000) );
  INV_X1 U17925 ( .A(n16000), .ZN(n16002) );
  AOI21_X1 U17926 ( .B1(n18395), .B2(n16002), .A(n16001), .ZN(n16003) );
  AOI211_X1 U17927 ( .C1(n16006), .C2(n16005), .A(n16004), .B(n16003), .ZN(
        n21378) );
  NAND2_X1 U17928 ( .A1(n21790), .A2(n18393), .ZN(n16007) );
  OAI211_X1 U17929 ( .C1(n16009), .C2(n16008), .A(n21378), .B(n16007), .ZN(
        n21803) );
  NOR2_X1 U17930 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21836), .ZN(n19253) );
  INV_X1 U17931 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21852) );
  INV_X1 U17932 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21841) );
  NAND2_X1 U17933 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18276) );
  NOR2_X1 U17934 ( .A1(n21841), .A2(n18276), .ZN(n17677) );
  INV_X1 U17935 ( .A(n17677), .ZN(n21834) );
  NOR2_X1 U17936 ( .A1(n21852), .A2(n21834), .ZN(n17664) );
  AOI211_X2 U17937 ( .C1(n21826), .C2(n21803), .A(n19253), .B(n17664), .ZN(
        n21362) );
  MUX2_X1 U17938 ( .A(n16010), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n21362), .Z(P3_U3284) );
  XOR2_X1 U17939 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n16011), .Z(n16014)
         );
  MUX2_X1 U17940 ( .A(n18972), .B(n16012), .S(n17044), .Z(n16013) );
  OAI21_X1 U17941 ( .B1(n16014), .B2(n17034), .A(n16013), .ZN(P2_U2882) );
  NAND2_X1 U17942 ( .A1(n15444), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n16016) );
  NAND2_X1 U17943 ( .A1(n17765), .A2(n17044), .ZN(n16015) );
  OAI211_X1 U17944 ( .C1(n19974), .C2(n17034), .A(n16016), .B(n16015), .ZN(
        P2_U2883) );
  INV_X1 U17945 ( .A(n17769), .ZN(n16020) );
  NOR2_X1 U17946 ( .A1(n19134), .A2(n16017), .ZN(n16019) );
  AOI21_X1 U17947 ( .B1(n16020), .B2(n16019), .A(n19201), .ZN(n16018) );
  OAI21_X1 U17948 ( .B1(n16020), .B2(n16019), .A(n16018), .ZN(n16028) );
  AOI22_X1 U17949 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19158), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19159), .ZN(n16021) );
  OAI211_X1 U17950 ( .C1(n19111), .C2(n17863), .A(n16021), .B(n19068), .ZN(
        n16022) );
  AOI21_X1 U17951 ( .B1(n19118), .B2(n16023), .A(n16022), .ZN(n16024) );
  OAI21_X1 U17952 ( .B1(n16025), .B2(n19144), .A(n16024), .ZN(n16026) );
  AOI21_X1 U17953 ( .B1(n17765), .B2(n19131), .A(n16026), .ZN(n16027) );
  OAI211_X1 U17954 ( .C1(n19974), .C2(n16973), .A(n16028), .B(n16027), .ZN(
        P2_U2851) );
  NAND2_X1 U17955 ( .A1(n16029), .A2(n14287), .ZN(n16031) );
  INV_X1 U17956 ( .A(n16031), .ZN(n16030) );
  NAND2_X1 U17957 ( .A1(n16030), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16131) );
  INV_X1 U17958 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16090) );
  NAND2_X1 U17959 ( .A1(n16031), .A2(n16090), .ZN(n16105) );
  NAND2_X1 U17960 ( .A1(n16131), .A2(n16105), .ZN(n16077) );
  NAND2_X1 U17961 ( .A1(n16033), .A2(n16032), .ZN(n16034) );
  NAND2_X1 U17962 ( .A1(n16049), .A2(n16034), .ZN(n19081) );
  INV_X1 U17963 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17428) );
  OAI21_X1 U17964 ( .B1(n19081), .B2(n16060), .A(n17428), .ZN(n17204) );
  NAND2_X1 U17965 ( .A1(n17295), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16036) );
  NAND2_X1 U17966 ( .A1(n16036), .A2(n16035), .ZN(n16037) );
  AND4_X1 U17967 ( .A1(n17204), .A2(n16039), .A3(n16038), .A4(n16037), .ZN(
        n16040) );
  INV_X1 U17968 ( .A(n19081), .ZN(n16043) );
  AND2_X1 U17969 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16042) );
  NAND2_X1 U17970 ( .A1(n16043), .A2(n16042), .ZN(n17203) );
  XNOR2_X1 U17971 ( .A(n16049), .B(n16048), .ZN(n19088) );
  NAND2_X1 U17972 ( .A1(n19088), .A2(n14287), .ZN(n17191) );
  NAND2_X1 U17973 ( .A1(n16051), .A2(n16050), .ZN(n16052) );
  AND2_X1 U17974 ( .A1(n16056), .A2(n16052), .ZN(n16053) );
  AOI21_X1 U17975 ( .B1(n16053), .B2(n14287), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17180) );
  INV_X1 U17976 ( .A(n16053), .ZN(n19107) );
  NAND2_X1 U17977 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16054) );
  XNOR2_X1 U17978 ( .A(n16056), .B(n16055), .ZN(n19116) );
  NAND2_X1 U17979 ( .A1(n19116), .A2(n14287), .ZN(n17169) );
  INV_X1 U17980 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16057) );
  XNOR2_X1 U17981 ( .A(n16059), .B(n16058), .ZN(n16061) );
  INV_X1 U17982 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17365) );
  OAI21_X1 U17983 ( .B1(n16061), .B2(n16060), .A(n17365), .ZN(n16063) );
  INV_X1 U17984 ( .A(n16061), .ZN(n19128) );
  AND2_X1 U17985 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16062) );
  NAND2_X1 U17986 ( .A1(n19128), .A2(n16062), .ZN(n16075) );
  INV_X1 U17987 ( .A(n16064), .ZN(n16065) );
  XNOR2_X1 U17988 ( .A(n16066), .B(n16065), .ZN(n16937) );
  NAND2_X1 U17989 ( .A1(n16937), .A2(n14287), .ZN(n16074) );
  INV_X1 U17990 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17377) );
  NAND2_X1 U17991 ( .A1(n16074), .A2(n17377), .ZN(n17163) );
  NAND2_X1 U17992 ( .A1(n16069), .A2(n16068), .ZN(n16070) );
  INV_X1 U17993 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17141) );
  INV_X1 U17994 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17345) );
  XNOR2_X1 U17995 ( .A(n16072), .B(n16071), .ZN(n19157) );
  INV_X1 U17996 ( .A(n17131), .ZN(n16073) );
  INV_X1 U17997 ( .A(n16075), .ZN(n16076) );
  INV_X1 U17998 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16080) );
  NAND2_X2 U17999 ( .A1(n17176), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17177) );
  NOR2_X1 U18000 ( .A1(n17365), .A2(n17377), .ZN(n17364) );
  INV_X1 U18001 ( .A(n17364), .ZN(n16082) );
  OR2_X1 U18002 ( .A1(n16082), .A2(n16057), .ZN(n16078) );
  INV_X1 U18003 ( .A(n17132), .ZN(n17140) );
  AOI21_X1 U18004 ( .B1(n17140), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16079) );
  NAND2_X1 U18005 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16112) );
  NOR2_X1 U18006 ( .A1(n16079), .A2(n16142), .ZN(n16102) );
  INV_X1 U18007 ( .A(n17413), .ZN(n17400) );
  INV_X1 U18008 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16081) );
  NOR2_X1 U18009 ( .A1(n16081), .A2(n16080), .ZN(n17389) );
  NAND3_X1 U18010 ( .A1(n17400), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n17389), .ZN(n17382) );
  NOR2_X1 U18011 ( .A1(n17382), .A2(n16082), .ZN(n16113) );
  NAND2_X1 U18012 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16113), .ZN(
        n17344) );
  XNOR2_X1 U18013 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16083) );
  NAND2_X1 U18014 ( .A1(n19047), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16096) );
  OAI21_X1 U18015 ( .B1(n17344), .B2(n16083), .A(n16096), .ZN(n16092) );
  INV_X1 U18016 ( .A(n16113), .ZN(n16160) );
  NOR2_X1 U18017 ( .A1(n16160), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17356) );
  NOR2_X1 U18018 ( .A1(n17579), .A2(n16084), .ZN(n17450) );
  OR2_X1 U18019 ( .A1(n16085), .A2(n17450), .ZN(n17561) );
  INV_X1 U18020 ( .A(n17422), .ZN(n16086) );
  NOR2_X1 U18021 ( .A1(n17581), .A2(n16086), .ZN(n16087) );
  NOR2_X1 U18022 ( .A1(n17561), .A2(n16087), .ZN(n17429) );
  AND2_X1 U18023 ( .A1(n17429), .A2(n17581), .ZN(n16088) );
  OR2_X1 U18024 ( .A1(n16088), .A2(n17364), .ZN(n16089) );
  INV_X1 U18025 ( .A(n17389), .ZN(n17399) );
  AOI21_X1 U18026 ( .B1(n17429), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16088), .ZN(n17416) );
  AOI211_X1 U18027 ( .C1(n19186), .C2(n17399), .A(n16057), .B(n17416), .ZN(
        n17391) );
  OR2_X1 U18028 ( .A1(n17391), .A2(n16088), .ZN(n17378) );
  NAND2_X1 U18029 ( .A1(n16089), .A2(n17378), .ZN(n17358) );
  NOR2_X1 U18030 ( .A1(n17356), .A2(n17358), .ZN(n17346) );
  NOR2_X1 U18031 ( .A1(n17346), .A2(n16090), .ZN(n16091) );
  AOI211_X1 U18032 ( .C1(n19189), .C2(n17053), .A(n16092), .B(n16091), .ZN(
        n16093) );
  OAI21_X1 U18033 ( .B1(n16980), .B2(n19184), .A(n16093), .ZN(n16094) );
  AOI21_X1 U18034 ( .B1(n16102), .B2(n17628), .A(n16094), .ZN(n16095) );
  OAI21_X1 U18035 ( .B1(n16104), .B2(n19182), .A(n16095), .ZN(P2_U3017) );
  OAI21_X1 U18036 ( .B1(n17762), .B2(n16097), .A(n16096), .ZN(n16098) );
  AOI21_X1 U18037 ( .B1(n17754), .B2(n16099), .A(n16098), .ZN(n16100) );
  OAI21_X1 U18038 ( .B1(n16980), .B2(n17773), .A(n16100), .ZN(n16101) );
  AOI21_X1 U18039 ( .B1(n16102), .B2(n17782), .A(n16101), .ZN(n16103) );
  OAI21_X1 U18040 ( .B1(n16104), .B2(n17774), .A(n16103), .ZN(P2_U2985) );
  NAND2_X1 U18041 ( .A1(n16106), .A2(n16105), .ZN(n16134) );
  NAND2_X1 U18042 ( .A1(n16134), .A2(n16131), .ZN(n16111) );
  AOI21_X1 U18043 ( .B1(n16108), .B2(n14287), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16133) );
  AND2_X1 U18044 ( .A1(n14287), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16107) );
  NAND2_X1 U18045 ( .A1(n16108), .A2(n16107), .ZN(n16132) );
  INV_X1 U18046 ( .A(n16132), .ZN(n16109) );
  NOR2_X1 U18047 ( .A1(n16133), .A2(n16109), .ZN(n16110) );
  XNOR2_X1 U18048 ( .A(n16111), .B(n16110), .ZN(n16130) );
  NAND2_X1 U18049 ( .A1(n16124), .A2(n17628), .ZN(n16123) );
  NOR2_X1 U18050 ( .A1(n16112), .A2(n17141), .ZN(n16116) );
  NAND2_X1 U18051 ( .A1(n16116), .A2(n16113), .ZN(n16114) );
  NOR2_X1 U18052 ( .A1(n16114), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16121) );
  NAND2_X1 U18053 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16116), .ZN(
        n16159) );
  AOI21_X1 U18054 ( .B1(n16159), .B2(n19186), .A(n17358), .ZN(n16156) );
  OR2_X1 U18055 ( .A1(n16156), .A2(n11430), .ZN(n16117) );
  NAND2_X1 U18056 ( .A1(n19047), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n16126) );
  NAND2_X1 U18057 ( .A1(n16119), .A2(n16118), .ZN(n16120) );
  OAI211_X1 U18058 ( .C1(n16130), .C2(n19182), .A(n16123), .B(n16122), .ZN(
        P2_U3016) );
  NAND2_X1 U18059 ( .A1(n16124), .A2(n17782), .ZN(n16129) );
  NAND2_X1 U18060 ( .A1(n17780), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16125) );
  OAI211_X1 U18061 ( .C1(n17790), .C2(n16913), .A(n16126), .B(n16125), .ZN(
        n16127) );
  AOI21_X1 U18062 ( .B1(n16414), .B2(n17784), .A(n16127), .ZN(n16128) );
  OAI211_X1 U18063 ( .C1(n16130), .C2(n17774), .A(n16129), .B(n16128), .ZN(
        P2_U2984) );
  OAI21_X2 U18064 ( .B1(n16134), .B2(n16133), .A(n11856), .ZN(n16141) );
  NOR2_X1 U18065 ( .A1(n16135), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n16138) );
  MUX2_X1 U18066 ( .A(n16138), .B(n16137), .S(n16136), .Z(n16918) );
  NAND2_X1 U18067 ( .A1(n16918), .A2(n14287), .ZN(n16139) );
  XNOR2_X1 U18068 ( .A(n16139), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16140) );
  XNOR2_X1 U18069 ( .A(n16141), .B(n16140), .ZN(n16176) );
  XNOR2_X1 U18070 ( .A(n16143), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16168) );
  AOI22_X1 U18071 ( .A1(n13164), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n16148) );
  NAND2_X1 U18072 ( .A1(n16146), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n16147) );
  OAI211_X1 U18073 ( .C1(n16149), .C2(n16155), .A(n16148), .B(n16147), .ZN(
        n16150) );
  NAND2_X1 U18074 ( .A1(n16169), .A2(n17633), .ZN(n16165) );
  AOI222_X1 U18075 ( .A1(n13394), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n13577), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n13595), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n16152) );
  INV_X1 U18076 ( .A(n16152), .ZN(n16153) );
  OR2_X1 U18077 ( .A1(n16156), .A2(n16155), .ZN(n16158) );
  INV_X1 U18078 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n17903) );
  NOR2_X1 U18079 ( .A1(n19068), .A2(n17903), .ZN(n16170) );
  INV_X1 U18080 ( .A(n16170), .ZN(n16157) );
  NAND2_X1 U18081 ( .A1(n16158), .A2(n16157), .ZN(n16162) );
  NOR3_X1 U18082 ( .A1(n16160), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16159), .ZN(n16161) );
  NAND2_X1 U18083 ( .A1(n16165), .A2(n16164), .ZN(n16166) );
  AOI21_X1 U18084 ( .B1(n16168), .B2(n17628), .A(n16166), .ZN(n16167) );
  OAI21_X1 U18085 ( .B1(n16176), .B2(n19182), .A(n16167), .ZN(P2_U3015) );
  NAND2_X1 U18086 ( .A1(n16168), .A2(n17782), .ZN(n16175) );
  AOI21_X1 U18087 ( .B1(n17780), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16170), .ZN(n16171) );
  OAI21_X1 U18088 ( .B1(n17790), .B2(n16172), .A(n16171), .ZN(n16173) );
  AOI21_X1 U18089 ( .B1(n16169), .B2(n17784), .A(n16173), .ZN(n16174) );
  OAI211_X1 U18090 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n16178), .A(n16177), 
        .B(n22441), .ZN(n16181) );
  NAND2_X1 U18091 ( .A1(n16179), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n16180) );
  OAI211_X1 U18092 ( .C1(n16182), .C2(n22430), .A(n16181), .B(n16180), .ZN(
        P1_U3477) );
  NAND2_X1 U18093 ( .A1(n20462), .A2(n22069), .ZN(n16189) );
  AOI22_X1 U18094 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n22030), .B1(n22034), 
        .B2(n22031), .ZN(n16183) );
  OAI21_X1 U18095 ( .B1(n22203), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n16183), .ZN(n16187) );
  INV_X1 U18096 ( .A(n16184), .ZN(n16185) );
  OAI22_X1 U18097 ( .A1(n22208), .A2(n16185), .B1(n22201), .B2(n11742), .ZN(
        n16186) );
  AOI211_X1 U18098 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n22206), .A(
        n16187), .B(n16186), .ZN(n16188) );
  OAI211_X1 U18099 ( .C1(n22050), .C2(n22430), .A(n16189), .B(n16188), .ZN(
        P1_U2839) );
  AOI22_X1 U18100 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16193) );
  AOI22_X1 U18101 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16192) );
  AOI22_X1 U18102 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16191) );
  AOI22_X1 U18103 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16190) );
  NAND4_X1 U18104 ( .A1(n16193), .A2(n16192), .A3(n16191), .A4(n16190), .ZN(
        n16200) );
  AOI22_X1 U18105 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16198) );
  AOI22_X1 U18106 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16234), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16197) );
  AOI22_X1 U18107 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16196) );
  AOI22_X1 U18108 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16195) );
  NAND4_X1 U18109 ( .A1(n16198), .A2(n16197), .A3(n16196), .A4(n16195), .ZN(
        n16199) );
  OR2_X1 U18110 ( .A1(n16200), .A2(n16199), .ZN(n17043) );
  AOI22_X1 U18111 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16205) );
  AOI22_X1 U18112 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16234), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16204) );
  AOI22_X1 U18113 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16203) );
  AOI22_X1 U18114 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16202) );
  NAND4_X1 U18115 ( .A1(n16205), .A2(n16204), .A3(n16203), .A4(n16202), .ZN(
        n16221) );
  INV_X1 U18116 ( .A(n13369), .ZN(n16209) );
  INV_X1 U18117 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16208) );
  INV_X1 U18118 ( .A(n16232), .ZN(n16207) );
  INV_X1 U18119 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16206) );
  OAI22_X1 U18120 ( .A1(n16209), .A2(n16208), .B1(n16207), .B2(n16206), .ZN(
        n16220) );
  INV_X1 U18121 ( .A(n16210), .ZN(n16215) );
  INV_X1 U18122 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16214) );
  INV_X1 U18123 ( .A(n16211), .ZN(n16213) );
  INV_X1 U18124 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16212) );
  OAI22_X1 U18125 ( .A1(n16215), .A2(n16214), .B1(n16213), .B2(n16212), .ZN(
        n16219) );
  AOI22_X1 U18126 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16217) );
  AOI22_X1 U18127 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16216) );
  NAND2_X1 U18128 ( .A1(n16217), .A2(n16216), .ZN(n16218) );
  NOR4_X1 U18129 ( .A1(n16221), .A2(n16220), .A3(n16219), .A4(n16218), .ZN(
        n17038) );
  AOI22_X1 U18130 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16225) );
  AOI22_X1 U18131 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16224) );
  AOI22_X1 U18132 ( .A1(n13344), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16223) );
  AOI22_X1 U18133 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16222) );
  NAND4_X1 U18134 ( .A1(n16225), .A2(n16224), .A3(n16223), .A4(n16222), .ZN(
        n16231) );
  AOI22_X1 U18135 ( .A1(n16194), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16239), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16229) );
  AOI22_X1 U18136 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16234), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16228) );
  AOI22_X1 U18137 ( .A1(n16241), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16242), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16227) );
  AOI22_X1 U18138 ( .A1(n16240), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16226) );
  NAND4_X1 U18139 ( .A1(n16229), .A2(n16228), .A3(n16227), .A4(n16226), .ZN(
        n16230) );
  OR2_X1 U18140 ( .A1(n16231), .A2(n16230), .ZN(n17028) );
  AOI22_X1 U18141 ( .A1(n16210), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16232), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16238) );
  AOI22_X1 U18142 ( .A1(n13369), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16211), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16237) );
  AOI22_X1 U18143 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11159), .B1(
        n13344), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16236) );
  AOI22_X1 U18144 ( .A1(n13446), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16235) );
  NAND4_X1 U18145 ( .A1(n16238), .A2(n16237), .A3(n16236), .A4(n16235), .ZN(
        n16248) );
  AOI22_X1 U18146 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n16239), .B1(
        n16194), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16246) );
  AOI22_X1 U18147 ( .A1(n13460), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13447), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16245) );
  AOI22_X1 U18148 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n16241), .B1(
        n16240), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16244) );
  AOI22_X1 U18149 ( .A1(n16242), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13368), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16243) );
  NAND4_X1 U18150 ( .A1(n16246), .A2(n16245), .A3(n16244), .A4(n16243), .ZN(
        n16247) );
  NOR2_X1 U18151 ( .A1(n16248), .A2(n16247), .ZN(n16266) );
  AOI22_X1 U18152 ( .A1(n13021), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11193), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16256) );
  AND2_X1 U18153 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16250) );
  OR2_X1 U18154 ( .A1(n16250), .A2(n16249), .ZN(n16396) );
  INV_X1 U18155 ( .A(n16396), .ZN(n16352) );
  NAND2_X1 U18156 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n16252) );
  NAND2_X1 U18157 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n16251) );
  AND3_X1 U18158 ( .A1(n16352), .A2(n16252), .A3(n16251), .ZN(n16255) );
  AOI22_X1 U18159 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16254) );
  AOI22_X1 U18160 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16253) );
  NAND4_X1 U18161 ( .A1(n16256), .A2(n16255), .A3(n16254), .A4(n16253), .ZN(
        n16265) );
  AOI22_X1 U18162 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16399), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16263) );
  AOI22_X1 U18163 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16262) );
  NAND2_X1 U18164 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n16258) );
  NAND2_X1 U18165 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n16257) );
  AND3_X1 U18166 ( .A1(n16258), .A2(n16396), .A3(n16257), .ZN(n16261) );
  AOI22_X1 U18167 ( .A1(n11194), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16260) );
  NAND4_X1 U18168 ( .A1(n16263), .A2(n16262), .A3(n16261), .A4(n16260), .ZN(
        n16264) );
  NAND2_X1 U18169 ( .A1(n16265), .A2(n16264), .ZN(n16267) );
  XNOR2_X1 U18170 ( .A(n16266), .B(n16267), .ZN(n17021) );
  INV_X1 U18171 ( .A(n16266), .ZN(n16269) );
  INV_X1 U18172 ( .A(n16267), .ZN(n16268) );
  NAND2_X1 U18173 ( .A1(n16269), .A2(n16268), .ZN(n16285) );
  AOI22_X1 U18174 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11196), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16275) );
  NAND2_X1 U18175 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n16271) );
  NAND2_X1 U18176 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n16270) );
  AND3_X1 U18177 ( .A1(n16352), .A2(n16271), .A3(n16270), .ZN(n16274) );
  AOI22_X1 U18178 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16273) );
  AOI22_X1 U18179 ( .A1(n13021), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16272) );
  NAND4_X1 U18180 ( .A1(n16275), .A2(n16274), .A3(n16273), .A4(n16272), .ZN(
        n16283) );
  AOI22_X1 U18181 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11195), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16281) );
  AOI22_X1 U18182 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16280) );
  NAND2_X1 U18183 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n16277) );
  NAND2_X1 U18184 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n16276) );
  AND3_X1 U18185 ( .A1(n16277), .A2(n16396), .A3(n16276), .ZN(n16279) );
  AOI22_X1 U18186 ( .A1(n13021), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16278) );
  NAND4_X1 U18187 ( .A1(n16281), .A2(n16280), .A3(n16279), .A4(n16278), .ZN(
        n16282) );
  NAND2_X1 U18188 ( .A1(n16283), .A2(n16282), .ZN(n16287) );
  INV_X1 U18189 ( .A(n16285), .ZN(n16284) );
  NAND2_X1 U18190 ( .A1(n16347), .A2(n16284), .ZN(n16286) );
  NOR2_X1 U18191 ( .A1(n16285), .A2(n16287), .ZN(n16309) );
  AOI22_X1 U18192 ( .A1(n16287), .A2(n16286), .B1(n16309), .B2(n11178), .ZN(
        n17014) );
  INV_X1 U18193 ( .A(n16309), .ZN(n16303) );
  AOI22_X1 U18194 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11193), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16294) );
  NAND2_X1 U18195 ( .A1(n16386), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n16289) );
  NAND2_X1 U18196 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n16288) );
  AND3_X1 U18197 ( .A1(n16352), .A2(n16289), .A3(n16288), .ZN(n16293) );
  AOI22_X1 U18198 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16292) );
  AOI22_X1 U18199 ( .A1(n13021), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16291) );
  NAND4_X1 U18200 ( .A1(n16294), .A2(n16293), .A3(n16292), .A4(n16291), .ZN(
        n16302) );
  AOI22_X1 U18201 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11193), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16300) );
  AOI22_X1 U18202 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16299) );
  NAND2_X1 U18203 ( .A1(n16386), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n16296) );
  NAND2_X1 U18204 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n16295) );
  AND3_X1 U18205 ( .A1(n16296), .A2(n16396), .A3(n16295), .ZN(n16298) );
  AOI22_X1 U18206 ( .A1(n13021), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16297) );
  NAND4_X1 U18207 ( .A1(n16300), .A2(n16299), .A3(n16298), .A4(n16297), .ZN(
        n16301) );
  AND2_X1 U18208 ( .A1(n16302), .A2(n16301), .ZN(n16308) );
  XNOR2_X1 U18209 ( .A(n16303), .B(n16308), .ZN(n16304) );
  NAND2_X1 U18210 ( .A1(n16304), .A2(n16347), .ZN(n16307) );
  INV_X1 U18211 ( .A(n16308), .ZN(n16306) );
  NOR2_X1 U18212 ( .A1(n11178), .A2(n16306), .ZN(n17009) );
  NAND2_X1 U18213 ( .A1(n17010), .A2(n17009), .ZN(n17008) );
  NAND2_X1 U18214 ( .A1(n16309), .A2(n16308), .ZN(n16325) );
  INV_X1 U18215 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20086) );
  AOI22_X1 U18216 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11193), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16315) );
  NAND2_X1 U18217 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n16311) );
  NAND2_X1 U18218 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n16310) );
  AND3_X1 U18219 ( .A1(n16352), .A2(n16311), .A3(n16310), .ZN(n16314) );
  AOI22_X1 U18220 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16313) );
  AOI22_X1 U18221 ( .A1(n13021), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16312) );
  NAND4_X1 U18222 ( .A1(n16315), .A2(n16314), .A3(n16313), .A4(n16312), .ZN(
        n16323) );
  AOI22_X1 U18223 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11190), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16321) );
  AOI22_X1 U18224 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16320) );
  NAND2_X1 U18225 ( .A1(n16386), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n16317) );
  NAND2_X1 U18226 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n16316) );
  AND3_X1 U18227 ( .A1(n16317), .A2(n16396), .A3(n16316), .ZN(n16319) );
  AOI22_X1 U18228 ( .A1(n13021), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16318) );
  NAND4_X1 U18229 ( .A1(n16321), .A2(n16320), .A3(n16319), .A4(n16318), .ZN(
        n16322) );
  NAND2_X1 U18230 ( .A1(n16323), .A2(n16322), .ZN(n16327) );
  AOI21_X1 U18231 ( .B1(n16325), .B2(n16327), .A(n16324), .ZN(n16326) );
  OR2_X1 U18232 ( .A1(n16325), .A2(n16327), .ZN(n16346) );
  INV_X1 U18233 ( .A(n16327), .ZN(n16328) );
  NAND2_X1 U18234 ( .A1(n13109), .A2(n16328), .ZN(n17003) );
  NOR2_X2 U18235 ( .A1(n17004), .A2(n17003), .ZN(n17002) );
  NOR2_X2 U18236 ( .A1(n17002), .A2(n16330), .ZN(n16366) );
  INV_X1 U18237 ( .A(n16346), .ZN(n16348) );
  AOI22_X1 U18238 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11190), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16336) );
  NAND2_X1 U18239 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n16332) );
  NAND2_X1 U18240 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n16331) );
  AND3_X1 U18241 ( .A1(n16352), .A2(n16332), .A3(n16331), .ZN(n16335) );
  AOI22_X1 U18242 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16334) );
  AOI22_X1 U18243 ( .A1(n16399), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16333) );
  NAND4_X1 U18244 ( .A1(n16336), .A2(n16335), .A3(n16334), .A4(n16333), .ZN(
        n16344) );
  AOI22_X1 U18245 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11189), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16342) );
  AOI22_X1 U18246 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16341) );
  NAND2_X1 U18247 ( .A1(n16386), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n16338) );
  NAND2_X1 U18248 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n16337) );
  AND3_X1 U18249 ( .A1(n16338), .A2(n16396), .A3(n16337), .ZN(n16340) );
  AOI22_X1 U18250 ( .A1(n16399), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16339) );
  NAND4_X1 U18251 ( .A1(n16342), .A2(n16341), .A3(n16340), .A4(n16339), .ZN(
        n16343) );
  NAND2_X1 U18252 ( .A1(n16344), .A2(n16343), .ZN(n16345) );
  INV_X1 U18253 ( .A(n16345), .ZN(n16349) );
  OR2_X1 U18254 ( .A1(n16346), .A2(n16345), .ZN(n16983) );
  OAI211_X1 U18255 ( .C1(n16348), .C2(n16349), .A(n16347), .B(n16983), .ZN(
        n16365) );
  AND2_X1 U18256 ( .A1(n13109), .A2(n16349), .ZN(n16994) );
  AOI22_X1 U18257 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11191), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16356) );
  NAND2_X1 U18258 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n16351) );
  NAND2_X1 U18259 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n16350) );
  AND3_X1 U18260 ( .A1(n16352), .A2(n16351), .A3(n16350), .ZN(n16355) );
  AOI22_X1 U18261 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16354) );
  AOI22_X1 U18262 ( .A1(n16399), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16353) );
  NAND4_X1 U18263 ( .A1(n16356), .A2(n16355), .A3(n16354), .A4(n16353), .ZN(
        n16364) );
  AOI22_X1 U18264 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11192), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16362) );
  AOI22_X1 U18265 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16361) );
  NAND2_X1 U18266 ( .A1(n16386), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n16358) );
  NAND2_X1 U18267 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n16357) );
  AND3_X1 U18268 ( .A1(n16358), .A2(n16396), .A3(n16357), .ZN(n16360) );
  AOI22_X1 U18269 ( .A1(n13021), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16359) );
  NAND4_X1 U18270 ( .A1(n16362), .A2(n16361), .A3(n16360), .A4(n16359), .ZN(
        n16363) );
  AND2_X1 U18271 ( .A1(n16364), .A2(n16363), .ZN(n16984) );
  INV_X1 U18272 ( .A(n16983), .ZN(n16367) );
  NAND3_X1 U18273 ( .A1(n16367), .A2(n16984), .A3(n11178), .ZN(n16977) );
  AOI22_X1 U18274 ( .A1(n11194), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16370) );
  NAND2_X1 U18275 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n16369) );
  NAND2_X1 U18276 ( .A1(n16376), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n16368) );
  NAND4_X1 U18277 ( .A1(n16370), .A2(n16396), .A3(n16369), .A4(n16368), .ZN(
        n16383) );
  AOI22_X1 U18278 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16399), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16372) );
  AOI22_X1 U18279 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16371) );
  NAND2_X1 U18280 ( .A1(n16372), .A2(n16371), .ZN(n16382) );
  INV_X1 U18281 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16373) );
  NOR2_X1 U18282 ( .A1(n16374), .A2(n16373), .ZN(n16375) );
  AOI211_X1 U18283 ( .C1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .C2(n16376), .A(
        n16396), .B(n16375), .ZN(n16380) );
  AOI22_X1 U18284 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16379) );
  AOI22_X1 U18285 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13321), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16378) );
  AOI22_X1 U18286 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11193), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16377) );
  NAND4_X1 U18287 ( .A1(n16380), .A2(n16379), .A3(n16378), .A4(n16377), .ZN(
        n16381) );
  OAI21_X1 U18288 ( .B1(n16383), .B2(n16382), .A(n16381), .ZN(n16976) );
  AOI22_X1 U18289 ( .A1(n16385), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16389) );
  NAND2_X1 U18290 ( .A1(n16386), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n16388) );
  NAND2_X1 U18291 ( .A1(n13321), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n16387) );
  NAND4_X1 U18292 ( .A1(n16389), .A2(n16388), .A3(n16387), .A4(n16396), .ZN(
        n16407) );
  AOI22_X1 U18293 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11195), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16392) );
  AOI22_X1 U18294 ( .A1(n16390), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16391) );
  NAND2_X1 U18295 ( .A1(n16392), .A2(n16391), .ZN(n16406) );
  NOR2_X1 U18296 ( .A1(n16394), .A2(n16393), .ZN(n16395) );
  AOI211_X1 U18297 ( .C1(n13321), .C2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n16396), .B(n16395), .ZN(n16404) );
  AOI22_X1 U18298 ( .A1(n16398), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16397), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16403) );
  AOI22_X1 U18299 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n16390), .B1(
        n16399), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16402) );
  AOI22_X1 U18300 ( .A1(n11196), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16384), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16401) );
  NAND4_X1 U18301 ( .A1(n16404), .A2(n16403), .A3(n16402), .A4(n16401), .ZN(
        n16405) );
  OAI21_X1 U18302 ( .B1(n16407), .B2(n16406), .A(n16405), .ZN(n16408) );
  XNOR2_X1 U18303 ( .A(n16409), .B(n16408), .ZN(n16417) );
  INV_X1 U18304 ( .A(n20225), .ZN(n17105) );
  AOI22_X1 U18305 ( .A1(n20223), .A2(n19693), .B1(n20221), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n16411) );
  NAND2_X1 U18306 ( .A1(n20224), .A2(BUF1_REG_30__SCAN_IN), .ZN(n16410) );
  OAI211_X1 U18307 ( .C1(n17105), .C2(n21231), .A(n16411), .B(n16410), .ZN(
        n16412) );
  AOI21_X1 U18308 ( .B1(n16115), .B2(n20169), .A(n16412), .ZN(n16413) );
  OAI21_X1 U18309 ( .B1(n16417), .B2(n20228), .A(n16413), .ZN(P2_U2889) );
  NAND2_X1 U18310 ( .A1(n15444), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n16416) );
  NAND2_X1 U18311 ( .A1(n16414), .A2(n17044), .ZN(n16415) );
  OAI211_X1 U18312 ( .C1(n16417), .C2(n17034), .A(n16416), .B(n16415), .ZN(
        P2_U2857) );
  OR2_X1 U18313 ( .A1(n16418), .A2(n16421), .ZN(n16427) );
  NAND2_X1 U18314 ( .A1(n22810), .A2(n16419), .ZN(n16426) );
  NAND2_X1 U18315 ( .A1(n16421), .A2(n16420), .ZN(n16425) );
  NAND2_X1 U18316 ( .A1(n16423), .A2(n16422), .ZN(n16424) );
  NAND4_X1 U18317 ( .A1(n16427), .A2(n16426), .A3(n16425), .A4(n16424), .ZN(
        n17734) );
  OR2_X1 U18318 ( .A1(n16428), .A2(n22261), .ZN(n16429) );
  NAND2_X1 U18319 ( .A1(n16429), .A2(n22253), .ZN(n21854) );
  AND2_X1 U18320 ( .A1(n16430), .A2(n21854), .ZN(n17735) );
  NOR2_X1 U18321 ( .A1(n17735), .A2(n22234), .ZN(n22218) );
  MUX2_X1 U18322 ( .A(P1_MORE_REG_SCAN_IN), .B(n17734), .S(n22218), .Z(
        P1_U3484) );
  INV_X1 U18323 ( .A(n16678), .ZN(n16599) );
  INV_X1 U18324 ( .A(n16434), .ZN(n16448) );
  OR2_X1 U18325 ( .A1(n16455), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16447) );
  NAND2_X1 U18326 ( .A1(n16451), .A2(n16435), .ZN(n16439) );
  INV_X1 U18327 ( .A(n16436), .ZN(n16437) );
  NAND2_X1 U18328 ( .A1(n16465), .A2(n16437), .ZN(n16438) );
  NAND2_X1 U18329 ( .A1(n16439), .A2(n16438), .ZN(n16442) );
  INV_X1 U18330 ( .A(n16440), .ZN(n16441) );
  INV_X1 U18331 ( .A(n16674), .ZN(n16443) );
  OAI22_X1 U18332 ( .A1(n16676), .A2(n22152), .B1(n22203), .B2(n16443), .ZN(
        n16444) );
  AOI21_X1 U18333 ( .B1(n22166), .B2(P1_EBX_REG_30__SCAN_IN), .A(n16444), .ZN(
        n16445) );
  OAI21_X1 U18334 ( .B1(n16815), .B2(n22208), .A(n16445), .ZN(n16446) );
  AOI21_X1 U18335 ( .B1(n16448), .B2(n16447), .A(n16446), .ZN(n16449) );
  OAI21_X1 U18336 ( .B1(n16599), .B2(n22209), .A(n16449), .ZN(P1_U2810) );
  OAI21_X1 U18337 ( .B1(n16465), .B2(n16452), .A(n16451), .ZN(n16560) );
  INV_X1 U18338 ( .A(n16560), .ZN(n16826) );
  AOI22_X1 U18339 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n22206), .B1(
        n22187), .B2(n16453), .ZN(n16454) );
  OAI21_X1 U18340 ( .B1(n22201), .B2(n16561), .A(n16454), .ZN(n16458) );
  AOI22_X1 U18341 ( .A1(n11375), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(n22200), .ZN(n16456) );
  AOI211_X1 U18342 ( .C1(n16826), .C2(n22165), .A(n16458), .B(n16457), .ZN(
        n16459) );
  OAI21_X1 U18343 ( .B1(n16450), .B2(n22209), .A(n16459), .ZN(P1_U2811) );
  INV_X1 U18344 ( .A(n16460), .ZN(n16461) );
  AOI21_X1 U18345 ( .B1(n16462), .B2(n16461), .A(n13649), .ZN(n16691) );
  NOR2_X1 U18346 ( .A1(n16482), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16471) );
  NOR2_X1 U18347 ( .A1(n16478), .A2(n16463), .ZN(n16464) );
  NAND3_X1 U18348 ( .A1(n16482), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n22200), 
        .ZN(n16469) );
  OAI22_X1 U18349 ( .A1(n16466), .A2(n22152), .B1(n22203), .B2(n16689), .ZN(
        n16467) );
  AOI21_X1 U18350 ( .B1(n22166), .B2(P1_EBX_REG_28__SCAN_IN), .A(n16467), .ZN(
        n16468) );
  OAI211_X1 U18351 ( .C1(n21984), .C2(n22208), .A(n16469), .B(n16468), .ZN(
        n16470) );
  AOI211_X1 U18352 ( .C1(n16691), .C2(n22172), .A(n16471), .B(n16470), .ZN(
        n16472) );
  INV_X1 U18353 ( .A(n16472), .ZN(P1_U2812) );
  AOI21_X1 U18354 ( .B1(n16474), .B2(n16486), .A(n16460), .ZN(n16700) );
  INV_X1 U18355 ( .A(n16700), .ZN(n16608) );
  INV_X1 U18356 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n16475) );
  OAI22_X1 U18357 ( .A1(n16509), .A2(n21976), .B1(n22189), .B2(n16475), .ZN(
        n16483) );
  NOR2_X1 U18358 ( .A1(n16488), .A2(n16476), .ZN(n16477) );
  OR2_X1 U18359 ( .A1(n16478), .A2(n16477), .ZN(n16829) );
  AOI22_X1 U18360 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n22206), .B1(
        n22187), .B2(n16696), .ZN(n16480) );
  NAND2_X1 U18361 ( .A1(n22166), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n16479) );
  OAI211_X1 U18362 ( .C1(n16829), .C2(n22208), .A(n16480), .B(n16479), .ZN(
        n16481) );
  AOI21_X1 U18363 ( .B1(n16483), .B2(n16482), .A(n16481), .ZN(n16484) );
  OAI21_X1 U18364 ( .B1(n16608), .B2(n22209), .A(n16484), .ZN(P1_U2813) );
  OAI21_X1 U18365 ( .B1(n16485), .B2(n16487), .A(n16486), .ZN(n16612) );
  INV_X1 U18366 ( .A(n16612), .ZN(n16706) );
  NOR2_X1 U18367 ( .A1(n16509), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n16497) );
  INV_X1 U18368 ( .A(n16488), .ZN(n16491) );
  NAND2_X1 U18369 ( .A1(n16505), .A2(n16489), .ZN(n16490) );
  NAND2_X1 U18370 ( .A1(n16491), .A2(n16490), .ZN(n21966) );
  NAND3_X1 U18371 ( .A1(n16509), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n22200), 
        .ZN(n16495) );
  OAI22_X1 U18372 ( .A1(n16492), .A2(n22152), .B1(n22203), .B2(n16704), .ZN(
        n16493) );
  AOI21_X1 U18373 ( .B1(n22166), .B2(P1_EBX_REG_26__SCAN_IN), .A(n16493), .ZN(
        n16494) );
  OAI211_X1 U18374 ( .C1(n21966), .C2(n22208), .A(n16495), .B(n16494), .ZN(
        n16496) );
  AOI211_X1 U18375 ( .C1(n16706), .C2(n22172), .A(n16497), .B(n16496), .ZN(
        n16498) );
  INV_X1 U18376 ( .A(n16498), .ZN(P1_U2814) );
  INV_X1 U18377 ( .A(n16485), .ZN(n16500) );
  OAI21_X1 U18378 ( .B1(n16501), .B2(n16499), .A(n16500), .ZN(n16712) );
  INV_X1 U18379 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20429) );
  INV_X1 U18380 ( .A(n22215), .ZN(n16502) );
  OAI21_X1 U18381 ( .B1(n22189), .B2(n20429), .A(n16502), .ZN(n16510) );
  NAND2_X1 U18382 ( .A1(n20479), .A2(n16503), .ZN(n16504) );
  NAND2_X1 U18383 ( .A1(n16505), .A2(n16504), .ZN(n21991) );
  AOI22_X1 U18384 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n22206), .B1(
        n22187), .B2(n16715), .ZN(n16507) );
  NAND2_X1 U18385 ( .A1(n22166), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n16506) );
  OAI211_X1 U18386 ( .C1(n21991), .C2(n22208), .A(n16507), .B(n16506), .ZN(
        n16508) );
  AOI21_X1 U18387 ( .B1(n16510), .B2(n16509), .A(n16508), .ZN(n16511) );
  OAI21_X1 U18388 ( .B1(n16712), .B2(n22209), .A(n16511), .ZN(P1_U2815) );
  INV_X1 U18389 ( .A(n16512), .ZN(n16514) );
  INV_X1 U18390 ( .A(n16513), .ZN(n16572) );
  AOI21_X1 U18391 ( .B1(n16514), .B2(n11203), .A(n16572), .ZN(n20547) );
  INV_X1 U18392 ( .A(n20547), .ZN(n16634) );
  INV_X1 U18393 ( .A(n16515), .ZN(n16517) );
  NOR3_X1 U18394 ( .A1(n22112), .A2(n16517), .A3(n16516), .ZN(n16536) );
  AOI211_X1 U18395 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(n16536), .A(n22189), 
        .B(n16526), .ZN(n16525) );
  INV_X1 U18396 ( .A(n16518), .ZN(n16520) );
  INV_X1 U18397 ( .A(n16575), .ZN(n16519) );
  AOI21_X1 U18398 ( .B1(n16520), .B2(n16519), .A(n16567), .ZN(n21937) );
  INV_X1 U18399 ( .A(n21937), .ZN(n16523) );
  OAI22_X1 U18400 ( .A1(n20550), .A2(n22203), .B1(n20475), .B2(n22201), .ZN(
        n16521) );
  AOI21_X1 U18401 ( .B1(n22206), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16521), .ZN(n16522) );
  OAI21_X1 U18402 ( .B1(n16523), .B2(n22208), .A(n16522), .ZN(n16524) );
  AOI211_X1 U18403 ( .C1(n16527), .C2(n16526), .A(n16525), .B(n16524), .ZN(
        n16528) );
  OAI21_X1 U18404 ( .B1(n16634), .B2(n22209), .A(n16528), .ZN(P1_U2818) );
  OR2_X1 U18405 ( .A1(n16529), .A2(n16546), .ZN(n16544) );
  AND2_X1 U18406 ( .A1(n16544), .A2(n16530), .ZN(n16532) );
  OR2_X1 U18407 ( .A1(n16532), .A2(n16531), .ZN(n20539) );
  OAI21_X1 U18408 ( .B1(n16535), .B2(n16534), .A(n16533), .ZN(n16542) );
  NOR2_X1 U18409 ( .A1(n22189), .A2(n16536), .ZN(n22177) );
  NAND2_X1 U18410 ( .A1(n11264), .A2(n16537), .ZN(n16538) );
  NAND2_X1 U18411 ( .A1(n11277), .A2(n16538), .ZN(n21924) );
  OAI22_X1 U18412 ( .A1(n20543), .A2(n22203), .B1(n20486), .B2(n22201), .ZN(
        n16539) );
  AOI21_X1 U18413 ( .B1(n22206), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16539), .ZN(n16540) );
  OAI21_X1 U18414 ( .B1(n21924), .B2(n22208), .A(n16540), .ZN(n16541) );
  AOI21_X1 U18415 ( .B1(n16542), .B2(n22177), .A(n16541), .ZN(n16543) );
  OAI21_X1 U18416 ( .B1(n20539), .B2(n22209), .A(n16543), .ZN(P1_U2820) );
  INV_X1 U18417 ( .A(n16544), .ZN(n16545) );
  AOI21_X1 U18418 ( .B1(n16546), .B2(n16529), .A(n16545), .ZN(n16736) );
  INV_X1 U18419 ( .A(n16736), .ZN(n16646) );
  NAND2_X1 U18420 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n22121), .ZN(n22140) );
  NOR2_X1 U18421 ( .A1(n22139), .A2(n22140), .ZN(n22141) );
  NAND2_X1 U18422 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n22141), .ZN(n22157) );
  INV_X1 U18423 ( .A(n22157), .ZN(n22150) );
  NAND2_X1 U18424 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n22150), .ZN(n22176) );
  AND2_X1 U18425 ( .A1(n22176), .A2(n22200), .ZN(n22171) );
  AOI221_X1 U18426 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), .C1(n16548), .C2(n16547), .A(n22176), .ZN(n16555) );
  OR2_X1 U18427 ( .A1(n16550), .A2(n16549), .ZN(n16551) );
  NAND2_X1 U18428 ( .A1(n11264), .A2(n16551), .ZN(n21936) );
  AOI21_X1 U18429 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n22206), .A(
        n22170), .ZN(n16553) );
  AOI22_X1 U18430 ( .A1(n16739), .A2(n22187), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n22166), .ZN(n16552) );
  OAI211_X1 U18431 ( .C1(n22208), .C2(n21936), .A(n16553), .B(n16552), .ZN(
        n16554) );
  AOI211_X1 U18432 ( .C1(n22171), .C2(P1_REIP_REG_19__SCAN_IN), .A(n16555), 
        .B(n16554), .ZN(n16556) );
  OAI21_X1 U18433 ( .B1(n16646), .B2(n22209), .A(n16556), .ZN(P1_U2821) );
  INV_X1 U18434 ( .A(n16804), .ZN(n16558) );
  OAI22_X1 U18435 ( .A1(n16558), .A2(n20480), .B1(n16557), .B2(n20493), .ZN(
        P1_U2841) );
  OAI222_X1 U18436 ( .A1(n16559), .A2(n20493), .B1(n20480), .B2(n16815), .C1(
        n20483), .C2(n16599), .ZN(P1_U2842) );
  OAI222_X1 U18437 ( .A1(n16561), .A2(n20493), .B1(n20480), .B2(n16560), .C1(
        n16450), .C2(n20483), .ZN(P1_U2843) );
  INV_X1 U18438 ( .A(n16691), .ZN(n16605) );
  OAI222_X1 U18439 ( .A1(n16562), .A2(n20493), .B1(n20483), .B2(n16605), .C1(
        n20480), .C2(n21984), .ZN(P1_U2844) );
  INV_X1 U18440 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n16563) );
  OAI222_X1 U18441 ( .A1(n16563), .A2(n20493), .B1(n20480), .B2(n16829), .C1(
        n16608), .C2(n20483), .ZN(P1_U2845) );
  OAI222_X1 U18442 ( .A1(n16564), .A2(n20493), .B1(n20480), .B2(n21966), .C1(
        n16612), .C2(n20483), .ZN(P1_U2846) );
  OAI222_X1 U18443 ( .A1(n16565), .A2(n20493), .B1(n20480), .B2(n21991), .C1(
        n16712), .C2(n20483), .ZN(P1_U2847) );
  OR2_X1 U18444 ( .A1(n16567), .A2(n16566), .ZN(n16568) );
  NAND2_X1 U18445 ( .A1(n20477), .A2(n16568), .ZN(n22192) );
  INV_X1 U18446 ( .A(n16569), .ZN(n16571) );
  INV_X1 U18447 ( .A(n16570), .ZN(n16617) );
  OAI21_X1 U18448 ( .B1(n16572), .B2(n16571), .A(n16617), .ZN(n22193) );
  OAI222_X1 U18449 ( .A1(n22192), .A2(n20480), .B1(n20493), .B2(n22198), .C1(
        n22193), .C2(n20483), .ZN(P1_U2849) );
  OAI21_X1 U18450 ( .B1(n16573), .B2(n16531), .A(n11203), .ZN(n22182) );
  AND2_X1 U18451 ( .A1(n11277), .A2(n16574), .ZN(n16576) );
  OR2_X1 U18452 ( .A1(n16576), .A2(n16575), .ZN(n22186) );
  OAI22_X1 U18453 ( .A1(n22186), .A2(n20480), .B1(n22180), .B2(n20493), .ZN(
        n16577) );
  INV_X1 U18454 ( .A(n16577), .ZN(n16578) );
  OAI21_X1 U18455 ( .B1(n22182), .B2(n20483), .A(n16578), .ZN(P1_U2851) );
  OAI222_X1 U18456 ( .A1(n21936), .A2(n20480), .B1(n20493), .B2(n16579), .C1(
        n16646), .C2(n20483), .ZN(P1_U2853) );
  NAND2_X1 U18457 ( .A1(n16580), .A2(n16581), .ZN(n16582) );
  NAND2_X1 U18458 ( .A1(n16583), .A2(n16582), .ZN(n22163) );
  NOR2_X1 U18459 ( .A1(n16585), .A2(n16586), .ZN(n16587) );
  OR2_X1 U18460 ( .A1(n16584), .A2(n16587), .ZN(n22156) );
  OAI222_X1 U18461 ( .A1(n22163), .A2(n20480), .B1(n20493), .B2(n22151), .C1(
        n22156), .C2(n20483), .ZN(P1_U2855) );
  NOR2_X1 U18462 ( .A1(n16588), .A2(n16591), .ZN(n16589) );
  NAND2_X1 U18463 ( .A1(n16659), .A2(n16589), .ZN(n16660) );
  AOI22_X1 U18464 ( .A1(n11350), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n16653), .ZN(n16593) );
  OAI211_X1 U18465 ( .C1(n15140), .C2(n16660), .A(n16594), .B(n16593), .ZN(
        P1_U2873) );
  INV_X1 U18466 ( .A(n16660), .ZN(n16654) );
  AOI22_X1 U18467 ( .A1(n16654), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n16653), .ZN(n16598) );
  NOR3_X4 U18468 ( .A1(n16653), .A2(n16596), .A3(n16595), .ZN(n16664) );
  AOI22_X1 U18469 ( .A1(n16664), .A2(n22397), .B1(n11350), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n16597) );
  OAI211_X1 U18470 ( .C1(n16599), .C2(n16667), .A(n16598), .B(n16597), .ZN(
        P1_U2874) );
  OAI22_X1 U18471 ( .A1(n16660), .A2(n13670), .B1(n22393), .B2(n16659), .ZN(
        n16600) );
  INV_X1 U18472 ( .A(n16600), .ZN(n16602) );
  AOI22_X1 U18473 ( .A1(n16664), .A2(n22390), .B1(n11350), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n16601) );
  OAI211_X1 U18474 ( .C1(n16450), .C2(n16667), .A(n16602), .B(n16601), .ZN(
        P1_U2875) );
  AOI22_X1 U18475 ( .A1(n16654), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n16653), .ZN(n16604) );
  AOI22_X1 U18476 ( .A1(n16664), .A2(n22382), .B1(n11350), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n16603) );
  OAI211_X1 U18477 ( .C1(n16605), .C2(n16667), .A(n16604), .B(n16603), .ZN(
        P1_U2876) );
  AOI22_X1 U18478 ( .A1(n16654), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n16653), .ZN(n16607) );
  AOI22_X1 U18479 ( .A1(n16664), .A2(n22375), .B1(n11350), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16606) );
  OAI211_X1 U18480 ( .C1(n16608), .C2(n16667), .A(n16607), .B(n16606), .ZN(
        P1_U2877) );
  OAI22_X1 U18481 ( .A1(n16660), .A2(n22556), .B1(n22371), .B2(n16659), .ZN(
        n16609) );
  INV_X1 U18482 ( .A(n16609), .ZN(n16611) );
  AOI22_X1 U18483 ( .A1(n16664), .A2(n22368), .B1(n11350), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n16610) );
  OAI211_X1 U18484 ( .C1(n16612), .C2(n16667), .A(n16611), .B(n16610), .ZN(
        P1_U2878) );
  AOI22_X1 U18485 ( .A1(n16654), .A2(DATAI_25_), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n16653), .ZN(n16615) );
  AOI22_X1 U18486 ( .A1(n16664), .A2(n16613), .B1(n11350), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n16614) );
  OAI211_X1 U18487 ( .C1(n16712), .C2(n16667), .A(n16615), .B(n16614), .ZN(
        P1_U2879) );
  AND2_X1 U18488 ( .A1(n16617), .A2(n16616), .ZN(n16618) );
  INV_X1 U18489 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n16619) );
  OAI22_X1 U18490 ( .A1(n16660), .A2(n22413), .B1(n16619), .B2(n16659), .ZN(
        n16620) );
  INV_X1 U18491 ( .A(n16620), .ZN(n16623) );
  AOI22_X1 U18492 ( .A1(n16664), .A2(n16621), .B1(n11350), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16622) );
  OAI211_X1 U18493 ( .C1(n22210), .C2(n16667), .A(n16623), .B(n16622), .ZN(
        P1_U2880) );
  OAI22_X1 U18494 ( .A1(n16660), .A2(n16624), .B1(n22354), .B2(n16659), .ZN(
        n16625) );
  INV_X1 U18495 ( .A(n16625), .ZN(n16628) );
  AOI22_X1 U18496 ( .A1(n16664), .A2(n16626), .B1(n11350), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16627) );
  OAI211_X1 U18497 ( .C1(n22193), .C2(n16667), .A(n16628), .B(n16627), .ZN(
        P1_U2881) );
  OAI22_X1 U18498 ( .A1(n16660), .A2(n16629), .B1(n22348), .B2(n16659), .ZN(
        n16630) );
  INV_X1 U18499 ( .A(n16630), .ZN(n16633) );
  AOI22_X1 U18500 ( .A1(n16664), .A2(n16631), .B1(n11350), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16632) );
  OAI211_X1 U18501 ( .C1(n16634), .C2(n16667), .A(n16633), .B(n16632), .ZN(
        P1_U2882) );
  AOI22_X1 U18502 ( .A1(n16654), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n16653), .ZN(n16637) );
  AOI22_X1 U18503 ( .A1(n16664), .A2(n16635), .B1(n11350), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n16636) );
  OAI211_X1 U18504 ( .C1(n22182), .C2(n16667), .A(n16637), .B(n16636), .ZN(
        P1_U2883) );
  OAI22_X1 U18505 ( .A1(n16660), .A2(n22633), .B1(n22336), .B2(n16659), .ZN(
        n16638) );
  INV_X1 U18506 ( .A(n16638), .ZN(n16640) );
  INV_X1 U18507 ( .A(n22334), .ZN(n22625) );
  AOI22_X1 U18508 ( .A1(n16664), .A2(n22625), .B1(n11350), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16639) );
  OAI211_X1 U18509 ( .C1(n20539), .C2(n16667), .A(n16640), .B(n16639), .ZN(
        P1_U2884) );
  OAI22_X1 U18510 ( .A1(n16660), .A2(n16641), .B1(n22330), .B2(n16659), .ZN(
        n16642) );
  INV_X1 U18511 ( .A(n16642), .ZN(n16645) );
  AOI22_X1 U18512 ( .A1(n16664), .A2(n16643), .B1(n11350), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n16644) );
  OAI211_X1 U18513 ( .C1(n16646), .C2(n16667), .A(n16645), .B(n16644), .ZN(
        P1_U2885) );
  OR2_X1 U18514 ( .A1(n16584), .A2(n16647), .ZN(n16648) );
  AND2_X1 U18515 ( .A1(n16529), .A2(n16648), .ZN(n22173) );
  INV_X1 U18516 ( .A(n22173), .ZN(n16652) );
  OAI22_X1 U18517 ( .A1(n16660), .A2(n22558), .B1(n22324), .B2(n16659), .ZN(
        n16649) );
  INV_X1 U18518 ( .A(n16649), .ZN(n16651) );
  AOI22_X1 U18519 ( .A1(n16664), .A2(n22555), .B1(n11350), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16650) );
  OAI211_X1 U18520 ( .C1(n16652), .C2(n16667), .A(n16651), .B(n16650), .ZN(
        P1_U2886) );
  AOI22_X1 U18521 ( .A1(n16654), .A2(DATAI_17_), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16653), .ZN(n16656) );
  AOI22_X1 U18522 ( .A1(n16664), .A2(n22315), .B1(n11350), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n16655) );
  OAI211_X1 U18523 ( .C1(n22156), .C2(n16667), .A(n16656), .B(n16655), .ZN(
        P1_U2887) );
  AOI21_X1 U18524 ( .B1(n16658), .B2(n16657), .A(n16585), .ZN(n22146) );
  INV_X1 U18525 ( .A(n22146), .ZN(n16668) );
  OAI22_X1 U18526 ( .A1(n16660), .A2(n22422), .B1(n22311), .B2(n16659), .ZN(
        n16661) );
  INV_X1 U18527 ( .A(n16661), .ZN(n16666) );
  INV_X1 U18528 ( .A(n22410), .ZN(n16663) );
  AOI22_X1 U18529 ( .A1(n16664), .A2(n16663), .B1(n11350), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n16665) );
  OAI211_X1 U18530 ( .C1(n16668), .C2(n16667), .A(n16666), .B(n16665), .ZN(
        P1_U2888) );
  NAND2_X1 U18531 ( .A1(n16669), .A2(n16823), .ZN(n16671) );
  NAND3_X1 U18532 ( .A1(n16672), .A2(n16671), .A3(n16670), .ZN(n16673) );
  INV_X1 U18533 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16809) );
  XNOR2_X1 U18534 ( .A(n16673), .B(n16809), .ZN(n16819) );
  NAND2_X1 U18535 ( .A1(n20520), .A2(n16674), .ZN(n16675) );
  NAND2_X1 U18536 ( .A1(n22170), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16806) );
  OAI211_X1 U18537 ( .C1(n16676), .C2(n20506), .A(n16675), .B(n16806), .ZN(
        n16677) );
  AOI21_X1 U18538 ( .B1(n16678), .B2(n20557), .A(n16677), .ZN(n16679) );
  OAI21_X1 U18539 ( .B1(n16819), .B2(n22216), .A(n16679), .ZN(P1_U2969) );
  NAND2_X1 U18540 ( .A1(n16680), .A2(n16681), .ZN(n16686) );
  NOR2_X1 U18541 ( .A1(n16682), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16683) );
  MUX2_X1 U18542 ( .A(n16683), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n20552), .Z(n16684) );
  NAND2_X1 U18543 ( .A1(n11861), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16717) );
  OAI211_X1 U18544 ( .C1(n16686), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16684), .B(n16717), .ZN(n16685) );
  AOI21_X1 U18545 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n16686), .A(
        n16685), .ZN(n16687) );
  XNOR2_X1 U18546 ( .A(n16687), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n21977) );
  NAND2_X1 U18547 ( .A1(n21999), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n21978) );
  NAND2_X1 U18548 ( .A1(n20551), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16688) );
  OAI211_X1 U18549 ( .C1(n20561), .C2(n16689), .A(n21978), .B(n16688), .ZN(
        n16690) );
  AOI21_X1 U18550 ( .B1(n16691), .B2(n20557), .A(n16690), .ZN(n16692) );
  OAI21_X1 U18551 ( .B1(n22216), .B2(n21977), .A(n16692), .ZN(P1_U2971) );
  NAND2_X1 U18552 ( .A1(n12929), .A2(n16693), .ZN(n16695) );
  XNOR2_X1 U18553 ( .A(n20552), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16694) );
  XNOR2_X1 U18554 ( .A(n16695), .B(n16694), .ZN(n16835) );
  NAND2_X1 U18555 ( .A1(n20520), .A2(n16696), .ZN(n16697) );
  NAND2_X1 U18556 ( .A1(n21999), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16830) );
  OAI211_X1 U18557 ( .C1(n20506), .C2(n16698), .A(n16697), .B(n16830), .ZN(
        n16699) );
  AOI21_X1 U18558 ( .B1(n16700), .B2(n20557), .A(n16699), .ZN(n16701) );
  OAI21_X1 U18559 ( .B1(n16835), .B2(n22216), .A(n16701), .ZN(P1_U2972) );
  OAI21_X1 U18560 ( .B1(n11789), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12929), .ZN(n21965) );
  AOI22_X1 U18561 ( .A1(n20551), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n21999), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n16703) );
  OAI21_X1 U18562 ( .B1(n20561), .B2(n16704), .A(n16703), .ZN(n16705) );
  AOI21_X1 U18563 ( .B1(n16706), .B2(n20557), .A(n16705), .ZN(n16707) );
  OAI21_X1 U18564 ( .B1(n22216), .B2(n21965), .A(n16707), .ZN(P1_U2973) );
  OAI21_X1 U18565 ( .B1(n16680), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n21969), .ZN(n16709) );
  NAND3_X1 U18566 ( .A1(n16709), .A2(n16708), .A3(n16717), .ZN(n16710) );
  XNOR2_X1 U18567 ( .A(n16710), .B(n21997), .ZN(n21990) );
  OAI22_X1 U18568 ( .A1(n20506), .A2(n16711), .B1(n21975), .B2(n20429), .ZN(
        n16714) );
  NOR2_X1 U18569 ( .A1(n16712), .A2(n20538), .ZN(n16713) );
  AOI211_X1 U18570 ( .C1(n20520), .C2(n16715), .A(n16714), .B(n16713), .ZN(
        n16716) );
  OAI21_X1 U18571 ( .B1(n22216), .B2(n21990), .A(n16716), .ZN(P1_U2974) );
  OAI21_X1 U18572 ( .B1(n11861), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16717), .ZN(n16718) );
  XOR2_X1 U18573 ( .A(n16718), .B(n16680), .Z(n22001) );
  OAI22_X1 U18574 ( .A1(n20506), .A2(n16719), .B1(n21975), .B2(n22191), .ZN(
        n16721) );
  NOR2_X1 U18575 ( .A1(n22193), .A2(n20538), .ZN(n16720) );
  AOI211_X1 U18576 ( .C1(n20520), .C2(n22188), .A(n16721), .B(n16720), .ZN(
        n16722) );
  OAI21_X1 U18577 ( .B1(n22001), .B2(n22216), .A(n16722), .ZN(P1_U2976) );
  INV_X1 U18578 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21932) );
  NAND3_X1 U18579 ( .A1(n16723), .A2(n14530), .A3(n21932), .ZN(n16727) );
  AND2_X1 U18580 ( .A1(n20552), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16724) );
  NAND2_X1 U18581 ( .A1(n16734), .A2(n16724), .ZN(n20534) );
  INV_X1 U18582 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16725) );
  NAND2_X1 U18583 ( .A1(n11861), .A2(n16725), .ZN(n16726) );
  AOI22_X1 U18584 ( .A1(n16727), .A2(n21944), .B1(n20534), .B2(n16726), .ZN(
        n16728) );
  XNOR2_X1 U18585 ( .A(n16728), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21952) );
  INV_X1 U18586 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n16729) );
  OAI22_X1 U18587 ( .A1(n20506), .A2(n16730), .B1(n16729), .B2(n21975), .ZN(
        n16732) );
  NOR2_X1 U18588 ( .A1(n22182), .A2(n20538), .ZN(n16731) );
  AOI211_X1 U18589 ( .C1(n20520), .C2(n22178), .A(n16732), .B(n16731), .ZN(
        n16733) );
  OAI21_X1 U18590 ( .B1(n22216), .B2(n21952), .A(n16733), .ZN(P1_U2978) );
  OR3_X1 U18591 ( .A1(n16734), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n20552), .ZN(n20533) );
  NAND2_X1 U18592 ( .A1(n20534), .A2(n20533), .ZN(n16735) );
  XNOR2_X1 U18593 ( .A(n16735), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21931) );
  NAND2_X1 U18594 ( .A1(n16736), .A2(n20557), .ZN(n16741) );
  OAI22_X1 U18595 ( .A1(n20506), .A2(n16737), .B1(n16548), .B2(n21975), .ZN(
        n16738) );
  AOI21_X1 U18596 ( .B1(n20520), .B2(n16739), .A(n16738), .ZN(n16740) );
  OAI211_X1 U18597 ( .C1(n21931), .C2(n22216), .A(n16741), .B(n16740), .ZN(
        P1_U2980) );
  NAND2_X1 U18598 ( .A1(n20551), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16742) );
  OAI211_X1 U18599 ( .C1(n20561), .C2(n22168), .A(n16743), .B(n16742), .ZN(
        n16744) );
  AOI21_X1 U18600 ( .B1(n22173), .B2(n20557), .A(n16744), .ZN(n16745) );
  OAI21_X1 U18601 ( .B1(n22216), .B2(n16746), .A(n16745), .ZN(P1_U2981) );
  NOR2_X1 U18602 ( .A1(n11861), .A2(n21911), .ZN(n20528) );
  NAND2_X1 U18603 ( .A1(n20528), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16751) );
  INV_X1 U18604 ( .A(n16747), .ZN(n16838) );
  NAND2_X1 U18605 ( .A1(n16748), .A2(n16838), .ZN(n16760) );
  AOI21_X1 U18606 ( .B1(n11861), .B2(n16749), .A(n16760), .ZN(n16750) );
  MUX2_X1 U18607 ( .A(n16751), .B(n20526), .S(n16750), .Z(n16753) );
  XNOR2_X1 U18608 ( .A(n16753), .B(n16752), .ZN(n21899) );
  NAND2_X1 U18609 ( .A1(n22170), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n21898) );
  OAI21_X1 U18610 ( .B1(n20506), .B2(n22153), .A(n21898), .ZN(n16755) );
  NOR2_X1 U18611 ( .A1(n22156), .A2(n20538), .ZN(n16754) );
  AOI211_X1 U18612 ( .C1(n20520), .C2(n22155), .A(n16755), .B(n16754), .ZN(
        n16756) );
  OAI21_X1 U18613 ( .B1(n21899), .B2(n22216), .A(n16756), .ZN(P1_U2982) );
  AOI21_X1 U18614 ( .B1(n16758), .B2(n16757), .A(n20552), .ZN(n16759) );
  NOR2_X1 U18615 ( .A1(n16760), .A2(n16759), .ZN(n20525) );
  XNOR2_X1 U18616 ( .A(n20552), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16761) );
  XNOR2_X1 U18617 ( .A(n20525), .B(n16761), .ZN(n21896) );
  NAND2_X1 U18618 ( .A1(n21896), .A2(n20556), .ZN(n16765) );
  OAI22_X1 U18619 ( .A1(n20506), .A2(n16762), .B1(n21975), .B2(n22139), .ZN(
        n16763) );
  AOI21_X1 U18620 ( .B1(n20520), .B2(n22131), .A(n16763), .ZN(n16764) );
  OAI211_X1 U18621 ( .C1(n20538), .C2(n16766), .A(n16765), .B(n16764), .ZN(
        P1_U2984) );
  INV_X1 U18622 ( .A(n16768), .ZN(n16769) );
  AOI21_X1 U18623 ( .B1(n16767), .B2(n16770), .A(n16769), .ZN(n20517) );
  AND2_X1 U18624 ( .A1(n16771), .A2(n16772), .ZN(n20516) );
  NAND2_X1 U18625 ( .A1(n20517), .A2(n20516), .ZN(n20515) );
  NAND2_X1 U18626 ( .A1(n20515), .A2(n16772), .ZN(n16774) );
  XNOR2_X1 U18627 ( .A(n16774), .B(n16773), .ZN(n21867) );
  INV_X1 U18628 ( .A(n21867), .ZN(n16780) );
  AOI22_X1 U18629 ( .A1(n20551), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n21999), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n16775) );
  OAI21_X1 U18630 ( .B1(n20561), .B2(n16776), .A(n16775), .ZN(n16777) );
  AOI21_X1 U18631 ( .B1(n16778), .B2(n20557), .A(n16777), .ZN(n16779) );
  OAI21_X1 U18632 ( .B1(n16780), .B2(n22216), .A(n16779), .ZN(P1_U2986) );
  NAND2_X1 U18633 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21946), .ZN(
        n16784) );
  NAND2_X1 U18634 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16781), .ZN(
        n21916) );
  INV_X1 U18635 ( .A(n21916), .ZN(n16783) );
  NAND2_X1 U18636 ( .A1(n16783), .A2(n16782), .ZN(n21917) );
  NOR2_X1 U18637 ( .A1(n16784), .A2(n21917), .ZN(n16789) );
  NOR2_X1 U18638 ( .A1(n21916), .A2(n16785), .ZN(n21921) );
  NAND3_X1 U18639 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21946), .A3(
        n21921), .ZN(n16792) );
  NOR2_X1 U18640 ( .A1(n16792), .A2(n16786), .ZN(n21959) );
  AOI21_X1 U18641 ( .B1(n16789), .B2(n21918), .A(n21959), .ZN(n21970) );
  NOR2_X1 U18642 ( .A1(n21970), .A2(n16787), .ZN(n21972) );
  NAND2_X1 U18643 ( .A1(n21972), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n21980) );
  NOR3_X1 U18644 ( .A1(n21980), .A2(n16808), .A3(n16823), .ZN(n16814) );
  NAND3_X1 U18645 ( .A1(n16814), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16894), .ZN(n16802) );
  AOI21_X1 U18646 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16789), .A(
        n16788), .ZN(n16790) );
  AOI211_X1 U18647 ( .C1(n16793), .C2(n16792), .A(n16791), .B(n16790), .ZN(
        n16794) );
  INV_X1 U18648 ( .A(n16794), .ZN(n22000) );
  AOI21_X1 U18649 ( .B1(n21969), .B2(n16798), .A(n22000), .ZN(n21998) );
  NAND2_X1 U18650 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21998), .ZN(
        n21971) );
  INV_X1 U18651 ( .A(n21971), .ZN(n16795) );
  NAND2_X1 U18652 ( .A1(n16795), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16796) );
  INV_X1 U18653 ( .A(n21940), .ZN(n16807) );
  AND2_X1 U18654 ( .A1(n16796), .A2(n16807), .ZN(n21986) );
  INV_X1 U18655 ( .A(n21986), .ZN(n16797) );
  NAND2_X1 U18656 ( .A1(n16797), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16813) );
  NAND2_X1 U18657 ( .A1(n16798), .A2(n16823), .ZN(n16810) );
  NAND2_X1 U18658 ( .A1(n16810), .A2(n12927), .ZN(n16799) );
  OAI211_X1 U18659 ( .C1(n16813), .C2(n16799), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16807), .ZN(n16800) );
  NAND3_X1 U18660 ( .A1(n16802), .A2(n16801), .A3(n16800), .ZN(n16803) );
  AOI21_X1 U18661 ( .B1(n16804), .B2(n21993), .A(n16803), .ZN(n16805) );
  INV_X1 U18662 ( .A(n16806), .ZN(n16812) );
  AOI21_X1 U18663 ( .B1(n16808), .B2(n16807), .A(n21986), .ZN(n16824) );
  AOI21_X1 U18664 ( .B1(n16824), .B2(n16810), .A(n16809), .ZN(n16811) );
  AOI211_X1 U18665 ( .C1(n16814), .C2(n16813), .A(n16812), .B(n16811), .ZN(
        n16818) );
  INV_X1 U18666 ( .A(n16815), .ZN(n16816) );
  NAND2_X1 U18667 ( .A1(n16816), .A2(n21993), .ZN(n16817) );
  OAI211_X1 U18668 ( .C1(n16819), .C2(n22010), .A(n16818), .B(n16817), .ZN(
        P1_U3001) );
  INV_X1 U18669 ( .A(n21980), .ZN(n16820) );
  NAND3_X1 U18670 ( .A1(n16820), .A2(n12927), .A3(n16823), .ZN(n16821) );
  OAI211_X1 U18671 ( .C1(n16824), .C2(n16823), .A(n16822), .B(n16821), .ZN(
        n16825) );
  AOI21_X1 U18672 ( .B1(n16826), .B2(n21993), .A(n16825), .ZN(n16827) );
  OAI21_X1 U18673 ( .B1(n16828), .B2(n22010), .A(n16827), .ZN(P1_U3002) );
  INV_X1 U18674 ( .A(n16829), .ZN(n16833) );
  NAND2_X1 U18675 ( .A1(n21986), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16831) );
  OAI211_X1 U18676 ( .C1(n21980), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16831), .B(n16830), .ZN(n16832) );
  AOI21_X1 U18677 ( .B1(n16833), .B2(n21993), .A(n16832), .ZN(n16834) );
  OAI21_X1 U18678 ( .B1(n16835), .B2(n22010), .A(n16834), .ZN(P1_U3004) );
  AOI21_X1 U18679 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n11861), .A(
        n16836), .ZN(n16842) );
  INV_X1 U18680 ( .A(n16767), .ZN(n16839) );
  AOI21_X1 U18681 ( .B1(n16839), .B2(n16838), .A(n16837), .ZN(n16840) );
  AOI21_X1 U18682 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n11861), .A(
        n16840), .ZN(n16841) );
  XOR2_X1 U18683 ( .A(n16842), .B(n16841), .Z(n20523) );
  OR4_X1 U18684 ( .A1(n16757), .A2(n16844), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n16843), .ZN(n16864) );
  INV_X1 U18685 ( .A(n16845), .ZN(n16846) );
  AOI21_X1 U18686 ( .B1(n16848), .B2(n16847), .A(n16846), .ZN(n22125) );
  NOR2_X1 U18687 ( .A1(n21975), .A2(n16849), .ZN(n16862) );
  INV_X1 U18688 ( .A(n16850), .ZN(n16855) );
  AOI21_X1 U18689 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16852), .A(
        n16851), .ZN(n16853) );
  AOI211_X1 U18690 ( .C1(n21918), .C2(n16855), .A(n16854), .B(n16853), .ZN(
        n16856) );
  OAI21_X1 U18691 ( .B1(n16858), .B2(n16857), .A(n16856), .ZN(n21865) );
  INV_X1 U18692 ( .A(n21865), .ZN(n16860) );
  AOI221_X1 U18693 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16860), 
        .C1(n16859), .C2(n16860), .A(n16758), .ZN(n16861) );
  AOI211_X1 U18694 ( .C1(n21993), .C2(n22125), .A(n16862), .B(n16861), .ZN(
        n16863) );
  OAI211_X1 U18695 ( .C1(n20523), .C2(n22010), .A(n16864), .B(n16863), .ZN(
        P1_U3017) );
  NOR2_X1 U18696 ( .A1(n16873), .A2(n16767), .ZN(n16865) );
  MUX2_X1 U18697 ( .A(n16873), .B(n16865), .S(n11861), .Z(n16866) );
  NAND3_X1 U18698 ( .A1(n16868), .A2(n16867), .A3(n21888), .ZN(n16871) );
  OAI21_X1 U18699 ( .B1(n16878), .B2(n21890), .A(n16876), .ZN(n21886) );
  NOR2_X1 U18700 ( .A1(n21975), .A2(n22114), .ZN(n20514) );
  NOR2_X1 U18701 ( .A1(n22009), .A2(n22101), .ZN(n16869) );
  AOI211_X1 U18702 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n21886), .A(
        n20514), .B(n16869), .ZN(n16870) );
  OAI211_X1 U18703 ( .C1(n20513), .C2(n22010), .A(n16871), .B(n16870), .ZN(
        P1_U3020) );
  INV_X1 U18704 ( .A(n16872), .ZN(n16875) );
  INV_X1 U18705 ( .A(n16873), .ZN(n16874) );
  OAI21_X1 U18706 ( .B1(n16875), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16874), .ZN(n20512) );
  OAI21_X1 U18707 ( .B1(n16878), .B2(n16877), .A(n16876), .ZN(n21881) );
  NAND4_X1 U18708 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n21888), .ZN(n21878) );
  AOI221_X1 U18709 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n11503), .C2(n16879), .A(
        n21878), .ZN(n16880) );
  AOI21_X1 U18710 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n21881), .A(
        n16880), .ZN(n16885) );
  OAI22_X1 U18711 ( .A1(n16882), .A2(n22009), .B1(n21975), .B2(n16881), .ZN(
        n16883) );
  INV_X1 U18712 ( .A(n16883), .ZN(n16884) );
  OAI211_X1 U18713 ( .C1(n20512), .C2(n22010), .A(n16885), .B(n16884), .ZN(
        P1_U3021) );
  INV_X1 U18714 ( .A(n16896), .ZN(n16886) );
  NAND3_X1 U18715 ( .A1(n16888), .A2(n16887), .A3(n16886), .ZN(n16889) );
  OAI21_X1 U18716 ( .B1(n16890), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n16889), .ZN(n16891) );
  AOI21_X1 U18717 ( .B1(n22500), .B2(n16892), .A(n16891), .ZN(n17721) );
  OAI22_X1 U18718 ( .A1(n16894), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16893), .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16902) );
  INV_X1 U18719 ( .A(n16902), .ZN(n16898) );
  NOR2_X1 U18720 ( .A1(n17744), .A2(n16895), .ZN(n16903) );
  INV_X1 U18721 ( .A(n22228), .ZN(n16909) );
  NOR3_X1 U18722 ( .A1(n16896), .A2(n15076), .A3(n16909), .ZN(n16897) );
  AOI21_X1 U18723 ( .B1(n16898), .B2(n16903), .A(n16897), .ZN(n16899) );
  OAI21_X1 U18724 ( .B1(n17721), .B2(n17669), .A(n16899), .ZN(n16900) );
  MUX2_X1 U18725 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16900), .S(
        n17674), .Z(P1_U3473) );
  INV_X1 U18726 ( .A(n16901), .ZN(n16904) );
  AOI22_X1 U18727 ( .A1(n16904), .A2(n22228), .B1(n16903), .B2(n16902), .ZN(
        n16905) );
  OAI21_X1 U18728 ( .B1(n16906), .B2(n17669), .A(n16905), .ZN(n16907) );
  MUX2_X1 U18729 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16907), .S(
        n17674), .Z(P1_U3472) );
  INV_X1 U18730 ( .A(n16908), .ZN(n16911) );
  OAI22_X1 U18731 ( .A1(n16911), .A2(n17669), .B1(n16910), .B2(n16909), .ZN(
        n16912) );
  MUX2_X1 U18732 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16912), .S(
        n17674), .Z(P1_U3469) );
  NAND3_X1 U18733 ( .A1(n16914), .A2(n16913), .A3(n19019), .ZN(n16922) );
  NOR2_X1 U18734 ( .A1(n16915), .A2(n16975), .ZN(n16917) );
  OAI22_X1 U18735 ( .A1(n12959), .A2(n19037), .B1(n17903), .B2(n19111), .ZN(
        n16916) );
  AOI211_X1 U18736 ( .C1(n19687), .C2(n19118), .A(n16917), .B(n16916), .ZN(
        n16921) );
  NAND2_X1 U18737 ( .A1(n16918), .A2(n19156), .ZN(n16920) );
  NAND2_X1 U18738 ( .A1(n16169), .A2(n19131), .ZN(n16919) );
  NAND4_X1 U18739 ( .A1(n16922), .A2(n16921), .A3(n16920), .A4(n16919), .ZN(
        P2_U2824) );
  NAND2_X1 U18740 ( .A1(n16924), .A2(n16925), .ZN(n16926) );
  NAND2_X1 U18741 ( .A1(n16923), .A2(n16926), .ZN(n17375) );
  NOR2_X1 U18742 ( .A1(n17090), .A2(n16928), .ZN(n16929) );
  OR2_X1 U18743 ( .A1(n16927), .A2(n16929), .ZN(n17086) );
  INV_X1 U18744 ( .A(n17086), .ZN(n17380) );
  AOI22_X1 U18745 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19159), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19155), .ZN(n16930) );
  OAI21_X1 U18746 ( .B1(n19108), .B2(n16931), .A(n16930), .ZN(n16932) );
  AOI21_X1 U18747 ( .B1(n17380), .B2(n19118), .A(n16932), .ZN(n16933) );
  OAI21_X1 U18748 ( .B1(n17375), .B2(n19163), .A(n16933), .ZN(n16936) );
  AOI211_X1 U18749 ( .C1(n16934), .C2(n17161), .A(n19201), .B(n19137), .ZN(
        n16935) );
  AOI211_X1 U18750 ( .C1(n19156), .C2(n16937), .A(n16936), .B(n16935), .ZN(
        n16938) );
  INV_X1 U18751 ( .A(n16938), .ZN(P2_U2830) );
  AOI211_X1 U18752 ( .C1(n16941), .C2(n16940), .A(n16939), .B(n19201), .ZN(
        n16942) );
  INV_X1 U18753 ( .A(n16942), .ZN(n16947) );
  AOI22_X1 U18754 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19159), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19155), .ZN(n16944) );
  NAND2_X1 U18755 ( .A1(n19158), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n16943) );
  OAI211_X1 U18756 ( .C1(n20022), .C2(n19161), .A(n16944), .B(n16943), .ZN(
        n16945) );
  AOI21_X1 U18757 ( .B1(n17045), .B2(n19131), .A(n16945), .ZN(n16946) );
  OAI211_X1 U18758 ( .C1(n19144), .C2(n16948), .A(n16947), .B(n16946), .ZN(
        P2_U2835) );
  NOR2_X1 U18759 ( .A1(n19201), .A2(n16949), .ZN(n19056) );
  INV_X1 U18760 ( .A(n16950), .ZN(n16956) );
  NOR2_X1 U18761 ( .A1(n19108), .A2(n13635), .ZN(n16953) );
  AOI22_X1 U18762 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19159), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19155), .ZN(n16951) );
  OAI211_X1 U18763 ( .C1(n19161), .C2(n20121), .A(n16951), .B(n19068), .ZN(
        n16952) );
  AOI211_X1 U18764 ( .C1(n16954), .C2(n19131), .A(n16953), .B(n16952), .ZN(
        n16955) );
  OAI21_X1 U18765 ( .B1(n16956), .B2(n19144), .A(n16955), .ZN(n16959) );
  INV_X1 U18766 ( .A(n16949), .ZN(n16957) );
  NOR3_X1 U18767 ( .A1(n16957), .A2(n19201), .A3(n16960), .ZN(n16958) );
  AOI211_X1 U18768 ( .C1(n19056), .C2(n16960), .A(n16959), .B(n16958), .ZN(
        n16961) );
  INV_X1 U18769 ( .A(n16961), .ZN(P2_U2837) );
  AOI211_X1 U18770 ( .C1(n17642), .C2(n16963), .A(n19134), .B(n16962), .ZN(
        n17649) );
  NAND2_X1 U18771 ( .A1(n17649), .A2(n19167), .ZN(n16972) );
  AOI22_X1 U18772 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19159), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19155), .ZN(n16964) );
  OAI21_X1 U18773 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19049), .A(
        n16964), .ZN(n16967) );
  NOR2_X1 U18774 ( .A1(n19144), .A2(n16965), .ZN(n16966) );
  AOI211_X1 U18775 ( .C1(n19118), .C2(n20168), .A(n16967), .B(n16966), .ZN(
        n16968) );
  OAI21_X1 U18776 ( .B1(n19108), .B2(n16969), .A(n16968), .ZN(n16970) );
  AOI21_X1 U18777 ( .B1(n17634), .B2(n19131), .A(n16970), .ZN(n16971) );
  OAI211_X1 U18778 ( .C1(n17799), .C2(n16973), .A(n16972), .B(n16971), .ZN(
        P2_U2854) );
  NAND2_X1 U18779 ( .A1(n16169), .A2(n17044), .ZN(n16974) );
  OAI21_X1 U18780 ( .B1(n17044), .B2(n16975), .A(n16974), .ZN(P2_U2856) );
  XNOR2_X1 U18781 ( .A(n16977), .B(n16976), .ZN(n16978) );
  XNOR2_X1 U18782 ( .A(n16979), .B(n16978), .ZN(n17055) );
  NOR2_X1 U18783 ( .A1(n16980), .A2(n15444), .ZN(n16981) );
  AOI21_X1 U18784 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n15444), .A(n16981), .ZN(
        n16982) );
  OAI21_X1 U18785 ( .B1(n17055), .B2(n17034), .A(n16982), .ZN(P2_U2858) );
  NAND2_X1 U18786 ( .A1(n11225), .A2(n16983), .ZN(n16985) );
  XNOR2_X1 U18787 ( .A(n16985), .B(n16984), .ZN(n17063) );
  OR2_X1 U18788 ( .A1(n16986), .A2(n16987), .ZN(n16988) );
  NAND2_X1 U18789 ( .A1(n16989), .A2(n16988), .ZN(n19164) );
  NOR2_X1 U18790 ( .A1(n19164), .A2(n15444), .ZN(n16990) );
  AOI21_X1 U18791 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15444), .A(n16990), .ZN(
        n16991) );
  OAI21_X1 U18792 ( .B1(n17063), .B2(n17034), .A(n16991), .ZN(P2_U2859) );
  NAND2_X1 U18793 ( .A1(n11225), .A2(n16992), .ZN(n16993) );
  XOR2_X1 U18794 ( .A(n16994), .B(n16993), .Z(n17073) );
  NOR2_X1 U18795 ( .A1(n16995), .A2(n16996), .ZN(n16997) );
  NOR2_X1 U18796 ( .A1(n19150), .A2(n15444), .ZN(n16998) );
  AOI21_X1 U18797 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15444), .A(n16998), .ZN(
        n16999) );
  OAI21_X1 U18798 ( .B1(n17073), .B2(n17034), .A(n16999), .ZN(P2_U2860) );
  AND2_X1 U18799 ( .A1(n16923), .A2(n17000), .ZN(n17001) );
  NOR2_X1 U18800 ( .A1(n16995), .A2(n17001), .ZN(n19132) );
  INV_X1 U18801 ( .A(n19132), .ZN(n17007) );
  AOI21_X1 U18802 ( .B1(n17004), .B2(n17003), .A(n17002), .ZN(n17074) );
  NAND2_X1 U18803 ( .A1(n17074), .A2(n17039), .ZN(n17006) );
  NAND2_X1 U18804 ( .A1(n15444), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n17005) );
  OAI211_X1 U18805 ( .C1(n17007), .C2(n15444), .A(n17006), .B(n17005), .ZN(
        P2_U2861) );
  OAI21_X1 U18806 ( .B1(n17010), .B2(n17009), .A(n17008), .ZN(n17089) );
  NAND2_X1 U18807 ( .A1(n15444), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n17012) );
  OR2_X1 U18808 ( .A1(n17375), .A2(n15444), .ZN(n17011) );
  OAI211_X1 U18809 ( .C1(n17089), .C2(n17034), .A(n17012), .B(n17011), .ZN(
        P2_U2862) );
  OAI21_X1 U18810 ( .B1(n17015), .B2(n17014), .A(n17013), .ZN(n17098) );
  OR2_X1 U18811 ( .A1(n17016), .A2(n17017), .ZN(n17018) );
  NAND2_X1 U18812 ( .A1(n16924), .A2(n17018), .ZN(n19117) );
  NOR2_X1 U18813 ( .A1(n19117), .A2(n15444), .ZN(n17019) );
  AOI21_X1 U18814 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15444), .A(n17019), .ZN(
        n17020) );
  OAI21_X1 U18815 ( .B1(n17098), .B2(n17034), .A(n17020), .ZN(P2_U2863) );
  XNOR2_X1 U18816 ( .A(n17027), .B(n17021), .ZN(n17110) );
  NOR2_X1 U18817 ( .A1(n17030), .A2(n17022), .ZN(n17023) );
  OR2_X1 U18818 ( .A1(n17016), .A2(n17023), .ZN(n19100) );
  NOR2_X1 U18819 ( .A1(n19100), .A2(n15444), .ZN(n17024) );
  AOI21_X1 U18820 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n15444), .A(n17024), .ZN(
        n17025) );
  OAI21_X1 U18821 ( .B1(n17110), .B2(n17034), .A(n17025), .ZN(P2_U2864) );
  OAI21_X1 U18822 ( .B1(n17026), .B2(n17028), .A(n17027), .ZN(n19923) );
  AND2_X1 U18823 ( .A1(n11223), .A2(n17029), .ZN(n17031) );
  OR2_X1 U18824 ( .A1(n17031), .A2(n17030), .ZN(n19089) );
  NOR2_X1 U18825 ( .A1(n19089), .A2(n15444), .ZN(n17032) );
  AOI21_X1 U18826 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n15444), .A(n17032), .ZN(
        n17033) );
  OAI21_X1 U18827 ( .B1(n19923), .B2(n17034), .A(n17033), .ZN(P2_U2865) );
  NAND2_X1 U18828 ( .A1(n17036), .A2(n17035), .ZN(n17037) );
  NAND2_X1 U18829 ( .A1(n11223), .A2(n17037), .ZN(n19076) );
  AOI21_X1 U18830 ( .B1(n17038), .B2(n17042), .A(n17026), .ZN(n17116) );
  NAND2_X1 U18831 ( .A1(n17116), .A2(n17039), .ZN(n17041) );
  NAND2_X1 U18832 ( .A1(n15444), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n17040) );
  OAI211_X1 U18833 ( .C1(n19076), .C2(n15444), .A(n17041), .B(n17040), .ZN(
        P2_U2866) );
  OAI21_X1 U18834 ( .B1(n16201), .B2(n17043), .A(n17042), .ZN(n20021) );
  NAND2_X1 U18835 ( .A1(n15444), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n17047) );
  NAND2_X1 U18836 ( .A1(n17045), .A2(n17044), .ZN(n17046) );
  OAI211_X1 U18837 ( .C1(n20021), .C2(n17034), .A(n17047), .B(n17046), .ZN(
        P2_U2867) );
  INV_X1 U18838 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n17051) );
  OAI22_X1 U18839 ( .A1(n17123), .A2(n19696), .B1(n17048), .B2(n19929), .ZN(
        n17049) );
  AOI21_X1 U18840 ( .B1(n20224), .B2(BUF1_REG_29__SCAN_IN), .A(n17049), .ZN(
        n17050) );
  OAI21_X1 U18841 ( .B1(n17105), .B2(n17051), .A(n17050), .ZN(n17052) );
  AOI21_X1 U18842 ( .B1(n17053), .B2(n20169), .A(n17052), .ZN(n17054) );
  OAI21_X1 U18843 ( .B1(n17055), .B2(n20228), .A(n17054), .ZN(P2_U2890) );
  INV_X1 U18844 ( .A(n19699), .ZN(n17056) );
  OAI22_X1 U18845 ( .A1(n17123), .A2(n17056), .B1(n14925), .B2(n19929), .ZN(
        n17057) );
  AOI21_X1 U18846 ( .B1(n20224), .B2(BUF1_REG_28__SCAN_IN), .A(n17057), .ZN(
        n17062) );
  NAND2_X1 U18847 ( .A1(n17067), .A2(n17058), .ZN(n17059) );
  AOI22_X1 U18848 ( .A1(n19160), .A2(n20169), .B1(n20225), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n17061) );
  OAI211_X1 U18849 ( .C1(n17063), .C2(n20228), .A(n17062), .B(n17061), .ZN(
        P2_U2891) );
  NAND2_X1 U18850 ( .A1(n17064), .A2(n17065), .ZN(n17066) );
  NAND2_X1 U18851 ( .A1(n17067), .A2(n17066), .ZN(n19154) );
  INV_X1 U18852 ( .A(n20169), .ZN(n20227) );
  AOI22_X1 U18853 ( .A1(n20223), .A2(n17068), .B1(n20221), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U18854 ( .A1(n20225), .A2(BUF2_REG_27__SCAN_IN), .B1(n20224), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n17069) );
  OAI211_X1 U18855 ( .C1(n19154), .C2(n20227), .A(n17070), .B(n17069), .ZN(
        n17071) );
  INV_X1 U18856 ( .A(n17071), .ZN(n17072) );
  OAI21_X1 U18857 ( .B1(n17073), .B2(n20228), .A(n17072), .ZN(P2_U2892) );
  INV_X1 U18858 ( .A(n17074), .ZN(n17082) );
  INV_X1 U18859 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17076) );
  INV_X1 U18860 ( .A(n20224), .ZN(n17103) );
  INV_X1 U18861 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n17075) );
  OAI22_X1 U18862 ( .A1(n17105), .A2(n17076), .B1(n17103), .B2(n17075), .ZN(
        n17080) );
  OR2_X1 U18863 ( .A1(n16927), .A2(n17077), .ZN(n17078) );
  NAND2_X1 U18864 ( .A1(n17064), .A2(n17078), .ZN(n19129) );
  OAI22_X1 U18865 ( .A1(n19129), .A2(n20227), .B1(n14923), .B2(n19929), .ZN(
        n17079) );
  AOI211_X1 U18866 ( .C1(n20223), .C2(n19705), .A(n17080), .B(n17079), .ZN(
        n17081) );
  OAI21_X1 U18867 ( .B1(n17082), .B2(n20228), .A(n17081), .ZN(P2_U2893) );
  AOI22_X1 U18868 ( .A1(n20223), .A2(n17083), .B1(n20221), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U18869 ( .A1(n20225), .A2(BUF2_REG_25__SCAN_IN), .B1(n20224), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n17084) );
  OAI211_X1 U18870 ( .C1(n17086), .C2(n20227), .A(n17085), .B(n17084), .ZN(
        n17087) );
  INV_X1 U18871 ( .A(n17087), .ZN(n17088) );
  OAI21_X1 U18872 ( .B1(n17089), .B2(n20228), .A(n17088), .ZN(P2_U2894) );
  INV_X1 U18873 ( .A(n19712), .ZN(n17095) );
  AOI21_X1 U18874 ( .B1(n17091), .B2(n17101), .A(n17090), .ZN(n19119) );
  INV_X1 U18875 ( .A(n19119), .ZN(n17093) );
  OAI22_X1 U18876 ( .A1(n17093), .A2(n20227), .B1(n17092), .B2(n19929), .ZN(
        n17094) );
  AOI21_X1 U18877 ( .B1(n20223), .B2(n17095), .A(n17094), .ZN(n17097) );
  AOI22_X1 U18878 ( .A1(n20225), .A2(BUF2_REG_24__SCAN_IN), .B1(n20224), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n17096) );
  OAI211_X1 U18879 ( .C1(n17098), .C2(n20228), .A(n17097), .B(n17096), .ZN(
        P2_U2895) );
  INV_X1 U18880 ( .A(n19721), .ZN(n17108) );
  NAND2_X1 U18881 ( .A1(n17409), .A2(n17099), .ZN(n17100) );
  NAND2_X1 U18882 ( .A1(n17101), .A2(n17100), .ZN(n19101) );
  OAI22_X1 U18883 ( .A1(n19101), .A2(n20227), .B1(n17102), .B2(n19929), .ZN(
        n17107) );
  INV_X1 U18884 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n17104) );
  OAI22_X1 U18885 ( .A1(n17105), .A2(n17104), .B1(n17103), .B2(n20610), .ZN(
        n17106) );
  AOI211_X1 U18886 ( .C1(n20223), .C2(n17108), .A(n17107), .B(n17106), .ZN(
        n17109) );
  OAI21_X1 U18887 ( .B1(n17110), .B2(n20228), .A(n17109), .ZN(P2_U2896) );
  AOI22_X1 U18888 ( .A1(n20225), .A2(BUF2_REG_21__SCAN_IN), .B1(n20224), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n17114) );
  NOR2_X1 U18889 ( .A1(n11267), .A2(n17111), .ZN(n17112) );
  OR2_X1 U18890 ( .A1(n17411), .A2(n17112), .ZN(n19075) );
  INV_X1 U18891 ( .A(n19075), .ZN(n17425) );
  AOI22_X1 U18892 ( .A1(n17425), .A2(n20169), .B1(n20221), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n17113) );
  OAI211_X1 U18893 ( .C1(n19980), .C2(n17123), .A(n17114), .B(n17113), .ZN(
        n17115) );
  AOI21_X1 U18894 ( .B1(n17116), .B2(n20123), .A(n17115), .ZN(n17117) );
  INV_X1 U18895 ( .A(n17117), .ZN(P2_U2898) );
  AOI22_X1 U18896 ( .A1(n20225), .A2(BUF2_REG_19__SCAN_IN), .B1(n20224), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n17122) );
  NAND2_X1 U18897 ( .A1(n14392), .A2(n17118), .ZN(n17119) );
  NAND2_X1 U18898 ( .A1(n17120), .A2(n17119), .ZN(n17439) );
  INV_X1 U18899 ( .A(n17439), .ZN(n19062) );
  AOI22_X1 U18900 ( .A1(n20169), .A2(n19062), .B1(n20221), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n17121) );
  OAI211_X1 U18901 ( .C1(n20077), .C2(n17123), .A(n17122), .B(n17121), .ZN(
        n17124) );
  AOI21_X1 U18902 ( .B1(n17125), .B2(n20123), .A(n17124), .ZN(n17126) );
  INV_X1 U18903 ( .A(n17126), .ZN(P2_U2900) );
  XNOR2_X1 U18904 ( .A(n17132), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17351) );
  NOR2_X1 U18905 ( .A1(n19164), .A2(n17773), .ZN(n17135) );
  NAND2_X1 U18906 ( .A1(n19047), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n17343) );
  NAND2_X1 U18907 ( .A1(n17780), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17133) );
  OAI211_X1 U18908 ( .C1(n17790), .C2(n19169), .A(n17343), .B(n17133), .ZN(
        n17134) );
  AOI211_X1 U18909 ( .C1(n17351), .C2(n17782), .A(n17135), .B(n17134), .ZN(
        n17136) );
  OAI21_X1 U18910 ( .B1(n17353), .B2(n17774), .A(n17136), .ZN(P2_U2986) );
  NAND2_X1 U18911 ( .A1(n11241), .A2(n17137), .ZN(n17138) );
  XNOR2_X1 U18912 ( .A(n17138), .B(n17141), .ZN(n17363) );
  INV_X1 U18913 ( .A(n17139), .ZN(n17146) );
  AOI21_X1 U18914 ( .B1(n17141), .B2(n17146), .A(n17140), .ZN(n17361) );
  NOR2_X1 U18915 ( .A1(n19068), .A2(n17895), .ZN(n17354) );
  NOR2_X1 U18916 ( .A1(n17790), .A2(n19148), .ZN(n17142) );
  AOI211_X1 U18917 ( .C1(n17780), .C2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17354), .B(n17142), .ZN(n17143) );
  OAI21_X1 U18918 ( .B1(n19150), .B2(n17773), .A(n17143), .ZN(n17144) );
  AOI21_X1 U18919 ( .B1(n17361), .B2(n17782), .A(n17144), .ZN(n17145) );
  OAI21_X1 U18920 ( .B1(n17774), .B2(n17363), .A(n17145), .ZN(P2_U2987) );
  NOR2_X1 U18921 ( .A1(n17177), .A2(n16057), .ZN(n17171) );
  NAND2_X1 U18922 ( .A1(n17171), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17157) );
  INV_X1 U18923 ( .A(n17157), .ZN(n17147) );
  OAI21_X1 U18924 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17147), .A(
        n17146), .ZN(n17374) );
  NOR2_X1 U18925 ( .A1(n19068), .A2(n17892), .ZN(n17366) );
  AOI21_X1 U18926 ( .B1(n17780), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17366), .ZN(n17148) );
  OAI21_X1 U18927 ( .B1(n17790), .B2(n19133), .A(n17148), .ZN(n17149) );
  AOI21_X1 U18928 ( .B1(n19132), .B2(n17784), .A(n17149), .ZN(n17156) );
  OAI21_X1 U18929 ( .B1(n17150), .B2(n17162), .A(n17163), .ZN(n17152) );
  INV_X1 U18930 ( .A(n17127), .ZN(n17153) );
  NAND2_X1 U18931 ( .A1(n17371), .A2(n17785), .ZN(n17155) );
  OAI211_X1 U18932 ( .C1(n17374), .C2(n17770), .A(n17156), .B(n17155), .ZN(
        P2_U2988) );
  OAI21_X1 U18933 ( .B1(n17171), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17157), .ZN(n17388) );
  NAND2_X1 U18934 ( .A1(n19047), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n17376) );
  OAI21_X1 U18935 ( .B1(n17762), .B2(n17158), .A(n17376), .ZN(n17160) );
  NOR2_X1 U18936 ( .A1(n17375), .A2(n17773), .ZN(n17159) );
  AOI211_X1 U18937 ( .C1(n17754), .C2(n17161), .A(n17160), .B(n17159), .ZN(
        n17167) );
  INV_X1 U18938 ( .A(n17162), .ZN(n17164) );
  NAND2_X1 U18939 ( .A1(n17164), .A2(n17163), .ZN(n17165) );
  XNOR2_X1 U18940 ( .A(n17150), .B(n17165), .ZN(n17385) );
  NAND2_X1 U18941 ( .A1(n17385), .A2(n17785), .ZN(n17166) );
  OAI211_X1 U18942 ( .C1(n17388), .C2(n17770), .A(n17167), .B(n17166), .ZN(
        P2_U2989) );
  XNOR2_X1 U18943 ( .A(n17169), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17170) );
  XNOR2_X1 U18944 ( .A(n17168), .B(n17170), .ZN(n17398) );
  AOI21_X1 U18945 ( .B1(n16057), .B2(n17177), .A(n17171), .ZN(n17396) );
  NOR2_X1 U18946 ( .A1(n19068), .A2(n17888), .ZN(n17393) );
  NOR2_X1 U18947 ( .A1(n17790), .A2(n19121), .ZN(n17172) );
  AOI211_X1 U18948 ( .C1(n17780), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n17393), .B(n17172), .ZN(n17173) );
  OAI21_X1 U18949 ( .B1(n19117), .B2(n17773), .A(n17173), .ZN(n17174) );
  AOI21_X1 U18950 ( .B1(n17396), .B2(n17782), .A(n17174), .ZN(n17175) );
  OAI21_X1 U18951 ( .B1(n17398), .B2(n17774), .A(n17175), .ZN(P2_U2990) );
  OAI21_X1 U18952 ( .B1(n17176), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17177), .ZN(n17408) );
  INV_X1 U18953 ( .A(n17178), .ZN(n17179) );
  NOR2_X1 U18954 ( .A1(n17180), .A2(n17179), .ZN(n17181) );
  XNOR2_X1 U18955 ( .A(n17182), .B(n17181), .ZN(n17406) );
  NAND2_X1 U18956 ( .A1(n19047), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n17401) );
  OAI21_X1 U18957 ( .B1(n17762), .B2(n17183), .A(n17401), .ZN(n17184) );
  AOI21_X1 U18958 ( .B1(n17754), .B2(n19106), .A(n17184), .ZN(n17185) );
  OAI21_X1 U18959 ( .B1(n19100), .B2(n17773), .A(n17185), .ZN(n17186) );
  AOI21_X1 U18960 ( .B1(n17406), .B2(n17785), .A(n17186), .ZN(n17187) );
  OAI21_X1 U18961 ( .B1(n17408), .B2(n17770), .A(n17187), .ZN(P2_U2991) );
  INV_X1 U18962 ( .A(n17188), .ZN(n17190) );
  INV_X1 U18963 ( .A(n17176), .ZN(n17189) );
  OAI21_X1 U18964 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17190), .A(
        n17189), .ZN(n17421) );
  XOR2_X1 U18965 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17191), .Z(
        n17192) );
  XNOR2_X1 U18966 ( .A(n17193), .B(n17192), .ZN(n17419) );
  NAND2_X1 U18967 ( .A1(n19047), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n17412) );
  OAI21_X1 U18968 ( .B1(n17762), .B2(n17194), .A(n17412), .ZN(n17195) );
  AOI21_X1 U18969 ( .B1(n17754), .B2(n19094), .A(n17195), .ZN(n17196) );
  OAI21_X1 U18970 ( .B1(n19089), .B2(n17773), .A(n17196), .ZN(n17197) );
  AOI21_X1 U18971 ( .B1(n17419), .B2(n17785), .A(n17197), .ZN(n17198) );
  OAI21_X1 U18972 ( .B1(n17421), .B2(n17770), .A(n17198), .ZN(P2_U2992) );
  OAI21_X1 U18973 ( .B1(n17199), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n17188), .ZN(n17435) );
  NAND2_X1 U18974 ( .A1(n19047), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n17423) );
  OAI21_X1 U18975 ( .B1(n17762), .B2(n17200), .A(n17423), .ZN(n17202) );
  NOR2_X1 U18976 ( .A1(n19076), .A2(n17773), .ZN(n17201) );
  AOI211_X1 U18977 ( .C1(n17754), .C2(n19080), .A(n17202), .B(n17201), .ZN(
        n17211) );
  NAND2_X1 U18978 ( .A1(n17204), .A2(n17203), .ZN(n17209) );
  AOI22_X1 U18979 ( .A1(n17207), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n11477), .B2(n17206), .ZN(n17208) );
  XOR2_X1 U18980 ( .A(n17209), .B(n17208), .Z(n17432) );
  NAND2_X1 U18981 ( .A1(n17432), .A2(n17785), .ZN(n17210) );
  OAI211_X1 U18982 ( .C1(n17435), .C2(n17770), .A(n17211), .B(n17210), .ZN(
        P2_U2993) );
  XNOR2_X1 U18983 ( .A(n17212), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17447) );
  INV_X1 U18984 ( .A(n17213), .ZN(n17214) );
  AOI21_X1 U18985 ( .B1(n17216), .B2(n17215), .A(n17214), .ZN(n17220) );
  NAND2_X1 U18986 ( .A1(n17218), .A2(n17217), .ZN(n17219) );
  XNOR2_X1 U18987 ( .A(n17220), .B(n17219), .ZN(n17445) );
  NAND2_X1 U18988 ( .A1(n19047), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n17437) );
  OAI21_X1 U18989 ( .B1(n17762), .B2(n17221), .A(n17437), .ZN(n17222) );
  AOI21_X1 U18990 ( .B1(n17754), .B2(n19066), .A(n17222), .ZN(n17223) );
  OAI21_X1 U18991 ( .B1(n17436), .B2(n17773), .A(n17223), .ZN(n17224) );
  AOI21_X1 U18992 ( .B1(n17445), .B2(n17785), .A(n17224), .ZN(n17225) );
  OAI21_X1 U18993 ( .B1(n17447), .B2(n17770), .A(n17225), .ZN(P2_U2995) );
  AND2_X1 U18994 ( .A1(n17227), .A2(n17226), .ZN(n17244) );
  NAND2_X1 U18995 ( .A1(n17244), .A2(n17243), .ZN(n17245) );
  NAND2_X1 U18996 ( .A1(n17245), .A2(n17228), .ZN(n17232) );
  NAND2_X1 U18997 ( .A1(n17230), .A2(n17229), .ZN(n17231) );
  XNOR2_X1 U18998 ( .A(n17232), .B(n17231), .ZN(n17457) );
  INV_X1 U18999 ( .A(n17457), .ZN(n17238) );
  OAI211_X1 U19000 ( .C1(n11359), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n17782), .B(n17233), .ZN(n17237) );
  NAND2_X1 U19001 ( .A1(n19040), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n17454) );
  NAND2_X1 U19002 ( .A1(n17780), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17234) );
  OAI211_X1 U19003 ( .C1(n17790), .C2(n19057), .A(n17454), .B(n17234), .ZN(
        n17235) );
  AOI21_X1 U19004 ( .B1(n19046), .B2(n17784), .A(n17235), .ZN(n17236) );
  OAI211_X1 U19005 ( .C1(n17238), .C2(n17774), .A(n17237), .B(n17236), .ZN(
        P2_U2997) );
  OAI211_X1 U19006 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n11239), .A(
        n17448), .B(n17782), .ZN(n17249) );
  INV_X1 U19007 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17242) );
  INV_X1 U19008 ( .A(n17239), .ZN(n17240) );
  NAND2_X1 U19009 ( .A1(n17754), .A2(n17240), .ZN(n17241) );
  NAND2_X1 U19010 ( .A1(n19047), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n17467) );
  OAI211_X1 U19011 ( .C1(n17762), .C2(n17242), .A(n17241), .B(n17467), .ZN(
        n17247) );
  NOR2_X1 U19012 ( .A1(n17244), .A2(n17243), .ZN(n17465) );
  INV_X1 U19013 ( .A(n17245), .ZN(n17464) );
  NOR3_X1 U19014 ( .A1(n17465), .A2(n17464), .A3(n17774), .ZN(n17246) );
  AOI211_X1 U19015 ( .C1(n17466), .C2(n17784), .A(n17247), .B(n17246), .ZN(
        n17248) );
  NAND2_X1 U19016 ( .A1(n17249), .A2(n17248), .ZN(P2_U2998) );
  INV_X1 U19017 ( .A(n11239), .ZN(n17458) );
  OAI21_X1 U19018 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17250), .A(
        n17458), .ZN(n17488) );
  NAND2_X1 U19019 ( .A1(n17252), .A2(n17251), .ZN(n17258) );
  INV_X1 U19020 ( .A(n17275), .ZN(n17254) );
  INV_X1 U19021 ( .A(n17272), .ZN(n17253) );
  OAI21_X1 U19022 ( .B1(n17254), .B2(n17253), .A(n17273), .ZN(n17266) );
  AND2_X1 U19023 ( .A1(n17256), .A2(n17255), .ZN(n17265) );
  NAND2_X1 U19024 ( .A1(n17266), .A2(n17265), .ZN(n17264) );
  NAND2_X1 U19025 ( .A1(n17264), .A2(n17256), .ZN(n17257) );
  XOR2_X1 U19026 ( .A(n17258), .B(n17257), .Z(n17486) );
  NAND2_X1 U19027 ( .A1(n19047), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n17477) );
  OAI21_X1 U19028 ( .B1(n17762), .B2(n19038), .A(n17477), .ZN(n17259) );
  AOI21_X1 U19029 ( .B1(n17754), .B2(n19034), .A(n17259), .ZN(n17260) );
  OAI21_X1 U19030 ( .B1(n19041), .B2(n17773), .A(n17260), .ZN(n17261) );
  AOI21_X1 U19031 ( .B1(n17486), .B2(n17785), .A(n17261), .ZN(n17262) );
  OAI21_X1 U19032 ( .B1(n17488), .B2(n17770), .A(n17262), .ZN(P2_U2999) );
  OAI21_X1 U19033 ( .B1(n17276), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17263), .ZN(n17502) );
  OAI21_X1 U19034 ( .B1(n17266), .B2(n17265), .A(n17264), .ZN(n17499) );
  NOR2_X1 U19035 ( .A1(n17493), .A2(n17773), .ZN(n17270) );
  NAND2_X1 U19036 ( .A1(n19047), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n17492) );
  NAND2_X1 U19037 ( .A1(n17780), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17267) );
  OAI211_X1 U19038 ( .C1(n17790), .C2(n17268), .A(n17492), .B(n17267), .ZN(
        n17269) );
  AOI211_X1 U19039 ( .C1(n17499), .C2(n17785), .A(n17270), .B(n17269), .ZN(
        n17271) );
  OAI21_X1 U19040 ( .B1(n17502), .B2(n17770), .A(n17271), .ZN(P2_U3000) );
  NAND2_X1 U19041 ( .A1(n17273), .A2(n17272), .ZN(n17274) );
  XNOR2_X1 U19042 ( .A(n17275), .B(n17274), .ZN(n17515) );
  AOI21_X1 U19043 ( .B1(n17504), .B2(n17516), .A(n17276), .ZN(n17503) );
  NAND2_X1 U19044 ( .A1(n17503), .A2(n17782), .ZN(n17282) );
  NAND2_X1 U19045 ( .A1(n19047), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n17506) );
  OAI21_X1 U19046 ( .B1(n17762), .B2(n17277), .A(n17506), .ZN(n17279) );
  NOR2_X1 U19047 ( .A1(n19027), .A2(n17773), .ZN(n17278) );
  AOI211_X1 U19048 ( .C1(n17280), .C2(n17754), .A(n17279), .B(n17278), .ZN(
        n17281) );
  OAI211_X1 U19049 ( .C1(n17774), .C2(n17515), .A(n17282), .B(n17281), .ZN(
        P2_U3001) );
  NAND2_X1 U19050 ( .A1(n11471), .A2(n17284), .ZN(n17286) );
  XOR2_X1 U19051 ( .A(n17286), .B(n17285), .Z(n17529) );
  NAND2_X1 U19052 ( .A1(n11811), .A2(n17523), .ZN(n17517) );
  NAND3_X1 U19053 ( .A1(n17517), .A2(n17782), .A3(n17516), .ZN(n17293) );
  NAND2_X1 U19054 ( .A1(n19047), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n17518) );
  OAI21_X1 U19055 ( .B1(n17762), .B2(n17288), .A(n17518), .ZN(n17291) );
  NOR2_X1 U19056 ( .A1(n17790), .A2(n17289), .ZN(n17290) );
  AOI211_X1 U19057 ( .C1(n17784), .C2(n17520), .A(n17291), .B(n17290), .ZN(
        n17292) );
  OAI211_X1 U19058 ( .C1(n17774), .C2(n17529), .A(n17293), .B(n17292), .ZN(
        P2_U3002) );
  INV_X1 U19059 ( .A(n17295), .ZN(n17296) );
  NOR2_X1 U19060 ( .A1(n17297), .A2(n17296), .ZN(n17298) );
  XNOR2_X1 U19061 ( .A(n17294), .B(n17298), .ZN(n17543) );
  AOI21_X1 U19062 ( .B1(n17533), .B2(n17304), .A(n17287), .ZN(n17530) );
  NAND2_X1 U19063 ( .A1(n17530), .A2(n17782), .ZN(n17303) );
  NAND2_X1 U19064 ( .A1(n19047), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U19065 ( .B1(n17762), .B2(n11682), .A(n17535), .ZN(n17301) );
  NOR2_X1 U19066 ( .A1(n17790), .A2(n17299), .ZN(n17300) );
  AOI211_X1 U19067 ( .C1(n17784), .C2(n17534), .A(n17301), .B(n17300), .ZN(
        n17302) );
  OAI211_X1 U19068 ( .C1(n17543), .C2(n17774), .A(n17303), .B(n17302), .ZN(
        P2_U3003) );
  OAI21_X1 U19069 ( .B1(n17315), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17304), .ZN(n17555) );
  NAND2_X1 U19070 ( .A1(n17327), .A2(n17322), .ZN(n17307) );
  NAND2_X1 U19071 ( .A1(n11311), .A2(n17305), .ZN(n17306) );
  XNOR2_X1 U19072 ( .A(n17307), .B(n17306), .ZN(n17552) );
  OAI22_X1 U19073 ( .A1(n17762), .A2(n11681), .B1(n17308), .B2(n19068), .ZN(
        n17309) );
  AOI21_X1 U19074 ( .B1(n17784), .B2(n17310), .A(n17309), .ZN(n17311) );
  OAI21_X1 U19075 ( .B1(n17790), .B2(n17312), .A(n17311), .ZN(n17313) );
  AOI21_X1 U19076 ( .B1(n17552), .B2(n17785), .A(n17313), .ZN(n17314) );
  OAI21_X1 U19077 ( .B1(n17555), .B2(n17770), .A(n17314), .ZN(P2_U3004) );
  INV_X1 U19078 ( .A(n17315), .ZN(n17557) );
  NAND2_X1 U19079 ( .A1(n17316), .A2(n17532), .ZN(n17556) );
  NAND3_X1 U19080 ( .A1(n17557), .A2(n17782), .A3(n17556), .ZN(n17331) );
  INV_X1 U19081 ( .A(n17317), .ZN(n19010) );
  OAI22_X1 U19082 ( .A1(n17318), .A2(n17762), .B1(n17790), .B2(n19010), .ZN(
        n17319) );
  AOI21_X1 U19083 ( .B1(n19047), .B2(P2_REIP_REG_9__SCAN_IN), .A(n17319), .ZN(
        n17330) );
  INV_X1 U19084 ( .A(n17322), .ZN(n17326) );
  AND2_X1 U19085 ( .A1(n17321), .A2(n17320), .ZN(n17325) );
  AND2_X1 U19086 ( .A1(n17323), .A2(n17322), .ZN(n17324) );
  OAI22_X1 U19087 ( .A1(n17327), .A2(n17326), .B1(n17325), .B2(n17324), .ZN(
        n17568) );
  OR2_X1 U19088 ( .A1(n17568), .A2(n17774), .ZN(n17329) );
  INV_X1 U19089 ( .A(n17559), .ZN(n19011) );
  NAND2_X1 U19090 ( .A1(n17784), .A2(n19011), .ZN(n17328) );
  NAND4_X1 U19091 ( .A1(n17331), .A2(n17330), .A3(n17329), .A4(n17328), .ZN(
        P2_U3005) );
  NAND2_X1 U19092 ( .A1(n17332), .A2(n17333), .ZN(n17574) );
  INV_X1 U19093 ( .A(n17573), .ZN(n17335) );
  AND2_X1 U19094 ( .A1(n17573), .A2(n17333), .ZN(n17334) );
  OAI22_X1 U19095 ( .A1(n17574), .A2(n17335), .B1(n17334), .B2(n17332), .ZN(
        n17609) );
  NAND2_X1 U19096 ( .A1(n17336), .A2(n17337), .ZN(n17595) );
  NAND3_X1 U19097 ( .A1(n11814), .A2(n17782), .A3(n17595), .ZN(n17342) );
  NOR2_X1 U19098 ( .A1(n17773), .A2(n19000), .ZN(n17340) );
  OAI22_X1 U19099 ( .A1(n17338), .A2(n17762), .B1(n18999), .B2(n19068), .ZN(
        n17339) );
  AOI211_X1 U19100 ( .C1(n18995), .C2(n17754), .A(n17340), .B(n17339), .ZN(
        n17341) );
  OAI211_X1 U19101 ( .C1(n17774), .C2(n17609), .A(n17342), .B(n17341), .ZN(
        P2_U3007) );
  OAI21_X1 U19102 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17344), .A(
        n17343), .ZN(n17348) );
  NOR2_X1 U19103 ( .A1(n17346), .A2(n17345), .ZN(n17347) );
  AOI211_X1 U19104 ( .C1(n19189), .C2(n19160), .A(n17348), .B(n17347), .ZN(
        n17349) );
  OAI21_X1 U19105 ( .B1(n19164), .B2(n19184), .A(n17349), .ZN(n17350) );
  AOI21_X1 U19106 ( .B1(n17351), .B2(n17628), .A(n17350), .ZN(n17352) );
  INV_X1 U19107 ( .A(n17354), .ZN(n17355) );
  OAI21_X1 U19108 ( .B1(n19154), .B2(n17622), .A(n17355), .ZN(n17357) );
  AOI211_X1 U19109 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n17358), .A(
        n17357), .B(n17356), .ZN(n17359) );
  OAI21_X1 U19110 ( .B1(n19150), .B2(n19184), .A(n17359), .ZN(n17360) );
  AOI21_X1 U19111 ( .B1(n17361), .B2(n17628), .A(n17360), .ZN(n17362) );
  OAI21_X1 U19112 ( .B1(n19182), .B2(n17363), .A(n17362), .ZN(P2_U3019) );
  AOI211_X1 U19113 ( .C1(n17377), .C2(n17365), .A(n17364), .B(n17382), .ZN(
        n17370) );
  INV_X1 U19114 ( .A(n17378), .ZN(n17367) );
  AOI21_X1 U19115 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17367), .A(
        n17366), .ZN(n17368) );
  OAI21_X1 U19116 ( .B1(n19129), .B2(n17622), .A(n17368), .ZN(n17369) );
  AOI211_X1 U19117 ( .C1(n19132), .C2(n17633), .A(n17370), .B(n17369), .ZN(
        n17373) );
  NAND2_X1 U19118 ( .A1(n17371), .A2(n17636), .ZN(n17372) );
  OAI211_X1 U19119 ( .C1(n17374), .C2(n19193), .A(n17373), .B(n17372), .ZN(
        P2_U3020) );
  INV_X1 U19120 ( .A(n17375), .ZN(n17384) );
  OAI21_X1 U19121 ( .B1(n17378), .B2(n17377), .A(n17376), .ZN(n17379) );
  AOI21_X1 U19122 ( .B1(n17380), .B2(n19189), .A(n17379), .ZN(n17381) );
  OAI21_X1 U19123 ( .B1(n17382), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17381), .ZN(n17383) );
  AOI21_X1 U19124 ( .B1(n17384), .B2(n17633), .A(n17383), .ZN(n17387) );
  NAND2_X1 U19125 ( .A1(n17385), .A2(n17636), .ZN(n17386) );
  OAI211_X1 U19126 ( .C1(n17388), .C2(n19193), .A(n17387), .B(n17386), .ZN(
        P2_U3021) );
  AOI21_X1 U19127 ( .B1(n17400), .B2(n17389), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17390) );
  NOR2_X1 U19128 ( .A1(n17391), .A2(n17390), .ZN(n17392) );
  AOI211_X1 U19129 ( .C1(n19189), .C2(n19119), .A(n17393), .B(n17392), .ZN(
        n17394) );
  OAI21_X1 U19130 ( .B1(n19184), .B2(n19117), .A(n17394), .ZN(n17395) );
  AOI21_X1 U19131 ( .B1(n17396), .B2(n17628), .A(n17395), .ZN(n17397) );
  OAI21_X1 U19132 ( .B1(n17398), .B2(n19182), .A(n17397), .ZN(P2_U3022) );
  OAI211_X1 U19133 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17400), .B(n17399), .ZN(
        n17402) );
  OAI211_X1 U19134 ( .C1(n17622), .C2(n19101), .A(n17402), .B(n17401), .ZN(
        n17403) );
  AOI21_X1 U19135 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17416), .A(
        n17403), .ZN(n17404) );
  OAI21_X1 U19136 ( .B1(n19100), .B2(n19184), .A(n17404), .ZN(n17405) );
  AOI21_X1 U19137 ( .B1(n17406), .B2(n17636), .A(n17405), .ZN(n17407) );
  OAI21_X1 U19138 ( .B1(n17408), .B2(n19193), .A(n17407), .ZN(P2_U3023) );
  OAI21_X1 U19139 ( .B1(n17411), .B2(n17410), .A(n17409), .ZN(n19090) );
  OAI21_X1 U19140 ( .B1(n17622), .B2(n19090), .A(n17412), .ZN(n17415) );
  NOR2_X1 U19141 ( .A1(n17413), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17414) );
  AOI211_X1 U19142 ( .C1(n17416), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n17415), .B(n17414), .ZN(n17417) );
  OAI21_X1 U19143 ( .B1(n19089), .B2(n19184), .A(n17417), .ZN(n17418) );
  AOI21_X1 U19144 ( .B1(n17419), .B2(n17636), .A(n17418), .ZN(n17420) );
  OAI21_X1 U19145 ( .B1(n17421), .B2(n19193), .A(n17420), .ZN(P2_U3024) );
  INV_X1 U19146 ( .A(n19076), .ZN(n17431) );
  OR3_X1 U19147 ( .A1(n17563), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n17422), .ZN(n17427) );
  INV_X1 U19148 ( .A(n17423), .ZN(n17424) );
  AOI21_X1 U19149 ( .B1(n19189), .B2(n17425), .A(n17424), .ZN(n17426) );
  OAI211_X1 U19150 ( .C1(n17429), .C2(n17428), .A(n17427), .B(n17426), .ZN(
        n17430) );
  AOI21_X1 U19151 ( .B1(n17431), .B2(n17633), .A(n17430), .ZN(n17434) );
  NAND2_X1 U19152 ( .A1(n17432), .A2(n17636), .ZN(n17433) );
  OAI211_X1 U19153 ( .C1(n17435), .C2(n19193), .A(n17434), .B(n17433), .ZN(
        P2_U3025) );
  INV_X1 U19154 ( .A(n17436), .ZN(n19063) );
  OAI211_X1 U19155 ( .C1(n17622), .C2(n17439), .A(n17438), .B(n17437), .ZN(
        n17440) );
  AOI21_X1 U19156 ( .B1(n19063), .B2(n17633), .A(n17440), .ZN(n17441) );
  OAI21_X1 U19157 ( .B1(n17443), .B2(n17442), .A(n17441), .ZN(n17444) );
  AOI21_X1 U19158 ( .B1(n17445), .B2(n17636), .A(n17444), .ZN(n17446) );
  OAI21_X1 U19159 ( .B1(n17447), .B2(n19193), .A(n17446), .ZN(P2_U3027) );
  INV_X1 U19160 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17473) );
  OAI21_X1 U19161 ( .B1(n17628), .B2(n17585), .A(n17448), .ZN(n17453) );
  AOI21_X1 U19162 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17449), .A(
        n17579), .ZN(n17451) );
  NOR3_X1 U19163 ( .A1(n17452), .A2(n17451), .A3(n17450), .ZN(n17479) );
  NAND2_X1 U19164 ( .A1(n17453), .A2(n17479), .ZN(n17463) );
  AOI21_X1 U19165 ( .B1(n17473), .B2(n19186), .A(n17463), .ZN(n17462) );
  NAND2_X1 U19166 ( .A1(n19046), .A2(n17633), .ZN(n17455) );
  OAI211_X1 U19167 ( .C1(n17622), .C2(n19061), .A(n17455), .B(n17454), .ZN(
        n17456) );
  AOI21_X1 U19168 ( .B1(n17457), .B2(n17636), .A(n17456), .ZN(n17460) );
  OAI22_X1 U19169 ( .A1(n17458), .A2(n19193), .B1(n17478), .B2(n17484), .ZN(
        n17471) );
  NAND3_X1 U19170 ( .A1(n17471), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17461), .ZN(n17459) );
  OAI211_X1 U19171 ( .C1(n17462), .C2(n17461), .A(n17460), .B(n17459), .ZN(
        P2_U3029) );
  INV_X1 U19172 ( .A(n17463), .ZN(n17474) );
  NOR3_X1 U19173 ( .A1(n17465), .A2(n17464), .A3(n19182), .ZN(n17470) );
  NAND2_X1 U19174 ( .A1(n17466), .A2(n17633), .ZN(n17468) );
  OAI211_X1 U19175 ( .C1(n17622), .C2(n20226), .A(n17468), .B(n17467), .ZN(
        n17469) );
  AOI211_X1 U19176 ( .C1(n17471), .C2(n17473), .A(n17470), .B(n17469), .ZN(
        n17472) );
  OAI21_X1 U19177 ( .B1(n17474), .B2(n17473), .A(n17472), .ZN(P2_U3030) );
  OR2_X1 U19178 ( .A1(n15803), .A2(n17475), .ZN(n17476) );
  NAND2_X1 U19179 ( .A1(n17476), .A2(n15787), .ZN(n19692) );
  OAI21_X1 U19180 ( .B1(n17622), .B2(n19692), .A(n17477), .ZN(n17481) );
  NOR2_X1 U19181 ( .A1(n17479), .A2(n17478), .ZN(n17480) );
  AOI211_X1 U19182 ( .C1(n17482), .C2(n17633), .A(n17481), .B(n17480), .ZN(
        n17483) );
  OAI21_X1 U19183 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17484), .A(
        n17483), .ZN(n17485) );
  AOI21_X1 U19184 ( .B1(n17486), .B2(n17636), .A(n17485), .ZN(n17487) );
  OAI21_X1 U19185 ( .B1(n17488), .B2(n19193), .A(n17487), .ZN(P2_U3031) );
  OR3_X1 U19186 ( .A1(n17563), .A2(n17532), .A3(n17547), .ZN(n17537) );
  OR2_X1 U19187 ( .A1(n17537), .A2(n17533), .ZN(n17494) );
  INV_X1 U19188 ( .A(n17494), .ZN(n17505) );
  NAND2_X1 U19189 ( .A1(n17505), .A2(n17523), .ZN(n17522) );
  AOI21_X1 U19190 ( .B1(n17489), .B2(n19186), .A(n17561), .ZN(n17524) );
  NAND2_X1 U19191 ( .A1(n17522), .A2(n17524), .ZN(n17512) );
  INV_X1 U19192 ( .A(n19695), .ZN(n17490) );
  NAND2_X1 U19193 ( .A1(n19189), .A2(n17490), .ZN(n17491) );
  OAI211_X1 U19194 ( .C1(n17493), .C2(n19184), .A(n17492), .B(n17491), .ZN(
        n17498) );
  AOI21_X1 U19195 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17496), .A(
        n17504), .ZN(n17495) );
  AOI211_X1 U19196 ( .C1(n17504), .C2(n17496), .A(n17495), .B(n17494), .ZN(
        n17497) );
  AOI211_X1 U19197 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17512), .A(
        n17498), .B(n17497), .ZN(n17501) );
  NAND2_X1 U19198 ( .A1(n17499), .A2(n17636), .ZN(n17500) );
  OAI211_X1 U19199 ( .C1(n17502), .C2(n19193), .A(n17501), .B(n17500), .ZN(
        P2_U3032) );
  NAND2_X1 U19200 ( .A1(n17503), .A2(n17628), .ZN(n17514) );
  NAND3_X1 U19201 ( .A1(n17505), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n17504), .ZN(n17507) );
  OAI211_X1 U19202 ( .C1(n19027), .C2(n19184), .A(n17507), .B(n17506), .ZN(
        n17511) );
  INV_X1 U19203 ( .A(n15804), .ZN(n17508) );
  OAI21_X1 U19204 ( .B1(n15923), .B2(n17509), .A(n17508), .ZN(n19698) );
  NOR2_X1 U19205 ( .A1(n19698), .A2(n17622), .ZN(n17510) );
  AOI211_X1 U19206 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n17512), .A(
        n17511), .B(n17510), .ZN(n17513) );
  OAI211_X1 U19207 ( .C1(n17515), .C2(n19182), .A(n17514), .B(n17513), .ZN(
        P2_U3033) );
  NAND3_X1 U19208 ( .A1(n17517), .A2(n17628), .A3(n17516), .ZN(n17528) );
  INV_X1 U19209 ( .A(n17518), .ZN(n17519) );
  AOI21_X1 U19210 ( .B1(n17520), .B2(n17633), .A(n17519), .ZN(n17521) );
  OAI211_X1 U19211 ( .C1(n17524), .C2(n17523), .A(n17522), .B(n17521), .ZN(
        n17525) );
  AOI21_X1 U19212 ( .B1(n17526), .B2(n19189), .A(n17525), .ZN(n17527) );
  OAI211_X1 U19213 ( .C1(n17529), .C2(n19182), .A(n17528), .B(n17527), .ZN(
        P2_U3034) );
  NAND2_X1 U19214 ( .A1(n17530), .A2(n17628), .ZN(n17542) );
  INV_X1 U19215 ( .A(n19704), .ZN(n17540) );
  INV_X1 U19216 ( .A(n17563), .ZN(n17531) );
  NAND3_X1 U19217 ( .A1(n17531), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17547), .ZN(n17546) );
  AOI21_X1 U19218 ( .B1(n17532), .B2(n19186), .A(n17561), .ZN(n17548) );
  AOI21_X1 U19219 ( .B1(n17546), .B2(n17548), .A(n17533), .ZN(n17539) );
  NAND2_X1 U19220 ( .A1(n17534), .A2(n17633), .ZN(n17536) );
  OAI211_X1 U19221 ( .C1(n17537), .C2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17536), .B(n17535), .ZN(n17538) );
  AOI211_X1 U19222 ( .C1(n17540), .C2(n19189), .A(n17539), .B(n17538), .ZN(
        n17541) );
  OAI211_X1 U19223 ( .C1(n17543), .C2(n19182), .A(n17542), .B(n17541), .ZN(
        P2_U3035) );
  NOR2_X1 U19224 ( .A1(n19184), .A2(n17544), .ZN(n17550) );
  NAND2_X1 U19225 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19047), .ZN(n17545) );
  OAI211_X1 U19226 ( .C1(n17548), .C2(n17547), .A(n17546), .B(n17545), .ZN(
        n17549) );
  AOI211_X1 U19227 ( .C1(n17551), .C2(n19189), .A(n17550), .B(n17549), .ZN(
        n17554) );
  NAND2_X1 U19228 ( .A1(n17552), .A2(n17636), .ZN(n17553) );
  OAI211_X1 U19229 ( .C1(n17555), .C2(n19193), .A(n17554), .B(n17553), .ZN(
        P2_U3036) );
  NAND3_X1 U19230 ( .A1(n17557), .A2(n17628), .A3(n17556), .ZN(n17567) );
  OAI21_X1 U19231 ( .B1(n15838), .B2(n17558), .A(n15811), .ZN(n19710) );
  INV_X1 U19232 ( .A(n19710), .ZN(n17565) );
  OAI22_X1 U19233 ( .A1(n19184), .A2(n17559), .B1(n13200), .B2(n19068), .ZN(
        n17560) );
  AOI21_X1 U19234 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17561), .A(
        n17560), .ZN(n17562) );
  OAI21_X1 U19235 ( .B1(n17563), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17562), .ZN(n17564) );
  AOI21_X1 U19236 ( .B1(n17565), .B2(n19189), .A(n17564), .ZN(n17566) );
  OAI211_X1 U19237 ( .C1(n17568), .C2(n19182), .A(n17567), .B(n17566), .ZN(
        P2_U3037) );
  AOI21_X1 U19238 ( .B1(n11257), .B2(n17572), .A(n17571), .ZN(n17781) );
  INV_X1 U19239 ( .A(n17781), .ZN(n17594) );
  NAND2_X1 U19240 ( .A1(n17574), .A2(n17573), .ZN(n17578) );
  NAND2_X1 U19241 ( .A1(n17576), .A2(n17575), .ZN(n17577) );
  XNOR2_X1 U19242 ( .A(n17578), .B(n17577), .ZN(n17786) );
  INV_X1 U19243 ( .A(n17613), .ZN(n17580) );
  OAI22_X1 U19244 ( .A1(n17581), .A2(n17580), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17579), .ZN(n17582) );
  INV_X1 U19245 ( .A(n17582), .ZN(n17583) );
  NAND2_X1 U19246 ( .A1(n17584), .A2(n17583), .ZN(n17617) );
  AOI21_X1 U19247 ( .B1(n17585), .B2(n17616), .A(n17617), .ZN(n17599) );
  OAI21_X1 U19248 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n17606), .ZN(n17586) );
  OAI22_X1 U19249 ( .A1(n19068), .A2(n15841), .B1(n17587), .B2(n17586), .ZN(
        n17588) );
  AOI21_X1 U19250 ( .B1(n17633), .B2(n17783), .A(n17588), .ZN(n17590) );
  NAND2_X1 U19251 ( .A1(n19189), .A2(n19711), .ZN(n17589) );
  OAI211_X1 U19252 ( .C1(n17599), .C2(n17591), .A(n17590), .B(n17589), .ZN(
        n17592) );
  AOI21_X1 U19253 ( .B1(n17786), .B2(n17636), .A(n17592), .ZN(n17593) );
  OAI21_X1 U19254 ( .B1(n17594), .B2(n19193), .A(n17593), .ZN(P2_U3038) );
  NAND3_X1 U19255 ( .A1(n11814), .A2(n17628), .A3(n17595), .ZN(n17608) );
  INV_X1 U19256 ( .A(n19000), .ZN(n17597) );
  NOR2_X1 U19257 ( .A1(n18999), .A2(n19068), .ZN(n17596) );
  AOI21_X1 U19258 ( .B1(n17633), .B2(n17597), .A(n17596), .ZN(n17598) );
  OAI21_X1 U19259 ( .B1(n17599), .B2(n17605), .A(n17598), .ZN(n17604) );
  OAI21_X1 U19260 ( .B1(n17602), .B2(n17601), .A(n17600), .ZN(n19716) );
  NOR2_X1 U19261 ( .A1(n19716), .A2(n17622), .ZN(n17603) );
  AOI211_X1 U19262 ( .C1(n17606), .C2(n17605), .A(n17604), .B(n17603), .ZN(
        n17607) );
  OAI211_X1 U19263 ( .C1(n17609), .C2(n19182), .A(n17608), .B(n17607), .ZN(
        P2_U3039) );
  XNOR2_X1 U19264 ( .A(n17610), .B(n17611), .ZN(n17775) );
  OR3_X1 U19265 ( .A1(n17612), .A2(n17771), .A3(n19193), .ZN(n17626) );
  NOR2_X1 U19266 ( .A1(n17614), .A2(n17613), .ZN(n17615) );
  NAND2_X1 U19267 ( .A1(n17616), .A2(n17615), .ZN(n17619) );
  NAND2_X1 U19268 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17617), .ZN(
        n17618) );
  OAI211_X1 U19269 ( .C1(n19068), .C2(n13185), .A(n17619), .B(n17618), .ZN(
        n17624) );
  XNOR2_X1 U19270 ( .A(n17621), .B(n17620), .ZN(n19931) );
  NOR2_X1 U19271 ( .A1(n19931), .A2(n17622), .ZN(n17623) );
  AOI211_X1 U19272 ( .C1(n18990), .C2(n17633), .A(n17624), .B(n17623), .ZN(
        n17625) );
  OAI211_X1 U19273 ( .C1(n17775), .C2(n19182), .A(n17626), .B(n17625), .ZN(
        P2_U3040) );
  NAND2_X1 U19274 ( .A1(n17628), .A2(n17627), .ZN(n17630) );
  OAI211_X1 U19275 ( .C1(n17631), .C2(n14719), .A(n17630), .B(n17629), .ZN(
        n17632) );
  AOI21_X1 U19276 ( .B1(n17634), .B2(n17633), .A(n17632), .ZN(n17640) );
  AOI22_X1 U19277 ( .A1(n17636), .A2(n17635), .B1(n19189), .B2(n20168), .ZN(
        n17639) );
  OAI211_X1 U19278 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19186), .B(n17637), .ZN(n17638) );
  NAND3_X1 U19279 ( .A1(n17640), .A2(n17639), .A3(n17638), .ZN(P2_U3045) );
  NOR2_X1 U19280 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17803) );
  AOI22_X1 U19281 ( .A1(n19134), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n17642), .B2(n19032), .ZN(n17648) );
  AOI22_X1 U19282 ( .A1(n17643), .A2(n17803), .B1(P2_STATE2_REG_1__SCAN_IN), 
        .B2(n17648), .ZN(n17644) );
  OAI21_X1 U19283 ( .B1(n19732), .B2(n17659), .A(n17644), .ZN(n17647) );
  OAI22_X1 U19284 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19876), .B1(n17645), 
        .B2(n19219), .ZN(n17646) );
  AOI21_X1 U19285 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17689), .A(n17646), .ZN(
        n17660) );
  MUX2_X1 U19286 ( .A(n17647), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n17660), .Z(P2_U3601) );
  NOR2_X1 U19287 ( .A1(n17648), .A2(n13265), .ZN(n17653) );
  AOI21_X1 U19288 ( .B1(n19134), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n17649), .ZN(n17655) );
  AOI222_X1 U19289 ( .A1(n17803), .A2(n17650), .B1(n17653), .B2(n17655), .C1(
        n19745), .C2(n19211), .ZN(n17652) );
  NAND2_X1 U19290 ( .A1(n17660), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17651) );
  OAI21_X1 U19291 ( .B1(n17660), .B2(n17652), .A(n17651), .ZN(P2_U3600) );
  INV_X1 U19292 ( .A(n17653), .ZN(n17656) );
  INV_X1 U19293 ( .A(n17803), .ZN(n19196) );
  OAI222_X1 U19294 ( .A1(n17659), .A2(n17805), .B1(n17656), .B2(n17655), .C1(
        n19196), .C2(n17654), .ZN(n17657) );
  MUX2_X1 U19295 ( .A(n17657), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n17660), .Z(P2_U3599) );
  OAI22_X1 U19296 ( .A1(n19768), .A2(n17659), .B1(n17658), .B2(n19196), .ZN(
        n17661) );
  INV_X1 U19297 ( .A(n17660), .ZN(n19180) );
  MUX2_X1 U19298 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17661), .S(
        n19180), .Z(P2_U3596) );
  NAND2_X1 U19299 ( .A1(n21806), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19286) );
  INV_X1 U19300 ( .A(n19286), .ZN(n19251) );
  OR2_X1 U19301 ( .A1(n17662), .A2(n18348), .ZN(n18277) );
  NAND2_X1 U19302 ( .A1(n21314), .A2(n20629), .ZN(n21843) );
  NAND2_X1 U19303 ( .A1(n21802), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21842) );
  INV_X1 U19304 ( .A(n21842), .ZN(n21358) );
  AOI21_X1 U19305 ( .B1(n21843), .B2(n18276), .A(n21358), .ZN(n17663) );
  INV_X1 U19306 ( .A(n17663), .ZN(n19252) );
  NAND2_X1 U19307 ( .A1(n21841), .A2(n19252), .ZN(n19586) );
  INV_X1 U19308 ( .A(n19586), .ZN(n19536) );
  AOI211_X1 U19309 ( .C1(n17677), .C2(n18277), .A(n19536), .B(n17664), .ZN(
        n18837) );
  AND2_X1 U19310 ( .A1(n21836), .A2(n18276), .ZN(n20633) );
  INV_X1 U19311 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n22243) );
  NOR2_X1 U19312 ( .A1(n21314), .A2(n22243), .ZN(n18700) );
  INV_X1 U19313 ( .A(n18700), .ZN(n18791) );
  NAND2_X1 U19314 ( .A1(n20633), .A2(n18791), .ZN(n17666) );
  NOR2_X1 U19315 ( .A1(n21809), .A2(n21815), .ZN(n19249) );
  AOI21_X1 U19316 ( .B1(n21836), .B2(n17666), .A(n19249), .ZN(n17665) );
  NOR3_X1 U19317 ( .A1(n19251), .A2(n18837), .A3(n17665), .ZN(n18836) );
  NAND3_X1 U19318 ( .A1(n20629), .A2(n21836), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19310) );
  INV_X1 U19319 ( .A(n19310), .ZN(n19289) );
  NAND2_X1 U19320 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17667) );
  AOI21_X1 U19321 ( .B1(n17667), .B2(n17666), .A(n18837), .ZN(n18838) );
  NOR2_X1 U19322 ( .A1(n19310), .A2(n19586), .ZN(n18834) );
  OAI22_X1 U19323 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19289), .B1(
        n18838), .B2(n18834), .ZN(n17668) );
  AOI22_X1 U19324 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18836), .B1(
        n17668), .B2(n21815), .ZN(P3_U2865) );
  OR3_X1 U19325 ( .A1(n17671), .A2(n17670), .A3(n17669), .ZN(n17672) );
  OAI21_X1 U19326 ( .B1(n17674), .B2(n17673), .A(n17672), .ZN(P1_U3468) );
  OAI21_X1 U19327 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n22250), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18914) );
  NAND2_X1 U19328 ( .A1(n22298), .A2(n18914), .ZN(n17676) );
  INV_X1 U19329 ( .A(n17676), .ZN(n22246) );
  NOR2_X1 U19330 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n22247) );
  OAI21_X1 U19331 ( .B1(BS16), .B2(n22247), .A(n22246), .ZN(n22244) );
  OAI21_X1 U19332 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n22246), .A(n22244), 
        .ZN(n17675) );
  INV_X1 U19333 ( .A(n17675), .ZN(P3_U3280) );
  AND2_X1 U19334 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17676), .ZN(P3_U3028) );
  AND2_X1 U19335 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17676), .ZN(P3_U3027) );
  AND2_X1 U19336 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17676), .ZN(P3_U3026) );
  AND2_X1 U19337 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17676), .ZN(P3_U3025) );
  AND2_X1 U19338 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17676), .ZN(P3_U3024) );
  AND2_X1 U19339 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17676), .ZN(P3_U3023) );
  AND2_X1 U19340 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17676), .ZN(P3_U3022) );
  AND2_X1 U19341 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17676), .ZN(P3_U3021) );
  AND2_X1 U19342 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17676), .ZN(
        P3_U3020) );
  AND2_X1 U19343 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17676), .ZN(
        P3_U3019) );
  AND2_X1 U19344 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17676), .ZN(
        P3_U3018) );
  AND2_X1 U19345 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17676), .ZN(
        P3_U3017) );
  AND2_X1 U19346 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17676), .ZN(
        P3_U3016) );
  AND2_X1 U19347 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17676), .ZN(
        P3_U3015) );
  AND2_X1 U19348 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17676), .ZN(
        P3_U3014) );
  AND2_X1 U19349 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17676), .ZN(
        P3_U3013) );
  AND2_X1 U19350 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17676), .ZN(
        P3_U3012) );
  AND2_X1 U19351 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17676), .ZN(
        P3_U3011) );
  AND2_X1 U19352 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17676), .ZN(
        P3_U3010) );
  AND2_X1 U19353 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17676), .ZN(
        P3_U3009) );
  AND2_X1 U19354 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17676), .ZN(
        P3_U3008) );
  AND2_X1 U19355 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17676), .ZN(
        P3_U3007) );
  AND2_X1 U19356 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17676), .ZN(
        P3_U3006) );
  AND2_X1 U19357 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17676), .ZN(
        P3_U3005) );
  AND2_X1 U19358 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17676), .ZN(
        P3_U3004) );
  AND2_X1 U19359 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17676), .ZN(
        P3_U3003) );
  AND2_X1 U19360 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17676), .ZN(
        P3_U3002) );
  AND2_X1 U19361 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17676), .ZN(
        P3_U3001) );
  AND2_X1 U19362 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17676), .ZN(
        P3_U3000) );
  AND2_X1 U19363 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17676), .ZN(
        P3_U2999) );
  AOI21_X1 U19364 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17678)
         );
  NOR4_X1 U19365 ( .A1(n21314), .A2(n21841), .A3(n22297), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n21786) );
  AOI211_X1 U19366 ( .C1(n18791), .C2(n17678), .A(n17677), .B(n21786), .ZN(
        P3_U2998) );
  AND2_X1 U19367 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18837), .ZN(
        P3_U2867) );
  NAND2_X1 U19368 ( .A1(n21841), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18827) );
  NAND2_X1 U19369 ( .A1(n21826), .A2(n21793), .ZN(n20639) );
  NAND2_X1 U19370 ( .A1(n21371), .A2(n17680), .ZN(n17679) );
  AND2_X1 U19371 ( .A1(n18903), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NOR2_X1 U19372 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21843), .ZN(n18274) );
  NOR2_X1 U19373 ( .A1(n18274), .A2(n20682), .ZN(n17683) );
  INV_X1 U19374 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18863) );
  NOR2_X1 U19375 ( .A1(n17682), .A2(n17681), .ZN(n18394) );
  INV_X1 U19376 ( .A(n18394), .ZN(n20631) );
  AOI22_X1 U19377 ( .A1(n17683), .A2(n18863), .B1(n20682), .B2(n20631), .ZN(
        P3_U3298) );
  INV_X1 U19378 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18862) );
  NAND2_X1 U19379 ( .A1(n19589), .A2(n20682), .ZN(n21113) );
  INV_X1 U19380 ( .A(n21113), .ZN(n20721) );
  AOI21_X1 U19381 ( .B1(n17683), .B2(n18862), .A(n20721), .ZN(P3_U3299) );
  NOR2_X1 U19382 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17685), .ZN(n22280) );
  AOI22_X1 U19383 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n22280), .B1(n17685), 
        .B2(n17684), .ZN(n17687) );
  INV_X1 U19384 ( .A(n17687), .ZN(n22242) );
  NOR2_X1 U19385 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n22273) );
  OAI21_X1 U19386 ( .B1(BS16), .B2(n22273), .A(n22242), .ZN(n22240) );
  OAI21_X1 U19387 ( .B1(n22242), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n22240), 
        .ZN(n17686) );
  INV_X1 U19388 ( .A(n17686), .ZN(P2_U3591) );
  AND2_X1 U19389 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17687), .ZN(P2_U3208) );
  AND2_X1 U19390 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17687), .ZN(P2_U3207) );
  INV_X1 U19391 ( .A(n22242), .ZN(n17688) );
  AND2_X1 U19392 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17688), .ZN(P2_U3206) );
  AND2_X1 U19393 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17687), .ZN(P2_U3205) );
  AND2_X1 U19394 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17688), .ZN(P2_U3204) );
  AND2_X1 U19395 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17687), .ZN(P2_U3203) );
  AND2_X1 U19396 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17688), .ZN(P2_U3202) );
  AND2_X1 U19397 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17687), .ZN(P2_U3201) );
  AND2_X1 U19398 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17688), .ZN(
        P2_U3200) );
  AND2_X1 U19399 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17687), .ZN(
        P2_U3199) );
  AND2_X1 U19400 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17687), .ZN(
        P2_U3198) );
  AND2_X1 U19401 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17688), .ZN(
        P2_U3197) );
  AND2_X1 U19402 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17688), .ZN(
        P2_U3196) );
  AND2_X1 U19403 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17688), .ZN(
        P2_U3195) );
  AND2_X1 U19404 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17688), .ZN(
        P2_U3194) );
  AND2_X1 U19405 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17688), .ZN(
        P2_U3193) );
  AND2_X1 U19406 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17687), .ZN(
        P2_U3192) );
  AND2_X1 U19407 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17687), .ZN(
        P2_U3191) );
  AND2_X1 U19408 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17687), .ZN(
        P2_U3190) );
  AND2_X1 U19409 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17687), .ZN(
        P2_U3189) );
  AND2_X1 U19410 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17687), .ZN(
        P2_U3188) );
  AND2_X1 U19411 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17687), .ZN(
        P2_U3187) );
  AND2_X1 U19412 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17688), .ZN(
        P2_U3186) );
  AND2_X1 U19413 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17688), .ZN(
        P2_U3185) );
  AND2_X1 U19414 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17688), .ZN(
        P2_U3184) );
  AND2_X1 U19415 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17688), .ZN(
        P2_U3183) );
  AND2_X1 U19416 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17688), .ZN(
        P2_U3182) );
  AND2_X1 U19417 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17688), .ZN(
        P2_U3181) );
  AND2_X1 U19418 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17688), .ZN(
        P2_U3180) );
  AND2_X1 U19419 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17688), .ZN(
        P2_U3179) );
  OAI221_X1 U19420 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(
        P2_STATEBS16_REG_SCAN_IN), .C1(n17752), .C2(n19213), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n17691) );
  AOI21_X1 U19421 ( .B1(n17691), .B2(n17690), .A(n17689), .ZN(P2_U3178) );
  NAND2_X1 U19422 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n17752), .ZN(n18963) );
  NAND2_X1 U19423 ( .A1(n17692), .A2(n18963), .ZN(n19214) );
  NAND2_X1 U19424 ( .A1(n17693), .A2(n19214), .ZN(n19725) );
  OAI221_X1 U19425 ( .B1(n14245), .B2(n19205), .C1(n19203), .C2(n19205), .A(
        n20234), .ZN(n17809) );
  NOR2_X1 U19426 ( .A1(n17695), .A2(n17809), .ZN(P2_U3047) );
  AND2_X1 U19427 ( .A1(n17836), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19428 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17699) );
  NOR4_X1 U19429 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17698) );
  NOR4_X1 U19430 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17697) );
  NOR4_X1 U19431 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17696) );
  NAND4_X1 U19432 ( .A1(n17699), .A2(n17698), .A3(n17697), .A4(n17696), .ZN(
        n17705) );
  NOR4_X1 U19433 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17703) );
  AOI211_X1 U19434 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17702) );
  NOR4_X1 U19435 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17701) );
  NOR4_X1 U19436 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17700) );
  NAND4_X1 U19437 ( .A1(n17703), .A2(n17702), .A3(n17701), .A4(n17700), .ZN(
        n17704) );
  NOR2_X1 U19438 ( .A1(n17705), .A2(n17704), .ZN(n17819) );
  INV_X1 U19439 ( .A(n17819), .ZN(n17817) );
  NOR2_X1 U19440 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17817), .ZN(n17812) );
  OR3_X1 U19441 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17816) );
  INV_X1 U19442 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17706) );
  AOI22_X1 U19443 ( .A1(n17812), .A2(n17816), .B1(n17817), .B2(n17706), .ZN(
        P2_U2821) );
  INV_X1 U19444 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17707) );
  AOI22_X1 U19445 ( .A1(n17812), .A2(n13343), .B1(n17817), .B2(n17707), .ZN(
        P2_U2820) );
  INV_X1 U19446 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17709) );
  NAND2_X1 U19447 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n22259), .ZN(n22806) );
  INV_X1 U19448 ( .A(n22806), .ZN(n22805) );
  AND2_X1 U19449 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n22266), .ZN(n17750) );
  OR2_X1 U19450 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n22270) );
  AOI21_X1 U19451 ( .B1(n17708), .B2(n22270), .A(n17710), .ZN(n22237) );
  AOI21_X1 U19452 ( .B1(n17709), .B2(n17710), .A(n22237), .ZN(P1_U3464) );
  AND2_X1 U19453 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n17710), .ZN(P1_U3193) );
  AND2_X1 U19454 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n17710), .ZN(P1_U3192) );
  AND2_X1 U19455 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n17710), .ZN(P1_U3191) );
  AND2_X1 U19456 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n17710), .ZN(P1_U3190) );
  AND2_X1 U19457 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n17710), .ZN(P1_U3189) );
  AND2_X1 U19458 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n17710), .ZN(P1_U3188) );
  AND2_X1 U19459 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n17710), .ZN(P1_U3187) );
  AND2_X1 U19460 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n17710), .ZN(P1_U3186) );
  AND2_X1 U19461 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n17710), .ZN(
        P1_U3185) );
  AND2_X1 U19462 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n17710), .ZN(
        P1_U3184) );
  AND2_X1 U19463 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n17710), .ZN(
        P1_U3183) );
  AND2_X1 U19464 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n17710), .ZN(
        P1_U3182) );
  AND2_X1 U19465 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n17710), .ZN(
        P1_U3181) );
  AND2_X1 U19466 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n17710), .ZN(
        P1_U3180) );
  AND2_X1 U19467 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n17710), .ZN(
        P1_U3179) );
  AND2_X1 U19468 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n17710), .ZN(
        P1_U3178) );
  AND2_X1 U19469 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n17710), .ZN(
        P1_U3177) );
  AND2_X1 U19470 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n17710), .ZN(
        P1_U3176) );
  AND2_X1 U19471 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n17710), .ZN(
        P1_U3175) );
  AND2_X1 U19472 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n17710), .ZN(
        P1_U3174) );
  AND2_X1 U19473 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n17710), .ZN(
        P1_U3173) );
  AND2_X1 U19474 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n17710), .ZN(
        P1_U3172) );
  AND2_X1 U19475 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n17710), .ZN(
        P1_U3171) );
  AND2_X1 U19476 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n17710), .ZN(
        P1_U3170) );
  AND2_X1 U19477 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n17710), .ZN(
        P1_U3169) );
  AND2_X1 U19478 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n17710), .ZN(
        P1_U3168) );
  AND2_X1 U19479 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n17710), .ZN(
        P1_U3167) );
  AND2_X1 U19480 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n17710), .ZN(
        P1_U3166) );
  AND2_X1 U19481 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n17710), .ZN(
        P1_U3165) );
  AND2_X1 U19482 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n17710), .ZN(
        P1_U3164) );
  NAND2_X1 U19483 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21855), .ZN(n22223) );
  OAI21_X1 U19484 ( .B1(n22253), .B2(n22223), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n22222) );
  AOI21_X1 U19485 ( .B1(n17711), .B2(n22225), .A(n22222), .ZN(n17746) );
  INV_X1 U19486 ( .A(n17712), .ZN(n17717) );
  OR3_X1 U19487 ( .A1(n17715), .A2(n17714), .A3(n17713), .ZN(n17716) );
  OAI221_X1 U19488 ( .B1(n17718), .B2(n17717), .C1(n17718), .C2(n22254), .A(
        n17716), .ZN(n17745) );
  NOR3_X1 U19489 ( .A1(n17720), .A2(n17719), .A3(n22485), .ZN(n17723) );
  NAND2_X1 U19490 ( .A1(n17723), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n17725) );
  OAI22_X1 U19491 ( .A1(n17723), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n17722), .B2(n17721), .ZN(n17724) );
  NAND2_X1 U19492 ( .A1(n17725), .A2(n17724), .ZN(n17726) );
  AOI222_X1 U19493 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17727), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17726), .C1(n17727), 
        .C2(n17726), .ZN(n17730) );
  OR2_X1 U19494 ( .A1(n17730), .A2(n12668), .ZN(n17729) );
  NAND2_X1 U19495 ( .A1(n17729), .A2(n17728), .ZN(n17732) );
  NAND2_X1 U19496 ( .A1(n17730), .A2(n12668), .ZN(n17731) );
  NAND2_X1 U19497 ( .A1(n17732), .A2(n17731), .ZN(n17741) );
  NOR2_X1 U19498 ( .A1(n17734), .A2(n17733), .ZN(n17737) );
  OAI21_X1 U19499 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n17735), .ZN(n17736) );
  NAND4_X1 U19500 ( .A1(n17739), .A2(n17738), .A3(n17737), .A4(n17736), .ZN(
        n17740) );
  AOI21_X1 U19501 ( .B1(n17741), .B2(n17748), .A(n17740), .ZN(n22235) );
  INV_X1 U19502 ( .A(n22235), .ZN(n17742) );
  AOI221_X1 U19503 ( .B1(n22225), .B2(n17744), .C1(n17742), .C2(n17744), .A(
        n17745), .ZN(n22227) );
  NOR2_X1 U19504 ( .A1(n22227), .A2(n22225), .ZN(n22226) );
  OAI211_X1 U19505 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n22253), .A(n22226), 
        .B(n17743), .ZN(n22231) );
  AOI22_X1 U19506 ( .A1(n17746), .A2(n17745), .B1(n17744), .B2(n22231), .ZN(
        P1_U3162) );
  NOR2_X1 U19507 ( .A1(n17748), .A2(n17747), .ZN(P1_U3032) );
  AND2_X1 U19508 ( .A1(n20393), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AOI21_X1 U19509 ( .B1(n17750), .B2(n17749), .A(n22805), .ZN(P1_U2802) );
  INV_X1 U19510 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17854) );
  OAI22_X1 U19511 ( .A1(n18968), .A2(n17854), .B1(n17752), .B2(n17751), .ZN(
        P2_U2816) );
  AOI22_X1 U19512 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19047), .B1(n17754), 
        .B2(n17753), .ZN(n17761) );
  NAND3_X1 U19513 ( .A1(n15556), .A2(n17755), .A3(n17782), .ZN(n17756) );
  OAI21_X1 U19514 ( .B1(n17773), .B2(n17757), .A(n17756), .ZN(n17758) );
  AOI21_X1 U19515 ( .B1(n17759), .B2(n17785), .A(n17758), .ZN(n17760) );
  OAI211_X1 U19516 ( .C1(n17763), .C2(n17762), .A(n17761), .B(n17760), .ZN(
        P2_U3011) );
  AOI22_X1 U19517 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17780), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19040), .ZN(n17768) );
  AOI222_X1 U19518 ( .A1(n17766), .A2(n17785), .B1(n17784), .B2(n17765), .C1(
        n17764), .C2(n17782), .ZN(n17767) );
  OAI211_X1 U19519 ( .C1(n17790), .C2(n17769), .A(n17768), .B(n17767), .ZN(
        P2_U3010) );
  AOI22_X1 U19520 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17780), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19040), .ZN(n17779) );
  NOR3_X1 U19521 ( .A1(n17612), .A2(n17771), .A3(n17770), .ZN(n17777) );
  OAI22_X1 U19522 ( .A1(n17775), .A2(n17774), .B1(n17773), .B2(n17772), .ZN(
        n17776) );
  NOR2_X1 U19523 ( .A1(n17777), .A2(n17776), .ZN(n17778) );
  OAI211_X1 U19524 ( .C1(n17790), .C2(n18988), .A(n17779), .B(n17778), .ZN(
        P2_U3008) );
  AOI22_X1 U19525 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17780), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19040), .ZN(n17788) );
  AOI222_X1 U19526 ( .A1(n17786), .A2(n17785), .B1(n17784), .B2(n17783), .C1(
        n17782), .C2(n17781), .ZN(n17787) );
  OAI211_X1 U19527 ( .C1(n17790), .C2(n17789), .A(n17788), .B(n17787), .ZN(
        P2_U3006) );
  INV_X1 U19528 ( .A(n17809), .ZN(n17811) );
  NAND3_X1 U19529 ( .A1(n17791), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n17792) );
  OAI21_X1 U19530 ( .B1(n19732), .B2(n18965), .A(n17792), .ZN(n17793) );
  AOI21_X1 U19531 ( .B1(n19891), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17793), 
        .ZN(n17794) );
  OAI22_X1 U19532 ( .A1(n19891), .A2(n17809), .B1(n17811), .B2(n17794), .ZN(
        P2_U3605) );
  AND2_X1 U19533 ( .A1(n19745), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19723) );
  NAND2_X1 U19534 ( .A1(n17805), .A2(n19723), .ZN(n19862) );
  OR2_X1 U19535 ( .A1(n19723), .A2(n19908), .ZN(n17800) );
  NAND2_X1 U19536 ( .A1(n17800), .A2(n19196), .ZN(n17807) );
  AOI22_X1 U19537 ( .A1(n17807), .A2(n19845), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n17795), .ZN(n17796) );
  OAI21_X1 U19538 ( .B1(n19862), .B2(n19908), .A(n17796), .ZN(n17797) );
  INV_X1 U19539 ( .A(n17797), .ZN(n17798) );
  AOI22_X1 U19540 ( .A1(n17811), .A2(n19766), .B1(n17798), .B2(n17809), .ZN(
        P2_U3603) );
  NAND2_X1 U19541 ( .A1(n17799), .A2(n22239), .ZN(n17802) );
  INV_X1 U19542 ( .A(n17800), .ZN(n17801) );
  AOI222_X1 U19543 ( .A1(n17803), .A2(n19745), .B1(n17802), .B2(n17801), .C1(
        n20168), .C2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17804) );
  AOI22_X1 U19544 ( .A1(n17811), .A2(n19889), .B1(n17804), .B2(n17809), .ZN(
        P2_U3604) );
  NAND2_X1 U19545 ( .A1(n19824), .A2(n19723), .ZN(n19814) );
  NAND2_X1 U19546 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19790), .ZN(n19776) );
  NAND2_X1 U19547 ( .A1(n19814), .A2(n19776), .ZN(n17808) );
  INV_X1 U19548 ( .A(n17806), .ZN(n20070) );
  AOI222_X1 U19549 ( .A1(n17808), .A2(n19880), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20070), .C1(n17807), .C2(n19863), .ZN(n17810) );
  AOI22_X1 U19550 ( .A1(n17811), .A2(n19777), .B1(n17810), .B2(n17809), .ZN(
        P2_U3602) );
  INV_X1 U19551 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22241) );
  NAND2_X1 U19552 ( .A1(n17812), .A2(n22241), .ZN(n17815) );
  INV_X1 U19553 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n17857) );
  OAI21_X1 U19554 ( .B1(n17857), .B2(n13343), .A(n17819), .ZN(n17813) );
  OAI21_X1 U19555 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17819), .A(n17813), 
        .ZN(n17814) );
  OAI221_X1 U19556 ( .B1(n17815), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17815), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17814), .ZN(P2_U2822) );
  INV_X1 U19557 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17818) );
  OAI221_X1 U19558 ( .B1(n17819), .B2(n17818), .C1(n17817), .C2(n17816), .A(
        n17815), .ZN(P2_U2823) );
  OAI22_X1 U19559 ( .A1(n22278), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n17907), .ZN(n17820) );
  INV_X1 U19560 ( .A(n17820), .ZN(P2_U3611) );
  INV_X1 U19561 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17821) );
  AOI22_X1 U19562 ( .A1(n17907), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17821), 
        .B2(n22278), .ZN(P2_U3608) );
  AOI21_X1 U19563 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n22242), .ZN(n17822) );
  INV_X1 U19564 ( .A(n17822), .ZN(P2_U2815) );
  INV_X1 U19565 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n17825) );
  AOI22_X1 U19566 ( .A1(n17851), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17824) );
  OAI21_X1 U19567 ( .B1(n17825), .B2(n17853), .A(n17824), .ZN(P2_U2951) );
  INV_X1 U19568 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17827) );
  AOI22_X1 U19569 ( .A1(n17851), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17826) );
  OAI21_X1 U19570 ( .B1(n17827), .B2(n17853), .A(n17826), .ZN(P2_U2950) );
  INV_X1 U19571 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17829) );
  AOI22_X1 U19572 ( .A1(n17851), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17836), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17828) );
  OAI21_X1 U19573 ( .B1(n17829), .B2(n17853), .A(n17828), .ZN(P2_U2949) );
  INV_X1 U19574 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17831) );
  AOI22_X1 U19575 ( .A1(n17841), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17836), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17830) );
  OAI21_X1 U19576 ( .B1(n17831), .B2(n17853), .A(n17830), .ZN(P2_U2948) );
  INV_X1 U19577 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17833) );
  AOI22_X1 U19578 ( .A1(n17851), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17836), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17832) );
  OAI21_X1 U19579 ( .B1(n17833), .B2(n17853), .A(n17832), .ZN(P2_U2947) );
  INV_X1 U19580 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n17835) );
  AOI22_X1 U19581 ( .A1(n17841), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17836), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17834) );
  OAI21_X1 U19582 ( .B1(n17835), .B2(n17853), .A(n17834), .ZN(P2_U2946) );
  INV_X1 U19583 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19930) );
  AOI22_X1 U19584 ( .A1(n17841), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17836), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17837) );
  OAI21_X1 U19585 ( .B1(n19930), .B2(n17853), .A(n17837), .ZN(P2_U2945) );
  AOI22_X1 U19586 ( .A1(n17841), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17838) );
  OAI21_X1 U19587 ( .B1(n19715), .B2(n17853), .A(n17838), .ZN(P2_U2944) );
  INV_X1 U19588 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19713) );
  AOI22_X1 U19589 ( .A1(n17841), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17839) );
  OAI21_X1 U19590 ( .B1(n19713), .B2(n17853), .A(n17839), .ZN(P2_U2943) );
  INV_X1 U19591 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19709) );
  AOI22_X1 U19592 ( .A1(n17851), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17840) );
  OAI21_X1 U19593 ( .B1(n19709), .B2(n17853), .A(n17840), .ZN(P2_U2942) );
  AOI22_X1 U19594 ( .A1(n17841), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17842) );
  OAI21_X1 U19595 ( .B1(n17843), .B2(n17853), .A(n17842), .ZN(P2_U2941) );
  INV_X1 U19596 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19703) );
  AOI22_X1 U19597 ( .A1(n17851), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17844) );
  OAI21_X1 U19598 ( .B1(n19703), .B2(n17853), .A(n17844), .ZN(P2_U2940) );
  AOI22_X1 U19599 ( .A1(n17851), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17845) );
  OAI21_X1 U19600 ( .B1(n17846), .B2(n17853), .A(n17845), .ZN(P2_U2939) );
  INV_X1 U19601 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19697) );
  AOI22_X1 U19602 ( .A1(n17851), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17847) );
  OAI21_X1 U19603 ( .B1(n19697), .B2(n17853), .A(n17847), .ZN(P2_U2938) );
  AOI22_X1 U19604 ( .A1(n17851), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17848) );
  OAI21_X1 U19605 ( .B1(n17849), .B2(n17853), .A(n17848), .ZN(P2_U2937) );
  AOI22_X1 U19606 ( .A1(n17851), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17850), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17852) );
  OAI21_X1 U19607 ( .B1(n19691), .B2(n17853), .A(n17852), .ZN(P2_U2936) );
  INV_X1 U19608 ( .A(P2_D_C_N_REG_SCAN_IN), .ZN(n17856) );
  AOI21_X1 U19609 ( .B1(P2_STATE_REG_1__SCAN_IN), .B2(n17854), .A(n22273), 
        .ZN(n17855) );
  OAI22_X1 U19610 ( .A1(n17907), .A2(n17856), .B1(P2_STATE_REG_0__SCAN_IN), 
        .B2(n17855), .ZN(P2_U2817) );
  OAI222_X1 U19611 ( .A1(n17904), .A2(n17859), .B1(n17858), .B2(n17907), .C1(
        n17857), .C2(n17900), .ZN(P2_U3212) );
  INV_X1 U19612 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n17860) );
  OAI222_X1 U19613 ( .A1(n17904), .A2(n17861), .B1(n17860), .B2(n17907), .C1(
        n17859), .C2(n17900), .ZN(P2_U3213) );
  INV_X1 U19614 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n17862) );
  OAI222_X1 U19615 ( .A1(n17904), .A2(n17863), .B1(n17862), .B2(n17907), .C1(
        n17861), .C2(n17900), .ZN(P2_U3214) );
  INV_X1 U19616 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n17864) );
  OAI222_X1 U19617 ( .A1(n17904), .A2(n18971), .B1(n17864), .B2(n17907), .C1(
        n17863), .C2(n17900), .ZN(P2_U3215) );
  INV_X1 U19618 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n17865) );
  OAI222_X1 U19619 ( .A1(n17904), .A2(n13185), .B1(n17865), .B2(n17907), .C1(
        n18971), .C2(n17900), .ZN(P2_U3216) );
  INV_X1 U19620 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n17866) );
  OAI222_X1 U19621 ( .A1(n17904), .A2(n18999), .B1(n17866), .B2(n17907), .C1(
        n13185), .C2(n17900), .ZN(P2_U3217) );
  INV_X1 U19622 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n17867) );
  OAI222_X1 U19623 ( .A1(n17904), .A2(n15841), .B1(n17867), .B2(n17907), .C1(
        n18999), .C2(n17900), .ZN(P2_U3218) );
  INV_X1 U19624 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n17868) );
  OAI222_X1 U19625 ( .A1(n17904), .A2(n13200), .B1(n17868), .B2(n17907), .C1(
        n15841), .C2(n17900), .ZN(P2_U3219) );
  INV_X1 U19626 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n17869) );
  OAI222_X1 U19627 ( .A1(n17900), .A2(n13200), .B1(n17869), .B2(n17907), .C1(
        n17308), .C2(n17904), .ZN(P2_U3220) );
  INV_X1 U19628 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n17870) );
  OAI222_X1 U19629 ( .A1(n17900), .A2(n17308), .B1(n17870), .B2(n17907), .C1(
        n17872), .C2(n17904), .ZN(P2_U3221) );
  INV_X1 U19630 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n17871) );
  OAI222_X1 U19631 ( .A1(n17900), .A2(n17872), .B1(n17871), .B2(n17907), .C1(
        n13531), .C2(n17904), .ZN(P2_U3222) );
  INV_X1 U19632 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n17873) );
  INV_X1 U19633 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19015) );
  OAI222_X1 U19634 ( .A1(n17900), .A2(n13531), .B1(n17873), .B2(n17907), .C1(
        n19015), .C2(n17904), .ZN(P2_U3223) );
  INV_X1 U19635 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n17874) );
  OAI222_X1 U19636 ( .A1(n17900), .A2(n19015), .B1(n17874), .B2(n17907), .C1(
        n13218), .C2(n17904), .ZN(P2_U3224) );
  INV_X1 U19637 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n17875) );
  OAI222_X1 U19638 ( .A1(n17900), .A2(n13218), .B1(n17875), .B2(n17907), .C1(
        n13224), .C2(n17904), .ZN(P2_U3225) );
  INV_X1 U19639 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n17876) );
  OAI222_X1 U19640 ( .A1(n17900), .A2(n13224), .B1(n17876), .B2(n17907), .C1(
        n17878), .C2(n17904), .ZN(P2_U3226) );
  INV_X1 U19641 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n17877) );
  OAI222_X1 U19642 ( .A1(n17900), .A2(n17878), .B1(n17877), .B2(n17907), .C1(
        n17880), .C2(n17904), .ZN(P2_U3227) );
  INV_X1 U19643 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n17879) );
  OAI222_X1 U19644 ( .A1(n17900), .A2(n17880), .B1(n17879), .B2(n17907), .C1(
        n13238), .C2(n17904), .ZN(P2_U3228) );
  INV_X1 U19645 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n17881) );
  OAI222_X1 U19646 ( .A1(n17904), .A2(n19070), .B1(n17881), .B2(n17907), .C1(
        n13238), .C2(n17900), .ZN(P2_U3229) );
  INV_X1 U19647 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n17882) );
  INV_X1 U19648 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n17883) );
  OAI222_X1 U19649 ( .A1(n17900), .A2(n19070), .B1(n17882), .B2(n17907), .C1(
        n17883), .C2(n17904), .ZN(P2_U3230) );
  INV_X1 U19650 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n17884) );
  OAI222_X1 U19651 ( .A1(n17904), .A2(n19083), .B1(n17884), .B2(n17907), .C1(
        n17883), .C2(n17900), .ZN(P2_U3231) );
  INV_X1 U19652 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n17885) );
  OAI222_X1 U19653 ( .A1(n17904), .A2(n13255), .B1(n17885), .B2(n17907), .C1(
        n19083), .C2(n17900), .ZN(P2_U3232) );
  INV_X1 U19654 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n17886) );
  OAI222_X1 U19655 ( .A1(n17904), .A2(n19110), .B1(n17886), .B2(n17907), .C1(
        n13255), .C2(n17900), .ZN(P2_U3233) );
  INV_X1 U19656 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n17887) );
  OAI222_X1 U19657 ( .A1(n17904), .A2(n17888), .B1(n17887), .B2(n17907), .C1(
        n19110), .C2(n17900), .ZN(P2_U3234) );
  INV_X1 U19658 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n17889) );
  OAI222_X1 U19659 ( .A1(n17904), .A2(n17891), .B1(n17889), .B2(n17907), .C1(
        n17888), .C2(n17900), .ZN(P2_U3235) );
  INV_X1 U19660 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n17890) );
  OAI222_X1 U19661 ( .A1(n17900), .A2(n17891), .B1(n17890), .B2(n17907), .C1(
        n17892), .C2(n17904), .ZN(P2_U3236) );
  INV_X1 U19662 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n17893) );
  OAI222_X1 U19663 ( .A1(n17904), .A2(n17895), .B1(n17893), .B2(n17907), .C1(
        n17892), .C2(n17900), .ZN(P2_U3237) );
  INV_X1 U19664 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n17894) );
  INV_X1 U19665 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n17897) );
  OAI222_X1 U19666 ( .A1(n17900), .A2(n17895), .B1(n17894), .B2(n17907), .C1(
        n17897), .C2(n17904), .ZN(P2_U3238) );
  INV_X1 U19667 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n17896) );
  OAI222_X1 U19668 ( .A1(n17900), .A2(n17897), .B1(n17896), .B2(n17907), .C1(
        n17899), .C2(n17904), .ZN(P2_U3239) );
  INV_X1 U19669 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n17898) );
  INV_X1 U19670 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n17901) );
  OAI222_X1 U19671 ( .A1(n17900), .A2(n17899), .B1(n17898), .B2(n17907), .C1(
        n17901), .C2(n17904), .ZN(P2_U3240) );
  INV_X1 U19672 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n17902) );
  OAI222_X1 U19673 ( .A1(n17904), .A2(n17903), .B1(n17902), .B2(n17907), .C1(
        n17901), .C2(n17900), .ZN(P2_U3241) );
  OAI22_X1 U19674 ( .A1(n22278), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n17907), .ZN(n17905) );
  INV_X1 U19675 ( .A(n17905), .ZN(P2_U3588) );
  OAI22_X1 U19676 ( .A1(n22278), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n17907), .ZN(n17906) );
  INV_X1 U19677 ( .A(n17906), .ZN(P2_U3587) );
  MUX2_X1 U19678 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n22278), .Z(P2_U3586) );
  OAI22_X1 U19679 ( .A1(n22278), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n17907), .ZN(n17908) );
  INV_X1 U19680 ( .A(n17908), .ZN(P2_U3585) );
  NOR2_X1 U19681 ( .A1(n17909), .A2(n18269), .ZN(n17933) );
  INV_X1 U19682 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20714) );
  NAND2_X1 U19683 ( .A1(n17910), .A2(n18270), .ZN(n17912) );
  NOR2_X1 U19684 ( .A1(n20714), .A2(n17912), .ZN(n17914) );
  AOI21_X1 U19685 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18268), .A(n17914), .ZN(
        n17911) );
  OAI22_X1 U19686 ( .A1(n17933), .A2(n17911), .B1(n19452), .B2(n18248), .ZN(
        P3_U2699) );
  INV_X1 U19687 ( .A(n17912), .ZN(n17916) );
  AOI21_X1 U19688 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18268), .A(n17916), .ZN(
        n17913) );
  INV_X1 U19689 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19494) );
  OAI22_X1 U19690 ( .A1(n17914), .A2(n17913), .B1(n19494), .B2(n18248), .ZN(
        P3_U2700) );
  OAI221_X1 U19691 ( .B1(n18267), .B2(n18265), .C1(n21219), .C2(n18265), .A(
        n20704), .ZN(n17915) );
  INV_X1 U19692 ( .A(n17915), .ZN(n17917) );
  AOI211_X1 U19693 ( .C1(n18271), .C2(n19534), .A(n17917), .B(n17916), .ZN(
        P3_U2701) );
  AOI22_X1 U19694 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17921) );
  AOI22_X1 U19695 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17920) );
  AOI22_X1 U19696 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17919) );
  AOI22_X1 U19697 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17918) );
  NAND4_X1 U19698 ( .A1(n17921), .A2(n17920), .A3(n17919), .A4(n17918), .ZN(
        n17927) );
  AOI22_X1 U19699 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17925) );
  AOI22_X1 U19700 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11160), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17924) );
  AOI22_X1 U19701 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17923) );
  AOI22_X1 U19702 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17922) );
  NAND4_X1 U19703 ( .A1(n17925), .A2(n17924), .A3(n17923), .A4(n17922), .ZN(
        n17926) );
  NOR2_X1 U19704 ( .A1(n17927), .A2(n17926), .ZN(n21293) );
  OAI21_X1 U19705 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17932), .A(n18033), .ZN(
        n17928) );
  AOI22_X1 U19706 ( .A1(n18271), .A2(n21293), .B1(n17928), .B2(n18268), .ZN(
        P3_U2695) );
  AOI21_X1 U19707 ( .B1(n20768), .B2(n17929), .A(n18271), .ZN(n17930) );
  INV_X1 U19708 ( .A(n17930), .ZN(n17931) );
  INV_X1 U19709 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19331) );
  OAI22_X1 U19710 ( .A1(n17932), .A2(n17931), .B1(n19331), .B2(n18248), .ZN(
        P3_U2696) );
  NAND2_X1 U19711 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17933), .ZN(n17936) );
  NAND3_X1 U19712 ( .A1(n17936), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n18268), .ZN(
        n17934) );
  OAI221_X1 U19713 ( .B1(n17936), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n18248), 
        .C2(n19371), .A(n17934), .ZN(P3_U2697) );
  AOI21_X1 U19714 ( .B1(n18273), .B2(n17935), .A(P3_EBX_REG_5__SCAN_IN), .ZN(
        n17938) );
  NAND2_X1 U19715 ( .A1(n18268), .A2(n17936), .ZN(n17937) );
  OAI22_X1 U19716 ( .A1(n17938), .A2(n17937), .B1(n19411), .B2(n18248), .ZN(
        P3_U2698) );
  INV_X1 U19717 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n20899) );
  NAND2_X1 U19718 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .ZN(n18038) );
  NOR2_X1 U19719 ( .A1(n18038), .A2(n17939), .ZN(n17963) );
  NAND2_X1 U19720 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17963), .ZN(n17950) );
  NAND2_X1 U19721 ( .A1(n18268), .A2(n17950), .ZN(n17964) );
  AOI22_X1 U19722 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17949) );
  AOI22_X1 U19723 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17948) );
  AOI22_X1 U19724 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17940) );
  OAI21_X1 U19725 ( .B1(n14959), .B2(n19686), .A(n17940), .ZN(n17946) );
  AOI22_X1 U19726 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17944) );
  AOI22_X1 U19727 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17943) );
  AOI22_X1 U19728 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17942) );
  AOI22_X1 U19729 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17941) );
  NAND4_X1 U19730 ( .A1(n17944), .A2(n17943), .A3(n17942), .A4(n17941), .ZN(
        n17945) );
  AOI211_X1 U19731 ( .C1(n11180), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n17946), .B(n17945), .ZN(n17947) );
  NAND3_X1 U19732 ( .A1(n17949), .A2(n17948), .A3(n17947), .ZN(n21269) );
  NOR3_X1 U19733 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n21179), .A3(n17950), .ZN(
        n17951) );
  AOI21_X1 U19734 ( .B1(n18271), .B2(n21269), .A(n17951), .ZN(n17952) );
  OAI21_X1 U19735 ( .B1(n20899), .B2(n17964), .A(n17952), .ZN(P3_U2687) );
  AOI22_X1 U19736 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17956) );
  AOI22_X1 U19737 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17955) );
  AOI22_X1 U19738 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17954) );
  AOI22_X1 U19739 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17953) );
  NAND4_X1 U19740 ( .A1(n17956), .A2(n17955), .A3(n17954), .A4(n17953), .ZN(
        n17962) );
  AOI22_X1 U19741 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11161), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17960) );
  AOI22_X1 U19742 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17959) );
  AOI22_X1 U19743 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17958) );
  AOI22_X1 U19744 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15006), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17957) );
  NAND4_X1 U19745 ( .A1(n17960), .A2(n17959), .A3(n17958), .A4(n17957), .ZN(
        n17961) );
  NOR2_X1 U19746 ( .A1(n17962), .A2(n17961), .ZN(n21286) );
  NOR2_X1 U19747 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17963), .ZN(n17965) );
  OAI22_X1 U19748 ( .A1(n21286), .A2(n18248), .B1(n17965), .B2(n17964), .ZN(
        P3_U2688) );
  INV_X1 U19749 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20853) );
  AOI22_X1 U19750 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17975) );
  AOI22_X1 U19751 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17974) );
  AOI22_X1 U19752 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17966) );
  OAI21_X1 U19753 ( .B1(n18010), .B2(n19411), .A(n17966), .ZN(n17972) );
  AOI22_X1 U19754 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17970) );
  AOI22_X1 U19755 ( .A1(n11160), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17969) );
  AOI22_X1 U19756 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17968) );
  AOI22_X1 U19757 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17967) );
  NAND4_X1 U19758 ( .A1(n17970), .A2(n17969), .A3(n17968), .A4(n17967), .ZN(
        n17971) );
  AOI211_X1 U19759 ( .C1(n11175), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n17972), .B(n17971), .ZN(n17973) );
  NAND3_X1 U19760 ( .A1(n17975), .A2(n17974), .A3(n17973), .ZN(n21123) );
  NAND2_X1 U19761 ( .A1(n18271), .A2(n21123), .ZN(n17976) );
  OAI221_X1 U19762 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17978), .C1(n20853), 
        .C2(n17977), .A(n17976), .ZN(P3_U2690) );
  AOI22_X1 U19763 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17983) );
  AOI22_X1 U19764 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17982) );
  AOI22_X1 U19765 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17981) );
  AOI22_X1 U19766 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17980) );
  NAND4_X1 U19767 ( .A1(n17983), .A2(n17982), .A3(n17981), .A4(n17980), .ZN(
        n17989) );
  AOI22_X1 U19768 ( .A1(n14985), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18323), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17987) );
  AOI22_X1 U19769 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17986) );
  AOI22_X1 U19770 ( .A1(n11160), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17985) );
  AOI22_X1 U19771 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15006), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17984) );
  NAND4_X1 U19772 ( .A1(n17987), .A2(n17986), .A3(n17985), .A4(n17984), .ZN(
        n17988) );
  NOR2_X1 U19773 ( .A1(n17989), .A2(n17988), .ZN(n21127) );
  NOR2_X1 U19774 ( .A1(n18271), .A2(n17990), .ZN(n18005) );
  NOR2_X1 U19775 ( .A1(n21179), .A2(n17991), .ZN(n17993) );
  INV_X1 U19776 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17992) );
  AOI22_X1 U19777 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18005), .B1(n17993), 
        .B2(n17992), .ZN(n17994) );
  OAI21_X1 U19778 ( .B1(n21127), .B2(n18268), .A(n17994), .ZN(P3_U2691) );
  AOI22_X1 U19779 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17998) );
  AOI22_X1 U19780 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11161), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17997) );
  AOI22_X1 U19781 ( .A1(n18321), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17996) );
  AOI22_X1 U19782 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17995) );
  NAND4_X1 U19783 ( .A1(n17998), .A2(n17997), .A3(n17996), .A4(n17995), .ZN(
        n18004) );
  AOI22_X1 U19784 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18002) );
  AOI22_X1 U19785 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18001) );
  AOI22_X1 U19786 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18000) );
  AOI22_X1 U19787 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18323), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17999) );
  NAND4_X1 U19788 ( .A1(n18002), .A2(n18001), .A3(n18000), .A4(n17999), .ZN(
        n18003) );
  NOR2_X1 U19789 ( .A1(n18004), .A2(n18003), .ZN(n21132) );
  OAI21_X1 U19790 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n18006), .A(n18005), .ZN(
        n18007) );
  OAI21_X1 U19791 ( .B1(n21132), .B2(n18268), .A(n18007), .ZN(P3_U2692) );
  NAND2_X1 U19792 ( .A1(n21219), .A2(n18008), .ZN(n18021) );
  NOR2_X1 U19793 ( .A1(n18271), .A2(n18008), .ZN(n18034) );
  AOI22_X1 U19794 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18019) );
  AOI22_X1 U19795 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18018) );
  AOI22_X1 U19796 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18009) );
  OAI21_X1 U19797 ( .B1(n18010), .B2(n19534), .A(n18009), .ZN(n18016) );
  AOI22_X1 U19798 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18014) );
  AOI22_X1 U19799 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18013) );
  AOI22_X1 U19800 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18012) );
  AOI22_X1 U19801 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18011) );
  NAND4_X1 U19802 ( .A1(n18014), .A2(n18013), .A3(n18012), .A4(n18011), .ZN(
        n18015) );
  AOI211_X1 U19803 ( .C1(n11173), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n18016), .B(n18015), .ZN(n18017) );
  NAND3_X1 U19804 ( .A1(n18019), .A2(n18018), .A3(n18017), .ZN(n21136) );
  AOI22_X1 U19805 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18034), .B1(n18271), 
        .B2(n21136), .ZN(n18020) );
  OAI21_X1 U19806 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18021), .A(n18020), .ZN(
        P3_U2693) );
  AOI22_X1 U19807 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n11170), .ZN(n18025) );
  AOI22_X1 U19808 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n15006), .ZN(n18024) );
  AOI22_X1 U19809 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18023) );
  AOI22_X1 U19810 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18324), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n11172), .ZN(n18022) );
  NAND4_X1 U19811 ( .A1(n18025), .A2(n18024), .A3(n18023), .A4(n18022), .ZN(
        n18032) );
  AOI22_X1 U19812 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18255), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n18348), .ZN(n18030) );
  AOI22_X1 U19813 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11160), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n11171), .ZN(n18029) );
  AOI22_X1 U19814 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18028) );
  AOI22_X1 U19815 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18027) );
  NAND4_X1 U19816 ( .A1(n18030), .A2(n18029), .A3(n18028), .A4(n18027), .ZN(
        n18031) );
  NOR2_X1 U19817 ( .A1(n18032), .A2(n18031), .ZN(n21143) );
  INV_X1 U19818 ( .A(n18033), .ZN(n18035) );
  OAI21_X1 U19819 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18035), .A(n18034), .ZN(
        n18036) );
  OAI21_X1 U19820 ( .B1(n21143), .B2(n18268), .A(n18036), .ZN(P3_U2694) );
  INV_X1 U19821 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21099) );
  INV_X1 U19822 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n18234) );
  INV_X1 U19823 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20913) );
  INV_X1 U19824 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20877) );
  NAND4_X1 U19825 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(P3_EBX_REG_9__SCAN_IN), .ZN(n18037)
         );
  NOR4_X1 U19826 ( .A1(n20899), .A2(n20877), .A3(n18038), .A4(n18037), .ZN(
        n18039) );
  NAND4_X1 U19827 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(n18040), .A4(n18039), .ZN(n18263) );
  NOR2_X1 U19828 ( .A1(n20913), .A2(n18263), .ZN(n18262) );
  NAND2_X1 U19829 ( .A1(n18273), .A2(n18262), .ZN(n18233) );
  NAND2_X1 U19830 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18247), .ZN(n18246) );
  INV_X1 U19831 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n21070) );
  INV_X1 U19832 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n18042) );
  INV_X1 U19833 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20961) );
  NAND4_X1 U19834 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(P3_EBX_REG_24__SCAN_IN), .ZN(n18041)
         );
  NOR4_X1 U19835 ( .A1(n21070), .A2(n18042), .A3(n20961), .A4(n18041), .ZN(
        n18043) );
  NAND4_X1 U19836 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n18145), .A4(n18043), .ZN(n18046) );
  NOR2_X1 U19837 ( .A1(n21099), .A2(n18046), .ZN(n18144) );
  NAND2_X1 U19838 ( .A1(n18268), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n18045) );
  NAND2_X1 U19839 ( .A1(n18144), .A2(n21219), .ZN(n18044) );
  OAI22_X1 U19840 ( .A1(n18144), .A2(n18045), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n18044), .ZN(P3_U2672) );
  NAND2_X1 U19841 ( .A1(n21099), .A2(n18046), .ZN(n18047) );
  NAND2_X1 U19842 ( .A1(n18047), .A2(n18268), .ZN(n18143) );
  AOI22_X1 U19843 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18048), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18052) );
  AOI22_X1 U19844 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18051) );
  AOI22_X1 U19845 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18050) );
  AOI22_X1 U19846 ( .A1(n18321), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18049) );
  NAND4_X1 U19847 ( .A1(n18052), .A2(n18051), .A3(n18050), .A4(n18049), .ZN(
        n18058) );
  AOI22_X1 U19848 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18056) );
  AOI22_X1 U19849 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18055) );
  AOI22_X1 U19850 ( .A1(n14985), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11161), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18054) );
  AOI22_X1 U19851 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18053) );
  NAND4_X1 U19852 ( .A1(n18056), .A2(n18055), .A3(n18054), .A4(n18053), .ZN(
        n18057) );
  NOR2_X1 U19853 ( .A1(n18058), .A2(n18057), .ZN(n18165) );
  AOI22_X1 U19854 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11161), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18062) );
  AOI22_X1 U19855 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18061) );
  AOI22_X1 U19856 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18060) );
  AOI22_X1 U19857 ( .A1(n18321), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18059) );
  NAND4_X1 U19858 ( .A1(n18062), .A2(n18061), .A3(n18060), .A4(n18059), .ZN(
        n18068) );
  AOI22_X1 U19859 ( .A1(n14985), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18066) );
  AOI22_X1 U19860 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18065) );
  AOI22_X1 U19861 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18064) );
  AOI22_X1 U19862 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18063) );
  NAND4_X1 U19863 ( .A1(n18066), .A2(n18065), .A3(n18064), .A4(n18063), .ZN(
        n18067) );
  NOR2_X1 U19864 ( .A1(n18068), .A2(n18067), .ZN(n18159) );
  AOI22_X1 U19865 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18072) );
  AOI22_X1 U19866 ( .A1(n14985), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18323), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18071) );
  AOI22_X1 U19867 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18070) );
  AOI22_X1 U19868 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18069) );
  NAND4_X1 U19869 ( .A1(n18072), .A2(n18071), .A3(n18070), .A4(n18069), .ZN(
        n18078) );
  AOI22_X1 U19870 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18076) );
  AOI22_X1 U19871 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18075) );
  AOI22_X1 U19872 ( .A1(n11161), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18074) );
  AOI22_X1 U19873 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18073) );
  NAND4_X1 U19874 ( .A1(n18076), .A2(n18075), .A3(n18074), .A4(n18073), .ZN(
        n18077) );
  NOR2_X1 U19875 ( .A1(n18078), .A2(n18077), .ZN(n18180) );
  AOI22_X1 U19876 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18082) );
  AOI22_X1 U19877 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18081) );
  AOI22_X1 U19878 ( .A1(n20722), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18080) );
  AOI22_X1 U19879 ( .A1(n11160), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18079) );
  NAND4_X1 U19880 ( .A1(n18082), .A2(n18081), .A3(n18080), .A4(n18079), .ZN(
        n18088) );
  AOI22_X1 U19881 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18086) );
  AOI22_X1 U19882 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18085) );
  AOI22_X1 U19883 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18084) );
  AOI22_X1 U19884 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14984), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18083) );
  NAND4_X1 U19885 ( .A1(n18086), .A2(n18085), .A3(n18084), .A4(n18083), .ZN(
        n18087) );
  NOR2_X1 U19886 ( .A1(n18088), .A2(n18087), .ZN(n18190) );
  AOI22_X1 U19887 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18092) );
  AOI22_X1 U19888 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18091) );
  AOI22_X1 U19889 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18090) );
  AOI22_X1 U19890 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18089) );
  NAND4_X1 U19891 ( .A1(n18092), .A2(n18091), .A3(n18090), .A4(n18089), .ZN(
        n18098) );
  AOI22_X1 U19892 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18096) );
  AOI22_X1 U19893 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18095) );
  AOI22_X1 U19894 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18094) );
  AOI22_X1 U19895 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18093) );
  NAND4_X1 U19896 ( .A1(n18096), .A2(n18095), .A3(n18094), .A4(n18093), .ZN(
        n18097) );
  NOR2_X1 U19897 ( .A1(n18098), .A2(n18097), .ZN(n18191) );
  NOR2_X1 U19898 ( .A1(n18190), .A2(n18191), .ZN(n18189) );
  AOI22_X1 U19899 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n11171), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18255), .ZN(n18109) );
  AOI22_X1 U19900 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n18366), .ZN(n18108) );
  INV_X1 U19901 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19580) );
  AOI22_X1 U19902 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18324), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18100) );
  OAI21_X1 U19903 ( .B1(n11852), .B2(n19580), .A(n18100), .ZN(n18106) );
  AOI22_X1 U19904 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n11170), .ZN(n18104) );
  AOI22_X1 U19905 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11167), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18103) );
  AOI22_X1 U19906 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18102) );
  AOI22_X1 U19907 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20722), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n11172), .ZN(n18101) );
  NAND4_X1 U19908 ( .A1(n18104), .A2(n18103), .A3(n18102), .A4(n18101), .ZN(
        n18105) );
  AOI211_X1 U19909 ( .C1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .C2(n11173), .A(
        n18106), .B(n18105), .ZN(n18107) );
  NAND3_X1 U19910 ( .A1(n18109), .A2(n18108), .A3(n18107), .ZN(n18185) );
  NAND2_X1 U19911 ( .A1(n18189), .A2(n18185), .ZN(n18184) );
  NOR2_X1 U19912 ( .A1(n18180), .A2(n18184), .ZN(n18179) );
  AOI22_X1 U19913 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18120) );
  AOI22_X1 U19914 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18119) );
  INV_X1 U19915 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18111) );
  AOI22_X1 U19916 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18110) );
  OAI21_X1 U19917 ( .B1(n18346), .B2(n18111), .A(n18110), .ZN(n18117) );
  AOI22_X1 U19918 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18115) );
  AOI22_X1 U19919 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18114) );
  AOI22_X1 U19920 ( .A1(n14985), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11160), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18113) );
  AOI22_X1 U19921 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18112) );
  NAND4_X1 U19922 ( .A1(n18115), .A2(n18114), .A3(n18113), .A4(n18112), .ZN(
        n18116) );
  AOI211_X1 U19923 ( .C1(n18323), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n18117), .B(n18116), .ZN(n18118) );
  NAND3_X1 U19924 ( .A1(n18120), .A2(n18119), .A3(n18118), .ZN(n18175) );
  NAND2_X1 U19925 ( .A1(n18179), .A2(n18175), .ZN(n18174) );
  NOR2_X1 U19926 ( .A1(n18159), .A2(n18174), .ZN(n18171) );
  AOI22_X1 U19927 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11160), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18131) );
  AOI22_X1 U19928 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18130) );
  AOI22_X1 U19929 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18121) );
  OAI21_X1 U19930 ( .B1(n11852), .B2(n19411), .A(n18121), .ZN(n18128) );
  AOI22_X1 U19931 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18126) );
  AOI22_X1 U19932 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18125) );
  AOI22_X1 U19933 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18124) );
  AOI22_X1 U19934 ( .A1(n18321), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18123) );
  NAND4_X1 U19935 ( .A1(n18126), .A2(n18125), .A3(n18124), .A4(n18123), .ZN(
        n18127) );
  AOI211_X1 U19936 ( .C1(n11174), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n18128), .B(n18127), .ZN(n18129) );
  NAND3_X1 U19937 ( .A1(n18131), .A2(n18130), .A3(n18129), .ZN(n18170) );
  NAND2_X1 U19938 ( .A1(n18171), .A2(n18170), .ZN(n18169) );
  NOR2_X1 U19939 ( .A1(n18165), .A2(n18169), .ZN(n18164) );
  AOI22_X1 U19940 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15006), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18135) );
  AOI22_X1 U19941 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18134) );
  AOI22_X1 U19942 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18133) );
  AOI22_X1 U19943 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18132) );
  NAND4_X1 U19944 ( .A1(n18135), .A2(n18134), .A3(n18133), .A4(n18132), .ZN(
        n18141) );
  AOI22_X1 U19945 ( .A1(n18323), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18139) );
  AOI22_X1 U19946 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18138) );
  AOI22_X1 U19947 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18137) );
  AOI22_X1 U19948 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18136) );
  NAND4_X1 U19949 ( .A1(n18139), .A2(n18138), .A3(n18137), .A4(n18136), .ZN(
        n18140) );
  NOR2_X1 U19950 ( .A1(n18141), .A2(n18140), .ZN(n18142) );
  XOR2_X1 U19951 ( .A(n18164), .B(n18142), .Z(n21232) );
  OAI22_X1 U19952 ( .A1(n18144), .A2(n18143), .B1(n21232), .B2(n18248), .ZN(
        P3_U2673) );
  NAND2_X1 U19953 ( .A1(n21219), .A2(n18145), .ZN(n18158) );
  NOR2_X1 U19954 ( .A1(n18271), .A2(n18145), .ZN(n18218) );
  AOI22_X1 U19955 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18149) );
  AOI22_X1 U19956 ( .A1(n18323), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15006), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18148) );
  AOI22_X1 U19957 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18147) );
  AOI22_X1 U19958 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18146) );
  NAND4_X1 U19959 ( .A1(n18149), .A2(n18148), .A3(n18147), .A4(n18146), .ZN(
        n18155) );
  AOI22_X1 U19960 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18153) );
  AOI22_X1 U19961 ( .A1(n11161), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18152) );
  AOI22_X1 U19962 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18151) );
  AOI22_X1 U19963 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18150) );
  NAND4_X1 U19964 ( .A1(n18153), .A2(n18152), .A3(n18151), .A4(n18150), .ZN(
        n18154) );
  NOR2_X1 U19965 ( .A1(n18155), .A2(n18154), .ZN(n21182) );
  INV_X1 U19966 ( .A(n21182), .ZN(n18156) );
  AOI22_X1 U19967 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18218), .B1(n18271), 
        .B2(n18156), .ZN(n18157) );
  OAI21_X1 U19968 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18158), .A(n18157), .ZN(
        P3_U2682) );
  INV_X1 U19969 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n21012) );
  INV_X1 U19970 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20989) );
  NOR2_X1 U19971 ( .A1(n20961), .A2(n18158), .ZN(n18195) );
  NAND2_X1 U19972 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18195), .ZN(n18188) );
  NAND2_X1 U19973 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n18194), .ZN(n18178) );
  NOR2_X1 U19974 ( .A1(n21012), .A2(n18178), .ZN(n18183) );
  NAND2_X1 U19975 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n18177), .ZN(n18173) );
  INV_X1 U19976 ( .A(n18173), .ZN(n18162) );
  AOI21_X1 U19977 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18268), .A(n18177), .ZN(
        n18161) );
  AOI21_X1 U19978 ( .B1(n18159), .B2(n18174), .A(n18171), .ZN(n21246) );
  INV_X1 U19979 ( .A(n21246), .ZN(n18160) );
  OAI22_X1 U19980 ( .A1(n18162), .A2(n18161), .B1(n18160), .B2(n18248), .ZN(
        P3_U2676) );
  NAND2_X1 U19981 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18162), .ZN(n18168) );
  NAND2_X1 U19982 ( .A1(n18268), .A2(n18173), .ZN(n18163) );
  OAI21_X1 U19983 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n18269), .A(n18163), .ZN(
        n18166) );
  AOI21_X1 U19984 ( .B1(n18165), .B2(n18169), .A(n18164), .ZN(n21237) );
  AOI22_X1 U19985 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n18166), .B1(n21237), 
        .B2(n18271), .ZN(n18167) );
  OAI21_X1 U19986 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n18168), .A(n18167), .ZN(
        P3_U2674) );
  OAI21_X1 U19987 ( .B1(n18171), .B2(n18170), .A(n18169), .ZN(n21245) );
  NAND3_X1 U19988 ( .A1(n18173), .A2(P3_EBX_REG_28__SCAN_IN), .A3(n18268), 
        .ZN(n18172) );
  OAI221_X1 U19989 ( .B1(n18173), .B2(P3_EBX_REG_28__SCAN_IN), .C1(n18248), 
        .C2(n21245), .A(n18172), .ZN(P3_U2675) );
  AOI21_X1 U19990 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18268), .A(n18183), .ZN(
        n18176) );
  OAI21_X1 U19991 ( .B1(n18179), .B2(n18175), .A(n18174), .ZN(n21228) );
  OAI22_X1 U19992 ( .A1(n18177), .A2(n18176), .B1(n21228), .B2(n18248), .ZN(
        P3_U2677) );
  INV_X1 U19993 ( .A(n18178), .ZN(n18187) );
  AOI21_X1 U19994 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18268), .A(n18187), .ZN(
        n18182) );
  AOI21_X1 U19995 ( .B1(n18180), .B2(n18184), .A(n18179), .ZN(n21216) );
  INV_X1 U19996 ( .A(n21216), .ZN(n18181) );
  OAI22_X1 U19997 ( .A1(n18183), .A2(n18182), .B1(n18181), .B2(n18248), .ZN(
        P3_U2678) );
  AOI21_X1 U19998 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18268), .A(n18194), .ZN(
        n18186) );
  OAI21_X1 U19999 ( .B1(n18189), .B2(n18185), .A(n18184), .ZN(n21260) );
  OAI22_X1 U20000 ( .A1(n18187), .A2(n18186), .B1(n21260), .B2(n18248), .ZN(
        P3_U2679) );
  INV_X1 U20001 ( .A(n18188), .ZN(n18207) );
  AOI21_X1 U20002 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18248), .A(n18207), .ZN(
        n18193) );
  AOI21_X1 U20003 ( .B1(n18191), .B2(n18190), .A(n18189), .ZN(n21261) );
  INV_X1 U20004 ( .A(n21261), .ZN(n18192) );
  OAI22_X1 U20005 ( .A1(n18194), .A2(n18193), .B1(n18248), .B2(n18192), .ZN(
        P3_U2680) );
  AOI21_X1 U20006 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18268), .A(n18195), .ZN(
        n18206) );
  AOI22_X1 U20007 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18199) );
  AOI22_X1 U20008 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18198) );
  AOI22_X1 U20009 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11160), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18197) );
  AOI22_X1 U20010 ( .A1(n18321), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18196) );
  NAND4_X1 U20011 ( .A1(n18199), .A2(n18198), .A3(n18197), .A4(n18196), .ZN(
        n18205) );
  AOI22_X1 U20012 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18203) );
  AOI22_X1 U20013 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18202) );
  AOI22_X1 U20014 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18323), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18201) );
  AOI22_X1 U20015 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18200) );
  NAND4_X1 U20016 ( .A1(n18203), .A2(n18202), .A3(n18201), .A4(n18200), .ZN(
        n18204) );
  NOR2_X1 U20017 ( .A1(n18205), .A2(n18204), .ZN(n21194) );
  OAI22_X1 U20018 ( .A1(n18207), .A2(n18206), .B1(n21194), .B2(n18248), .ZN(
        P3_U2681) );
  AOI22_X1 U20019 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18217) );
  AOI22_X1 U20020 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U20021 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18208) );
  OAI21_X1 U20022 ( .B1(n14959), .B2(n19452), .A(n18208), .ZN(n18214) );
  AOI22_X1 U20023 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18212) );
  AOI22_X1 U20024 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15006), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18211) );
  AOI22_X1 U20025 ( .A1(n11161), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18210) );
  AOI22_X1 U20026 ( .A1(n18323), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18209) );
  NAND4_X1 U20027 ( .A1(n18212), .A2(n18211), .A3(n18210), .A4(n18209), .ZN(
        n18213) );
  AOI211_X1 U20028 ( .C1(n11174), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n18214), .B(n18213), .ZN(n18215) );
  NAND3_X1 U20029 ( .A1(n18217), .A2(n18216), .A3(n18215), .ZN(n21186) );
  INV_X1 U20030 ( .A(n21186), .ZN(n18221) );
  OAI21_X1 U20031 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18219), .A(n18218), .ZN(
        n18220) );
  OAI21_X1 U20032 ( .B1(n18221), .B2(n18268), .A(n18220), .ZN(P3_U2683) );
  AOI22_X1 U20033 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18232) );
  AOI22_X1 U20034 ( .A1(n18323), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18231) );
  AOI22_X1 U20035 ( .A1(n18321), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18222) );
  OAI21_X1 U20036 ( .B1(n14959), .B2(n19534), .A(n18222), .ZN(n18229) );
  AOI22_X1 U20037 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18227) );
  AOI22_X1 U20038 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18226) );
  AOI22_X1 U20039 ( .A1(n11161), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18225) );
  AOI22_X1 U20040 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18224) );
  NAND4_X1 U20041 ( .A1(n18227), .A2(n18226), .A3(n18225), .A4(n18224), .ZN(
        n18228) );
  AOI211_X1 U20042 ( .C1(n14984), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n18229), .B(n18228), .ZN(n18230) );
  NAND3_X1 U20043 ( .A1(n18232), .A2(n18231), .A3(n18230), .ZN(n21204) );
  AOI21_X1 U20044 ( .B1(n18234), .B2(n18233), .A(n18247), .ZN(n18235) );
  MUX2_X1 U20045 ( .A(n21204), .B(n18235), .S(n18268), .Z(P3_U2685) );
  AOI22_X1 U20046 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18239) );
  AOI22_X1 U20047 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18238) );
  AOI22_X1 U20048 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U20049 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18236) );
  NAND4_X1 U20050 ( .A1(n18239), .A2(n18238), .A3(n18237), .A4(n18236), .ZN(
        n18245) );
  AOI22_X1 U20051 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18243) );
  AOI22_X1 U20052 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18242) );
  AOI22_X1 U20053 ( .A1(n18323), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18241) );
  AOI22_X1 U20054 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18240) );
  NAND4_X1 U20055 ( .A1(n18243), .A2(n18242), .A3(n18241), .A4(n18240), .ZN(
        n18244) );
  NOR2_X1 U20056 ( .A1(n18245), .A2(n18244), .ZN(n21203) );
  OAI21_X1 U20057 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18247), .A(n18246), .ZN(
        n18249) );
  AOI22_X1 U20058 ( .A1(n18271), .A2(n21203), .B1(n18249), .B2(n18248), .ZN(
        P3_U2684) );
  AOI22_X1 U20059 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18348), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n11170), .ZN(n18253) );
  AOI22_X1 U20060 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18252) );
  AOI22_X1 U20061 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18366), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n11172), .ZN(n18251) );
  AOI22_X1 U20062 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n20722), .ZN(n18250) );
  NAND4_X1 U20063 ( .A1(n18253), .A2(n18252), .A3(n18251), .A4(n18250), .ZN(
        n18261) );
  AOI22_X1 U20064 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18323), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18259) );
  AOI22_X1 U20065 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11163), .B1(
        n11160), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18258) );
  AOI22_X1 U20066 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U20067 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18256) );
  NAND4_X1 U20068 ( .A1(n18259), .A2(n18258), .A3(n18257), .A4(n18256), .ZN(
        n18260) );
  NOR2_X1 U20069 ( .A1(n18261), .A2(n18260), .ZN(n21215) );
  AOI211_X1 U20070 ( .C1(n20913), .C2(n18263), .A(n18262), .B(n18269), .ZN(
        n18264) );
  AOI21_X1 U20071 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18265), .A(n18264), .ZN(
        n18266) );
  OAI21_X1 U20072 ( .B1(n21215), .B2(n18268), .A(n18266), .ZN(P3_U2686) );
  OAI21_X1 U20073 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n18267), .ZN(n20688) );
  INV_X1 U20074 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20694) );
  OAI222_X1 U20075 ( .A1(n20688), .A2(n18269), .B1(n20694), .B2(n18273), .C1(
        n19580), .C2(n18268), .ZN(P3_U2702) );
  INV_X1 U20076 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n20695) );
  AOI22_X1 U20077 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18271), .B1(
        n18270), .B2(n20695), .ZN(n18272) );
  OAI21_X1 U20078 ( .B1(n18273), .B2(n20695), .A(n18272), .ZN(P3_U2703) );
  INV_X1 U20079 ( .A(n18274), .ZN(n18427) );
  OAI21_X1 U20080 ( .B1(n21798), .B2(n20639), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18275) );
  OAI21_X1 U20081 ( .B1(n18427), .B2(n21841), .A(n18275), .ZN(P3_U2634) );
  NOR2_X1 U20082 ( .A1(n20633), .A2(n18837), .ZN(n18279) );
  AOI21_X1 U20083 ( .B1(n21852), .B2(n18277), .A(n18276), .ZN(n21839) );
  NOR2_X1 U20084 ( .A1(n21839), .A2(n19251), .ZN(n18278) );
  OAI22_X1 U20085 ( .A1(n21806), .A2(n18279), .B1(n18837), .B2(n18278), .ZN(
        P3_U2863) );
  AOI22_X1 U20086 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18289) );
  AOI22_X1 U20087 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18288) );
  AOI22_X1 U20088 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18280) );
  OAI21_X1 U20089 ( .B1(n18346), .B2(n19331), .A(n18280), .ZN(n18286) );
  AOI22_X1 U20090 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18284) );
  AOI22_X1 U20091 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18283) );
  AOI22_X1 U20092 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18282) );
  AOI22_X1 U20093 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18281) );
  NAND4_X1 U20094 ( .A1(n18284), .A2(n18283), .A3(n18282), .A4(n18281), .ZN(
        n18285) );
  AOI211_X1 U20095 ( .C1(n18347), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n18286), .B(n18285), .ZN(n18287) );
  NAND3_X1 U20096 ( .A1(n18289), .A2(n18288), .A3(n18287), .ZN(n18400) );
  AOI22_X1 U20097 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18293) );
  AOI22_X1 U20098 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18292) );
  AOI22_X1 U20099 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18291) );
  AOI22_X1 U20100 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18290) );
  NAND4_X1 U20101 ( .A1(n18293), .A2(n18292), .A3(n18291), .A4(n18290), .ZN(
        n18299) );
  AOI22_X1 U20102 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18297) );
  AOI22_X1 U20103 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18296) );
  AOI22_X1 U20104 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18295) );
  AOI22_X1 U20105 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18294) );
  NAND4_X1 U20106 ( .A1(n18297), .A2(n18296), .A3(n18295), .A4(n18294), .ZN(
        n18298) );
  AOI22_X1 U20107 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18303) );
  AOI22_X1 U20108 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18302) );
  AOI22_X1 U20109 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18301) );
  AOI22_X1 U20110 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18300) );
  NAND4_X1 U20111 ( .A1(n18303), .A2(n18302), .A3(n18301), .A4(n18300), .ZN(
        n18309) );
  AOI22_X1 U20112 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18307) );
  AOI22_X1 U20113 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18335), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18306) );
  AOI22_X1 U20114 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18305) );
  AOI22_X1 U20115 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18304) );
  NAND4_X1 U20116 ( .A1(n18307), .A2(n18306), .A3(n18305), .A4(n18304), .ZN(
        n18308) );
  AOI22_X1 U20117 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18319) );
  AOI22_X1 U20118 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18318) );
  AOI22_X1 U20119 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18310) );
  OAI21_X1 U20120 ( .B1(n18346), .B2(n19534), .A(n18310), .ZN(n18316) );
  AOI22_X1 U20121 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18314) );
  AOI22_X1 U20122 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18313) );
  AOI22_X1 U20123 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18312) );
  AOI22_X1 U20124 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18323), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18311) );
  NAND4_X1 U20125 ( .A1(n18314), .A2(n18313), .A3(n18312), .A4(n18311), .ZN(
        n18315) );
  AOI211_X1 U20126 ( .C1(n11180), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n18316), .B(n18315), .ZN(n18317) );
  AOI22_X1 U20127 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n11163), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18333) );
  AOI22_X1 U20128 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18320), .B1(
        n11173), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18332) );
  AOI22_X1 U20129 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18321), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n18366), .ZN(n18322) );
  OAI21_X1 U20130 ( .B1(n19580), .B2(n18346), .A(n18322), .ZN(n18330) );
  AOI22_X1 U20131 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11161), .B1(
        n18323), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18328) );
  AOI22_X1 U20132 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18327) );
  AOI22_X1 U20133 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18324), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n11170), .ZN(n18326) );
  AOI22_X1 U20134 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n18348), .ZN(n18325) );
  NAND4_X1 U20135 ( .A1(n18328), .A2(n18327), .A3(n18326), .A4(n18325), .ZN(
        n18329) );
  AOI22_X1 U20136 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18344) );
  AOI22_X1 U20137 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18343) );
  AOI22_X1 U20138 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18334) );
  OAI21_X1 U20139 ( .B1(n18346), .B2(n19452), .A(n18334), .ZN(n18341) );
  AOI22_X1 U20140 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U20141 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18338) );
  AOI22_X1 U20142 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18337) );
  AOI22_X1 U20143 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18336) );
  NAND4_X1 U20144 ( .A1(n18339), .A2(n18338), .A3(n18337), .A4(n18336), .ZN(
        n18340) );
  AOI211_X1 U20145 ( .C1(n11167), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n18341), .B(n18340), .ZN(n18342) );
  NAND3_X1 U20146 ( .A1(n18344), .A2(n18343), .A3(n18342), .ZN(n21161) );
  NAND2_X1 U20147 ( .A1(n18359), .A2(n21161), .ZN(n18358) );
  AOI22_X1 U20148 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18366), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18357) );
  AOI22_X1 U20149 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18356) );
  AOI22_X1 U20150 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18345) );
  OAI21_X1 U20151 ( .B1(n18346), .B2(n19371), .A(n18345), .ZN(n18354) );
  AOI22_X1 U20152 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18352) );
  AOI22_X1 U20153 ( .A1(n11180), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18335), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18351) );
  AOI22_X1 U20154 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18350) );
  AOI22_X1 U20155 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18349) );
  NAND4_X1 U20156 ( .A1(n18352), .A2(n18351), .A3(n18350), .A4(n18349), .ZN(
        n18353) );
  AOI211_X1 U20157 ( .C1(n18254), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n18354), .B(n18353), .ZN(n18355) );
  NAND3_X1 U20158 ( .A1(n18357), .A2(n18356), .A3(n18355), .ZN(n21152) );
  XOR2_X1 U20159 ( .A(n21156), .B(n18358), .Z(n18383) );
  XOR2_X1 U20160 ( .A(n21161), .B(n18359), .Z(n18360) );
  NAND2_X1 U20161 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18360), .ZN(
        n18382) );
  XOR2_X1 U20162 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n18360), .Z(
        n18788) );
  NOR2_X1 U20163 ( .A1(n18361), .A2(n18412), .ZN(n18363) );
  NAND2_X1 U20164 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18365), .ZN(
        n18379) );
  NAND2_X1 U20165 ( .A1(n21301), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18378) );
  XNOR2_X1 U20166 ( .A(n18412), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18818) );
  AOI22_X1 U20167 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18370) );
  AOI22_X1 U20168 ( .A1(n18324), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18369) );
  AOI22_X1 U20169 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n20722), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18368) );
  AOI22_X1 U20170 ( .A1(n11173), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18367) );
  NAND4_X1 U20171 ( .A1(n18370), .A2(n18369), .A3(n18368), .A4(n18367), .ZN(
        n18377) );
  AOI22_X1 U20172 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18375) );
  AOI22_X1 U20173 ( .A1(n11167), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18348), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18374) );
  AOI22_X1 U20174 ( .A1(n18371), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U20175 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18372) );
  NAND4_X1 U20176 ( .A1(n18375), .A2(n18374), .A3(n18373), .A4(n18372), .ZN(
        n18376) );
  INV_X1 U20177 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21532) );
  NOR2_X1 U20178 ( .A1(n18826), .A2(n21532), .ZN(n18825) );
  NAND2_X1 U20179 ( .A1(n18818), .A2(n18825), .ZN(n18817) );
  NAND2_X1 U20180 ( .A1(n18378), .A2(n18817), .ZN(n18811) );
  NAND2_X1 U20181 ( .A1(n18812), .A2(n18811), .ZN(n18810) );
  NAND2_X1 U20182 ( .A1(n18379), .A2(n18810), .ZN(n18380) );
  NAND2_X1 U20183 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18380), .ZN(
        n18381) );
  INV_X1 U20184 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21443) );
  XNOR2_X1 U20185 ( .A(n21443), .B(n18380), .ZN(n18797) );
  XOR2_X1 U20186 ( .A(n21165), .B(n18408), .Z(n18796) );
  NAND2_X1 U20187 ( .A1(n18797), .A2(n18796), .ZN(n18795) );
  NAND2_X1 U20188 ( .A1(n18383), .A2(n18384), .ZN(n18385) );
  NAND2_X1 U20189 ( .A1(n18385), .A2(n18777), .ZN(n18765) );
  XOR2_X1 U20190 ( .A(n21152), .B(n18386), .Z(n18387) );
  XOR2_X1 U20191 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n18387), .Z(
        n18766) );
  NAND2_X1 U20192 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18387), .ZN(
        n18388) );
  AOI21_X1 U20193 ( .B1(n21655), .B2(n18389), .A(n18640), .ZN(n18391) );
  NAND2_X1 U20194 ( .A1(n18391), .A2(n18453), .ZN(n18392) );
  NAND2_X1 U20195 ( .A1(n21649), .A2(n18737), .ZN(n18698) );
  INV_X1 U20196 ( .A(n21826), .ZN(n21847) );
  OR2_X1 U20197 ( .A1(n20684), .A2(n18395), .ZN(n21319) );
  NAND2_X2 U20198 ( .A1(n21367), .A2(n21628), .ZN(n21795) );
  INV_X1 U20199 ( .A(n18397), .ZN(n18398) );
  AOI21_X1 U20200 ( .B1(n18399), .B2(n18398), .A(n21797), .ZN(n21794) );
  NOR2_X1 U20201 ( .A1(n21165), .A2(n18405), .ZN(n18416) );
  NAND2_X1 U20202 ( .A1(n18416), .A2(n21161), .ZN(n18403) );
  NOR2_X1 U20203 ( .A1(n21156), .A2(n18403), .ZN(n18402) );
  NAND2_X1 U20204 ( .A1(n18402), .A2(n21152), .ZN(n18401) );
  NOR2_X1 U20205 ( .A1(n21655), .A2(n18401), .ZN(n18425) );
  XOR2_X1 U20206 ( .A(n21655), .B(n18401), .Z(n18757) );
  XOR2_X1 U20207 ( .A(n21152), .B(n18402), .Z(n18419) );
  XOR2_X1 U20208 ( .A(n21156), .B(n18403), .Z(n18404) );
  NAND2_X1 U20209 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18404), .ZN(
        n18418) );
  XOR2_X1 U20210 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n18404), .Z(
        n18775) );
  XOR2_X1 U20211 ( .A(n21165), .B(n18405), .Z(n18406) );
  NAND2_X1 U20212 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18406), .ZN(
        n18414) );
  XOR2_X1 U20213 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18406), .Z(
        n18802) );
  OAI21_X1 U20214 ( .B1(n18826), .B2(n18408), .A(n18407), .ZN(n18409) );
  NAND2_X1 U20215 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18409), .ZN(
        n18413) );
  XNOR2_X1 U20216 ( .A(n18364), .B(n18409), .ZN(n18809) );
  AOI21_X1 U20217 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18412), .A(
        n11540), .ZN(n18411) );
  NOR2_X1 U20218 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18412), .ZN(
        n18410) );
  AOI221_X1 U20219 ( .B1(n11540), .B2(n18412), .C1(n18411), .C2(n21532), .A(
        n18410), .ZN(n18808) );
  NAND2_X1 U20220 ( .A1(n18809), .A2(n18808), .ZN(n18807) );
  NAND2_X1 U20221 ( .A1(n18413), .A2(n18807), .ZN(n18801) );
  NAND2_X1 U20222 ( .A1(n18802), .A2(n18801), .ZN(n18800) );
  NAND2_X1 U20223 ( .A1(n18414), .A2(n18800), .ZN(n18415) );
  NAND2_X1 U20224 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18415), .ZN(
        n18417) );
  INV_X1 U20225 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21444) );
  XNOR2_X1 U20226 ( .A(n21444), .B(n18415), .ZN(n18785) );
  XOR2_X1 U20227 ( .A(n21161), .B(n18416), .Z(n18784) );
  NAND2_X1 U20228 ( .A1(n18785), .A2(n18784), .ZN(n18783) );
  NAND2_X1 U20229 ( .A1(n18417), .A2(n18783), .ZN(n18774) );
  NAND2_X1 U20230 ( .A1(n18775), .A2(n18774), .ZN(n18773) );
  NAND2_X1 U20231 ( .A1(n18419), .A2(n18420), .ZN(n18421) );
  INV_X1 U20232 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21479) );
  NAND2_X1 U20233 ( .A1(n18425), .A2(n18422), .ZN(n18426) );
  INV_X1 U20234 ( .A(n18422), .ZN(n18424) );
  NAND2_X1 U20235 ( .A1(n18425), .A2(n18424), .ZN(n18423) );
  INV_X1 U20236 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21783) );
  INV_X1 U20237 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21762) );
  NOR2_X1 U20238 ( .A1(n21783), .A2(n21762), .ZN(n21493) );
  INV_X1 U20239 ( .A(n21493), .ZN(n21499) );
  INV_X1 U20240 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18707) );
  NOR2_X1 U20241 ( .A1(n21499), .A2(n18707), .ZN(n21488) );
  NAND2_X1 U20242 ( .A1(n21488), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n21508) );
  INV_X1 U20243 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21754) );
  NOR2_X1 U20244 ( .A1(n21508), .A2(n21754), .ZN(n21518) );
  NAND2_X1 U20245 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21518), .ZN(
        n21539) );
  INV_X1 U20246 ( .A(n18493), .ZN(n18673) );
  INV_X1 U20247 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21743) );
  INV_X1 U20248 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21738) );
  NOR2_X1 U20249 ( .A1(n21743), .A2(n21738), .ZN(n21719) );
  INV_X1 U20250 ( .A(n21719), .ZN(n21717) );
  INV_X1 U20251 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21529) );
  NAND2_X1 U20252 ( .A1(n21721), .A2(n21518), .ZN(n18691) );
  NOR2_X2 U20253 ( .A1(n21529), .A2(n18691), .ZN(n21542) );
  NAND2_X1 U20254 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21542), .ZN(
        n18494) );
  INV_X1 U20255 ( .A(n18494), .ZN(n21530) );
  INV_X1 U20256 ( .A(n18746), .ZN(n18645) );
  NOR2_X2 U20257 ( .A1(n21529), .A2(n18683), .ZN(n21546) );
  NAND2_X1 U20258 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21546), .ZN(
        n18495) );
  INV_X1 U20259 ( .A(n18495), .ZN(n21718) );
  OAI22_X1 U20260 ( .A1(n21530), .A2(n18645), .B1(n21718), .B2(n18832), .ZN(
        n18468) );
  AOI21_X1 U20261 ( .B1(n18673), .B2(n21717), .A(n18468), .ZN(n18678) );
  INV_X1 U20262 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18566) );
  INV_X1 U20263 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18740) );
  NOR2_X1 U20264 ( .A1(n18740), .A2(n18752), .ZN(n18739) );
  NAND2_X1 U20265 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20845) );
  NAND2_X1 U20266 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18461) );
  INV_X1 U20267 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20693) );
  NOR2_X1 U20268 ( .A1(n18429), .A2(n20693), .ZN(n18670) );
  AOI21_X4 U20269 ( .B1(n20633), .B2(n21841), .A(n21850), .ZN(n18815) );
  AOI21_X1 U20270 ( .B1(n18700), .B2(n18429), .A(n18815), .ZN(n18675) );
  OAI21_X1 U20271 ( .B1(n18670), .B2(n18827), .A(n18675), .ZN(n18445) );
  INV_X2 U20272 ( .A(n19584), .ZN(n19585) );
  AOI21_X1 U20273 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18671), .A(
        n19585), .ZN(n18471) );
  NOR3_X1 U20274 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18471), .A3(
        n18429), .ZN(n18446) );
  NOR2_X1 U20275 ( .A1(n18427), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18728) );
  INV_X1 U20276 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21735) );
  NAND3_X2 U20277 ( .A1(n22243), .A2(n18828), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18620) );
  INV_X1 U20278 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18428) );
  NAND2_X1 U20279 ( .A1(n11266), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18444) );
  OAI21_X1 U20280 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18670), .A(
        n18444), .ZN(n20924) );
  OAI22_X1 U20281 ( .A1(n11165), .A2(n21735), .B1(n18620), .B2(n20924), .ZN(
        n18430) );
  AOI211_X1 U20282 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18445), .A(
        n18446), .B(n18430), .ZN(n18441) );
  NAND2_X1 U20283 ( .A1(n21649), .A2(n18566), .ZN(n18523) );
  OAI21_X1 U20284 ( .B1(n21649), .B2(n18566), .A(n18523), .ZN(n18439) );
  NOR2_X1 U20285 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18713) );
  AND2_X1 U20286 ( .A1(n18713), .A2(n18707), .ZN(n18431) );
  NAND2_X1 U20287 ( .A1(n18432), .A2(n21754), .ZN(n18433) );
  NOR2_X2 U20288 ( .A1(n18475), .A2(n18433), .ZN(n18454) );
  NOR2_X1 U20289 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18434) );
  AOI21_X1 U20290 ( .B1(n18454), .B2(n18434), .A(n18640), .ZN(n18435) );
  INV_X1 U20291 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21545) );
  NOR2_X1 U20292 ( .A1(n21545), .A2(n21539), .ZN(n21382) );
  INV_X1 U20293 ( .A(n21382), .ZN(n21731) );
  NOR2_X1 U20294 ( .A1(n18492), .A2(n21717), .ZN(n18442) );
  INV_X1 U20295 ( .A(n18435), .ZN(n18438) );
  XOR2_X1 U20296 ( .A(n18439), .B(n11593), .Z(n21733) );
  NOR2_X1 U20297 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21717), .ZN(
        n21732) );
  AOI22_X1 U20298 ( .A1(n18745), .A2(n21733), .B1(n18673), .B2(n21732), .ZN(
        n18440) );
  OAI211_X1 U20299 ( .C1(n18678), .C2(n18566), .A(n18441), .B(n18440), .ZN(
        P3_U2812) );
  NAND2_X1 U20300 ( .A1(n21719), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n21383) );
  INV_X1 U20301 ( .A(n21383), .ZN(n21380) );
  NAND2_X1 U20302 ( .A1(n21380), .A2(n18673), .ZN(n18526) );
  INV_X1 U20303 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21706) );
  NAND3_X1 U20304 ( .A1(n21380), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n21530), .ZN(n21695) );
  NAND3_X1 U20305 ( .A1(n21380), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n21718), .ZN(n21698) );
  AOI22_X1 U20306 ( .A1(n18746), .A2(n21695), .B1(n18820), .B2(n21698), .ZN(
        n18530) );
  NAND3_X1 U20307 ( .A1(n18640), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18442), .ZN(n18524) );
  OAI21_X1 U20308 ( .B1(n11593), .B2(n18523), .A(n18524), .ZN(n18443) );
  XOR2_X1 U20309 ( .A(n18443), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n21703) );
  INV_X1 U20310 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18936) );
  NOR2_X1 U20311 ( .A1(n11165), .A2(n18936), .ZN(n21702) );
  INV_X1 U20312 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20928) );
  NOR2_X1 U20313 ( .A1(n18515), .A2(n20693), .ZN(n18497) );
  AOI21_X1 U20314 ( .B1(n20928), .B2(n18444), .A(n18497), .ZN(n20927) );
  OAI21_X1 U20315 ( .B1(n18446), .B2(n18445), .A(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18448) );
  INV_X1 U20316 ( .A(n18471), .ZN(n18630) );
  NAND3_X1 U20317 ( .A1(n11266), .A2(n20928), .A3(n18630), .ZN(n18447) );
  OAI211_X1 U20318 ( .C1(n11641), .C2(n18620), .A(n18448), .B(n18447), .ZN(
        n18449) );
  AOI211_X1 U20319 ( .C1(n18745), .C2(n21703), .A(n21702), .B(n18449), .ZN(
        n18450) );
  OAI221_X1 U20320 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18526), 
        .C1(n21706), .C2(n18530), .A(n18450), .ZN(P3_U2811) );
  NOR2_X1 U20321 ( .A1(n18451), .A2(n20693), .ZN(n18684) );
  AOI21_X1 U20322 ( .B1(n18700), .B2(n18451), .A(n18815), .ZN(n18688) );
  OAI21_X1 U20323 ( .B1(n18684), .B2(n18827), .A(n18688), .ZN(n18466) );
  INV_X1 U20324 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18457) );
  INV_X1 U20325 ( .A(n18684), .ZN(n18452) );
  NOR2_X1 U20326 ( .A1(n18457), .A2(n18452), .ZN(n20874) );
  AOI21_X1 U20327 ( .B1(n18457), .B2(n18452), .A(n20874), .ZN(n20876) );
  AOI22_X1 U20328 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18466), .B1(
        n18672), .B2(n20876), .ZN(n18460) );
  INV_X1 U20329 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21477) );
  NOR2_X1 U20330 ( .A1(n21477), .A2(n21479), .ZN(n21381) );
  AND3_X1 U20331 ( .A1(n18453), .A2(n18640), .A3(n21381), .ZN(n18722) );
  NAND2_X1 U20332 ( .A1(n21518), .A2(n18722), .ZN(n18692) );
  INV_X1 U20333 ( .A(n18698), .ZN(n18455) );
  NAND2_X1 U20334 ( .A1(n18455), .A2(n18454), .ZN(n18693) );
  AOI22_X1 U20335 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18692), .B1(
        n18693), .B2(n21529), .ZN(n18456) );
  XOR2_X1 U20336 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18456), .Z(
        n21538) );
  NOR2_X1 U20337 ( .A1(n18471), .A2(n18451), .ZN(n18462) );
  AOI22_X1 U20338 ( .A1(n18745), .A2(n21538), .B1(n18462), .B2(n18457), .ZN(
        n18459) );
  NAND2_X1 U20339 ( .A1(n18728), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n21547) );
  OAI21_X1 U20340 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n11252), .A(
        n18468), .ZN(n18458) );
  NAND4_X1 U20341 ( .A1(n18460), .A2(n18459), .A3(n21547), .A4(n18458), .ZN(
        P3_U2815) );
  NAND2_X1 U20342 ( .A1(n18674), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20914) );
  OAI21_X1 U20343 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20874), .A(
        n20914), .ZN(n20887) );
  OAI211_X1 U20344 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18462), .B(n18461), .ZN(n18464) );
  NAND2_X1 U20345 ( .A1(n21780), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18463) );
  OAI211_X1 U20346 ( .C1(n18620), .C2(n20887), .A(n18464), .B(n18463), .ZN(
        n18465) );
  AOI21_X1 U20347 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18466), .A(
        n18465), .ZN(n18470) );
  AOI22_X1 U20348 ( .A1(n18640), .A2(n21743), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21649), .ZN(n18467) );
  XNOR2_X1 U20349 ( .A(n18492), .B(n18467), .ZN(n21745) );
  AOI22_X1 U20350 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18468), .B1(
        n18745), .B2(n21745), .ZN(n18469) );
  OAI211_X1 U20351 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18493), .A(
        n18470), .B(n18469), .ZN(P3_U2814) );
  NAND2_X1 U20352 ( .A1(n21488), .A2(n18432), .ZN(n21517) );
  NOR2_X1 U20353 ( .A1(n18471), .A2(n18472), .ZN(n18481) );
  INV_X1 U20354 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20843) );
  NOR2_X1 U20355 ( .A1(n18472), .A2(n20693), .ZN(n18701) );
  INV_X1 U20356 ( .A(n18827), .ZN(n18535) );
  AOI21_X1 U20357 ( .B1(n18700), .B2(n18472), .A(n18535), .ZN(n18473) );
  OAI21_X1 U20358 ( .B1(n18701), .B2(n18473), .A(n18828), .ZN(n18484) );
  INV_X1 U20359 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20840) );
  NAND2_X1 U20360 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18701), .ZN(
        n20850) );
  OAI21_X1 U20361 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18701), .A(
        n20850), .ZN(n20838) );
  OAI22_X1 U20362 ( .A1(n11165), .A2(n20840), .B1(n18620), .B2(n20838), .ZN(
        n18474) );
  AOI221_X1 U20363 ( .B1(n18481), .B2(n20843), .C1(n18484), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18474), .ZN(n18479) );
  INV_X1 U20364 ( .A(n21491), .ZN(n21379) );
  NOR2_X1 U20365 ( .A1(n21508), .A2(n21379), .ZN(n21506) );
  NOR2_X1 U20366 ( .A1(n21489), .A2(n21508), .ZN(n21514) );
  OAI22_X1 U20367 ( .A1(n21506), .A2(n18832), .B1(n21514), .B2(n18645), .ZN(
        n18488) );
  NAND2_X1 U20368 ( .A1(n21649), .A2(n18475), .ZN(n18485) );
  OAI221_X1 U20369 ( .B1(n21649), .B2(n21488), .C1(n21649), .C2(n18476), .A(
        n18485), .ZN(n18477) );
  XOR2_X1 U20370 ( .A(n18432), .B(n18477), .Z(n21505) );
  AOI22_X1 U20371 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18488), .B1(
        n18745), .B2(n21505), .ZN(n18478) );
  OAI211_X1 U20372 ( .C1(n18733), .C2(n21517), .A(n18479), .B(n18478), .ZN(
        P3_U2818) );
  OR2_X1 U20373 ( .A1(n21508), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n21761) );
  INV_X1 U20374 ( .A(n20850), .ZN(n18480) );
  NAND2_X1 U20375 ( .A1(n18687), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18685) );
  OAI21_X1 U20376 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18480), .A(
        n18685), .ZN(n20848) );
  OAI211_X1 U20377 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18481), .B(n20845), .ZN(n18482) );
  NAND2_X1 U20378 ( .A1(n21780), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n21759) );
  OAI211_X1 U20379 ( .C1(n18620), .C2(n20848), .A(n18482), .B(n21759), .ZN(
        n18483) );
  AOI21_X1 U20380 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18484), .A(
        n18483), .ZN(n18490) );
  OAI22_X1 U20381 ( .A1(n18640), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n18708), .B2(n21508), .ZN(n18486) );
  NAND2_X1 U20382 ( .A1(n18486), .A2(n18485), .ZN(n18487) );
  XOR2_X1 U20383 ( .A(n18487), .B(n21754), .Z(n21758) );
  AOI22_X1 U20384 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18488), .B1(
        n18745), .B2(n21758), .ZN(n18489) );
  OAI211_X1 U20385 ( .C1(n18733), .C2(n21761), .A(n18490), .B(n18489), .ZN(
        P3_U2817) );
  INV_X1 U20386 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18565) );
  NOR2_X1 U20387 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18523), .ZN(
        n18491) );
  INV_X1 U20388 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21707) );
  NAND2_X1 U20389 ( .A1(n18491), .A2(n21707), .ZN(n18510) );
  NOR2_X1 U20390 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18510), .ZN(
        n18531) );
  NAND2_X1 U20391 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21392) );
  INV_X1 U20392 ( .A(n21392), .ZN(n21387) );
  NAND2_X1 U20393 ( .A1(n21387), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21551) );
  OR2_X1 U20394 ( .A1(n21383), .A2(n21551), .ZN(n18496) );
  NOR2_X1 U20395 ( .A1(n18496), .A2(n18492), .ZN(n18560) );
  INV_X1 U20396 ( .A(n18522), .ZN(n18563) );
  OAI21_X1 U20397 ( .B1(n18531), .B2(n18560), .A(n18563), .ZN(n18532) );
  XNOR2_X1 U20398 ( .A(n18565), .B(n18532), .ZN(n21556) );
  NOR2_X1 U20399 ( .A1(n18496), .A2(n18493), .ZN(n18572) );
  NOR2_X2 U20400 ( .A1(n18496), .A2(n18494), .ZN(n21388) );
  OAI22_X1 U20401 ( .A1(n21388), .A2(n18645), .B1(n21389), .B2(n18832), .ZN(
        n18512) );
  INV_X1 U20402 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18517) );
  INV_X1 U20403 ( .A(n18497), .ZN(n18516) );
  AOI21_X1 U20404 ( .B1(n18535), .B2(n18516), .A(n18815), .ZN(n18498) );
  OAI21_X1 U20405 ( .B1(n18499), .B2(n18791), .A(n18498), .ZN(n18521) );
  AOI21_X1 U20406 ( .B1(n18671), .B2(n18517), .A(n18521), .ZN(n18507) );
  INV_X1 U20407 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18503) );
  NAND3_X1 U20408 ( .A1(n18499), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18500) );
  NOR2_X1 U20409 ( .A1(n18534), .A2(n20693), .ZN(n18537) );
  AOI21_X1 U20410 ( .B1(n18503), .B2(n18500), .A(n18537), .ZN(n20970) );
  INV_X1 U20411 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20957) );
  NAND2_X1 U20412 ( .A1(n18499), .A2(n18630), .ZN(n18508) );
  AOI221_X1 U20413 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n18503), .C2(n20957), .A(
        n18508), .ZN(n18501) );
  AOI21_X1 U20414 ( .B1(n20970), .B2(n18672), .A(n18501), .ZN(n18502) );
  NAND2_X1 U20415 ( .A1(n21780), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21558) );
  OAI211_X1 U20416 ( .C1(n18507), .C2(n18503), .A(n18502), .B(n21558), .ZN(
        n18504) );
  AOI221_X1 U20417 ( .B1(n18572), .B2(n18565), .C1(n18512), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18504), .ZN(n18505) );
  OAI21_X1 U20418 ( .B1(n18682), .B2(n21556), .A(n18505), .ZN(P3_U2808) );
  INV_X1 U20419 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21554) );
  NAND2_X1 U20420 ( .A1(n21387), .A2(n21554), .ZN(n21398) );
  NAND2_X1 U20421 ( .A1(n18499), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18506) );
  XOR2_X1 U20422 ( .A(n20957), .B(n18506), .Z(n20956) );
  NAND2_X1 U20423 ( .A1(n21780), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n21396) );
  OAI221_X1 U20424 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18508), .C1(
        n20957), .C2(n18507), .A(n21396), .ZN(n18509) );
  AOI21_X1 U20425 ( .B1(n18672), .B2(n20956), .A(n18509), .ZN(n18514) );
  OAI22_X1 U20426 ( .A1(n21392), .A2(n18524), .B1(n11593), .B2(n18510), .ZN(
        n18511) );
  XNOR2_X1 U20427 ( .A(n21554), .B(n18511), .ZN(n21395) );
  AOI22_X1 U20428 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18512), .B1(
        n18745), .B2(n21395), .ZN(n18513) );
  OAI211_X1 U20429 ( .C1(n18526), .C2(n21398), .A(n18514), .B(n18513), .ZN(
        P3_U2809) );
  OAI21_X1 U20430 ( .B1(n18515), .B2(n19584), .A(n18517), .ZN(n18520) );
  INV_X1 U20431 ( .A(n18671), .ZN(n18518) );
  AOI22_X1 U20432 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18499), .B1(
        n18517), .B2(n18516), .ZN(n20943) );
  AOI21_X1 U20433 ( .B1(n18620), .B2(n18518), .A(n11642), .ZN(n18519) );
  INV_X1 U20434 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20950) );
  NOR2_X1 U20435 ( .A1(n11165), .A2(n20950), .ZN(n21711) );
  AOI211_X1 U20436 ( .C1(n18521), .C2(n18520), .A(n18519), .B(n21711), .ZN(
        n18529) );
  XOR2_X1 U20437 ( .A(n18525), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n21712) );
  INV_X1 U20438 ( .A(n18526), .ZN(n18624) );
  NAND2_X1 U20439 ( .A1(n21707), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21714) );
  INV_X1 U20440 ( .A(n21714), .ZN(n18527) );
  AOI22_X1 U20441 ( .A1(n18745), .A2(n21712), .B1(n18624), .B2(n18527), .ZN(
        n18528) );
  OAI211_X1 U20442 ( .C1(n18530), .C2(n21707), .A(n18529), .B(n18528), .ZN(
        P3_U2810) );
  INV_X1 U20443 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21679) );
  NAND2_X1 U20444 ( .A1(n18531), .A2(n18565), .ZN(n18562) );
  AOI221_X1 U20445 ( .B1(n21649), .B2(n18562), .C1(n18565), .C2(n18562), .A(
        n18532), .ZN(n18533) );
  XOR2_X1 U20446 ( .A(n21679), .B(n18533), .Z(n21685) );
  INV_X1 U20447 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20986) );
  NOR2_X1 U20448 ( .A1(n18555), .A2(n19584), .ZN(n18543) );
  INV_X1 U20449 ( .A(n18534), .ZN(n18542) );
  NAND2_X1 U20450 ( .A1(n21780), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n21683) );
  INV_X1 U20451 ( .A(n21683), .ZN(n18541) );
  INV_X1 U20452 ( .A(n18537), .ZN(n18536) );
  AOI211_X1 U20453 ( .C1(n18535), .C2(n18536), .A(n18815), .B(n18543), .ZN(
        n18553) );
  AND2_X1 U20454 ( .A1(n18555), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18577) );
  AOI21_X1 U20455 ( .B1(n20986), .B2(n18536), .A(n18577), .ZN(n20985) );
  NOR2_X1 U20456 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18518), .ZN(
        n18538) );
  AOI22_X1 U20457 ( .A1(n18672), .A2(n20985), .B1(n18538), .B2(n18537), .ZN(
        n18539) );
  OAI21_X1 U20458 ( .B1(n18553), .B2(n20986), .A(n18539), .ZN(n18540) );
  AOI211_X1 U20459 ( .C1(n18543), .C2(n18542), .A(n18541), .B(n18540), .ZN(
        n18551) );
  NOR2_X1 U20460 ( .A1(n21679), .A2(n18565), .ZN(n18544) );
  INV_X1 U20461 ( .A(n18544), .ZN(n18571) );
  NAND2_X1 U20462 ( .A1(n18544), .A2(n21388), .ZN(n21672) );
  NAND2_X1 U20463 ( .A1(n18746), .A2(n21672), .ZN(n18545) );
  OAI21_X1 U20464 ( .B1(n21676), .B2(n18832), .A(n18545), .ZN(n18573) );
  NAND2_X1 U20465 ( .A1(n18820), .A2(n18552), .ZN(n18547) );
  INV_X1 U20466 ( .A(n21388), .ZN(n18546) );
  OAI22_X1 U20467 ( .A1(n18548), .A2(n18547), .B1(n18546), .B2(n18545), .ZN(
        n18549) );
  AOI22_X1 U20468 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18573), .B1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18549), .ZN(n18550) );
  OAI211_X1 U20469 ( .C1(n18682), .C2(n21685), .A(n18551), .B(n18550), .ZN(
        P3_U2807) );
  INV_X1 U20470 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21562) );
  INV_X1 U20471 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21694) );
  XOR2_X1 U20472 ( .A(n21562), .B(n18588), .Z(n21568) );
  OAI21_X1 U20473 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18518), .A(
        n18553), .ZN(n18579) );
  INV_X1 U20474 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18556) );
  INV_X1 U20475 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18554) );
  NAND2_X1 U20476 ( .A1(n18555), .A2(n18630), .ZN(n18581) );
  AOI221_X1 U20477 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n18556), .C2(n18554), .A(
        n18581), .ZN(n18559) );
  INV_X1 U20478 ( .A(n11165), .ZN(n21780) );
  NAND2_X1 U20479 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18577), .ZN(
        n18576) );
  NOR2_X1 U20480 ( .A1(n18585), .A2(n20693), .ZN(n18619) );
  AOI21_X1 U20481 ( .B1(n18556), .B2(n18576), .A(n18619), .ZN(n21010) );
  AOI22_X1 U20482 ( .A1(n21780), .A2(P3_REIP_REG_25__SCAN_IN), .B1(n18672), 
        .B2(n21010), .ZN(n18557) );
  INV_X1 U20483 ( .A(n18557), .ZN(n18558) );
  AOI211_X1 U20484 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18579), .A(
        n18559), .B(n18558), .ZN(n18570) );
  NOR2_X1 U20485 ( .A1(n21694), .A2(n21672), .ZN(n18587) );
  XOR2_X1 U20486 ( .A(n18587), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n21569) );
  INV_X1 U20487 ( .A(n18560), .ZN(n18561) );
  OAI22_X1 U20488 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18562), .B1(
        n18561), .B2(n18571), .ZN(n18564) );
  NOR2_X1 U20489 ( .A1(n21551), .A2(n18565), .ZN(n21677) );
  NAND2_X1 U20490 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21677), .ZN(
        n18567) );
  OAI21_X1 U20491 ( .B1(n21649), .B2(n18614), .A(n18613), .ZN(n18568) );
  XOR2_X1 U20492 ( .A(n18568), .B(n21562), .Z(n21572) );
  AOI22_X1 U20493 ( .A1(n18746), .A2(n21569), .B1(n18745), .B2(n21572), .ZN(
        n18569) );
  OAI211_X1 U20494 ( .C1(n18832), .C2(n21568), .A(n18570), .B(n18569), .ZN(
        P3_U2805) );
  NOR2_X1 U20495 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18571), .ZN(
        n21688) );
  AOI22_X1 U20496 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18573), .B1(
        n21688), .B2(n18572), .ZN(n18584) );
  OAI21_X1 U20497 ( .B1(n18575), .B2(n21694), .A(n18574), .ZN(n21690) );
  OAI21_X1 U20498 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18577), .A(
        n18576), .ZN(n18578) );
  INV_X1 U20499 ( .A(n18578), .ZN(n21000) );
  AOI22_X1 U20500 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18579), .B1(
        n18672), .B2(n21000), .ZN(n18580) );
  NAND2_X1 U20501 ( .A1(n18728), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n21691) );
  OAI211_X1 U20502 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n18581), .A(
        n18580), .B(n21691), .ZN(n18582) );
  AOI21_X1 U20503 ( .B1(n21690), .B2(n18745), .A(n18582), .ZN(n18583) );
  NAND2_X1 U20504 ( .A1(n18584), .A2(n18583), .ZN(P3_U2806) );
  NAND2_X1 U20505 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18586) );
  NAND3_X1 U20506 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n21677), .ZN(n21563) );
  NOR2_X1 U20507 ( .A1(n18586), .A2(n21563), .ZN(n21604) );
  INV_X1 U20508 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21610) );
  NAND2_X1 U20509 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21610), .ZN(
        n21651) );
  INV_X1 U20510 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18617) );
  NOR2_X1 U20511 ( .A1(n18593), .A2(n20693), .ZN(n18604) );
  INV_X1 U20512 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n21050) );
  NOR2_X1 U20513 ( .A1(n18667), .A2(n20693), .ZN(n18633) );
  INV_X1 U20514 ( .A(n18633), .ZN(n18657) );
  OAI21_X1 U20515 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18604), .A(
        n18657), .ZN(n21066) );
  INV_X1 U20516 ( .A(n21066), .ZN(n21058) );
  INV_X1 U20517 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21598) );
  INV_X1 U20518 ( .A(n18586), .ZN(n18596) );
  NAND2_X1 U20519 ( .A1(n18596), .A2(n18587), .ZN(n18627) );
  INV_X1 U20520 ( .A(n18627), .ZN(n21590) );
  NAND2_X1 U20521 ( .A1(n18596), .A2(n18588), .ZN(n21576) );
  INV_X1 U20522 ( .A(n21576), .ZN(n18651) );
  OAI22_X1 U20523 ( .A1(n21590), .A2(n18645), .B1(n18651), .B2(n18832), .ZN(
        n18623) );
  NOR2_X1 U20524 ( .A1(n21598), .A2(n18623), .ZN(n18612) );
  AOI211_X1 U20525 ( .C1(n18645), .C2(n18832), .A(n18612), .B(n21610), .ZN(
        n18595) );
  NAND2_X1 U20526 ( .A1(n21050), .A2(n18630), .ZN(n18592) );
  NAND2_X1 U20527 ( .A1(n21780), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n21668) );
  AND3_X1 U20528 ( .A1(n11647), .A2(n18630), .A3(n18589), .ZN(n18605) );
  OAI22_X1 U20529 ( .A1(n18589), .A2(n18791), .B1(n18619), .B2(n18827), .ZN(
        n18590) );
  NOR2_X1 U20530 ( .A1(n18815), .A2(n18590), .ZN(n18616) );
  OAI21_X1 U20531 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18518), .A(
        n18616), .ZN(n18608) );
  OAI21_X1 U20532 ( .B1(n18605), .B2(n18608), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18591) );
  OAI211_X1 U20533 ( .C1(n18593), .C2(n18592), .A(n21668), .B(n18591), .ZN(
        n18594) );
  AOI211_X1 U20534 ( .C1(n18672), .C2(n21058), .A(n18595), .B(n18594), .ZN(
        n18603) );
  NOR2_X1 U20535 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18640), .ZN(
        n18637) );
  AOI21_X1 U20536 ( .B1(n18640), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18637), .ZN(n21665) );
  INV_X1 U20537 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21578) );
  AOI21_X1 U20538 ( .B1(n21578), .B2(n21562), .A(n18640), .ZN(n18597) );
  AND2_X2 U20539 ( .A1(n18599), .A2(n18598), .ZN(n18600) );
  OAI211_X1 U20540 ( .C1(n21665), .C2(n18601), .A(n18745), .B(n21647), .ZN(
        n18602) );
  OAI211_X1 U20541 ( .C1(n18649), .C2(n21651), .A(n18603), .B(n18602), .ZN(
        P3_U2802) );
  AND2_X1 U20542 ( .A1(n21598), .A2(n18649), .ZN(n18611) );
  NAND2_X1 U20543 ( .A1(n18589), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18618) );
  AOI21_X1 U20544 ( .B1(n11647), .B2(n18618), .A(n18604), .ZN(n21041) );
  INV_X1 U20545 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21035) );
  NOR2_X1 U20546 ( .A1(n11165), .A2(n21035), .ZN(n21595) );
  AOI211_X1 U20547 ( .C1(n18672), .C2(n21041), .A(n21595), .B(n18605), .ZN(
        n18610) );
  OAI21_X1 U20548 ( .B1(n18640), .B2(n18607), .A(n18606), .ZN(n21596) );
  AOI22_X1 U20549 ( .A1(n18745), .A2(n21596), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18608), .ZN(n18609) );
  OAI211_X1 U20550 ( .C1(n18612), .C2(n18611), .A(n18610), .B(n18609), .ZN(
        P3_U2803) );
  OAI221_X1 U20551 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21649), 
        .C1(n21562), .C2(n18614), .A(n18613), .ZN(n18615) );
  XOR2_X1 U20552 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n18615), .Z(
        n21587) );
  AOI221_X1 U20553 ( .B1(n18585), .B2(n18617), .C1(n19584), .C2(n18617), .A(
        n18616), .ZN(n18622) );
  OAI21_X1 U20554 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18619), .A(
        n18618), .ZN(n21029) );
  NAND2_X1 U20555 ( .A1(n21780), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n21585) );
  OAI221_X1 U20556 ( .B1(n21029), .B2(n18620), .C1(n21029), .C2(n18518), .A(
        n21585), .ZN(n18621) );
  AOI211_X1 U20557 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n18623), .A(
        n18622), .B(n18621), .ZN(n18626) );
  NOR2_X1 U20558 ( .A1(n21562), .A2(n21563), .ZN(n21581) );
  NAND3_X1 U20559 ( .A1(n18624), .A2(n21581), .A3(n21578), .ZN(n18625) );
  OAI211_X1 U20560 ( .C1(n21587), .C2(n18682), .A(n18626), .B(n18625), .ZN(
        P3_U2804) );
  INV_X1 U20561 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21646) );
  INV_X1 U20562 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21618) );
  INV_X1 U20563 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21630) );
  NOR2_X1 U20564 ( .A1(n21618), .A2(n21630), .ZN(n21637) );
  NAND2_X1 U20565 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21613) );
  NOR2_X1 U20566 ( .A1(n21613), .A2(n18627), .ZN(n21659) );
  NAND2_X1 U20567 ( .A1(n21637), .A2(n21659), .ZN(n18628) );
  XNOR2_X1 U20568 ( .A(n21646), .B(n18628), .ZN(n21643) );
  INV_X1 U20569 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n21097) );
  INV_X1 U20570 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21079) );
  NAND2_X1 U20571 ( .A1(n18656), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18629) );
  XOR2_X2 U20572 ( .A(n21097), .B(n18629), .Z(n21054) );
  NAND2_X1 U20573 ( .A1(n21780), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n21645) );
  INV_X1 U20574 ( .A(n21645), .ZN(n18636) );
  NAND2_X1 U20575 ( .A1(n18631), .A2(n18630), .ZN(n18648) );
  XNOR2_X1 U20576 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18634) );
  NOR2_X1 U20577 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18518), .ZN(
        n18663) );
  NAND2_X1 U20578 ( .A1(n19585), .A2(n18632), .ZN(n18666) );
  OAI211_X1 U20579 ( .C1(n18633), .C2(n18827), .A(n18828), .B(n18666), .ZN(
        n18655) );
  NOR2_X1 U20580 ( .A1(n18663), .A2(n18655), .ZN(n18647) );
  OAI22_X1 U20581 ( .A1(n18648), .A2(n18634), .B1(n18647), .B2(n21097), .ZN(
        n18635) );
  AOI211_X1 U20582 ( .C1(n21054), .C2(n18672), .A(n18636), .B(n18635), .ZN(
        n18644) );
  XNOR2_X1 U20583 ( .A(n18641), .B(n21646), .ZN(n21644) );
  NOR2_X1 U20584 ( .A1(n21613), .A2(n21576), .ZN(n21660) );
  NAND2_X1 U20585 ( .A1(n21637), .A2(n21660), .ZN(n18642) );
  XOR2_X1 U20586 ( .A(n18642), .B(n21646), .Z(n21640) );
  AOI22_X1 U20587 ( .A1(n18745), .A2(n21644), .B1(n18820), .B2(n21640), .ZN(
        n18643) );
  OAI211_X1 U20588 ( .C1(n21643), .C2(n18645), .A(n18644), .B(n18643), .ZN(
        P3_U2799) );
  AOI22_X1 U20589 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21664), .B1(
        n18658), .B2(n21618), .ZN(n18646) );
  XOR2_X1 U20590 ( .A(n21630), .B(n18646), .Z(n21636) );
  INV_X1 U20591 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n21083) );
  XNOR2_X1 U20592 ( .A(n18656), .B(n21083), .ZN(n21094) );
  INV_X1 U20593 ( .A(n11165), .ZN(n21537) );
  NAND2_X1 U20594 ( .A1(n21537), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n21635) );
  OAI221_X1 U20595 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18648), .C1(
        n21083), .C2(n18647), .A(n21635), .ZN(n18653) );
  NOR2_X1 U20596 ( .A1(n21613), .A2(n21618), .ZN(n21627) );
  INV_X1 U20597 ( .A(n21627), .ZN(n18650) );
  NAND2_X1 U20598 ( .A1(n21590), .A2(n21627), .ZN(n21600) );
  NAND2_X1 U20599 ( .A1(n18651), .A2(n21627), .ZN(n21599) );
  AOI22_X1 U20600 ( .A1(n18746), .A2(n21600), .B1(n18820), .B2(n21599), .ZN(
        n18661) );
  INV_X1 U20601 ( .A(n18661), .ZN(n18652) );
  OAI21_X1 U20602 ( .B1(n21636), .B2(n18682), .A(n18654), .ZN(P3_U2800) );
  AOI22_X1 U20603 ( .A1(n21780), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18655), .ZN(n18665) );
  AOI21_X1 U20604 ( .B1(n21079), .B2(n18657), .A(n18656), .ZN(n21069) );
  AOI211_X1 U20605 ( .C1(n21660), .C2(n18820), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n21659), .ZN(n18660) );
  OAI22_X1 U20606 ( .A1(n18661), .A2(n18660), .B1(n21621), .B2(n18682), .ZN(
        n18662) );
  AOI221_X1 U20607 ( .B1(n18672), .B2(n21069), .C1(n18663), .C2(n21069), .A(
        n18662), .ZN(n18664) );
  OAI211_X1 U20608 ( .C1(n18667), .C2(n18666), .A(n18665), .B(n18664), .ZN(
        P3_U2801) );
  AOI21_X1 U20609 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18669), .A(
        n18668), .ZN(n21742) );
  AOI21_X1 U20610 ( .B1(n11638), .B2(n20914), .A(n18670), .ZN(n20901) );
  NOR2_X2 U20611 ( .A1(n18672), .A2(n18671), .ZN(n18813) );
  INV_X1 U20612 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20907) );
  NOR2_X1 U20613 ( .A1(n11165), .A2(n20907), .ZN(n18680) );
  AOI21_X1 U20614 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18673), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18677) );
  AOI21_X1 U20615 ( .B1(n18674), .B2(n19585), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18676) );
  OAI22_X1 U20616 ( .A1(n18678), .A2(n18677), .B1(n18676), .B2(n18675), .ZN(
        n18679) );
  AOI211_X1 U20617 ( .C1(n20901), .C2(n18821), .A(n18680), .B(n18679), .ZN(
        n18681) );
  OAI21_X1 U20618 ( .B1(n21742), .B2(n18682), .A(n18681), .ZN(P3_U2813) );
  AOI21_X1 U20619 ( .B1(n21529), .B2(n18683), .A(n21546), .ZN(n21520) );
  INV_X1 U20620 ( .A(n21520), .ZN(n18697) );
  INV_X1 U20621 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18686) );
  AOI21_X1 U20622 ( .B1(n18686), .B2(n18685), .A(n18684), .ZN(n20861) );
  AOI21_X1 U20623 ( .B1(n18687), .B2(n19585), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18689) );
  NAND2_X1 U20624 ( .A1(n21780), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n21527) );
  OAI21_X1 U20625 ( .B1(n18689), .B2(n18688), .A(n21527), .ZN(n18690) );
  AOI21_X1 U20626 ( .B1(n20861), .B2(n18821), .A(n18690), .ZN(n18696) );
  AOI21_X1 U20627 ( .B1(n21529), .B2(n18691), .A(n21542), .ZN(n21521) );
  NAND2_X1 U20628 ( .A1(n18693), .A2(n18692), .ZN(n18694) );
  XOR2_X1 U20629 ( .A(n18694), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n21525) );
  AOI22_X1 U20630 ( .A1(n18746), .A2(n21521), .B1(n18745), .B2(n21525), .ZN(
        n18695) );
  OAI211_X1 U20631 ( .C1(n18832), .C2(n18697), .A(n18696), .B(n18695), .ZN(
        P3_U2816) );
  AOI22_X1 U20632 ( .A1(n18820), .A2(n21379), .B1(n18746), .B2(n21489), .ZN(
        n18732) );
  NOR2_X1 U20633 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18698), .ZN(
        n18723) );
  AOI22_X1 U20634 ( .A1(n21493), .A2(n18722), .B1(n18713), .B2(n18723), .ZN(
        n18699) );
  XOR2_X1 U20635 ( .A(n18707), .B(n18699), .Z(n21501) );
  AOI211_X1 U20636 ( .C1(n21499), .C2(n18707), .A(n18733), .B(n21488), .ZN(
        n18705) );
  NAND2_X1 U20637 ( .A1(n20835), .A2(n19585), .ZN(n18716) );
  NOR2_X1 U20638 ( .A1(n18815), .A2(n18700), .ZN(n18769) );
  INV_X1 U20639 ( .A(n18769), .ZN(n18822) );
  NAND3_X1 U20640 ( .A1(n18822), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n18716), .ZN(n18703) );
  INV_X1 U20641 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20826) );
  NAND2_X1 U20642 ( .A1(n20835), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18714) );
  AOI21_X1 U20643 ( .B1(n20826), .B2(n18714), .A(n18701), .ZN(n20822) );
  AOI22_X1 U20644 ( .A1(n21780), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n20822), 
        .B2(n18821), .ZN(n18702) );
  OAI211_X1 U20645 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18716), .A(
        n18703), .B(n18702), .ZN(n18704) );
  AOI211_X1 U20646 ( .C1(n18745), .C2(n21501), .A(n18705), .B(n18704), .ZN(
        n18706) );
  OAI21_X1 U20647 ( .B1(n18732), .B2(n18707), .A(n18706), .ZN(P3_U2819) );
  INV_X1 U20648 ( .A(n18708), .ZN(n18710) );
  AOI21_X1 U20649 ( .B1(n21649), .B2(n21783), .A(n18722), .ZN(n18709) );
  AOI21_X1 U20650 ( .B1(n21783), .B2(n18710), .A(n18709), .ZN(n18712) );
  AOI221_X1 U20651 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18722), .C1(
        n21783), .C2(n18723), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18711) );
  AOI21_X1 U20652 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18712), .A(
        n18711), .ZN(n21763) );
  NOR3_X1 U20653 ( .A1(n21493), .A2(n18713), .A3(n18733), .ZN(n18720) );
  INV_X1 U20654 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20793) );
  NAND2_X1 U20655 ( .A1(n18750), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n20777) );
  NOR2_X1 U20656 ( .A1(n20693), .A2(n20777), .ZN(n18751) );
  NAND2_X1 U20657 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18751), .ZN(
        n20789) );
  NOR2_X1 U20658 ( .A1(n20793), .A2(n20789), .ZN(n20797) );
  OAI21_X1 U20659 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20797), .A(
        n18714), .ZN(n20808) );
  NAND4_X1 U20660 ( .A1(n18715), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18739), .A4(n19585), .ZN(n18726) );
  NOR2_X1 U20661 ( .A1(n20793), .A2(n18726), .ZN(n18725) );
  OAI211_X1 U20662 ( .C1(n18725), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18822), .B(n18716), .ZN(n18718) );
  NAND2_X1 U20663 ( .A1(n21537), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18717) );
  OAI211_X1 U20664 ( .C1(n18813), .C2(n20808), .A(n18718), .B(n18717), .ZN(
        n18719) );
  AOI211_X1 U20665 ( .C1(n21763), .C2(n18745), .A(n18720), .B(n18719), .ZN(
        n18721) );
  OAI21_X1 U20666 ( .B1(n18732), .B2(n21762), .A(n18721), .ZN(P3_U2820) );
  NOR2_X1 U20667 ( .A1(n18723), .A2(n18722), .ZN(n18724) );
  XOR2_X1 U20668 ( .A(n18724), .B(n21783), .Z(n21778) );
  AOI211_X1 U20669 ( .C1(n18726), .C2(n20793), .A(n18769), .B(n18725), .ZN(
        n18730) );
  AOI21_X1 U20670 ( .B1(n20793), .B2(n20789), .A(n20797), .ZN(n18727) );
  INV_X1 U20671 ( .A(n18727), .ZN(n20798) );
  INV_X1 U20672 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20811) );
  OAI22_X1 U20673 ( .A1(n18813), .A2(n20798), .B1(n11165), .B2(n20811), .ZN(
        n18729) );
  AOI211_X1 U20674 ( .C1(n18745), .C2(n21778), .A(n18730), .B(n18729), .ZN(
        n18731) );
  OAI221_X1 U20675 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18733), .C1(
        n21783), .C2(n18732), .A(n18731), .ZN(P3_U2821) );
  OAI21_X1 U20676 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18735), .A(
        n18734), .ZN(n21483) );
  AOI21_X1 U20677 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21649), .A(
        n18736), .ZN(n18738) );
  XOR2_X1 U20678 ( .A(n18738), .B(n18737), .Z(n21487) );
  INV_X1 U20679 ( .A(n21487), .ZN(n18744) );
  OAI21_X1 U20680 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18751), .A(
        n20789), .ZN(n20779) );
  OAI21_X1 U20681 ( .B1(n18750), .B2(n18791), .A(n18828), .ZN(n18759) );
  AOI211_X1 U20682 ( .C1(n18740), .C2(n20777), .A(n18739), .B(n19584), .ZN(
        n18741) );
  AOI21_X1 U20683 ( .B1(n18759), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n18741), .ZN(n18742) );
  NAND2_X1 U20684 ( .A1(n21780), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n21485) );
  OAI211_X1 U20685 ( .C1(n18813), .C2(n20779), .A(n18742), .B(n21485), .ZN(
        n18743) );
  AOI221_X1 U20686 ( .B1(n18746), .B2(n21487), .C1(n18745), .C2(n18744), .A(
        n18743), .ZN(n18747) );
  OAI21_X1 U20687 ( .B1(n18832), .B2(n21483), .A(n18747), .ZN(P3_U2822) );
  OAI21_X1 U20688 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18749), .A(
        n18748), .ZN(n21475) );
  NAND2_X1 U20689 ( .A1(n18750), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20750) );
  AOI21_X1 U20690 ( .B1(n18752), .B2(n20750), .A(n18751), .ZN(n20764) );
  NAND3_X1 U20691 ( .A1(n18715), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n19585), .ZN(n18753) );
  INV_X1 U20692 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n21470) );
  OAI22_X1 U20693 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18753), .B1(
        n11165), .B2(n21470), .ZN(n18754) );
  AOI21_X1 U20694 ( .B1(n20764), .B2(n18821), .A(n18754), .ZN(n18761) );
  AOI21_X1 U20695 ( .B1(n18757), .B2(n18756), .A(n18755), .ZN(n18758) );
  XOR2_X1 U20696 ( .A(n18758), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n21473) );
  AOI22_X1 U20697 ( .A1(n18820), .A2(n21473), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18759), .ZN(n18760) );
  OAI211_X1 U20698 ( .C1(n18831), .C2(n21475), .A(n18761), .B(n18760), .ZN(
        P3_U2823) );
  OAI21_X1 U20699 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18763), .A(
        n18762), .ZN(n21457) );
  NAND2_X1 U20700 ( .A1(n18715), .A2(n19585), .ZN(n18767) );
  OAI21_X1 U20701 ( .B1(n18766), .B2(n18765), .A(n18764), .ZN(n21459) );
  OAI22_X1 U20702 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18767), .B1(
        n18831), .B2(n21459), .ZN(n18768) );
  AOI21_X1 U20703 ( .B1(n18728), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18768), .ZN(
        n18772) );
  AOI21_X1 U20704 ( .B1(n19585), .B2(n18715), .A(n18769), .ZN(n18781) );
  NAND2_X1 U20705 ( .A1(n18715), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20757) );
  INV_X1 U20706 ( .A(n20757), .ZN(n18770) );
  OAI21_X1 U20707 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18770), .A(
        n20750), .ZN(n20756) );
  INV_X1 U20708 ( .A(n20756), .ZN(n20751) );
  AOI22_X1 U20709 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18781), .B1(
        n20751), .B2(n18821), .ZN(n18771) );
  OAI211_X1 U20710 ( .C1(n18832), .C2(n21457), .A(n18772), .B(n18771), .ZN(
        P3_U2824) );
  OAI21_X1 U20711 ( .B1(n18775), .B2(n18774), .A(n18773), .ZN(n21448) );
  OAI21_X1 U20712 ( .B1(n18815), .B2(n18776), .A(n20745), .ZN(n18780) );
  NOR2_X1 U20713 ( .A1(n18776), .A2(n20693), .ZN(n20719) );
  OAI21_X1 U20714 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20719), .A(
        n20757), .ZN(n20739) );
  OAI21_X1 U20715 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18778), .A(
        n18777), .ZN(n21454) );
  OAI22_X1 U20716 ( .A1(n18813), .A2(n20739), .B1(n18831), .B2(n21454), .ZN(
        n18779) );
  AOI21_X1 U20717 ( .B1(n18781), .B2(n18780), .A(n18779), .ZN(n18782) );
  NAND2_X1 U20718 ( .A1(n21537), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21452) );
  OAI211_X1 U20719 ( .C1(n18832), .C2(n21448), .A(n18782), .B(n21452), .ZN(
        P3_U2825) );
  OAI21_X1 U20720 ( .B1(n18785), .B2(n18784), .A(n18783), .ZN(n21436) );
  NAND2_X1 U20721 ( .A1(n18792), .A2(n19585), .ZN(n18789) );
  OAI21_X1 U20722 ( .B1(n18788), .B2(n18787), .A(n18786), .ZN(n21442) );
  OAI22_X1 U20723 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18789), .B1(
        n18831), .B2(n21442), .ZN(n18790) );
  AOI21_X1 U20724 ( .B1(n18728), .B2(P3_REIP_REG_4__SCAN_IN), .A(n18790), .ZN(
        n18794) );
  OAI21_X1 U20725 ( .B1(n18792), .B2(n18791), .A(n18828), .ZN(n18805) );
  INV_X1 U20726 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20724) );
  NAND2_X1 U20727 ( .A1(n18792), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20728) );
  AOI21_X1 U20728 ( .B1(n20724), .B2(n20728), .A(n20719), .ZN(n20730) );
  AOI22_X1 U20729 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18805), .B1(
        n20730), .B2(n18821), .ZN(n18793) );
  OAI211_X1 U20730 ( .C1(n18832), .C2(n21436), .A(n18794), .B(n18793), .ZN(
        P3_U2826) );
  OAI21_X1 U20731 ( .B1(n18797), .B2(n18796), .A(n18795), .ZN(n21430) );
  NOR2_X1 U20732 ( .A1(n18815), .A2(n18798), .ZN(n18804) );
  NOR2_X1 U20733 ( .A1(n18798), .A2(n20693), .ZN(n18799) );
  OAI21_X1 U20734 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18799), .A(
        n20728), .ZN(n20709) );
  OAI21_X1 U20735 ( .B1(n18802), .B2(n18801), .A(n18800), .ZN(n21429) );
  OAI22_X1 U20736 ( .A1(n18813), .A2(n20709), .B1(n18832), .B2(n21429), .ZN(
        n18803) );
  AOI221_X1 U20737 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18805), .C1(
        n18804), .C2(n18805), .A(n18803), .ZN(n18806) );
  NAND2_X1 U20738 ( .A1(n21537), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n21432) );
  OAI211_X1 U20739 ( .C1(n18831), .C2(n21430), .A(n18806), .B(n21432), .ZN(
        P3_U2827) );
  OAI21_X1 U20740 ( .B1(n18809), .B2(n18808), .A(n18807), .ZN(n21418) );
  AOI22_X1 U20741 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20693), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18798), .ZN(n20699) );
  OAI21_X1 U20742 ( .B1(n18812), .B2(n18811), .A(n18810), .ZN(n21415) );
  OAI22_X1 U20743 ( .A1(n18813), .A2(n20699), .B1(n18831), .B2(n21415), .ZN(
        n18814) );
  AOI221_X1 U20744 ( .B1(n18815), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19585), .C2(n18798), .A(n18814), .ZN(n18816) );
  NAND2_X1 U20745 ( .A1(n21537), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n21422) );
  OAI211_X1 U20746 ( .C1(n18832), .C2(n21418), .A(n18816), .B(n21422), .ZN(
        P3_U2828) );
  OAI21_X1 U20747 ( .B1(n18818), .B2(n18825), .A(n18817), .ZN(n21408) );
  NAND2_X1 U20748 ( .A1(n21532), .A2(n18826), .ZN(n18819) );
  XNOR2_X1 U20749 ( .A(n18819), .B(n18818), .ZN(n21409) );
  AOI22_X1 U20750 ( .A1(n21780), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18820), 
        .B2(n21409), .ZN(n18824) );
  AOI22_X1 U20751 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18822), .B1(
        n18821), .B2(n20693), .ZN(n18823) );
  OAI211_X1 U20752 ( .C1(n18831), .C2(n21408), .A(n18824), .B(n18823), .ZN(
        P3_U2829) );
  AOI21_X1 U20753 ( .B1(n18826), .B2(n21532), .A(n18825), .ZN(n21405) );
  INV_X1 U20754 ( .A(n21405), .ZN(n21404) );
  NAND3_X1 U20755 ( .A1(n21314), .A2(n18828), .A3(n18827), .ZN(n18829) );
  AOI22_X1 U20756 ( .A1(n21780), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18829), .ZN(n18830) );
  OAI221_X1 U20757 ( .B1(n21405), .B2(n18832), .C1(n21404), .C2(n18831), .A(
        n18830), .ZN(P3_U2830) );
  INV_X1 U20758 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21818) );
  NAND2_X1 U20759 ( .A1(n19249), .A2(n21818), .ZN(n19285) );
  INV_X1 U20760 ( .A(n19285), .ZN(n19278) );
  NAND2_X1 U20761 ( .A1(n21815), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19275) );
  NAND2_X1 U20762 ( .A1(n21818), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19293) );
  NAND2_X1 U20763 ( .A1(n19275), .A2(n19293), .ZN(n18833) );
  AOI22_X1 U20764 ( .A1(n19278), .A2(n18838), .B1(n18834), .B2(n18833), .ZN(
        n18835) );
  OAI21_X1 U20765 ( .B1(n18836), .B2(n21818), .A(n18835), .ZN(P3_U2866) );
  NOR3_X1 U20766 ( .A1(n19289), .A2(n19251), .A3(n18837), .ZN(n18840) );
  INV_X1 U20767 ( .A(n18838), .ZN(n18839) );
  AOI22_X1 U20768 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18840), .B1(
        n18839), .B2(n21809), .ZN(P3_U2864) );
  NOR4_X1 U20769 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18844) );
  NOR4_X1 U20770 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18843) );
  NOR4_X1 U20771 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18842) );
  NOR4_X1 U20772 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18841) );
  NAND4_X1 U20773 ( .A1(n18844), .A2(n18843), .A3(n18842), .A4(n18841), .ZN(
        n18850) );
  NOR4_X1 U20774 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18848) );
  AOI211_X1 U20775 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18847) );
  NOR4_X1 U20776 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18846) );
  NOR4_X1 U20777 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18845) );
  NAND4_X1 U20778 ( .A1(n18848), .A2(n18847), .A3(n18846), .A4(n18845), .ZN(
        n18849) );
  NOR2_X1 U20779 ( .A1(n18850), .A2(n18849), .ZN(n18855) );
  INV_X1 U20780 ( .A(n18855), .ZN(n18858) );
  NOR2_X1 U20781 ( .A1(n18858), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18857) );
  INV_X1 U20782 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n21399) );
  INV_X1 U20783 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18953) );
  AOI22_X1 U20784 ( .A1(n18857), .A2(n21399), .B1(n18858), .B2(n18953), .ZN(
        P3_U3293) );
  NOR2_X1 U20785 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18854) );
  AOI21_X1 U20786 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n21399), .A(n18854), 
        .ZN(n18853) );
  INV_X1 U20787 ( .A(n18857), .ZN(n18861) );
  NOR2_X1 U20788 ( .A1(n18858), .A2(n21399), .ZN(n18851) );
  AOI22_X1 U20789 ( .A1(P3_BYTEENABLE_REG_2__SCAN_IN), .A2(n18858), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n18851), .ZN(n18852) );
  OAI21_X1 U20790 ( .B1(n18853), .B2(n18861), .A(n18852), .ZN(P3_U3292) );
  NOR2_X1 U20791 ( .A1(n18855), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18856)
         );
  NAND3_X1 U20792 ( .A1(n18855), .A2(n18854), .A3(n21399), .ZN(n18859) );
  OAI21_X1 U20793 ( .B1(n18857), .B2(n18856), .A(n18859), .ZN(P3_U2638) );
  NAND2_X1 U20794 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n18858), .ZN(n18860) );
  OAI211_X1 U20795 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(n18861), .A(n18860), 
        .B(n18859), .ZN(P3_U2639) );
  INV_X1 U20796 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18954) );
  AOI22_X1 U20797 ( .A1(n22252), .A2(n18862), .B1(n18954), .B2(n22298), .ZN(
        P3_U3297) );
  OAI22_X1 U20798 ( .A1(n22298), .A2(n18863), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n22252), .ZN(n18864) );
  INV_X1 U20799 ( .A(n18864), .ZN(P3_U3294) );
  AOI22_X1 U20800 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n22298), .B1(n22247), .B2(
        n22249), .ZN(n18865) );
  OAI21_X1 U20801 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n22298), .A(n18865), 
        .ZN(P3_U2635) );
  AOI22_X1 U20802 ( .A1(n21785), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18866) );
  OAI21_X1 U20803 ( .B1(n11420), .B2(n18887), .A(n18866), .ZN(P3_U2767) );
  INV_X1 U20804 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n21296) );
  AOI22_X1 U20805 ( .A1(n21785), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18867) );
  OAI21_X1 U20806 ( .B1(n21296), .B2(n18887), .A(n18867), .ZN(P3_U2766) );
  INV_X1 U20807 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n21170) );
  AOI22_X1 U20808 ( .A1(n21785), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18868) );
  OAI21_X1 U20809 ( .B1(n21170), .B2(n18887), .A(n18868), .ZN(P3_U2765) );
  INV_X1 U20810 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18870) );
  AOI22_X1 U20811 ( .A1(n21785), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18903), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18869) );
  OAI21_X1 U20812 ( .B1(n18870), .B2(n18887), .A(n18869), .ZN(P3_U2764) );
  INV_X1 U20813 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21147) );
  AOI22_X1 U20814 ( .A1(n21785), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18903), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18871) );
  OAI21_X1 U20815 ( .B1(n21147), .B2(n18887), .A(n18871), .ZN(P3_U2763) );
  INV_X1 U20816 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18873) );
  AOI22_X1 U20817 ( .A1(n21785), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18903), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18872) );
  OAI21_X1 U20818 ( .B1(n18873), .B2(n18887), .A(n18872), .ZN(P3_U2762) );
  INV_X1 U20819 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n21148) );
  AOI22_X1 U20820 ( .A1(n21785), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18903), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18874) );
  OAI21_X1 U20821 ( .B1(n21148), .B2(n18887), .A(n18874), .ZN(P3_U2761) );
  INV_X1 U20822 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18876) );
  AOI22_X1 U20823 ( .A1(n21785), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18875) );
  OAI21_X1 U20824 ( .B1(n18876), .B2(n18887), .A(n18875), .ZN(P3_U2760) );
  INV_X1 U20825 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21287) );
  AOI22_X1 U20826 ( .A1(n21785), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18877) );
  OAI21_X1 U20827 ( .B1(n21287), .B2(n18887), .A(n18877), .ZN(P3_U2759) );
  INV_X1 U20828 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n21141) );
  AOI22_X1 U20829 ( .A1(n18901), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18878) );
  OAI21_X1 U20830 ( .B1(n21141), .B2(n18887), .A(n18878), .ZN(P3_U2758) );
  INV_X1 U20831 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18880) );
  AOI22_X1 U20832 ( .A1(n18901), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18879) );
  OAI21_X1 U20833 ( .B1(n18880), .B2(n18887), .A(n18879), .ZN(P3_U2757) );
  INV_X1 U20834 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n21130) );
  AOI22_X1 U20835 ( .A1(n18901), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18881) );
  OAI21_X1 U20836 ( .B1(n21130), .B2(n18887), .A(n18881), .ZN(P3_U2756) );
  INV_X1 U20837 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18883) );
  AOI22_X1 U20838 ( .A1(n18901), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18882) );
  OAI21_X1 U20839 ( .B1(n18883), .B2(n18887), .A(n18882), .ZN(P3_U2755) );
  INV_X1 U20840 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20674) );
  AOI22_X1 U20841 ( .A1(n18901), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18884) );
  OAI21_X1 U20842 ( .B1(n20674), .B2(n18887), .A(n18884), .ZN(P3_U2754) );
  INV_X1 U20843 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20676) );
  AOI22_X1 U20844 ( .A1(n18901), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18885) );
  OAI21_X1 U20845 ( .B1(n20676), .B2(n18887), .A(n18885), .ZN(P3_U2753) );
  INV_X1 U20846 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21282) );
  AOI22_X1 U20847 ( .A1(n18901), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18886) );
  OAI21_X1 U20848 ( .B1(n21282), .B2(n18887), .A(n18886), .ZN(P3_U2752) );
  INV_X1 U20849 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18890) );
  NAND2_X1 U20850 ( .A1(n18888), .A2(n21115), .ZN(n18913) );
  AOI22_X1 U20851 ( .A1(n18901), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18889) );
  OAI21_X1 U20852 ( .B1(n18890), .B2(n18913), .A(n18889), .ZN(P3_U2751) );
  INV_X1 U20853 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n21205) );
  AOI22_X1 U20854 ( .A1(n18901), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18891) );
  OAI21_X1 U20855 ( .B1(n21205), .B2(n18913), .A(n18891), .ZN(P3_U2750) );
  INV_X1 U20856 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n21207) );
  AOI22_X1 U20857 ( .A1(n18901), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18892) );
  OAI21_X1 U20858 ( .B1(n21207), .B2(n18913), .A(n18892), .ZN(P3_U2749) );
  INV_X1 U20859 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18894) );
  AOI22_X1 U20860 ( .A1(n21785), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18903), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18893) );
  OAI21_X1 U20861 ( .B1(n18894), .B2(n18913), .A(n18893), .ZN(P3_U2748) );
  INV_X1 U20862 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18896) );
  AOI22_X1 U20863 ( .A1(n21785), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18903), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18895) );
  OAI21_X1 U20864 ( .B1(n18896), .B2(n18913), .A(n18895), .ZN(P3_U2747) );
  INV_X1 U20865 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21185) );
  AOI22_X1 U20866 ( .A1(n21785), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18903), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18897) );
  OAI21_X1 U20867 ( .B1(n21185), .B2(n18913), .A(n18897), .ZN(P3_U2746) );
  INV_X1 U20868 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18899) );
  AOI22_X1 U20869 ( .A1(n21785), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18903), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18898) );
  OAI21_X1 U20870 ( .B1(n18899), .B2(n18913), .A(n18898), .ZN(P3_U2745) );
  INV_X1 U20871 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n21263) );
  AOI22_X1 U20872 ( .A1(n21785), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18903), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18900) );
  OAI21_X1 U20873 ( .B1(n21263), .B2(n18913), .A(n18900), .ZN(P3_U2744) );
  INV_X1 U20874 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n21255) );
  AOI22_X1 U20875 ( .A1(n18901), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18902) );
  OAI21_X1 U20876 ( .B1(n21255), .B2(n18913), .A(n18902), .ZN(P3_U2743) );
  INV_X1 U20877 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n21220) );
  AOI22_X1 U20878 ( .A1(n21785), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18903), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18904) );
  OAI21_X1 U20879 ( .B1(n21220), .B2(n18913), .A(n18904), .ZN(P3_U2742) );
  INV_X1 U20880 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18906) );
  AOI22_X1 U20881 ( .A1(n21785), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18905) );
  OAI21_X1 U20882 ( .B1(n18906), .B2(n18913), .A(n18905), .ZN(P3_U2741) );
  INV_X1 U20883 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n21248) );
  AOI22_X1 U20884 ( .A1(n21785), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18907) );
  OAI21_X1 U20885 ( .B1(n21248), .B2(n18913), .A(n18907), .ZN(P3_U2740) );
  INV_X1 U20886 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18909) );
  AOI22_X1 U20887 ( .A1(n21785), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18908) );
  OAI21_X1 U20888 ( .B1(n18909), .B2(n18913), .A(n18908), .ZN(P3_U2739) );
  INV_X1 U20889 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20654) );
  AOI22_X1 U20890 ( .A1(n21785), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18910) );
  OAI21_X1 U20891 ( .B1(n20654), .B2(n18913), .A(n18910), .ZN(P3_U2738) );
  INV_X1 U20892 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n21236) );
  AOI22_X1 U20893 ( .A1(n21785), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18911), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18912) );
  OAI21_X1 U20894 ( .B1(n21236), .B2(n18913), .A(n18912), .ZN(P3_U2737) );
  NOR2_X1 U20895 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18914), .ZN(n18915) );
  NOR2_X1 U20896 ( .A1(n22252), .A2(n18915), .ZN(P3_U2633) );
  INV_X1 U20897 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18917) );
  INV_X1 U20898 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n22300) );
  NAND2_X1 U20899 ( .A1(n22300), .A2(n22252), .ZN(n18951) );
  INV_X1 U20900 ( .A(n18951), .ZN(n18946) );
  AOI22_X1 U20901 ( .A1(n18946), .A2(P3_REIP_REG_2__SCAN_IN), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n22298), .ZN(n18916) );
  OAI21_X1 U20902 ( .B1(n18948), .B2(n18917), .A(n18916), .ZN(P3_U3032) );
  INV_X1 U20903 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20705) );
  AOI22_X1 U20904 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18949), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n22298), .ZN(n18918) );
  OAI21_X1 U20905 ( .B1(n20705), .B2(n18951), .A(n18918), .ZN(P3_U3033) );
  AOI22_X1 U20906 ( .A1(n18946), .A2(P3_REIP_REG_4__SCAN_IN), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n22298), .ZN(n18919) );
  OAI21_X1 U20907 ( .B1(n18948), .B2(n20705), .A(n18919), .ZN(P3_U3034) );
  INV_X1 U20908 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20736) );
  AOI22_X1 U20909 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18949), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n22298), .ZN(n18920) );
  OAI21_X1 U20910 ( .B1(n20736), .B2(n18951), .A(n18920), .ZN(P3_U3035) );
  AOI22_X1 U20911 ( .A1(n18946), .A2(P3_REIP_REG_6__SCAN_IN), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n22298), .ZN(n18921) );
  OAI21_X1 U20912 ( .B1(n18948), .B2(n20736), .A(n18921), .ZN(P3_U3036) );
  AOI22_X1 U20913 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18949), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n22298), .ZN(n18922) );
  OAI21_X1 U20914 ( .B1(n21470), .B2(n18951), .A(n18922), .ZN(P3_U3037) );
  AOI22_X1 U20915 ( .A1(n18946), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n22298), .ZN(n18923) );
  OAI21_X1 U20916 ( .B1(n18948), .B2(n21470), .A(n18923), .ZN(P3_U3038) );
  INV_X1 U20917 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20792) );
  AOI22_X1 U20918 ( .A1(n18946), .A2(P3_REIP_REG_9__SCAN_IN), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n22298), .ZN(n18924) );
  OAI21_X1 U20919 ( .B1(n18948), .B2(n20792), .A(n18924), .ZN(P3_U3039) );
  AOI22_X1 U20920 ( .A1(n18946), .A2(P3_REIP_REG_10__SCAN_IN), .B1(
        P3_ADDRESS_REG_8__SCAN_IN), .B2(n22298), .ZN(n18925) );
  OAI21_X1 U20921 ( .B1(n18948), .B2(n20811), .A(n18925), .ZN(P3_U3040) );
  INV_X1 U20922 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n21503) );
  AOI22_X1 U20923 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18949), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n22298), .ZN(n18926) );
  OAI21_X1 U20924 ( .B1(n21503), .B2(n18951), .A(n18926), .ZN(P3_U3041) );
  AOI22_X1 U20925 ( .A1(n18946), .A2(P3_REIP_REG_12__SCAN_IN), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n22298), .ZN(n18927) );
  OAI21_X1 U20926 ( .B1(n18948), .B2(n21503), .A(n18927), .ZN(P3_U3042) );
  AOI22_X1 U20927 ( .A1(n18946), .A2(P3_REIP_REG_13__SCAN_IN), .B1(
        P3_ADDRESS_REG_11__SCAN_IN), .B2(n22298), .ZN(n18928) );
  OAI21_X1 U20928 ( .B1(n18948), .B2(n20840), .A(n18928), .ZN(P3_U3043) );
  INV_X1 U20929 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20865) );
  AOI22_X1 U20930 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n18949), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n22298), .ZN(n18929) );
  OAI21_X1 U20931 ( .B1(n20865), .B2(n18951), .A(n18929), .ZN(P3_U3044) );
  AOI22_X1 U20932 ( .A1(n18946), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n22298), .ZN(n18930) );
  OAI21_X1 U20933 ( .B1(n18948), .B2(n20865), .A(n18930), .ZN(P3_U3045) );
  INV_X1 U20934 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20884) );
  AOI22_X1 U20935 ( .A1(n18946), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(n22298), .ZN(n18931) );
  OAI21_X1 U20936 ( .B1(n18948), .B2(n20884), .A(n18931), .ZN(P3_U3046) );
  INV_X1 U20937 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n21751) );
  AOI22_X1 U20938 ( .A1(n18946), .A2(P3_REIP_REG_17__SCAN_IN), .B1(
        P3_ADDRESS_REG_15__SCAN_IN), .B2(n22298), .ZN(n18932) );
  OAI21_X1 U20939 ( .B1(n18948), .B2(n21751), .A(n18932), .ZN(P3_U3047) );
  AOI22_X1 U20940 ( .A1(n18946), .A2(P3_REIP_REG_18__SCAN_IN), .B1(
        P3_ADDRESS_REG_16__SCAN_IN), .B2(n22298), .ZN(n18933) );
  OAI21_X1 U20941 ( .B1(n18948), .B2(n20907), .A(n18933), .ZN(P3_U3048) );
  AOI22_X1 U20942 ( .A1(n18946), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_ADDRESS_REG_17__SCAN_IN), .B2(n22298), .ZN(n18934) );
  OAI21_X1 U20943 ( .B1(n18948), .B2(n21735), .A(n18934), .ZN(P3_U3049) );
  AOI22_X1 U20944 ( .A1(n18946), .A2(P3_REIP_REG_20__SCAN_IN), .B1(
        P3_ADDRESS_REG_18__SCAN_IN), .B2(n22298), .ZN(n18935) );
  OAI21_X1 U20945 ( .B1(n18948), .B2(n18936), .A(n18935), .ZN(P3_U3050) );
  AOI22_X1 U20946 ( .A1(n18946), .A2(P3_REIP_REG_21__SCAN_IN), .B1(
        P3_ADDRESS_REG_19__SCAN_IN), .B2(n22298), .ZN(n18937) );
  OAI21_X1 U20947 ( .B1(n18948), .B2(n20950), .A(n18937), .ZN(P3_U3051) );
  INV_X1 U20948 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20966) );
  AOI22_X1 U20949 ( .A1(n18946), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(n22298), .ZN(n18938) );
  OAI21_X1 U20950 ( .B1(n18948), .B2(n20966), .A(n18938), .ZN(P3_U3052) );
  INV_X1 U20951 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20977) );
  AOI22_X1 U20952 ( .A1(n18946), .A2(P3_REIP_REG_23__SCAN_IN), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n22298), .ZN(n18939) );
  OAI21_X1 U20953 ( .B1(n18948), .B2(n20977), .A(n18939), .ZN(P3_U3053) );
  INV_X1 U20954 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n21006) );
  AOI22_X1 U20955 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n18949), .B1(
        P3_ADDRESS_REG_22__SCAN_IN), .B2(n22298), .ZN(n18940) );
  OAI21_X1 U20956 ( .B1(n21006), .B2(n18951), .A(n18940), .ZN(P3_U3054) );
  AOI22_X1 U20957 ( .A1(n18946), .A2(P3_REIP_REG_25__SCAN_IN), .B1(
        P3_ADDRESS_REG_23__SCAN_IN), .B2(n22298), .ZN(n18941) );
  OAI21_X1 U20958 ( .B1(n18948), .B2(n21006), .A(n18941), .ZN(P3_U3055) );
  INV_X1 U20959 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21021) );
  AOI22_X1 U20960 ( .A1(n18946), .A2(P3_REIP_REG_26__SCAN_IN), .B1(
        P3_ADDRESS_REG_24__SCAN_IN), .B2(n22298), .ZN(n18942) );
  OAI21_X1 U20961 ( .B1(n18948), .B2(n21021), .A(n18942), .ZN(P3_U3056) );
  INV_X1 U20962 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21033) );
  AOI22_X1 U20963 ( .A1(n18946), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_ADDRESS_REG_25__SCAN_IN), .B2(n22298), .ZN(n18943) );
  OAI21_X1 U20964 ( .B1(n18948), .B2(n21033), .A(n18943), .ZN(P3_U3057) );
  AOI22_X1 U20965 ( .A1(n18946), .A2(P3_REIP_REG_28__SCAN_IN), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n22298), .ZN(n18944) );
  OAI21_X1 U20966 ( .B1(n18948), .B2(n21035), .A(n18944), .ZN(P3_U3058) );
  INV_X1 U20967 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21065) );
  AOI22_X1 U20968 ( .A1(n18946), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n22298), .ZN(n18945) );
  OAI21_X1 U20969 ( .B1(n18948), .B2(n21065), .A(n18945), .ZN(P3_U3059) );
  INV_X1 U20970 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21076) );
  AOI22_X1 U20971 ( .A1(n18946), .A2(P3_REIP_REG_30__SCAN_IN), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(n22298), .ZN(n18947) );
  OAI21_X1 U20972 ( .B1(n18948), .B2(n21076), .A(n18947), .ZN(P3_U3060) );
  INV_X1 U20973 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n21091) );
  AOI22_X1 U20974 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18949), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n22298), .ZN(n18950) );
  OAI21_X1 U20975 ( .B1(n21091), .B2(n18951), .A(n18950), .ZN(P3_U3061) );
  INV_X1 U20976 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18952) );
  AOI22_X1 U20977 ( .A1(n22252), .A2(n18953), .B1(n18952), .B2(n22298), .ZN(
        P3_U3277) );
  MUX2_X1 U20978 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .B(P3_BE_N_REG_1__SCAN_IN), .S(n22298), .Z(P3_U3276) );
  MUX2_X1 U20979 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .B(P3_BE_N_REG_2__SCAN_IN), .S(n22298), .Z(P3_U3275) );
  MUX2_X1 U20980 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .B(P3_BE_N_REG_3__SCAN_IN), .S(n22298), .Z(P3_U3274) );
  NOR4_X1 U20981 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18956)
         );
  NOR4_X1 U20982 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18954), .ZN(n18955) );
  NAND3_X1 U20983 ( .A1(n18956), .A2(n18955), .A3(U215), .ZN(U213) );
  NAND2_X1 U20984 ( .A1(n19213), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n18964) );
  INV_X1 U20985 ( .A(n18964), .ZN(n18962) );
  INV_X1 U20986 ( .A(n18957), .ZN(n22283) );
  OAI21_X1 U20987 ( .B1(n22283), .B2(n22239), .A(n18958), .ZN(n18960) );
  NAND3_X1 U20988 ( .A1(n22283), .A2(n20237), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18959) );
  MUX2_X1 U20989 ( .A(n18960), .B(n18959), .S(n11178), .Z(n18961) );
  OAI21_X1 U20990 ( .B1(n18962), .B2(n19214), .A(n18961), .ZN(n18970) );
  OAI22_X1 U20991 ( .A1(n18966), .A2(n18965), .B1(n18964), .B2(n18963), .ZN(
        n18967) );
  NOR2_X1 U20992 ( .A1(n18968), .A2(n18967), .ZN(n18969) );
  MUX2_X1 U20993 ( .A(n18970), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n18969), 
        .Z(P2_U3610) );
  OAI21_X1 U20994 ( .B1(n18971), .B2(n19111), .A(n19068), .ZN(n18975) );
  OAI22_X1 U20995 ( .A1(n19144), .A2(n18973), .B1(n19108), .B2(n18972), .ZN(
        n18974) );
  AOI211_X1 U20996 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19159), .A(
        n18975), .B(n18974), .ZN(n18982) );
  NAND2_X1 U20997 ( .A1(n19032), .A2(n18976), .ZN(n18977) );
  XNOR2_X1 U20998 ( .A(n18978), .B(n18977), .ZN(n18980) );
  AOI22_X1 U20999 ( .A1(n18980), .A2(n19167), .B1(n19131), .B2(n18979), .ZN(
        n18981) );
  OAI211_X1 U21000 ( .C1(n19161), .C2(n19978), .A(n18982), .B(n18981), .ZN(
        P2_U2850) );
  AOI21_X1 U21001 ( .B1(n19158), .B2(P2_EBX_REG_6__SCAN_IN), .A(n19047), .ZN(
        n18983) );
  INV_X1 U21002 ( .A(n18983), .ZN(n18986) );
  OAI22_X1 U21003 ( .A1(n19144), .A2(n18984), .B1(n13185), .B2(n19111), .ZN(
        n18985) );
  AOI211_X1 U21004 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19159), .A(
        n18986), .B(n18985), .ZN(n18993) );
  NOR2_X1 U21005 ( .A1(n19134), .A2(n18987), .ZN(n18989) );
  XNOR2_X1 U21006 ( .A(n18989), .B(n18988), .ZN(n18991) );
  AOI22_X1 U21007 ( .A1(n18991), .A2(n19167), .B1(n19131), .B2(n18990), .ZN(
        n18992) );
  OAI211_X1 U21008 ( .C1(n19161), .C2(n19931), .A(n18993), .B(n18992), .ZN(
        P2_U2849) );
  NAND2_X1 U21009 ( .A1(n19032), .A2(n18994), .ZN(n18996) );
  XOR2_X1 U21010 ( .A(n18996), .B(n18995), .Z(n19004) );
  AOI22_X1 U21011 ( .A1(n18997), .A2(n19156), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19159), .ZN(n18998) );
  OAI211_X1 U21012 ( .C1(n18999), .C2(n19111), .A(n18998), .B(n19068), .ZN(
        n19002) );
  OAI22_X1 U21013 ( .A1(n19716), .A2(n19161), .B1(n19163), .B2(n19000), .ZN(
        n19001) );
  AOI211_X1 U21014 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19158), .A(n19002), .B(
        n19001), .ZN(n19003) );
  OAI21_X1 U21015 ( .B1(n19004), .B2(n19201), .A(n19003), .ZN(P2_U2848) );
  OAI21_X1 U21016 ( .B1(n13200), .B2(n19111), .A(n19068), .ZN(n19007) );
  OAI22_X1 U21017 ( .A1(n19005), .A2(n19144), .B1(n19108), .B2(n13630), .ZN(
        n19006) );
  AOI211_X1 U21018 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19159), .A(
        n19007), .B(n19006), .ZN(n19014) );
  NAND2_X1 U21019 ( .A1(n19032), .A2(n19008), .ZN(n19009) );
  XOR2_X1 U21020 ( .A(n19010), .B(n19009), .Z(n19012) );
  AOI22_X1 U21021 ( .A1(n19012), .A2(n19167), .B1(n19011), .B2(n19131), .ZN(
        n19013) );
  OAI211_X1 U21022 ( .C1(n19710), .C2(n19161), .A(n19014), .B(n19013), .ZN(
        P2_U2846) );
  NOR2_X1 U21023 ( .A1(n19111), .A2(n19015), .ZN(n19024) );
  INV_X1 U21024 ( .A(n19016), .ZN(n19020) );
  INV_X1 U21025 ( .A(n19017), .ZN(n19018) );
  OAI211_X1 U21026 ( .C1(n19020), .C2(n19026), .A(n19019), .B(n19018), .ZN(
        n19022) );
  AOI22_X1 U21027 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19159), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19158), .ZN(n19021) );
  NAND3_X1 U21028 ( .A1(n19022), .A2(n19021), .A3(n19068), .ZN(n19023) );
  AOI211_X1 U21029 ( .C1(n19025), .C2(n19156), .A(n19024), .B(n19023), .ZN(
        n19030) );
  OAI22_X1 U21030 ( .A1(n19027), .A2(n19163), .B1(n19049), .B2(n19026), .ZN(
        n19028) );
  INV_X1 U21031 ( .A(n19028), .ZN(n19029) );
  OAI211_X1 U21032 ( .C1(n19698), .C2(n19161), .A(n19030), .B(n19029), .ZN(
        P2_U2842) );
  NAND2_X1 U21033 ( .A1(n19032), .A2(n19031), .ZN(n19033) );
  XOR2_X1 U21034 ( .A(n19034), .B(n19033), .Z(n19045) );
  AOI22_X1 U21035 ( .A1(n19035), .A2(n19156), .B1(P2_EBX_REG_15__SCAN_IN), 
        .B2(n19158), .ZN(n19036) );
  OAI21_X1 U21036 ( .B1(n19038), .B2(n19037), .A(n19036), .ZN(n19039) );
  AOI211_X1 U21037 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19155), .A(n19040), 
        .B(n19039), .ZN(n19044) );
  OAI22_X1 U21038 ( .A1(n19041), .A2(n19163), .B1(n19692), .B2(n19161), .ZN(
        n19042) );
  INV_X1 U21039 ( .A(n19042), .ZN(n19043) );
  OAI211_X1 U21040 ( .C1(n19201), .C2(n19045), .A(n19044), .B(n19043), .ZN(
        P2_U2840) );
  NAND2_X1 U21041 ( .A1(n19046), .A2(n19131), .ZN(n19052) );
  AOI21_X1 U21042 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19159), .A(
        n19047), .ZN(n19048) );
  OAI21_X1 U21043 ( .B1(n19049), .B2(n19057), .A(n19048), .ZN(n19050) );
  AOI21_X1 U21044 ( .B1(n19155), .B2(P2_REIP_REG_17__SCAN_IN), .A(n19050), 
        .ZN(n19051) );
  OAI211_X1 U21045 ( .C1(n19108), .C2(n19053), .A(n19052), .B(n19051), .ZN(
        n19054) );
  AOI21_X1 U21046 ( .B1(n19156), .B2(n19055), .A(n19054), .ZN(n19060) );
  OAI21_X1 U21047 ( .B1(n19058), .B2(n19057), .A(n19056), .ZN(n19059) );
  OAI211_X1 U21048 ( .C1(n19161), .C2(n19061), .A(n19060), .B(n19059), .ZN(
        P2_U2838) );
  AOI22_X1 U21049 ( .A1(n19063), .A2(n19131), .B1(n19062), .B2(n19118), .ZN(
        n19074) );
  AOI211_X1 U21050 ( .C1(n19066), .C2(n19065), .A(n19064), .B(n19201), .ZN(
        n19072) );
  AOI22_X1 U21051 ( .A1(n19067), .A2(n19156), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n19158), .ZN(n19069) );
  OAI211_X1 U21052 ( .C1(n19070), .C2(n19111), .A(n19069), .B(n19068), .ZN(
        n19071) );
  AOI211_X1 U21053 ( .C1(n19159), .C2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19072), .B(n19071), .ZN(n19073) );
  NAND2_X1 U21054 ( .A1(n19074), .A2(n19073), .ZN(P2_U2836) );
  OAI22_X1 U21055 ( .A1(n19076), .A2(n19163), .B1(n19075), .B2(n19161), .ZN(
        n19077) );
  INV_X1 U21056 ( .A(n19077), .ZN(n19087) );
  AOI211_X1 U21057 ( .C1(n19080), .C2(n19079), .A(n19078), .B(n19201), .ZN(
        n19085) );
  OAI222_X1 U21058 ( .A1(n19111), .A2(n19083), .B1(n19082), .B2(n19108), .C1(
        n19081), .C2(n19144), .ZN(n19084) );
  AOI211_X1 U21059 ( .C1(n19159), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n19085), .B(n19084), .ZN(n19086) );
  NAND2_X1 U21060 ( .A1(n19087), .A2(n19086), .ZN(P2_U2834) );
  AOI22_X1 U21061 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19159), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19155), .ZN(n19099) );
  AOI22_X1 U21062 ( .A1(n19088), .A2(n19156), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n19158), .ZN(n19098) );
  INV_X1 U21063 ( .A(n19089), .ZN(n19091) );
  INV_X1 U21064 ( .A(n19090), .ZN(n19924) );
  AOI22_X1 U21065 ( .A1(n19091), .A2(n19131), .B1(n19924), .B2(n19118), .ZN(
        n19097) );
  AOI21_X1 U21066 ( .B1(n19094), .B2(n19093), .A(n19092), .ZN(n19095) );
  NAND2_X1 U21067 ( .A1(n19167), .A2(n19095), .ZN(n19096) );
  NAND4_X1 U21068 ( .A1(n19099), .A2(n19098), .A3(n19097), .A4(n19096), .ZN(
        P2_U2833) );
  INV_X1 U21069 ( .A(n19100), .ZN(n19103) );
  INV_X1 U21070 ( .A(n19101), .ZN(n19102) );
  AOI22_X1 U21071 ( .A1(n19103), .A2(n19131), .B1(n19102), .B2(n19118), .ZN(
        n19115) );
  AOI211_X1 U21072 ( .C1(n19106), .C2(n19105), .A(n19104), .B(n19201), .ZN(
        n19113) );
  OAI222_X1 U21073 ( .A1(n19111), .A2(n19110), .B1(n19109), .B2(n19108), .C1(
        n19107), .C2(n19144), .ZN(n19112) );
  AOI211_X1 U21074 ( .C1(n19159), .C2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n19113), .B(n19112), .ZN(n19114) );
  NAND2_X1 U21075 ( .A1(n19115), .A2(n19114), .ZN(P2_U2832) );
  AOI22_X1 U21076 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19159), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19155), .ZN(n19127) );
  AOI22_X1 U21077 ( .A1(n19116), .A2(n19156), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n19158), .ZN(n19126) );
  INV_X1 U21078 ( .A(n19117), .ZN(n19120) );
  AOI22_X1 U21079 ( .A1(n19120), .A2(n19131), .B1(n19119), .B2(n19118), .ZN(
        n19125) );
  OR2_X1 U21080 ( .A1(n19121), .A2(n19134), .ZN(n19123) );
  OAI21_X1 U21081 ( .B1(n19134), .B2(n19104), .A(n19121), .ZN(n19122) );
  OAI211_X1 U21082 ( .C1(n19104), .C2(n19123), .A(n19167), .B(n19122), .ZN(
        n19124) );
  NAND4_X1 U21083 ( .A1(n19127), .A2(n19126), .A3(n19125), .A4(n19124), .ZN(
        P2_U2831) );
  AOI22_X1 U21084 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19159), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19155), .ZN(n19141) );
  AOI22_X1 U21085 ( .A1(n19128), .A2(n19156), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n19158), .ZN(n19140) );
  NOR2_X1 U21086 ( .A1(n19129), .A2(n19161), .ZN(n19130) );
  AOI21_X1 U21087 ( .B1(n19132), .B2(n19131), .A(n19130), .ZN(n19139) );
  OR2_X1 U21088 ( .A1(n19133), .A2(n19134), .ZN(n19136) );
  OAI21_X1 U21089 ( .B1(n19134), .B2(n19137), .A(n19133), .ZN(n19135) );
  OAI211_X1 U21090 ( .C1(n19137), .C2(n19136), .A(n19167), .B(n19135), .ZN(
        n19138) );
  NAND4_X1 U21091 ( .A1(n19141), .A2(n19140), .A3(n19139), .A4(n19138), .ZN(
        P2_U2829) );
  AOI22_X1 U21092 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19159), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19155), .ZN(n19143) );
  OAI21_X1 U21093 ( .B1(n11639), .B2(n19144), .A(n19143), .ZN(n19145) );
  AOI21_X1 U21094 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19158), .A(n19145), .ZN(
        n19153) );
  OAI211_X1 U21095 ( .C1(n19148), .C2(n19147), .A(n19146), .B(n19167), .ZN(
        n19149) );
  OAI21_X1 U21096 ( .B1(n19150), .B2(n19163), .A(n19149), .ZN(n19151) );
  INV_X1 U21097 ( .A(n19151), .ZN(n19152) );
  OAI211_X1 U21098 ( .C1(n19154), .C2(n19161), .A(n19153), .B(n19152), .ZN(
        P2_U2828) );
  AOI22_X1 U21099 ( .A1(n19157), .A2(n19156), .B1(n19155), .B2(
        P2_REIP_REG_28__SCAN_IN), .ZN(n19173) );
  AOI22_X1 U21100 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19159), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n19158), .ZN(n19172) );
  INV_X1 U21101 ( .A(n19160), .ZN(n19162) );
  OAI22_X1 U21102 ( .A1(n19164), .A2(n19163), .B1(n19162), .B2(n19161), .ZN(
        n19165) );
  INV_X1 U21103 ( .A(n19165), .ZN(n19171) );
  OAI211_X1 U21104 ( .C1(n19169), .C2(n19168), .A(n19167), .B(n19166), .ZN(
        n19170) );
  NAND4_X1 U21105 ( .A1(n19173), .A2(n19172), .A3(n19171), .A4(n19170), .ZN(
        P2_U2827) );
  INV_X1 U21106 ( .A(n19174), .ZN(n19176) );
  NOR4_X1 U21107 ( .A1(n13315), .A2(n19176), .A3(n11178), .A4(n19196), .ZN(
        n19177) );
  NAND2_X1 U21108 ( .A1(n19180), .A2(n19177), .ZN(n19178) );
  OAI21_X1 U21109 ( .B1(n19180), .B2(n19179), .A(n19178), .ZN(P2_U3595) );
  OAI22_X1 U21110 ( .A1(n19184), .A2(n19183), .B1(n19182), .B2(n19181), .ZN(
        n19188) );
  MUX2_X1 U21111 ( .A(n19186), .B(n19185), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n19187) );
  AOI211_X1 U21112 ( .C1(n19190), .C2(n19189), .A(n19188), .B(n19187), .ZN(
        n19192) );
  OAI211_X1 U21113 ( .C1(n19194), .C2(n19193), .A(n19192), .B(n19191), .ZN(
        P2_U3046) );
  NAND2_X1 U21114 ( .A1(n19210), .A2(n19195), .ZN(n19212) );
  NAND2_X1 U21115 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19213), .ZN(n19197) );
  OAI21_X1 U21116 ( .B1(n19197), .B2(n19196), .A(n19219), .ZN(n19200) );
  NAND2_X1 U21117 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n22274), .ZN(n19198) );
  AOI21_X1 U21118 ( .B1(n19204), .B2(n19212), .A(n19198), .ZN(n19199) );
  AOI21_X1 U21119 ( .B1(n19212), .B2(n19200), .A(n19199), .ZN(n19202) );
  NAND2_X1 U21120 ( .A1(n19202), .A2(n19201), .ZN(P2_U3177) );
  INV_X1 U21121 ( .A(n19203), .ZN(n19206) );
  OAI22_X1 U21122 ( .A1(n19206), .A2(n19205), .B1(n19204), .B2(n19213), .ZN(
        n19208) );
  OR2_X1 U21123 ( .A1(n19208), .A2(n19207), .ZN(n19209) );
  AOI21_X1 U21124 ( .B1(n19210), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n19209), 
        .ZN(n19217) );
  NOR2_X1 U21125 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19211), .ZN(n19215) );
  OAI22_X1 U21126 ( .A1(n19215), .A2(n19214), .B1(n19213), .B2(n19212), .ZN(
        n19216) );
  OAI211_X1 U21127 ( .C1(n19218), .C2(n19219), .A(n19217), .B(n19216), .ZN(
        P2_U3176) );
  NOR2_X1 U21128 ( .A1(n19220), .A2(n19219), .ZN(n19223) );
  MUX2_X1 U21129 ( .A(P2_MORE_REG_SCAN_IN), .B(n19221), .S(n19223), .Z(
        P2_U3609) );
  OAI21_X1 U21130 ( .B1(n19223), .B2(n14245), .A(n19222), .ZN(P2_U2819) );
  INV_X1 U21131 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20627) );
  INV_X1 U21132 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n21230) );
  AOI22_X1 U21133 ( .A1(n19581), .A2(n20627), .B1(n21230), .B2(U215), .ZN(U282) );
  OAI22_X1 U21134 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19581), .ZN(n19224) );
  INV_X1 U21135 ( .A(n19224), .ZN(U281) );
  OAI22_X1 U21136 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19581), .ZN(n19225) );
  INV_X1 U21137 ( .A(n19225), .ZN(U280) );
  OAI22_X1 U21138 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19581), .ZN(n19226) );
  INV_X1 U21139 ( .A(n19226), .ZN(U279) );
  OAI22_X1 U21140 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19581), .ZN(n19227) );
  INV_X1 U21141 ( .A(n19227), .ZN(U278) );
  OAI22_X1 U21142 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19581), .ZN(n19228) );
  INV_X1 U21143 ( .A(n19228), .ZN(U277) );
  OAI22_X1 U21144 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19581), .ZN(n19229) );
  INV_X1 U21145 ( .A(n19229), .ZN(U276) );
  OAI22_X1 U21146 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19581), .ZN(n19230) );
  INV_X1 U21147 ( .A(n19230), .ZN(U275) );
  OAI22_X1 U21148 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19581), .ZN(n19231) );
  INV_X1 U21149 ( .A(n19231), .ZN(U274) );
  OAI22_X1 U21150 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19581), .ZN(n19232) );
  INV_X1 U21151 ( .A(n19232), .ZN(U273) );
  OAI22_X1 U21152 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19581), .ZN(n19233) );
  INV_X1 U21153 ( .A(n19233), .ZN(U272) );
  OAI22_X1 U21154 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19581), .ZN(n19234) );
  INV_X1 U21155 ( .A(n19234), .ZN(U271) );
  OAI22_X1 U21156 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19247), .ZN(n19235) );
  INV_X1 U21157 ( .A(n19235), .ZN(U270) );
  OAI22_X1 U21158 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19581), .ZN(n19236) );
  INV_X1 U21159 ( .A(n19236), .ZN(U269) );
  OAI22_X1 U21160 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19247), .ZN(n19237) );
  INV_X1 U21161 ( .A(n19237), .ZN(U268) );
  OAI22_X1 U21162 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19581), .ZN(n19238) );
  INV_X1 U21163 ( .A(n19238), .ZN(U267) );
  OAI22_X1 U21164 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19247), .ZN(n19239) );
  INV_X1 U21165 ( .A(n19239), .ZN(U266) );
  OAI22_X1 U21166 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19581), .ZN(n19240) );
  INV_X1 U21167 ( .A(n19240), .ZN(U265) );
  OAI22_X1 U21168 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19247), .ZN(n19241) );
  INV_X1 U21169 ( .A(n19241), .ZN(U264) );
  OAI22_X1 U21170 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19247), .ZN(n19242) );
  INV_X1 U21171 ( .A(n19242), .ZN(U263) );
  OAI22_X1 U21172 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19247), .ZN(n19243) );
  INV_X1 U21173 ( .A(n19243), .ZN(U262) );
  OAI22_X1 U21174 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19247), .ZN(n19244) );
  INV_X1 U21175 ( .A(n19244), .ZN(U261) );
  OAI22_X1 U21176 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n19247), .ZN(n19245) );
  INV_X1 U21177 ( .A(n19245), .ZN(U260) );
  OAI22_X1 U21178 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19247), .ZN(n19246) );
  INV_X1 U21179 ( .A(n19246), .ZN(U259) );
  OAI22_X1 U21180 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19247), .ZN(n19248) );
  INV_X1 U21181 ( .A(n19248), .ZN(U258) );
  NAND3_X1 U21182 ( .A1(n21809), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19259) );
  NOR2_X2 U21183 ( .A1(n19259), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19605) );
  INV_X1 U21184 ( .A(n19605), .ZN(n19598) );
  NOR2_X1 U21185 ( .A1(n21230), .A2(n19584), .ZN(n19328) );
  INV_X1 U21186 ( .A(n19328), .ZN(n19297) );
  INV_X1 U21187 ( .A(n19259), .ZN(n19260) );
  NAND2_X1 U21188 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19260), .ZN(
        n19593) );
  INV_X1 U21189 ( .A(n19593), .ZN(n19682) );
  NAND2_X1 U21190 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19585), .ZN(n19308) );
  INV_X1 U21191 ( .A(n19308), .ZN(n19326) );
  NOR2_X1 U21192 ( .A1(n21836), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21829) );
  NAND2_X1 U21193 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19249), .ZN(
        n19250) );
  NOR2_X1 U21194 ( .A1(n21829), .A2(n19250), .ZN(n19587) );
  INV_X1 U21195 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21150) );
  NOR2_X2 U21196 ( .A1(n21150), .A2(n19586), .ZN(n19325) );
  AOI22_X1 U21197 ( .A1(n19682), .A2(n19326), .B1(n19587), .B2(n19325), .ZN(
        n19255) );
  INV_X1 U21198 ( .A(n19250), .ZN(n19318) );
  NOR2_X1 U21199 ( .A1(n19251), .A2(n19586), .ZN(n19276) );
  AOI22_X1 U21200 ( .A1(n19585), .A2(n19260), .B1(n19318), .B2(n19276), .ZN(
        n19590) );
  NAND2_X1 U21201 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19318), .ZN(
        n19569) );
  INV_X1 U21202 ( .A(n19569), .ZN(n19669) );
  NAND2_X1 U21203 ( .A1(n19253), .A2(n19252), .ZN(n19588) );
  NOR2_X2 U21204 ( .A1(n21219), .A2(n19588), .ZN(n19327) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19590), .B1(
        n19669), .B2(n19327), .ZN(n19254) );
  OAI211_X1 U21206 ( .C1(n19598), .C2(n19297), .A(n19255), .B(n19254), .ZN(
        P3_U2995) );
  NOR2_X1 U21207 ( .A1(n21809), .A2(n19275), .ZN(n19268) );
  NAND2_X1 U21208 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19268), .ZN(
        n19541) );
  INV_X1 U21209 ( .A(n19541), .ZN(n19610) );
  NAND2_X1 U21210 ( .A1(n21806), .A2(n19318), .ZN(n19675) );
  INV_X1 U21211 ( .A(n19675), .ZN(n19679) );
  NOR2_X1 U21212 ( .A1(n19682), .A2(n19679), .ZN(n19323) );
  NOR2_X1 U21213 ( .A1(n21829), .A2(n19323), .ZN(n19594) );
  AOI22_X1 U21214 ( .A1(n19328), .A2(n19610), .B1(n19325), .B2(n19594), .ZN(
        n19258) );
  NOR2_X1 U21215 ( .A1(n19605), .A2(n19610), .ZN(n19263) );
  OAI21_X1 U21216 ( .B1(n21836), .B2(n21806), .A(n19536), .ZN(n19322) );
  AOI221_X1 U21217 ( .B1(n19323), .B2(n19310), .C1(n19323), .C2(n19263), .A(
        n19322), .ZN(n19256) );
  INV_X1 U21218 ( .A(n19256), .ZN(n19595) );
  AOI22_X1 U21219 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19595), .B1(
        n19327), .B2(n19679), .ZN(n19257) );
  OAI211_X1 U21220 ( .C1(n19598), .C2(n19308), .A(n19258), .B(n19257), .ZN(
        P3_U2987) );
  INV_X1 U21221 ( .A(n19268), .ZN(n19267) );
  NOR2_X2 U21222 ( .A1(n19267), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19616) );
  INV_X1 U21223 ( .A(n19616), .ZN(n19603) );
  NOR2_X1 U21224 ( .A1(n21829), .A2(n19259), .ZN(n19599) );
  AOI22_X1 U21225 ( .A1(n19326), .A2(n19610), .B1(n19325), .B2(n19599), .ZN(
        n19262) );
  AOI22_X1 U21226 ( .A1(n19585), .A2(n19268), .B1(n19276), .B2(n19260), .ZN(
        n19600) );
  AOI22_X1 U21227 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19600), .B1(
        n19327), .B2(n19682), .ZN(n19261) );
  OAI211_X1 U21228 ( .C1(n19297), .C2(n19603), .A(n19262), .B(n19261), .ZN(
        P3_U2979) );
  NAND2_X1 U21229 ( .A1(n21809), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19298) );
  INV_X1 U21230 ( .A(n19622), .ZN(n19614) );
  NOR2_X1 U21231 ( .A1(n21829), .A2(n19263), .ZN(n19604) );
  AOI22_X1 U21232 ( .A1(n19326), .A2(n19616), .B1(n19325), .B2(n19604), .ZN(
        n19266) );
  NOR2_X1 U21233 ( .A1(n19616), .A2(n19622), .ZN(n19271) );
  OAI22_X1 U21234 ( .A1(n19584), .A2(n19271), .B1(n19322), .B2(n19263), .ZN(
        n19264) );
  INV_X1 U21235 ( .A(n19264), .ZN(n19606) );
  AOI22_X1 U21236 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19327), .ZN(n19265) );
  OAI211_X1 U21237 ( .C1(n19297), .C2(n19614), .A(n19266), .B(n19265), .ZN(
        P3_U2971) );
  NAND2_X1 U21238 ( .A1(n21809), .A2(n21806), .ZN(n21811) );
  NOR2_X2 U21239 ( .A1(n21811), .A2(n19275), .ZN(n19628) );
  INV_X1 U21240 ( .A(n19628), .ZN(n19620) );
  NOR2_X1 U21241 ( .A1(n21829), .A2(n19267), .ZN(n19609) );
  AOI22_X1 U21242 ( .A1(n19326), .A2(n19622), .B1(n19325), .B2(n19609), .ZN(
        n19270) );
  INV_X1 U21243 ( .A(n19275), .ZN(n19277) );
  AOI22_X1 U21244 ( .A1(n19585), .A2(n19277), .B1(n19276), .B2(n19268), .ZN(
        n19611) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19611), .B1(
        n19327), .B2(n19610), .ZN(n19269) );
  OAI211_X1 U21246 ( .C1(n19297), .C2(n19620), .A(n19270), .B(n19269), .ZN(
        P3_U2963) );
  NAND2_X1 U21247 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19278), .ZN(
        n19626) );
  INV_X1 U21248 ( .A(n19626), .ZN(n19634) );
  NOR2_X1 U21249 ( .A1(n21829), .A2(n19271), .ZN(n19615) );
  AOI22_X1 U21250 ( .A1(n19328), .A2(n19634), .B1(n19325), .B2(n19615), .ZN(
        n19274) );
  NAND2_X1 U21251 ( .A1(n19620), .A2(n19626), .ZN(n19282) );
  INV_X1 U21252 ( .A(n19282), .ZN(n19281) );
  OAI21_X1 U21253 ( .B1(n19281), .B2(n19310), .A(n19271), .ZN(n19272) );
  OAI211_X1 U21254 ( .C1(n19616), .C2(n21836), .A(n19536), .B(n19272), .ZN(
        n19617) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19617), .B1(
        n19327), .B2(n19616), .ZN(n19273) );
  OAI211_X1 U21256 ( .C1(n19308), .C2(n19620), .A(n19274), .B(n19273), .ZN(
        P3_U2955) );
  NAND2_X1 U21257 ( .A1(n21806), .A2(n19278), .ZN(n19632) );
  INV_X1 U21258 ( .A(n19632), .ZN(n19639) );
  INV_X1 U21259 ( .A(n21829), .ZN(n20681) );
  NAND2_X1 U21260 ( .A1(n21809), .A2(n20681), .ZN(n19315) );
  NOR2_X1 U21261 ( .A1(n19275), .A2(n19315), .ZN(n19621) );
  AOI22_X1 U21262 ( .A1(n19328), .A2(n19639), .B1(n19325), .B2(n19621), .ZN(
        n19280) );
  AND2_X1 U21263 ( .A1(n21809), .A2(n19276), .ZN(n19317) );
  AOI22_X1 U21264 ( .A1(n19585), .A2(n19278), .B1(n19277), .B2(n19317), .ZN(
        n19623) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19623), .B1(
        n19327), .B2(n19622), .ZN(n19279) );
  OAI211_X1 U21266 ( .C1(n19308), .C2(n19626), .A(n19280), .B(n19279), .ZN(
        P3_U2947) );
  NOR2_X2 U21267 ( .A1(n19298), .A2(n19293), .ZN(n19645) );
  INV_X1 U21268 ( .A(n19645), .ZN(n19554) );
  NOR2_X1 U21269 ( .A1(n21829), .A2(n19281), .ZN(n19627) );
  AOI22_X1 U21270 ( .A1(n19326), .A2(n19639), .B1(n19325), .B2(n19627), .ZN(
        n19284) );
  NAND2_X1 U21271 ( .A1(n19632), .A2(n19554), .ZN(n19290) );
  INV_X1 U21272 ( .A(n19322), .ZN(n19301) );
  AOI22_X1 U21273 ( .A1(n19585), .A2(n19290), .B1(n19301), .B2(n19282), .ZN(
        n19629) );
  AOI22_X1 U21274 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19629), .B1(
        n19327), .B2(n19628), .ZN(n19283) );
  OAI211_X1 U21275 ( .C1(n19297), .C2(n19554), .A(n19284), .B(n19283), .ZN(
        P3_U2939) );
  NOR2_X2 U21276 ( .A1(n21811), .A2(n19293), .ZN(n19651) );
  NOR2_X1 U21277 ( .A1(n21829), .A2(n19285), .ZN(n19633) );
  AOI22_X1 U21278 ( .A1(n19328), .A2(n19651), .B1(n19325), .B2(n19633), .ZN(
        n19288) );
  INV_X1 U21279 ( .A(n19293), .ZN(n19294) );
  AOI21_X1 U21280 ( .B1(n21809), .B2(n19310), .A(n19586), .ZN(n19304) );
  NAND3_X1 U21281 ( .A1(n19294), .A2(n19304), .A3(n19286), .ZN(n19635) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19635), .B1(
        n19327), .B2(n19634), .ZN(n19287) );
  OAI211_X1 U21283 ( .C1(n19308), .C2(n19554), .A(n19288), .B(n19287), .ZN(
        P3_U2931) );
  NOR2_X1 U21284 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19316) );
  INV_X1 U21285 ( .A(n19316), .ZN(n19314) );
  NOR2_X1 U21286 ( .A1(n21809), .A2(n19314), .ZN(n19305) );
  NAND2_X1 U21287 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19305), .ZN(
        n19649) );
  AND2_X1 U21288 ( .A1(n20681), .A2(n19290), .ZN(n19638) );
  AOI22_X1 U21289 ( .A1(n19326), .A2(n19651), .B1(n19325), .B2(n19638), .ZN(
        n19292) );
  INV_X1 U21290 ( .A(n19651), .ZN(n19643) );
  NAND2_X1 U21291 ( .A1(n19643), .A2(n19649), .ZN(n19300) );
  OAI221_X1 U21292 ( .B1(n19290), .B2(n19289), .C1(n19290), .C2(n19300), .A(
        n19301), .ZN(n19640) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19640), .B1(
        n19327), .B2(n19639), .ZN(n19291) );
  OAI211_X1 U21294 ( .C1(n19297), .C2(n19649), .A(n19292), .B(n19291), .ZN(
        P3_U2923) );
  NAND2_X1 U21295 ( .A1(n19305), .A2(n21806), .ZN(n19564) );
  INV_X1 U21296 ( .A(n19649), .ZN(n19657) );
  NOR2_X1 U21297 ( .A1(n19315), .A2(n19293), .ZN(n19644) );
  AOI22_X1 U21298 ( .A1(n19326), .A2(n19657), .B1(n19325), .B2(n19644), .ZN(
        n19296) );
  AOI22_X1 U21299 ( .A1(n19585), .A2(n19305), .B1(n19317), .B2(n19294), .ZN(
        n19646) );
  AOI22_X1 U21300 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19646), .B1(
        n19327), .B2(n19645), .ZN(n19295) );
  OAI211_X1 U21301 ( .C1(n19297), .C2(n19564), .A(n19296), .B(n19295), .ZN(
        P3_U2915) );
  INV_X1 U21302 ( .A(n19298), .ZN(n19299) );
  NAND2_X1 U21303 ( .A1(n19299), .A2(n19316), .ZN(n19660) );
  INV_X1 U21304 ( .A(n19660), .ZN(n19670) );
  AND2_X1 U21305 ( .A1(n20681), .A2(n19300), .ZN(n19650) );
  AOI22_X1 U21306 ( .A1(n19328), .A2(n19670), .B1(n19325), .B2(n19650), .ZN(
        n19303) );
  NAND2_X1 U21307 ( .A1(n19564), .A2(n19660), .ZN(n19309) );
  AOI22_X1 U21308 ( .A1(n19585), .A2(n19309), .B1(n19301), .B2(n19300), .ZN(
        n19652) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19652), .B1(
        n19327), .B2(n19651), .ZN(n19302) );
  OAI211_X1 U21310 ( .C1(n19308), .C2(n19564), .A(n19303), .B(n19302), .ZN(
        P3_U2907) );
  OAI211_X1 U21311 ( .C1(n19657), .C2(n21836), .A(n19316), .B(n19304), .ZN(
        n19656) );
  AND2_X1 U21312 ( .A1(n20681), .A2(n19305), .ZN(n19655) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19656), .B1(
        n19325), .B2(n19655), .ZN(n19307) );
  AOI22_X1 U21314 ( .A1(n19328), .A2(n19576), .B1(n19327), .B2(n19657), .ZN(
        n19306) );
  OAI211_X1 U21315 ( .C1(n19308), .C2(n19660), .A(n19307), .B(n19306), .ZN(
        P3_U2899) );
  INV_X1 U21316 ( .A(n19327), .ZN(n19321) );
  AND2_X1 U21317 ( .A1(n20681), .A2(n19309), .ZN(n19661) );
  AOI22_X1 U21318 ( .A1(n19326), .A2(n19576), .B1(n19325), .B2(n19661), .ZN(
        n19313) );
  INV_X1 U21319 ( .A(n19564), .ZN(n19662) );
  NOR2_X1 U21320 ( .A1(n19669), .A2(n19576), .ZN(n19324) );
  OAI22_X1 U21321 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19660), .B1(n19324), 
        .B2(n19310), .ZN(n19311) );
  OAI21_X1 U21322 ( .B1(n19662), .B2(n19311), .A(n19536), .ZN(n19663) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19663), .B1(
        n19328), .B2(n19669), .ZN(n19312) );
  OAI211_X1 U21324 ( .C1(n19321), .C2(n19564), .A(n19313), .B(n19312), .ZN(
        P3_U2891) );
  NOR2_X1 U21325 ( .A1(n19315), .A2(n19314), .ZN(n19668) );
  AOI22_X1 U21326 ( .A1(n19669), .A2(n19326), .B1(n19325), .B2(n19668), .ZN(
        n19320) );
  AOI22_X1 U21327 ( .A1(n19585), .A2(n19318), .B1(n19317), .B2(n19316), .ZN(
        n19671) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19671), .B1(
        n19328), .B2(n19679), .ZN(n19319) );
  OAI211_X1 U21329 ( .C1(n19321), .C2(n19660), .A(n19320), .B(n19319), .ZN(
        P3_U2883) );
  OAI22_X1 U21330 ( .A1(n19323), .A2(n19584), .B1(n19324), .B2(n19322), .ZN(
        n19685) );
  NOR2_X1 U21331 ( .A1(n21829), .A2(n19324), .ZN(n19677) );
  AOI22_X1 U21332 ( .A1(n19326), .A2(n19679), .B1(n19325), .B2(n19677), .ZN(
        n19330) );
  AOI22_X1 U21333 ( .A1(n19328), .A2(n19682), .B1(n19327), .B2(n19576), .ZN(
        n19329) );
  OAI211_X1 U21334 ( .C1(n19331), .C2(n19685), .A(n19330), .B(n19329), .ZN(
        P3_U2875) );
  OAI22_X1 U21335 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19581), .ZN(n19332) );
  INV_X1 U21336 ( .A(n19332), .ZN(U257) );
  INV_X1 U21337 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n21193) );
  NOR2_X1 U21338 ( .A1(n21193), .A2(n19584), .ZN(n19368) );
  INV_X1 U21339 ( .A(n19368), .ZN(n19359) );
  NAND2_X1 U21340 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19585), .ZN(n19364) );
  INV_X1 U21341 ( .A(n19364), .ZN(n19366) );
  NOR2_X2 U21342 ( .A1(n21199), .A2(n19586), .ZN(n19365) );
  AOI22_X1 U21343 ( .A1(n19605), .A2(n19366), .B1(n19587), .B2(n19365), .ZN(
        n19334) );
  NOR2_X2 U21344 ( .A1(n21180), .A2(n19588), .ZN(n19367) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19590), .B1(
        n19669), .B2(n19367), .ZN(n19333) );
  OAI211_X1 U21346 ( .C1(n19593), .C2(n19359), .A(n19334), .B(n19333), .ZN(
        P3_U2994) );
  AOI22_X1 U21347 ( .A1(n19610), .A2(n19366), .B1(n19594), .B2(n19365), .ZN(
        n19336) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19595), .B1(
        n19679), .B2(n19367), .ZN(n19335) );
  OAI211_X1 U21349 ( .C1(n19598), .C2(n19359), .A(n19336), .B(n19335), .ZN(
        P3_U2986) );
  AOI22_X1 U21350 ( .A1(n19616), .A2(n19366), .B1(n19599), .B2(n19365), .ZN(
        n19338) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19600), .B1(
        n19682), .B2(n19367), .ZN(n19337) );
  OAI211_X1 U21352 ( .C1(n19541), .C2(n19359), .A(n19338), .B(n19337), .ZN(
        P3_U2978) );
  AOI22_X1 U21353 ( .A1(n19616), .A2(n19368), .B1(n19604), .B2(n19365), .ZN(
        n19340) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19367), .ZN(n19339) );
  OAI211_X1 U21355 ( .C1(n19614), .C2(n19364), .A(n19340), .B(n19339), .ZN(
        P3_U2970) );
  AOI22_X1 U21356 ( .A1(n19628), .A2(n19366), .B1(n19609), .B2(n19365), .ZN(
        n19342) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19367), .ZN(n19341) );
  OAI211_X1 U21358 ( .C1(n19614), .C2(n19359), .A(n19342), .B(n19341), .ZN(
        P3_U2962) );
  AOI22_X1 U21359 ( .A1(n19634), .A2(n19366), .B1(n19615), .B2(n19365), .ZN(
        n19344) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19367), .ZN(n19343) );
  OAI211_X1 U21361 ( .C1(n19620), .C2(n19359), .A(n19344), .B(n19343), .ZN(
        P3_U2954) );
  AOI22_X1 U21362 ( .A1(n19639), .A2(n19366), .B1(n19621), .B2(n19365), .ZN(
        n19346) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19367), .ZN(n19345) );
  OAI211_X1 U21364 ( .C1(n19626), .C2(n19359), .A(n19346), .B(n19345), .ZN(
        P3_U2946) );
  AOI22_X1 U21365 ( .A1(n19645), .A2(n19366), .B1(n19627), .B2(n19365), .ZN(
        n19348) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19367), .ZN(n19347) );
  OAI211_X1 U21367 ( .C1(n19632), .C2(n19359), .A(n19348), .B(n19347), .ZN(
        P3_U2938) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19635), .B1(
        n19633), .B2(n19365), .ZN(n19350) );
  AOI22_X1 U21369 ( .A1(n19634), .A2(n19367), .B1(n19651), .B2(n19366), .ZN(
        n19349) );
  OAI211_X1 U21370 ( .C1(n19554), .C2(n19359), .A(n19350), .B(n19349), .ZN(
        P3_U2930) );
  AOI22_X1 U21371 ( .A1(n19657), .A2(n19366), .B1(n19638), .B2(n19365), .ZN(
        n19352) );
  AOI22_X1 U21372 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19367), .ZN(n19351) );
  OAI211_X1 U21373 ( .C1(n19643), .C2(n19359), .A(n19352), .B(n19351), .ZN(
        P3_U2922) );
  AOI22_X1 U21374 ( .A1(n19662), .A2(n19366), .B1(n19644), .B2(n19365), .ZN(
        n19354) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19367), .ZN(n19353) );
  OAI211_X1 U21376 ( .C1(n19649), .C2(n19359), .A(n19354), .B(n19353), .ZN(
        P3_U2914) );
  AOI22_X1 U21377 ( .A1(n19670), .A2(n19366), .B1(n19650), .B2(n19365), .ZN(
        n19356) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19652), .B1(
        n19651), .B2(n19367), .ZN(n19355) );
  OAI211_X1 U21379 ( .C1(n19564), .C2(n19359), .A(n19356), .B(n19355), .ZN(
        P3_U2906) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19656), .B1(
        n19655), .B2(n19365), .ZN(n19358) );
  AOI22_X1 U21381 ( .A1(n19657), .A2(n19367), .B1(n19576), .B2(n19366), .ZN(
        n19357) );
  OAI211_X1 U21382 ( .C1(n19660), .C2(n19359), .A(n19358), .B(n19357), .ZN(
        P3_U2898) );
  AOI22_X1 U21383 ( .A1(n19576), .A2(n19368), .B1(n19661), .B2(n19365), .ZN(
        n19361) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19367), .ZN(n19360) );
  OAI211_X1 U21385 ( .C1(n19569), .C2(n19364), .A(n19361), .B(n19360), .ZN(
        P3_U2890) );
  AOI22_X1 U21386 ( .A1(n19669), .A2(n19368), .B1(n19668), .B2(n19365), .ZN(
        n19363) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19367), .ZN(n19362) );
  OAI211_X1 U21388 ( .C1(n19675), .C2(n19364), .A(n19363), .B(n19362), .ZN(
        P3_U2882) );
  AOI22_X1 U21389 ( .A1(n19682), .A2(n19366), .B1(n19677), .B2(n19365), .ZN(
        n19370) );
  AOI22_X1 U21390 ( .A1(n19679), .A2(n19368), .B1(n19576), .B2(n19367), .ZN(
        n19369) );
  OAI211_X1 U21391 ( .C1(n19371), .C2(n19685), .A(n19370), .B(n19369), .ZN(
        P3_U2874) );
  OAI22_X1 U21392 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19581), .ZN(n19372) );
  INV_X1 U21393 ( .A(n19372), .ZN(U256) );
  NOR2_X1 U21394 ( .A1(n17051), .A2(n19584), .ZN(n19406) );
  INV_X1 U21395 ( .A(n19406), .ZN(n19404) );
  NAND2_X1 U21396 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n19585), .ZN(n19401) );
  INV_X1 U21397 ( .A(n19401), .ZN(n19408) );
  INV_X1 U21398 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21159) );
  NOR2_X2 U21399 ( .A1(n21159), .A2(n19586), .ZN(n19405) );
  AOI22_X1 U21400 ( .A1(n19682), .A2(n19408), .B1(n19587), .B2(n19405), .ZN(
        n19374) );
  NOR2_X2 U21401 ( .A1(n15979), .A2(n19588), .ZN(n19407) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19590), .B1(
        n19669), .B2(n19407), .ZN(n19373) );
  OAI211_X1 U21403 ( .C1(n19598), .C2(n19404), .A(n19374), .B(n19373), .ZN(
        P3_U2993) );
  AOI22_X1 U21404 ( .A1(n19605), .A2(n19408), .B1(n19594), .B2(n19405), .ZN(
        n19376) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19595), .B1(
        n19679), .B2(n19407), .ZN(n19375) );
  OAI211_X1 U21406 ( .C1(n19541), .C2(n19404), .A(n19376), .B(n19375), .ZN(
        P3_U2985) );
  AOI22_X1 U21407 ( .A1(n19616), .A2(n19406), .B1(n19599), .B2(n19405), .ZN(
        n19378) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19600), .B1(
        n19682), .B2(n19407), .ZN(n19377) );
  OAI211_X1 U21409 ( .C1(n19541), .C2(n19401), .A(n19378), .B(n19377), .ZN(
        P3_U2977) );
  AOI22_X1 U21410 ( .A1(n19622), .A2(n19406), .B1(n19604), .B2(n19405), .ZN(
        n19380) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19407), .ZN(n19379) );
  OAI211_X1 U21412 ( .C1(n19603), .C2(n19401), .A(n19380), .B(n19379), .ZN(
        P3_U2969) );
  AOI22_X1 U21413 ( .A1(n19628), .A2(n19406), .B1(n19609), .B2(n19405), .ZN(
        n19382) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19407), .ZN(n19381) );
  OAI211_X1 U21415 ( .C1(n19614), .C2(n19401), .A(n19382), .B(n19381), .ZN(
        P3_U2961) );
  AOI22_X1 U21416 ( .A1(n19628), .A2(n19408), .B1(n19615), .B2(n19405), .ZN(
        n19384) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19407), .ZN(n19383) );
  OAI211_X1 U21418 ( .C1(n19626), .C2(n19404), .A(n19384), .B(n19383), .ZN(
        P3_U2953) );
  AOI22_X1 U21419 ( .A1(n19634), .A2(n19408), .B1(n19621), .B2(n19405), .ZN(
        n19386) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19407), .ZN(n19385) );
  OAI211_X1 U21421 ( .C1(n19632), .C2(n19404), .A(n19386), .B(n19385), .ZN(
        P3_U2945) );
  AOI22_X1 U21422 ( .A1(n19639), .A2(n19408), .B1(n19627), .B2(n19405), .ZN(
        n19388) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19407), .ZN(n19387) );
  OAI211_X1 U21424 ( .C1(n19554), .C2(n19404), .A(n19388), .B(n19387), .ZN(
        P3_U2937) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19635), .B1(
        n19633), .B2(n19405), .ZN(n19390) );
  AOI22_X1 U21426 ( .A1(n19634), .A2(n19407), .B1(n19645), .B2(n19408), .ZN(
        n19389) );
  OAI211_X1 U21427 ( .C1(n19643), .C2(n19404), .A(n19390), .B(n19389), .ZN(
        P3_U2929) );
  AOI22_X1 U21428 ( .A1(n19651), .A2(n19408), .B1(n19638), .B2(n19405), .ZN(
        n19392) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19407), .ZN(n19391) );
  OAI211_X1 U21430 ( .C1(n19649), .C2(n19404), .A(n19392), .B(n19391), .ZN(
        P3_U2921) );
  AOI22_X1 U21431 ( .A1(n19657), .A2(n19408), .B1(n19644), .B2(n19405), .ZN(
        n19394) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19407), .ZN(n19393) );
  OAI211_X1 U21433 ( .C1(n19564), .C2(n19404), .A(n19394), .B(n19393), .ZN(
        P3_U2913) );
  AOI22_X1 U21434 ( .A1(n19670), .A2(n19406), .B1(n19650), .B2(n19405), .ZN(
        n19396) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19652), .B1(
        n19651), .B2(n19407), .ZN(n19395) );
  OAI211_X1 U21436 ( .C1(n19564), .C2(n19401), .A(n19396), .B(n19395), .ZN(
        P3_U2905) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19656), .B1(
        n19655), .B2(n19405), .ZN(n19398) );
  AOI22_X1 U21438 ( .A1(n19657), .A2(n19407), .B1(n19576), .B2(n19406), .ZN(
        n19397) );
  OAI211_X1 U21439 ( .C1(n19660), .C2(n19401), .A(n19398), .B(n19397), .ZN(
        P3_U2897) );
  INV_X1 U21440 ( .A(n19576), .ZN(n19667) );
  AOI22_X1 U21441 ( .A1(n19669), .A2(n19406), .B1(n19661), .B2(n19405), .ZN(
        n19400) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19407), .ZN(n19399) );
  OAI211_X1 U21443 ( .C1(n19667), .C2(n19401), .A(n19400), .B(n19399), .ZN(
        P3_U2889) );
  AOI22_X1 U21444 ( .A1(n19669), .A2(n19408), .B1(n19668), .B2(n19405), .ZN(
        n19403) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19407), .ZN(n19402) );
  OAI211_X1 U21446 ( .C1(n19675), .C2(n19404), .A(n19403), .B(n19402), .ZN(
        P3_U2881) );
  AOI22_X1 U21447 ( .A1(n19682), .A2(n19406), .B1(n19677), .B2(n19405), .ZN(
        n19410) );
  AOI22_X1 U21448 ( .A1(n19679), .A2(n19408), .B1(n19576), .B2(n19407), .ZN(
        n19409) );
  OAI211_X1 U21449 ( .C1(n19411), .C2(n19685), .A(n19410), .B(n19409), .ZN(
        P3_U2873) );
  OAI22_X1 U21450 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19581), .ZN(n19412) );
  INV_X1 U21451 ( .A(n19412), .ZN(U255) );
  INV_X1 U21452 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19413) );
  NOR2_X1 U21453 ( .A1(n19413), .A2(n19584), .ZN(n19447) );
  INV_X1 U21454 ( .A(n19447), .ZN(n19442) );
  NAND2_X1 U21455 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n19585), .ZN(n19445) );
  INV_X1 U21456 ( .A(n19445), .ZN(n19449) );
  INV_X1 U21457 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n21191) );
  NOR2_X2 U21458 ( .A1(n21191), .A2(n19586), .ZN(n19446) );
  AOI22_X1 U21459 ( .A1(n19682), .A2(n19449), .B1(n19587), .B2(n19446), .ZN(
        n19415) );
  NOR2_X2 U21460 ( .A1(n21364), .A2(n19588), .ZN(n19448) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19590), .B1(
        n19669), .B2(n19448), .ZN(n19414) );
  OAI211_X1 U21462 ( .C1(n19598), .C2(n19442), .A(n19415), .B(n19414), .ZN(
        P3_U2992) );
  AOI22_X1 U21463 ( .A1(n19605), .A2(n19449), .B1(n19594), .B2(n19446), .ZN(
        n19417) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19595), .B1(
        n19679), .B2(n19448), .ZN(n19416) );
  OAI211_X1 U21465 ( .C1(n19541), .C2(n19442), .A(n19417), .B(n19416), .ZN(
        P3_U2984) );
  AOI22_X1 U21466 ( .A1(n19610), .A2(n19449), .B1(n19599), .B2(n19446), .ZN(
        n19419) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19600), .B1(
        n19682), .B2(n19448), .ZN(n19418) );
  OAI211_X1 U21468 ( .C1(n19603), .C2(n19442), .A(n19419), .B(n19418), .ZN(
        P3_U2976) );
  AOI22_X1 U21469 ( .A1(n19616), .A2(n19449), .B1(n19604), .B2(n19446), .ZN(
        n19421) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19448), .ZN(n19420) );
  OAI211_X1 U21471 ( .C1(n19614), .C2(n19442), .A(n19421), .B(n19420), .ZN(
        P3_U2968) );
  AOI22_X1 U21472 ( .A1(n19628), .A2(n19447), .B1(n19609), .B2(n19446), .ZN(
        n19423) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19448), .ZN(n19422) );
  OAI211_X1 U21474 ( .C1(n19614), .C2(n19445), .A(n19423), .B(n19422), .ZN(
        P3_U2960) );
  AOI22_X1 U21475 ( .A1(n19628), .A2(n19449), .B1(n19615), .B2(n19446), .ZN(
        n19425) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19448), .ZN(n19424) );
  OAI211_X1 U21477 ( .C1(n19626), .C2(n19442), .A(n19425), .B(n19424), .ZN(
        P3_U2952) );
  AOI22_X1 U21478 ( .A1(n19634), .A2(n19449), .B1(n19621), .B2(n19446), .ZN(
        n19427) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19448), .ZN(n19426) );
  OAI211_X1 U21480 ( .C1(n19632), .C2(n19442), .A(n19427), .B(n19426), .ZN(
        P3_U2944) );
  AOI22_X1 U21481 ( .A1(n19645), .A2(n19447), .B1(n19627), .B2(n19446), .ZN(
        n19429) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19448), .ZN(n19428) );
  OAI211_X1 U21483 ( .C1(n19632), .C2(n19445), .A(n19429), .B(n19428), .ZN(
        P3_U2936) );
  AOI22_X1 U21484 ( .A1(n19645), .A2(n19449), .B1(n19633), .B2(n19446), .ZN(
        n19431) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19635), .B1(
        n19634), .B2(n19448), .ZN(n19430) );
  OAI211_X1 U21486 ( .C1(n19643), .C2(n19442), .A(n19431), .B(n19430), .ZN(
        P3_U2928) );
  AOI22_X1 U21487 ( .A1(n19657), .A2(n19447), .B1(n19638), .B2(n19446), .ZN(
        n19433) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19448), .ZN(n19432) );
  OAI211_X1 U21489 ( .C1(n19643), .C2(n19445), .A(n19433), .B(n19432), .ZN(
        P3_U2920) );
  AOI22_X1 U21490 ( .A1(n19662), .A2(n19447), .B1(n19644), .B2(n19446), .ZN(
        n19435) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19448), .ZN(n19434) );
  OAI211_X1 U21492 ( .C1(n19649), .C2(n19445), .A(n19435), .B(n19434), .ZN(
        P3_U2912) );
  AOI22_X1 U21493 ( .A1(n19670), .A2(n19447), .B1(n19650), .B2(n19446), .ZN(
        n19437) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19652), .B1(
        n19651), .B2(n19448), .ZN(n19436) );
  OAI211_X1 U21495 ( .C1(n19564), .C2(n19445), .A(n19437), .B(n19436), .ZN(
        P3_U2904) );
  AOI22_X1 U21496 ( .A1(n19576), .A2(n19447), .B1(n19655), .B2(n19446), .ZN(
        n19439) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19656), .B1(
        n19657), .B2(n19448), .ZN(n19438) );
  OAI211_X1 U21498 ( .C1(n19660), .C2(n19445), .A(n19439), .B(n19438), .ZN(
        P3_U2896) );
  AOI22_X1 U21499 ( .A1(n19576), .A2(n19449), .B1(n19661), .B2(n19446), .ZN(
        n19441) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19448), .ZN(n19440) );
  OAI211_X1 U21501 ( .C1(n19569), .C2(n19442), .A(n19441), .B(n19440), .ZN(
        P3_U2888) );
  AOI22_X1 U21502 ( .A1(n19679), .A2(n19447), .B1(n19668), .B2(n19446), .ZN(
        n19444) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19448), .ZN(n19443) );
  OAI211_X1 U21504 ( .C1(n19569), .C2(n19445), .A(n19444), .B(n19443), .ZN(
        P3_U2880) );
  AOI22_X1 U21505 ( .A1(n19682), .A2(n19447), .B1(n19677), .B2(n19446), .ZN(
        n19451) );
  AOI22_X1 U21506 ( .A1(n19679), .A2(n19449), .B1(n19576), .B2(n19448), .ZN(
        n19450) );
  OAI211_X1 U21507 ( .C1(n19452), .C2(n19685), .A(n19451), .B(n19450), .ZN(
        P3_U2872) );
  OAI22_X1 U21508 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19581), .ZN(n19453) );
  INV_X1 U21509 ( .A(n19453), .ZN(U254) );
  INV_X1 U21510 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19454) );
  NOR2_X1 U21511 ( .A1(n19584), .A2(n19454), .ZN(n19489) );
  INV_X1 U21512 ( .A(n19489), .ZN(n19487) );
  NAND2_X1 U21513 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19585), .ZN(n19482) );
  INV_X1 U21514 ( .A(n19482), .ZN(n19491) );
  INV_X1 U21515 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n21168) );
  NOR2_X2 U21516 ( .A1(n19586), .A2(n21168), .ZN(n19488) );
  AOI22_X1 U21517 ( .A1(n19605), .A2(n19491), .B1(n19587), .B2(n19488), .ZN(
        n19457) );
  NOR2_X2 U21518 ( .A1(n19455), .A2(n19588), .ZN(n19490) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19590), .B1(
        n19669), .B2(n19490), .ZN(n19456) );
  OAI211_X1 U21520 ( .C1(n19593), .C2(n19487), .A(n19457), .B(n19456), .ZN(
        P3_U2991) );
  AOI22_X1 U21521 ( .A1(n19610), .A2(n19491), .B1(n19594), .B2(n19488), .ZN(
        n19459) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19595), .B1(
        n19679), .B2(n19490), .ZN(n19458) );
  OAI211_X1 U21523 ( .C1(n19598), .C2(n19487), .A(n19459), .B(n19458), .ZN(
        P3_U2983) );
  AOI22_X1 U21524 ( .A1(n19610), .A2(n19489), .B1(n19599), .B2(n19488), .ZN(
        n19461) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19600), .B1(
        n19682), .B2(n19490), .ZN(n19460) );
  OAI211_X1 U21526 ( .C1(n19603), .C2(n19482), .A(n19461), .B(n19460), .ZN(
        P3_U2975) );
  AOI22_X1 U21527 ( .A1(n19616), .A2(n19489), .B1(n19604), .B2(n19488), .ZN(
        n19463) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19490), .ZN(n19462) );
  OAI211_X1 U21529 ( .C1(n19614), .C2(n19482), .A(n19463), .B(n19462), .ZN(
        P3_U2967) );
  AOI22_X1 U21530 ( .A1(n19628), .A2(n19491), .B1(n19609), .B2(n19488), .ZN(
        n19465) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19490), .ZN(n19464) );
  OAI211_X1 U21532 ( .C1(n19614), .C2(n19487), .A(n19465), .B(n19464), .ZN(
        P3_U2959) );
  AOI22_X1 U21533 ( .A1(n19628), .A2(n19489), .B1(n19615), .B2(n19488), .ZN(
        n19467) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19490), .ZN(n19466) );
  OAI211_X1 U21535 ( .C1(n19626), .C2(n19482), .A(n19467), .B(n19466), .ZN(
        P3_U2951) );
  AOI22_X1 U21536 ( .A1(n19639), .A2(n19491), .B1(n19621), .B2(n19488), .ZN(
        n19469) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19490), .ZN(n19468) );
  OAI211_X1 U21538 ( .C1(n19626), .C2(n19487), .A(n19469), .B(n19468), .ZN(
        P3_U2943) );
  AOI22_X1 U21539 ( .A1(n19639), .A2(n19489), .B1(n19627), .B2(n19488), .ZN(
        n19471) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19490), .ZN(n19470) );
  OAI211_X1 U21541 ( .C1(n19554), .C2(n19482), .A(n19471), .B(n19470), .ZN(
        P3_U2935) );
  AOI22_X1 U21542 ( .A1(n19645), .A2(n19489), .B1(n19633), .B2(n19488), .ZN(
        n19473) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19635), .B1(
        n19634), .B2(n19490), .ZN(n19472) );
  OAI211_X1 U21544 ( .C1(n19643), .C2(n19482), .A(n19473), .B(n19472), .ZN(
        P3_U2927) );
  AOI22_X1 U21545 ( .A1(n19657), .A2(n19491), .B1(n19638), .B2(n19488), .ZN(
        n19475) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19490), .ZN(n19474) );
  OAI211_X1 U21547 ( .C1(n19643), .C2(n19487), .A(n19475), .B(n19474), .ZN(
        P3_U2919) );
  AOI22_X1 U21548 ( .A1(n19657), .A2(n19489), .B1(n19644), .B2(n19488), .ZN(
        n19477) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19490), .ZN(n19476) );
  OAI211_X1 U21550 ( .C1(n19564), .C2(n19482), .A(n19477), .B(n19476), .ZN(
        P3_U2911) );
  AOI22_X1 U21551 ( .A1(n19662), .A2(n19489), .B1(n19650), .B2(n19488), .ZN(
        n19479) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19652), .B1(
        n19651), .B2(n19490), .ZN(n19478) );
  OAI211_X1 U21553 ( .C1(n19660), .C2(n19482), .A(n19479), .B(n19478), .ZN(
        P3_U2903) );
  AOI22_X1 U21554 ( .A1(n19670), .A2(n19489), .B1(n19655), .B2(n19488), .ZN(
        n19481) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19656), .B1(
        n19657), .B2(n19490), .ZN(n19480) );
  OAI211_X1 U21556 ( .C1(n19667), .C2(n19482), .A(n19481), .B(n19480), .ZN(
        P3_U2895) );
  AOI22_X1 U21557 ( .A1(n19669), .A2(n19491), .B1(n19661), .B2(n19488), .ZN(
        n19484) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19490), .ZN(n19483) );
  OAI211_X1 U21559 ( .C1(n19667), .C2(n19487), .A(n19484), .B(n19483), .ZN(
        P3_U2887) );
  AOI22_X1 U21560 ( .A1(n19679), .A2(n19491), .B1(n19668), .B2(n19488), .ZN(
        n19486) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19490), .ZN(n19485) );
  OAI211_X1 U21562 ( .C1(n19569), .C2(n19487), .A(n19486), .B(n19485), .ZN(
        P3_U2879) );
  AOI22_X1 U21563 ( .A1(n19679), .A2(n19489), .B1(n19677), .B2(n19488), .ZN(
        n19493) );
  AOI22_X1 U21564 ( .A1(n19682), .A2(n19491), .B1(n19576), .B2(n19490), .ZN(
        n19492) );
  OAI211_X1 U21565 ( .C1(n19494), .C2(n19685), .A(n19493), .B(n19492), .ZN(
        P3_U2871) );
  OAI22_X1 U21566 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19581), .ZN(n19495) );
  INV_X1 U21567 ( .A(n19495), .ZN(U253) );
  NOR2_X1 U21568 ( .A1(n17076), .A2(n19584), .ZN(n19531) );
  INV_X1 U21569 ( .A(n19531), .ZN(n19524) );
  NAND2_X1 U21570 ( .A1(n19585), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19527) );
  INV_X1 U21571 ( .A(n19527), .ZN(n19529) );
  INV_X1 U21572 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n21211) );
  NOR2_X2 U21573 ( .A1(n19586), .A2(n21211), .ZN(n19528) );
  AOI22_X1 U21574 ( .A1(n19682), .A2(n19529), .B1(n19587), .B2(n19528), .ZN(
        n19497) );
  NOR2_X2 U21575 ( .A1(n21369), .A2(n19588), .ZN(n19530) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19590), .B1(
        n19669), .B2(n19530), .ZN(n19496) );
  OAI211_X1 U21577 ( .C1(n19598), .C2(n19524), .A(n19497), .B(n19496), .ZN(
        P3_U2990) );
  AOI22_X1 U21578 ( .A1(n19610), .A2(n19531), .B1(n19594), .B2(n19528), .ZN(
        n19499) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19595), .B1(
        n19679), .B2(n19530), .ZN(n19498) );
  OAI211_X1 U21580 ( .C1(n19598), .C2(n19527), .A(n19499), .B(n19498), .ZN(
        P3_U2982) );
  AOI22_X1 U21581 ( .A1(n19610), .A2(n19529), .B1(n19599), .B2(n19528), .ZN(
        n19501) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19600), .B1(
        n19682), .B2(n19530), .ZN(n19500) );
  OAI211_X1 U21583 ( .C1(n19603), .C2(n19524), .A(n19501), .B(n19500), .ZN(
        P3_U2974) );
  AOI22_X1 U21584 ( .A1(n19622), .A2(n19531), .B1(n19604), .B2(n19528), .ZN(
        n19503) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19530), .ZN(n19502) );
  OAI211_X1 U21586 ( .C1(n19603), .C2(n19527), .A(n19503), .B(n19502), .ZN(
        P3_U2966) );
  AOI22_X1 U21587 ( .A1(n19628), .A2(n19531), .B1(n19609), .B2(n19528), .ZN(
        n19505) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19530), .ZN(n19504) );
  OAI211_X1 U21589 ( .C1(n19614), .C2(n19527), .A(n19505), .B(n19504), .ZN(
        P3_U2958) );
  AOI22_X1 U21590 ( .A1(n19628), .A2(n19529), .B1(n19615), .B2(n19528), .ZN(
        n19507) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19530), .ZN(n19506) );
  OAI211_X1 U21592 ( .C1(n19626), .C2(n19524), .A(n19507), .B(n19506), .ZN(
        P3_U2950) );
  AOI22_X1 U21593 ( .A1(n19639), .A2(n19531), .B1(n19621), .B2(n19528), .ZN(
        n19509) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19530), .ZN(n19508) );
  OAI211_X1 U21595 ( .C1(n19626), .C2(n19527), .A(n19509), .B(n19508), .ZN(
        P3_U2942) );
  AOI22_X1 U21596 ( .A1(n19639), .A2(n19529), .B1(n19627), .B2(n19528), .ZN(
        n19511) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19530), .ZN(n19510) );
  OAI211_X1 U21598 ( .C1(n19554), .C2(n19524), .A(n19511), .B(n19510), .ZN(
        P3_U2934) );
  AOI22_X1 U21599 ( .A1(n19645), .A2(n19529), .B1(n19633), .B2(n19528), .ZN(
        n19513) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19635), .B1(
        n19634), .B2(n19530), .ZN(n19512) );
  OAI211_X1 U21601 ( .C1(n19643), .C2(n19524), .A(n19513), .B(n19512), .ZN(
        P3_U2926) );
  AOI22_X1 U21602 ( .A1(n19651), .A2(n19529), .B1(n19638), .B2(n19528), .ZN(
        n19515) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19530), .ZN(n19514) );
  OAI211_X1 U21604 ( .C1(n19649), .C2(n19524), .A(n19515), .B(n19514), .ZN(
        P3_U2918) );
  AOI22_X1 U21605 ( .A1(n19657), .A2(n19529), .B1(n19644), .B2(n19528), .ZN(
        n19517) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19530), .ZN(n19516) );
  OAI211_X1 U21607 ( .C1(n19564), .C2(n19524), .A(n19517), .B(n19516), .ZN(
        P3_U2910) );
  AOI22_X1 U21608 ( .A1(n19662), .A2(n19529), .B1(n19650), .B2(n19528), .ZN(
        n19519) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19652), .B1(
        n19651), .B2(n19530), .ZN(n19518) );
  OAI211_X1 U21610 ( .C1(n19660), .C2(n19524), .A(n19519), .B(n19518), .ZN(
        P3_U2902) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19656), .B1(
        n19655), .B2(n19528), .ZN(n19521) );
  AOI22_X1 U21612 ( .A1(n19657), .A2(n19530), .B1(n19576), .B2(n19531), .ZN(
        n19520) );
  OAI211_X1 U21613 ( .C1(n19660), .C2(n19527), .A(n19521), .B(n19520), .ZN(
        P3_U2894) );
  AOI22_X1 U21614 ( .A1(n19576), .A2(n19529), .B1(n19661), .B2(n19528), .ZN(
        n19523) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19530), .ZN(n19522) );
  OAI211_X1 U21616 ( .C1(n19569), .C2(n19524), .A(n19523), .B(n19522), .ZN(
        P3_U2886) );
  AOI22_X1 U21617 ( .A1(n19679), .A2(n19531), .B1(n19668), .B2(n19528), .ZN(
        n19526) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19530), .ZN(n19525) );
  OAI211_X1 U21619 ( .C1(n19569), .C2(n19527), .A(n19526), .B(n19525), .ZN(
        P3_U2878) );
  AOI22_X1 U21620 ( .A1(n19679), .A2(n19529), .B1(n19677), .B2(n19528), .ZN(
        n19533) );
  AOI22_X1 U21621 ( .A1(n19682), .A2(n19531), .B1(n19576), .B2(n19530), .ZN(
        n19532) );
  OAI211_X1 U21622 ( .C1(n19534), .C2(n19685), .A(n19533), .B(n19532), .ZN(
        P3_U2870) );
  OAI22_X1 U21623 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19581), .ZN(n19535) );
  INV_X1 U21624 ( .A(n19535), .ZN(U252) );
  INV_X1 U21625 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n21224) );
  NOR2_X1 U21626 ( .A1(n21224), .A2(n19584), .ZN(n19577) );
  INV_X1 U21627 ( .A(n19577), .ZN(n19572) );
  NAND2_X1 U21628 ( .A1(n19585), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19563) );
  INV_X1 U21629 ( .A(n19563), .ZN(n19574) );
  AND2_X1 U21630 ( .A1(n19536), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19573) );
  AOI22_X1 U21631 ( .A1(n19682), .A2(n19574), .B1(n19587), .B2(n19573), .ZN(
        n19538) );
  NOR2_X2 U21632 ( .A1(n20684), .A2(n19588), .ZN(n19575) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19590), .B1(
        n19669), .B2(n19575), .ZN(n19537) );
  OAI211_X1 U21634 ( .C1(n19598), .C2(n19572), .A(n19538), .B(n19537), .ZN(
        P3_U2989) );
  AOI22_X1 U21635 ( .A1(n19605), .A2(n19574), .B1(n19594), .B2(n19573), .ZN(
        n19540) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19595), .B1(
        n19679), .B2(n19575), .ZN(n19539) );
  OAI211_X1 U21637 ( .C1(n19541), .C2(n19572), .A(n19540), .B(n19539), .ZN(
        P3_U2981) );
  AOI22_X1 U21638 ( .A1(n19610), .A2(n19574), .B1(n19599), .B2(n19573), .ZN(
        n19543) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19600), .B1(
        n19682), .B2(n19575), .ZN(n19542) );
  OAI211_X1 U21640 ( .C1(n19603), .C2(n19572), .A(n19543), .B(n19542), .ZN(
        P3_U2973) );
  AOI22_X1 U21641 ( .A1(n19616), .A2(n19574), .B1(n19604), .B2(n19573), .ZN(
        n19545) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19575), .ZN(n19544) );
  OAI211_X1 U21643 ( .C1(n19614), .C2(n19572), .A(n19545), .B(n19544), .ZN(
        P3_U2965) );
  AOI22_X1 U21644 ( .A1(n19622), .A2(n19574), .B1(n19609), .B2(n19573), .ZN(
        n19547) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19575), .ZN(n19546) );
  OAI211_X1 U21646 ( .C1(n19620), .C2(n19572), .A(n19547), .B(n19546), .ZN(
        P3_U2957) );
  AOI22_X1 U21647 ( .A1(n19634), .A2(n19577), .B1(n19615), .B2(n19573), .ZN(
        n19549) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19575), .ZN(n19548) );
  OAI211_X1 U21649 ( .C1(n19620), .C2(n19563), .A(n19549), .B(n19548), .ZN(
        P3_U2949) );
  AOI22_X1 U21650 ( .A1(n19639), .A2(n19577), .B1(n19621), .B2(n19573), .ZN(
        n19551) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19575), .ZN(n19550) );
  OAI211_X1 U21652 ( .C1(n19626), .C2(n19563), .A(n19551), .B(n19550), .ZN(
        P3_U2941) );
  AOI22_X1 U21653 ( .A1(n19639), .A2(n19574), .B1(n19627), .B2(n19573), .ZN(
        n19553) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19575), .ZN(n19552) );
  OAI211_X1 U21655 ( .C1(n19554), .C2(n19572), .A(n19553), .B(n19552), .ZN(
        P3_U2933) );
  AOI22_X1 U21656 ( .A1(n19645), .A2(n19574), .B1(n19633), .B2(n19573), .ZN(
        n19556) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19635), .B1(
        n19634), .B2(n19575), .ZN(n19555) );
  OAI211_X1 U21658 ( .C1(n19643), .C2(n19572), .A(n19556), .B(n19555), .ZN(
        P3_U2925) );
  AOI22_X1 U21659 ( .A1(n19651), .A2(n19574), .B1(n19638), .B2(n19573), .ZN(
        n19558) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19575), .ZN(n19557) );
  OAI211_X1 U21661 ( .C1(n19649), .C2(n19572), .A(n19558), .B(n19557), .ZN(
        P3_U2917) );
  AOI22_X1 U21662 ( .A1(n19662), .A2(n19577), .B1(n19644), .B2(n19573), .ZN(
        n19560) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19575), .ZN(n19559) );
  OAI211_X1 U21664 ( .C1(n19649), .C2(n19563), .A(n19560), .B(n19559), .ZN(
        P3_U2909) );
  AOI22_X1 U21665 ( .A1(n19670), .A2(n19577), .B1(n19650), .B2(n19573), .ZN(
        n19562) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19652), .B1(
        n19651), .B2(n19575), .ZN(n19561) );
  OAI211_X1 U21667 ( .C1(n19564), .C2(n19563), .A(n19562), .B(n19561), .ZN(
        P3_U2901) );
  AOI22_X1 U21668 ( .A1(n19670), .A2(n19574), .B1(n19655), .B2(n19573), .ZN(
        n19566) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19656), .B1(
        n19657), .B2(n19575), .ZN(n19565) );
  OAI211_X1 U21670 ( .C1(n19667), .C2(n19572), .A(n19566), .B(n19565), .ZN(
        P3_U2893) );
  AOI22_X1 U21671 ( .A1(n19576), .A2(n19574), .B1(n19661), .B2(n19573), .ZN(
        n19568) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19575), .ZN(n19567) );
  OAI211_X1 U21673 ( .C1(n19569), .C2(n19572), .A(n19568), .B(n19567), .ZN(
        P3_U2885) );
  AOI22_X1 U21674 ( .A1(n19669), .A2(n19574), .B1(n19668), .B2(n19573), .ZN(
        n19571) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19575), .ZN(n19570) );
  OAI211_X1 U21676 ( .C1(n19675), .C2(n19572), .A(n19571), .B(n19570), .ZN(
        P3_U2877) );
  AOI22_X1 U21677 ( .A1(n19679), .A2(n19574), .B1(n19677), .B2(n19573), .ZN(
        n19579) );
  AOI22_X1 U21678 ( .A1(n19682), .A2(n19577), .B1(n19576), .B2(n19575), .ZN(
        n19578) );
  OAI211_X1 U21679 ( .C1(n19580), .C2(n19685), .A(n19579), .B(n19578), .ZN(
        P3_U2869) );
  OAI22_X1 U21680 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19581), .ZN(n19582) );
  INV_X1 U21681 ( .A(n19582), .ZN(U251) );
  INV_X1 U21682 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19583) );
  NOR2_X1 U21683 ( .A1(n19584), .A2(n19583), .ZN(n19678) );
  INV_X1 U21684 ( .A(n19678), .ZN(n19666) );
  NAND2_X1 U21685 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19585), .ZN(n19674) );
  INV_X1 U21686 ( .A(n19674), .ZN(n19681) );
  INV_X1 U21687 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n21274) );
  NOR2_X2 U21688 ( .A1(n19586), .A2(n21274), .ZN(n19676) );
  AOI22_X1 U21689 ( .A1(n19605), .A2(n19681), .B1(n19587), .B2(n19676), .ZN(
        n19592) );
  NOR2_X2 U21690 ( .A1(n19589), .A2(n19588), .ZN(n19680) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19590), .B1(
        n19669), .B2(n19680), .ZN(n19591) );
  OAI211_X1 U21692 ( .C1(n19593), .C2(n19666), .A(n19592), .B(n19591), .ZN(
        P3_U2988) );
  AOI22_X1 U21693 ( .A1(n19610), .A2(n19681), .B1(n19594), .B2(n19676), .ZN(
        n19597) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19595), .B1(
        n19679), .B2(n19680), .ZN(n19596) );
  OAI211_X1 U21695 ( .C1(n19598), .C2(n19666), .A(n19597), .B(n19596), .ZN(
        P3_U2980) );
  AOI22_X1 U21696 ( .A1(n19610), .A2(n19678), .B1(n19599), .B2(n19676), .ZN(
        n19602) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19600), .B1(
        n19682), .B2(n19680), .ZN(n19601) );
  OAI211_X1 U21698 ( .C1(n19603), .C2(n19674), .A(n19602), .B(n19601), .ZN(
        P3_U2972) );
  AOI22_X1 U21699 ( .A1(n19616), .A2(n19678), .B1(n19604), .B2(n19676), .ZN(
        n19608) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19680), .ZN(n19607) );
  OAI211_X1 U21701 ( .C1(n19614), .C2(n19674), .A(n19608), .B(n19607), .ZN(
        P3_U2964) );
  AOI22_X1 U21702 ( .A1(n19628), .A2(n19681), .B1(n19609), .B2(n19676), .ZN(
        n19613) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19680), .ZN(n19612) );
  OAI211_X1 U21704 ( .C1(n19614), .C2(n19666), .A(n19613), .B(n19612), .ZN(
        P3_U2956) );
  AOI22_X1 U21705 ( .A1(n19634), .A2(n19681), .B1(n19615), .B2(n19676), .ZN(
        n19619) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19680), .ZN(n19618) );
  OAI211_X1 U21707 ( .C1(n19620), .C2(n19666), .A(n19619), .B(n19618), .ZN(
        P3_U2948) );
  AOI22_X1 U21708 ( .A1(n19639), .A2(n19681), .B1(n19621), .B2(n19676), .ZN(
        n19625) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19680), .ZN(n19624) );
  OAI211_X1 U21710 ( .C1(n19626), .C2(n19666), .A(n19625), .B(n19624), .ZN(
        P3_U2940) );
  AOI22_X1 U21711 ( .A1(n19645), .A2(n19681), .B1(n19627), .B2(n19676), .ZN(
        n19631) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19680), .ZN(n19630) );
  OAI211_X1 U21713 ( .C1(n19632), .C2(n19666), .A(n19631), .B(n19630), .ZN(
        P3_U2932) );
  AOI22_X1 U21714 ( .A1(n19645), .A2(n19678), .B1(n19633), .B2(n19676), .ZN(
        n19637) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19635), .B1(
        n19634), .B2(n19680), .ZN(n19636) );
  OAI211_X1 U21716 ( .C1(n19643), .C2(n19674), .A(n19637), .B(n19636), .ZN(
        P3_U2924) );
  AOI22_X1 U21717 ( .A1(n19657), .A2(n19681), .B1(n19638), .B2(n19676), .ZN(
        n19642) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19680), .ZN(n19641) );
  OAI211_X1 U21719 ( .C1(n19643), .C2(n19666), .A(n19642), .B(n19641), .ZN(
        P3_U2916) );
  AOI22_X1 U21720 ( .A1(n19662), .A2(n19681), .B1(n19644), .B2(n19676), .ZN(
        n19648) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19680), .ZN(n19647) );
  OAI211_X1 U21722 ( .C1(n19649), .C2(n19666), .A(n19648), .B(n19647), .ZN(
        P3_U2908) );
  AOI22_X1 U21723 ( .A1(n19662), .A2(n19678), .B1(n19650), .B2(n19676), .ZN(
        n19654) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19652), .B1(
        n19651), .B2(n19680), .ZN(n19653) );
  OAI211_X1 U21725 ( .C1(n19660), .C2(n19674), .A(n19654), .B(n19653), .ZN(
        P3_U2900) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19656), .B1(
        n19655), .B2(n19676), .ZN(n19659) );
  AOI22_X1 U21727 ( .A1(n19657), .A2(n19680), .B1(n19576), .B2(n19681), .ZN(
        n19658) );
  OAI211_X1 U21728 ( .C1(n19660), .C2(n19666), .A(n19659), .B(n19658), .ZN(
        P3_U2892) );
  AOI22_X1 U21729 ( .A1(n19669), .A2(n19681), .B1(n19661), .B2(n19676), .ZN(
        n19665) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19663), .B1(
        n19662), .B2(n19680), .ZN(n19664) );
  OAI211_X1 U21731 ( .C1(n19667), .C2(n19666), .A(n19665), .B(n19664), .ZN(
        P3_U2884) );
  AOI22_X1 U21732 ( .A1(n19669), .A2(n19678), .B1(n19668), .B2(n19676), .ZN(
        n19673) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19680), .ZN(n19672) );
  OAI211_X1 U21734 ( .C1(n19675), .C2(n19674), .A(n19673), .B(n19672), .ZN(
        P3_U2876) );
  AOI22_X1 U21735 ( .A1(n19679), .A2(n19678), .B1(n19677), .B2(n19676), .ZN(
        n19684) );
  AOI22_X1 U21736 ( .A1(n19682), .A2(n19681), .B1(n19576), .B2(n19680), .ZN(
        n19683) );
  OAI211_X1 U21737 ( .C1(n19686), .C2(n19685), .A(n19684), .B(n19683), .ZN(
        P3_U2868) );
  AOI22_X1 U21738 ( .A1(n19687), .A2(n20169), .B1(BUF2_REG_31__SCAN_IN), .B2(
        n20225), .ZN(n19689) );
  AOI22_X1 U21739 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n20221), .B1(n20224), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19688) );
  NAND2_X1 U21740 ( .A1(n19689), .A2(n19688), .ZN(P2_U2888) );
  OAI222_X1 U21741 ( .A1(n19692), .A2(n19979), .B1(n19691), .B2(n19929), .C1(
        n19690), .C2(n20176), .ZN(P2_U2904) );
  AOI22_X1 U21742 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n20221), .B1(n19693), 
        .B2(n19972), .ZN(n19694) );
  OAI21_X1 U21743 ( .B1(n19979), .B2(n19695), .A(n19694), .ZN(P2_U2905) );
  OAI222_X1 U21744 ( .A1(n19698), .A2(n19979), .B1(n19697), .B2(n19929), .C1(
        n20176), .C2(n19696), .ZN(P2_U2906) );
  AOI22_X1 U21745 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n20221), .B1(n19699), 
        .B2(n19972), .ZN(n19700) );
  OAI21_X1 U21746 ( .B1(n19979), .B2(n19701), .A(n19700), .ZN(P2_U2907) );
  OAI222_X1 U21747 ( .A1(n19704), .A2(n19979), .B1(n19703), .B2(n19929), .C1(
        n20176), .C2(n19702), .ZN(P2_U2908) );
  AOI22_X1 U21748 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n20221), .B1(n19705), 
        .B2(n19972), .ZN(n19706) );
  OAI21_X1 U21749 ( .B1(n19979), .B2(n19707), .A(n19706), .ZN(P2_U2909) );
  OAI222_X1 U21750 ( .A1(n19710), .A2(n19979), .B1(n19709), .B2(n19929), .C1(
        n20176), .C2(n19708), .ZN(P2_U2910) );
  INV_X1 U21751 ( .A(n19711), .ZN(n19714) );
  OAI222_X1 U21752 ( .A1(n19714), .A2(n19979), .B1(n19713), .B2(n19929), .C1(
        n20176), .C2(n19712), .ZN(P2_U2911) );
  OAI222_X1 U21753 ( .A1(n19716), .A2(n19979), .B1(n19715), .B2(n19929), .C1(
        n20176), .C2(n19721), .ZN(P2_U2912) );
  AOI22_X1 U21754 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20240), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20241), .ZN(n19921) );
  NAND3_X1 U21755 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19733) );
  NOR2_X1 U21756 ( .A1(n19719), .A2(n19777), .ZN(n20238) );
  OAI21_X1 U21757 ( .B1(n14161), .B2(n20238), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19720) );
  OAI21_X1 U21758 ( .B1(n19733), .B2(n19908), .A(n19720), .ZN(n20239) );
  NOR2_X2 U21759 ( .A1(n13338), .A2(n20236), .ZN(n19906) );
  AOI22_X1 U21760 ( .A1(n20239), .A2(n19722), .B1(n20238), .B2(n19906), .ZN(
        n19731) );
  INV_X1 U21761 ( .A(n19723), .ZN(n19724) );
  NOR2_X1 U21762 ( .A1(n19746), .A2(n19724), .ZN(n19729) );
  INV_X1 U21763 ( .A(n19733), .ZN(n19728) );
  AOI21_X1 U21764 ( .B1(n14161), .B2(n19911), .A(n20238), .ZN(n19726) );
  NAND2_X1 U21765 ( .A1(n19865), .A2(n19726), .ZN(n19727) );
  OAI211_X1 U21766 ( .C1(n19729), .C2(n19728), .A(n19914), .B(n19727), .ZN(
        n20242) );
  INV_X1 U21767 ( .A(n19860), .ZN(n19820) );
  NOR2_X2 U21768 ( .A1(n19746), .A2(n19820), .ZN(n20246) );
  AOI22_X1 U21769 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20240), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20241), .ZN(n19903) );
  INV_X1 U21770 ( .A(n19903), .ZN(n19907) );
  AOI22_X1 U21771 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20242), .B1(
        n20246), .B2(n19907), .ZN(n19730) );
  OAI211_X1 U21772 ( .C1(n19921), .C2(n20344), .A(n19731), .B(n19730), .ZN(
        P2_U3175) );
  INV_X1 U21773 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19742) );
  AOI21_X1 U21774 ( .B1(n14164), .B2(n19911), .A(n19910), .ZN(n19736) );
  NAND3_X1 U21775 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19889), .ZN(n19757) );
  NOR2_X1 U21776 ( .A1(n19891), .A2(n19757), .ZN(n20252) );
  NOR2_X1 U21777 ( .A1(n19823), .A2(n19860), .ZN(n19775) );
  OR2_X1 U21778 ( .A1(n19775), .A2(n22239), .ZN(n19877) );
  OAI21_X1 U21779 ( .B1(n19746), .B2(n19877), .A(n19880), .ZN(n19739) );
  NOR2_X1 U21780 ( .A1(n20252), .A2(n19739), .ZN(n19735) );
  NOR2_X1 U21781 ( .A1(n19733), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20245) );
  INV_X1 U21782 ( .A(n20245), .ZN(n19734) );
  OAI22_X1 U21783 ( .A1(n19736), .A2(n19735), .B1(n20234), .B2(n19734), .ZN(
        n20250) );
  NOR2_X2 U21784 ( .A1(n19746), .A2(n19884), .ZN(n20254) );
  AOI22_X1 U21785 ( .A1(n19907), .A2(n20254), .B1(n19906), .B2(n20245), .ZN(
        n19741) );
  NOR2_X1 U21786 ( .A1(n20252), .A2(n20245), .ZN(n19738) );
  OAI21_X1 U21787 ( .B1(n14164), .B2(n20245), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19737) );
  OAI21_X1 U21788 ( .B1(n19739), .B2(n19738), .A(n19737), .ZN(n20247) );
  INV_X1 U21789 ( .A(n19921), .ZN(n19900) );
  AOI22_X1 U21790 ( .A1(n19722), .A2(n20247), .B1(n20246), .B2(n19900), .ZN(
        n19740) );
  OAI211_X1 U21791 ( .C1(n19742), .C2(n20250), .A(n19741), .B(n19740), .ZN(
        P2_U3167) );
  INV_X1 U21792 ( .A(n20261), .ZN(n20258) );
  OAI21_X1 U21793 ( .B1(n14151), .B2(n20252), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19744) );
  OAI21_X1 U21794 ( .B1(n19757), .B2(n19908), .A(n19744), .ZN(n20253) );
  AOI22_X1 U21795 ( .A1(n20253), .A2(n19722), .B1(n19906), .B2(n20252), .ZN(
        n19752) );
  OR2_X1 U21796 ( .A1(n19745), .A2(n22239), .ZN(n19894) );
  OAI21_X1 U21797 ( .B1(n19746), .B2(n19894), .A(n19757), .ZN(n19750) );
  NAND2_X1 U21798 ( .A1(n14151), .A2(n19911), .ZN(n19748) );
  INV_X1 U21799 ( .A(n20252), .ZN(n19747) );
  NAND3_X1 U21800 ( .A1(n19748), .A2(n19747), .A3(n19908), .ZN(n19749) );
  NAND3_X1 U21801 ( .A1(n19750), .A2(n19914), .A3(n19749), .ZN(n20255) );
  AOI22_X1 U21802 ( .A1(n19900), .A2(n20254), .B1(n20255), .B2(
        P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n19751) );
  OAI211_X1 U21803 ( .C1(n19903), .C2(n20258), .A(n19752), .B(n19751), .ZN(
        P2_U3159) );
  INV_X1 U21804 ( .A(n19753), .ZN(n19755) );
  INV_X1 U21805 ( .A(n19754), .ZN(n19828) );
  NAND2_X1 U21806 ( .A1(n19755), .A2(n19828), .ZN(n19849) );
  INV_X1 U21807 ( .A(n19756), .ZN(n19759) );
  NOR2_X1 U21808 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19757), .ZN(
        n20259) );
  OAI21_X1 U21809 ( .B1(n14160), .B2(n20259), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19758) );
  OAI21_X1 U21810 ( .B1(n19849), .B2(n19759), .A(n19758), .ZN(n20260) );
  AOI22_X1 U21811 ( .A1(n20260), .A2(n19722), .B1(n19906), .B2(n20259), .ZN(
        n19765) );
  OAI21_X1 U21812 ( .B1(n20261), .B2(n20040), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19760) );
  OAI21_X1 U21813 ( .B1(n19849), .B2(n19777), .A(n19760), .ZN(n19763) );
  AOI211_X1 U21814 ( .C1(n14160), .C2(n19911), .A(n19880), .B(n20259), .ZN(
        n19761) );
  NOR2_X1 U21815 ( .A1(n20234), .A2(n19761), .ZN(n19762) );
  NAND2_X1 U21816 ( .A1(n19763), .A2(n19762), .ZN(n20262) );
  AOI22_X1 U21817 ( .A1(n20262), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n19900), .B2(n20261), .ZN(n19764) );
  OAI211_X1 U21818 ( .C1(n19903), .C2(n20270), .A(n19765), .B(n19764), .ZN(
        P2_U3151) );
  NAND3_X1 U21819 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19766), .ZN(n19774) );
  NOR2_X1 U21820 ( .A1(n19891), .A2(n19774), .ZN(n20265) );
  OAI21_X1 U21821 ( .B1(n14179), .B2(n20265), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19767) );
  OAI21_X1 U21822 ( .B1(n19774), .B2(n19908), .A(n19767), .ZN(n20266) );
  AOI22_X1 U21823 ( .A1(n20266), .A2(n19722), .B1(n19906), .B2(n20265), .ZN(
        n19773) );
  NAND2_X1 U21824 ( .A1(n19790), .A2(n19860), .ZN(n20193) );
  OAI21_X1 U21825 ( .B1(n19768), .B2(n19862), .A(n19774), .ZN(n19771) );
  AOI211_X1 U21826 ( .C1(n14179), .C2(n19911), .A(n19880), .B(n20265), .ZN(
        n19769) );
  NOR2_X1 U21827 ( .A1(n20234), .A2(n19769), .ZN(n19770) );
  NAND2_X1 U21828 ( .A1(n19771), .A2(n19770), .ZN(n20267) );
  AOI22_X1 U21829 ( .A1(n19907), .A2(n20272), .B1(n20267), .B2(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n19772) );
  OAI211_X1 U21830 ( .C1(n19921), .C2(n20270), .A(n19773), .B(n19772), .ZN(
        P2_U3143) );
  NOR2_X1 U21831 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19774), .ZN(
        n20271) );
  AOI22_X1 U21832 ( .A1(n19900), .A2(n20272), .B1(n19906), .B2(n20271), .ZN(
        n19789) );
  OR2_X1 U21833 ( .A1(n19776), .A2(n19775), .ZN(n19784) );
  NOR3_X1 U21834 ( .A1(n19777), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19795) );
  INV_X1 U21835 ( .A(n19795), .ZN(n19802) );
  NOR2_X1 U21836 ( .A1(n19891), .A2(n19802), .ZN(n20277) );
  NOR2_X1 U21837 ( .A1(n20271), .A2(n20277), .ZN(n19783) );
  NAND2_X1 U21838 ( .A1(n19784), .A2(n19783), .ZN(n19781) );
  INV_X1 U21839 ( .A(n14149), .ZN(n19779) );
  INV_X1 U21840 ( .A(n20271), .ZN(n19778) );
  OAI21_X1 U21841 ( .B1(n19779), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19778), 
        .ZN(n19780) );
  MUX2_X1 U21842 ( .A(n19781), .B(n19780), .S(n19908), .Z(n19782) );
  NAND2_X1 U21843 ( .A1(n19782), .A2(n19914), .ZN(n20274) );
  OAI21_X1 U21844 ( .B1(n14149), .B2(n20271), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19787) );
  INV_X1 U21845 ( .A(n19783), .ZN(n19785) );
  NAND3_X1 U21846 ( .A1(n19880), .A2(n19785), .A3(n19784), .ZN(n19786) );
  NAND2_X1 U21847 ( .A1(n19787), .A2(n19786), .ZN(n20273) );
  AOI22_X1 U21848 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20274), .B1(
        n19722), .B2(n20273), .ZN(n19788) );
  OAI211_X1 U21849 ( .C1(n19903), .C2(n20282), .A(n19789), .B(n19788), .ZN(
        P2_U3135) );
  INV_X1 U21850 ( .A(n19835), .ZN(n19887) );
  NAND2_X1 U21851 ( .A1(n19790), .A2(n19887), .ZN(n19803) );
  AOI22_X1 U21852 ( .A1(n19907), .A2(n20284), .B1(n19906), .B2(n20277), .ZN(
        n19800) );
  OAI21_X1 U21853 ( .B1(n19791), .B2(n19894), .A(n19880), .ZN(n19798) );
  NAND2_X1 U21854 ( .A1(n19796), .A2(n19911), .ZN(n19793) );
  INV_X1 U21855 ( .A(n20277), .ZN(n19792) );
  NAND3_X1 U21856 ( .A1(n19793), .A2(n19908), .A3(n19792), .ZN(n19794) );
  OAI211_X1 U21857 ( .C1(n19798), .C2(n19795), .A(n19914), .B(n19794), .ZN(
        n20279) );
  OAI21_X1 U21858 ( .B1(n19796), .B2(n20277), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19797) );
  OAI21_X1 U21859 ( .B1(n19798), .B2(n19802), .A(n19797), .ZN(n20278) );
  AOI22_X1 U21860 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20279), .B1(
        n19722), .B2(n20278), .ZN(n19799) );
  OAI211_X1 U21861 ( .C1(n19921), .C2(n20282), .A(n19800), .B(n19799), .ZN(
        P2_U3127) );
  NOR2_X1 U21862 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19802), .ZN(
        n20283) );
  AOI22_X1 U21863 ( .A1(n19900), .A2(n20284), .B1(n19906), .B2(n20283), .ZN(
        n19812) );
  AOI21_X1 U21864 ( .B1(n19803), .B2(n20294), .A(n22239), .ZN(n19804) );
  NOR2_X1 U21865 ( .A1(n19804), .A2(n19908), .ZN(n19807) );
  AOI21_X1 U21866 ( .B1(n14159), .B2(n19876), .A(n19910), .ZN(n19805) );
  AOI21_X1 U21867 ( .B1(n19807), .B2(n19815), .A(n19805), .ZN(n19806) );
  INV_X1 U21868 ( .A(n19807), .ZN(n19810) );
  OAI21_X1 U21869 ( .B1(n14159), .B2(n20283), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19809) );
  NOR2_X1 U21870 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20283), .ZN(n19808) );
  AOI22_X1 U21871 ( .A1(n19810), .A2(n19809), .B1(n19808), .B2(n19815), .ZN(
        n20285) );
  AOI22_X1 U21872 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20286), .B1(
        n19722), .B2(n20285), .ZN(n19811) );
  OAI211_X1 U21873 ( .C1(n19903), .C2(n20294), .A(n19812), .B(n19811), .ZN(
        P2_U3119) );
  NOR2_X1 U21874 ( .A1(n19889), .A2(n19847), .ZN(n19818) );
  INV_X1 U21875 ( .A(n19818), .ZN(n19825) );
  INV_X1 U21876 ( .A(n19815), .ZN(n20289) );
  OAI21_X1 U21877 ( .B1(n14163), .B2(n20289), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19813) );
  OAI21_X1 U21878 ( .B1(n19825), .B2(n19908), .A(n19813), .ZN(n20290) );
  AOI22_X1 U21879 ( .A1(n20290), .A2(n19722), .B1(n20289), .B2(n19906), .ZN(
        n19822) );
  INV_X1 U21880 ( .A(n19814), .ZN(n19819) );
  NAND2_X1 U21881 ( .A1(n14163), .A2(n19911), .ZN(n19816) );
  AOI21_X1 U21882 ( .B1(n19816), .B2(n19815), .A(n20234), .ZN(n19817) );
  OAI22_X1 U21883 ( .A1(n19819), .A2(n19818), .B1(n19910), .B2(n19817), .ZN(
        n20291) );
  NOR2_X2 U21884 ( .A1(n19836), .A2(n19820), .ZN(n20297) );
  AOI22_X1 U21885 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20291), .B1(
        n20297), .B2(n19907), .ZN(n19821) );
  OAI211_X1 U21886 ( .C1(n19921), .C2(n20294), .A(n19822), .B(n19821), .ZN(
        P2_U3111) );
  INV_X1 U21887 ( .A(n19873), .ZN(n19827) );
  NOR2_X1 U21888 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19825), .ZN(
        n20295) );
  OAI21_X1 U21889 ( .B1(n14153), .B2(n20295), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19826) );
  OAI21_X1 U21890 ( .B1(n19847), .B2(n19827), .A(n19826), .ZN(n20296) );
  AOI22_X1 U21891 ( .A1(n20296), .A2(n19722), .B1(n19906), .B2(n20295), .ZN(
        n19834) );
  OAI22_X1 U21892 ( .A1(n19836), .A2(n19877), .B1(n19847), .B2(n19828), .ZN(
        n19832) );
  NAND2_X1 U21893 ( .A1(n14153), .A2(n19911), .ZN(n19830) );
  INV_X1 U21894 ( .A(n20295), .ZN(n19829) );
  NAND3_X1 U21895 ( .A1(n19830), .A2(n19829), .A3(n19908), .ZN(n19831) );
  NAND3_X1 U21896 ( .A1(n19832), .A2(n19914), .A3(n19831), .ZN(n20298) );
  AOI22_X1 U21897 ( .A1(n20298), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n20297), .B2(n19900), .ZN(n19833) );
  OAI211_X1 U21898 ( .C1(n19903), .C2(n20306), .A(n19834), .B(n19833), .ZN(
        P2_U3103) );
  NOR3_X2 U21899 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19891), .A3(
        n19847), .ZN(n20301) );
  AOI22_X1 U21900 ( .A1(n20308), .A2(n19907), .B1(n19906), .B2(n20301), .ZN(
        n19844) );
  OAI21_X1 U21901 ( .B1(n19836), .B2(n19894), .A(n19880), .ZN(n19842) );
  NOR2_X1 U21902 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19847), .ZN(
        n19839) );
  AOI21_X1 U21903 ( .B1(n14152), .B2(n19911), .A(n20301), .ZN(n19837) );
  NAND2_X1 U21904 ( .A1(n19865), .A2(n19837), .ZN(n19838) );
  OAI211_X1 U21905 ( .C1(n19842), .C2(n19839), .A(n19914), .B(n19838), .ZN(
        n20303) );
  INV_X1 U21906 ( .A(n19839), .ZN(n19841) );
  OAI21_X1 U21907 ( .B1(n14152), .B2(n20301), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19840) );
  OAI21_X1 U21908 ( .B1(n19842), .B2(n19841), .A(n19840), .ZN(n20302) );
  AOI22_X1 U21909 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20303), .B1(
        n19722), .B2(n20302), .ZN(n19843) );
  OAI211_X1 U21910 ( .C1(n19921), .C2(n20306), .A(n19844), .B(n19843), .ZN(
        P2_U3095) );
  NOR2_X1 U21911 ( .A1(n19847), .A2(n19905), .ZN(n20307) );
  AOI22_X1 U21912 ( .A1(n20308), .A2(n19900), .B1(n19906), .B2(n20307), .ZN(
        n19859) );
  OAI21_X1 U21913 ( .B1(n20315), .B2(n20308), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19848) );
  NAND2_X1 U21914 ( .A1(n19848), .A2(n19880), .ZN(n19857) );
  NOR2_X1 U21915 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19849), .ZN(
        n19854) );
  INV_X1 U21916 ( .A(n14146), .ZN(n19852) );
  INV_X1 U21917 ( .A(n19911), .ZN(n19851) );
  OAI21_X1 U21918 ( .B1(n19880), .B2(n20307), .A(n19914), .ZN(n19850) );
  OAI21_X1 U21919 ( .B1(n19852), .B2(n19851), .A(n19850), .ZN(n19853) );
  INV_X1 U21920 ( .A(n19854), .ZN(n19856) );
  OAI21_X1 U21921 ( .B1(n14146), .B2(n20307), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19855) );
  AOI22_X1 U21922 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20310), .B1(
        n19722), .B2(n20309), .ZN(n19858) );
  OAI211_X1 U21923 ( .C1(n19903), .C2(n20313), .A(n19859), .B(n19858), .ZN(
        P2_U3087) );
  NOR2_X1 U21924 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19890) );
  INV_X1 U21925 ( .A(n19890), .ZN(n19904) );
  NOR2_X1 U21926 ( .A1(n19904), .A2(n19861), .ZN(n20314) );
  AOI22_X1 U21927 ( .A1(n20315), .A2(n19900), .B1(n20314), .B2(n19906), .ZN(
        n19871) );
  OAI21_X1 U21928 ( .B1(n19863), .B2(n19862), .A(n19880), .ZN(n19869) );
  NAND2_X1 U21929 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19890), .ZN(
        n19872) );
  INV_X1 U21930 ( .A(n19872), .ZN(n19867) );
  AOI21_X1 U21931 ( .B1(n14150), .B2(n19911), .A(n20314), .ZN(n19864) );
  NAND2_X1 U21932 ( .A1(n19865), .A2(n19864), .ZN(n19866) );
  OAI211_X1 U21933 ( .C1(n19869), .C2(n19867), .A(n19914), .B(n19866), .ZN(
        n20317) );
  OAI21_X1 U21934 ( .B1(n14150), .B2(n20314), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19868) );
  OAI21_X1 U21935 ( .B1(n19869), .B2(n19872), .A(n19868), .ZN(n20316) );
  AOI22_X1 U21936 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20317), .B1(
        n19722), .B2(n20316), .ZN(n19870) );
  OAI211_X1 U21937 ( .C1(n19903), .C2(n20326), .A(n19871), .B(n19870), .ZN(
        P2_U3079) );
  NOR2_X1 U21938 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19872), .ZN(
        n20320) );
  OAI21_X1 U21939 ( .B1(n14148), .B2(n20320), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19875) );
  AND2_X1 U21940 ( .A1(n19890), .A2(n19873), .ZN(n19878) );
  INV_X1 U21941 ( .A(n19878), .ZN(n19874) );
  NAND2_X1 U21942 ( .A1(n19875), .A2(n19874), .ZN(n20321) );
  AOI22_X1 U21943 ( .A1(n20321), .A2(n19722), .B1(n19906), .B2(n20320), .ZN(
        n19886) );
  AOI21_X1 U21944 ( .B1(n14148), .B2(n19876), .A(n20320), .ZN(n19882) );
  INV_X1 U21945 ( .A(n19877), .ZN(n19879) );
  AOI21_X1 U21946 ( .B1(n19888), .B2(n19879), .A(n19878), .ZN(n19881) );
  MUX2_X1 U21947 ( .A(n19882), .B(n19881), .S(n19880), .Z(n19883) );
  OR2_X1 U21948 ( .A1(n19883), .A2(n20234), .ZN(n20323) );
  NOR2_X2 U21949 ( .A1(n19895), .A2(n19884), .ZN(n20330) );
  AOI22_X1 U21950 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20323), .B1(
        n20330), .B2(n19907), .ZN(n19885) );
  OAI211_X1 U21951 ( .C1(n19921), .C2(n20326), .A(n19886), .B(n19885), .ZN(
        P2_U3071) );
  NAND2_X1 U21952 ( .A1(n19890), .A2(n19889), .ZN(n19893) );
  NOR3_X2 U21953 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19891), .A3(
        n19904), .ZN(n20328) );
  OAI21_X1 U21954 ( .B1(n14158), .B2(n20328), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19892) );
  OAI21_X1 U21955 ( .B1(n19893), .B2(n19908), .A(n19892), .ZN(n20329) );
  AOI22_X1 U21956 ( .A1(n20329), .A2(n19722), .B1(n19906), .B2(n20328), .ZN(
        n19902) );
  OAI22_X1 U21957 ( .A1(n19895), .A2(n19894), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19904), .ZN(n19899) );
  NAND2_X1 U21958 ( .A1(n14158), .A2(n19911), .ZN(n19897) );
  INV_X1 U21959 ( .A(n20328), .ZN(n19896) );
  NAND3_X1 U21960 ( .A1(n19897), .A2(n19896), .A3(n19908), .ZN(n19898) );
  NAND3_X1 U21961 ( .A1(n19899), .A2(n19914), .A3(n19898), .ZN(n20331) );
  AOI22_X1 U21962 ( .A1(n20331), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n20330), .B2(n19900), .ZN(n19901) );
  OAI211_X1 U21963 ( .C1(n19903), .C2(n20334), .A(n19902), .B(n19901), .ZN(
        P2_U3063) );
  INV_X1 U21964 ( .A(n20344), .ZN(n20215) );
  NOR2_X1 U21965 ( .A1(n19905), .A2(n19904), .ZN(n20335) );
  AOI22_X1 U21966 ( .A1(n19907), .A2(n20215), .B1(n19906), .B2(n20335), .ZN(
        n19920) );
  AOI21_X1 U21967 ( .B1(n20334), .B2(n20344), .A(n22239), .ZN(n19909) );
  NOR2_X1 U21968 ( .A1(n19909), .A2(n19908), .ZN(n19916) );
  INV_X1 U21969 ( .A(n20238), .ZN(n19913) );
  AOI21_X1 U21970 ( .B1(n14162), .B2(n19911), .A(n19910), .ZN(n19912) );
  AOI21_X1 U21971 ( .B1(n19916), .B2(n19913), .A(n19912), .ZN(n19915) );
  OAI21_X1 U21972 ( .B1(n20238), .B2(n20335), .A(n19916), .ZN(n19918) );
  OAI21_X1 U21973 ( .B1(n14162), .B2(n20335), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19917) );
  NAND2_X1 U21974 ( .A1(n19918), .A2(n19917), .ZN(n20340) );
  AOI22_X1 U21975 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n19722), .ZN(n19919) );
  OAI211_X1 U21976 ( .C1(n19921), .C2(n20334), .A(n19920), .B(n19919), .ZN(
        P2_U3055) );
  AOI22_X1 U21977 ( .A1(n20223), .A2(n19922), .B1(n20221), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n19928) );
  AOI22_X1 U21978 ( .A1(n20225), .A2(BUF2_REG_22__SCAN_IN), .B1(n20224), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n19927) );
  INV_X1 U21979 ( .A(n19923), .ZN(n19925) );
  AOI22_X1 U21980 ( .A1(n19925), .A2(n20123), .B1(n20169), .B2(n19924), .ZN(
        n19926) );
  NAND3_X1 U21981 ( .A1(n19928), .A2(n19927), .A3(n19926), .ZN(P2_U2897) );
  OAI222_X1 U21982 ( .A1(n19931), .A2(n19979), .B1(n19930), .B2(n19929), .C1(
        n20176), .C2(n19932), .ZN(P2_U2913) );
  AOI22_X1 U21983 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n20241), .B1(
        BUF1_REG_22__SCAN_IN), .B2(n20240), .ZN(n19964) );
  NOR2_X2 U21984 ( .A1(n14700), .A2(n20236), .ZN(n19967) );
  AOI22_X1 U21985 ( .A1(n20239), .A2(n19933), .B1(n20238), .B2(n19967), .ZN(
        n19935) );
  INV_X1 U21986 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n21231) );
  OAI22_X1 U21987 ( .A1(n21231), .A2(n20080), .B1(n20623), .B2(n20081), .ZN(
        n19961) );
  AOI22_X1 U21988 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20242), .B1(
        n20246), .B2(n19961), .ZN(n19934) );
  OAI211_X1 U21989 ( .C1(n19964), .C2(n20344), .A(n19935), .B(n19934), .ZN(
        P2_U3174) );
  INV_X1 U21990 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n19938) );
  AOI22_X1 U21991 ( .A1(n20254), .A2(n19961), .B1(n19967), .B2(n20245), .ZN(
        n19937) );
  AOI22_X1 U21992 ( .A1(n19933), .A2(n20247), .B1(n20246), .B2(n19968), .ZN(
        n19936) );
  OAI211_X1 U21993 ( .C1(n19938), .C2(n20250), .A(n19937), .B(n19936), .ZN(
        P2_U3166) );
  INV_X1 U21994 ( .A(n19961), .ZN(n19971) );
  AOI22_X1 U21995 ( .A1(n20253), .A2(n19933), .B1(n19967), .B2(n20252), .ZN(
        n19940) );
  AOI22_X1 U21996 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20255), .B1(
        n19968), .B2(n20254), .ZN(n19939) );
  OAI211_X1 U21997 ( .C1(n19971), .C2(n20258), .A(n19940), .B(n19939), .ZN(
        P2_U3158) );
  AOI22_X1 U21998 ( .A1(n20260), .A2(n19933), .B1(n19967), .B2(n20259), .ZN(
        n19942) );
  AOI22_X1 U21999 ( .A1(n20262), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n20261), .B2(n19968), .ZN(n19941) );
  OAI211_X1 U22000 ( .C1(n19971), .C2(n20270), .A(n19942), .B(n19941), .ZN(
        P2_U3150) );
  AOI22_X1 U22001 ( .A1(n20266), .A2(n19933), .B1(n19967), .B2(n20265), .ZN(
        n19944) );
  AOI22_X1 U22002 ( .A1(n20272), .A2(n19961), .B1(n20267), .B2(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n19943) );
  OAI211_X1 U22003 ( .C1(n19964), .C2(n20270), .A(n19944), .B(n19943), .ZN(
        P2_U3142) );
  AOI22_X1 U22004 ( .A1(n19968), .A2(n20272), .B1(n19967), .B2(n20271), .ZN(
        n19946) );
  AOI22_X1 U22005 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20274), .B1(
        n19933), .B2(n20273), .ZN(n19945) );
  OAI211_X1 U22006 ( .C1(n19971), .C2(n20282), .A(n19946), .B(n19945), .ZN(
        P2_U3134) );
  AOI22_X1 U22007 ( .A1(n20284), .A2(n19961), .B1(n19967), .B2(n20277), .ZN(
        n19948) );
  AOI22_X1 U22008 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20279), .B1(
        n19933), .B2(n20278), .ZN(n19947) );
  OAI211_X1 U22009 ( .C1(n19964), .C2(n20282), .A(n19948), .B(n19947), .ZN(
        P2_U3126) );
  AOI22_X1 U22010 ( .A1(n19968), .A2(n20284), .B1(n19967), .B2(n20283), .ZN(
        n19950) );
  AOI22_X1 U22011 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20286), .B1(
        n19933), .B2(n20285), .ZN(n19949) );
  OAI211_X1 U22012 ( .C1(n19971), .C2(n20294), .A(n19950), .B(n19949), .ZN(
        P2_U3118) );
  AOI22_X1 U22013 ( .A1(n20290), .A2(n19933), .B1(n20289), .B2(n19967), .ZN(
        n19952) );
  AOI22_X1 U22014 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20291), .B1(
        n20297), .B2(n19961), .ZN(n19951) );
  OAI211_X1 U22015 ( .C1(n19964), .C2(n20294), .A(n19952), .B(n19951), .ZN(
        P2_U3110) );
  AOI22_X1 U22016 ( .A1(n20296), .A2(n19933), .B1(n19967), .B2(n20295), .ZN(
        n19954) );
  AOI22_X1 U22017 ( .A1(n20298), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n20297), .B2(n19968), .ZN(n19953) );
  OAI211_X1 U22018 ( .C1(n19971), .C2(n20306), .A(n19954), .B(n19953), .ZN(
        P2_U3102) );
  AOI22_X1 U22019 ( .A1(n20308), .A2(n19961), .B1(n19967), .B2(n20301), .ZN(
        n19956) );
  AOI22_X1 U22020 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20303), .B1(
        n19933), .B2(n20302), .ZN(n19955) );
  OAI211_X1 U22021 ( .C1(n19964), .C2(n20306), .A(n19956), .B(n19955), .ZN(
        P2_U3094) );
  AOI22_X1 U22022 ( .A1(n20308), .A2(n19968), .B1(n19967), .B2(n20307), .ZN(
        n19958) );
  AOI22_X1 U22023 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20310), .B1(
        n19933), .B2(n20309), .ZN(n19957) );
  OAI211_X1 U22024 ( .C1(n19971), .C2(n20313), .A(n19958), .B(n19957), .ZN(
        P2_U3086) );
  AOI22_X1 U22025 ( .A1(n20315), .A2(n19968), .B1(n20314), .B2(n19967), .ZN(
        n19960) );
  AOI22_X1 U22026 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20317), .B1(
        n19933), .B2(n20316), .ZN(n19959) );
  OAI211_X1 U22027 ( .C1(n19971), .C2(n20326), .A(n19960), .B(n19959), .ZN(
        P2_U3078) );
  AOI22_X1 U22028 ( .A1(n20321), .A2(n19933), .B1(n19967), .B2(n20320), .ZN(
        n19963) );
  AOI22_X1 U22029 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20323), .B1(
        n20330), .B2(n19961), .ZN(n19962) );
  OAI211_X1 U22030 ( .C1(n19964), .C2(n20326), .A(n19963), .B(n19962), .ZN(
        P2_U3070) );
  AOI22_X1 U22031 ( .A1(n20329), .A2(n19933), .B1(n19967), .B2(n20328), .ZN(
        n19966) );
  AOI22_X1 U22032 ( .A1(n20331), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n20330), .B2(n19968), .ZN(n19965) );
  OAI211_X1 U22033 ( .C1(n19971), .C2(n20334), .A(n19966), .B(n19965), .ZN(
        P2_U3062) );
  INV_X1 U22034 ( .A(n20334), .ZN(n20338) );
  AOI22_X1 U22035 ( .A1(n20338), .A2(n19968), .B1(n19967), .B2(n20335), .ZN(
        n19970) );
  AOI22_X1 U22036 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n19933), .ZN(n19969) );
  OAI211_X1 U22037 ( .C1(n19971), .C2(n20344), .A(n19970), .B(n19969), .ZN(
        P2_U3054) );
  INV_X1 U22038 ( .A(n19980), .ZN(n19973) );
  AOI22_X1 U22039 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n20221), .B1(n19973), .B2(
        n19972), .ZN(n19977) );
  OR3_X1 U22040 ( .A1(n19975), .A2(n19974), .A3(n20228), .ZN(n19976) );
  OAI211_X1 U22041 ( .C1(n19979), .C2(n19978), .A(n19977), .B(n19976), .ZN(
        P2_U2914) );
  INV_X1 U22042 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n21181) );
  OAI22_X1 U22043 ( .A1(n21181), .A2(n20080), .B1(n20605), .B2(n20081), .ZN(
        n20011) );
  NOR2_X2 U22044 ( .A1(n19982), .A2(n20236), .ZN(n20015) );
  AOI22_X1 U22045 ( .A1(n20239), .A2(n19981), .B1(n20238), .B2(n20015), .ZN(
        n19984) );
  AOI22_X1 U22046 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20240), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20241), .ZN(n20014) );
  INV_X1 U22047 ( .A(n20014), .ZN(n20016) );
  AOI22_X1 U22048 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20242), .B1(
        n20246), .B2(n20016), .ZN(n19983) );
  OAI211_X1 U22049 ( .C1(n20019), .C2(n20344), .A(n19984), .B(n19983), .ZN(
        P2_U3173) );
  AOI22_X1 U22050 ( .A1(n20016), .A2(n20254), .B1(n20015), .B2(n20245), .ZN(
        n19986) );
  AOI22_X1 U22051 ( .A1(n19981), .A2(n20247), .B1(n20246), .B2(n20011), .ZN(
        n19985) );
  OAI211_X1 U22052 ( .C1(n16212), .C2(n20250), .A(n19986), .B(n19985), .ZN(
        P2_U3165) );
  AOI22_X1 U22053 ( .A1(n20253), .A2(n19981), .B1(n20015), .B2(n20252), .ZN(
        n19988) );
  AOI22_X1 U22054 ( .A1(n20255), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n20254), .B2(n20011), .ZN(n19987) );
  OAI211_X1 U22055 ( .C1(n20014), .C2(n20258), .A(n19988), .B(n19987), .ZN(
        P2_U3157) );
  AOI22_X1 U22056 ( .A1(n20260), .A2(n19981), .B1(n20015), .B2(n20259), .ZN(
        n19990) );
  AOI22_X1 U22057 ( .A1(n20262), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n20261), .B2(n20011), .ZN(n19989) );
  OAI211_X1 U22058 ( .C1(n20014), .C2(n20270), .A(n19990), .B(n19989), .ZN(
        P2_U3149) );
  AOI22_X1 U22059 ( .A1(n20266), .A2(n19981), .B1(n20015), .B2(n20265), .ZN(
        n19992) );
  AOI22_X1 U22060 ( .A1(n20016), .A2(n20272), .B1(n20267), .B2(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n19991) );
  OAI211_X1 U22061 ( .C1(n20019), .C2(n20270), .A(n19992), .B(n19991), .ZN(
        P2_U3141) );
  AOI22_X1 U22062 ( .A1(n20190), .A2(n20016), .B1(n20015), .B2(n20271), .ZN(
        n19994) );
  AOI22_X1 U22063 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20274), .B1(
        n19981), .B2(n20273), .ZN(n19993) );
  OAI211_X1 U22064 ( .C1(n20019), .C2(n20193), .A(n19994), .B(n19993), .ZN(
        P2_U3133) );
  AOI22_X1 U22065 ( .A1(n20016), .A2(n20284), .B1(n20015), .B2(n20277), .ZN(
        n19996) );
  AOI22_X1 U22066 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20279), .B1(
        n19981), .B2(n20278), .ZN(n19995) );
  OAI211_X1 U22067 ( .C1(n20019), .C2(n20282), .A(n19996), .B(n19995), .ZN(
        P2_U3125) );
  AOI22_X1 U22068 ( .A1(n20284), .A2(n20011), .B1(n20015), .B2(n20283), .ZN(
        n19998) );
  AOI22_X1 U22069 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20286), .B1(
        n19981), .B2(n20285), .ZN(n19997) );
  OAI211_X1 U22070 ( .C1(n20014), .C2(n20294), .A(n19998), .B(n19997), .ZN(
        P2_U3117) );
  AOI22_X1 U22071 ( .A1(n20290), .A2(n19981), .B1(n20289), .B2(n20015), .ZN(
        n20000) );
  AOI22_X1 U22072 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20291), .B1(
        n20297), .B2(n20016), .ZN(n19999) );
  OAI211_X1 U22073 ( .C1(n20019), .C2(n20294), .A(n20000), .B(n19999), .ZN(
        P2_U3109) );
  AOI22_X1 U22074 ( .A1(n20296), .A2(n19981), .B1(n20015), .B2(n20295), .ZN(
        n20002) );
  AOI22_X1 U22075 ( .A1(n20298), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n20297), .B2(n20011), .ZN(n20001) );
  OAI211_X1 U22076 ( .C1(n20014), .C2(n20306), .A(n20002), .B(n20001), .ZN(
        P2_U3101) );
  AOI22_X1 U22077 ( .A1(n20308), .A2(n20016), .B1(n20015), .B2(n20301), .ZN(
        n20004) );
  AOI22_X1 U22078 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20303), .B1(
        n19981), .B2(n20302), .ZN(n20003) );
  OAI211_X1 U22079 ( .C1(n20019), .C2(n20306), .A(n20004), .B(n20003), .ZN(
        P2_U3093) );
  AOI22_X1 U22080 ( .A1(n20308), .A2(n20011), .B1(n20015), .B2(n20307), .ZN(
        n20006) );
  AOI22_X1 U22081 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20310), .B1(
        n19981), .B2(n20309), .ZN(n20005) );
  OAI211_X1 U22082 ( .C1(n20014), .C2(n20313), .A(n20006), .B(n20005), .ZN(
        P2_U3085) );
  AOI22_X1 U22083 ( .A1(n20315), .A2(n20011), .B1(n20314), .B2(n20015), .ZN(
        n20008) );
  AOI22_X1 U22084 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20317), .B1(
        n19981), .B2(n20316), .ZN(n20007) );
  OAI211_X1 U22085 ( .C1(n20014), .C2(n20326), .A(n20008), .B(n20007), .ZN(
        P2_U3077) );
  AOI22_X1 U22086 ( .A1(n20321), .A2(n19981), .B1(n20015), .B2(n20320), .ZN(
        n20010) );
  AOI22_X1 U22087 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20323), .B1(
        n20330), .B2(n20016), .ZN(n20009) );
  OAI211_X1 U22088 ( .C1(n20019), .C2(n20326), .A(n20010), .B(n20009), .ZN(
        P2_U3069) );
  AOI22_X1 U22089 ( .A1(n20329), .A2(n19981), .B1(n20015), .B2(n20328), .ZN(
        n20013) );
  AOI22_X1 U22090 ( .A1(n20331), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n20330), .B2(n20011), .ZN(n20012) );
  OAI211_X1 U22091 ( .C1(n20014), .C2(n20334), .A(n20013), .B(n20012), .ZN(
        P2_U3061) );
  AOI22_X1 U22092 ( .A1(n20016), .A2(n20215), .B1(n20015), .B2(n20335), .ZN(
        n20018) );
  AOI22_X1 U22093 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n19981), .ZN(n20017) );
  OAI211_X1 U22094 ( .C1(n20019), .C2(n20334), .A(n20018), .B(n20017), .ZN(
        P2_U3053) );
  AOI22_X1 U22095 ( .A1(n20223), .A2(n20020), .B1(n20221), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n20027) );
  AOI22_X1 U22096 ( .A1(n20225), .A2(BUF2_REG_20__SCAN_IN), .B1(n20224), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n20026) );
  INV_X1 U22097 ( .A(n20021), .ZN(n20024) );
  INV_X1 U22098 ( .A(n20022), .ZN(n20023) );
  AOI22_X1 U22099 ( .A1(n20024), .A2(n20123), .B1(n20023), .B2(n20169), .ZN(
        n20025) );
  NAND3_X1 U22100 ( .A1(n20027), .A2(n20026), .A3(n20025), .ZN(P2_U2899) );
  AOI22_X1 U22101 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20240), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20241), .ZN(n20069) );
  NOR2_X2 U22102 ( .A1(n20030), .A2(n20236), .ZN(n20065) );
  AOI22_X1 U22103 ( .A1(n20239), .A2(n20029), .B1(n20238), .B2(n20065), .ZN(
        n20032) );
  AOI22_X1 U22104 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n20241), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n20240), .ZN(n20064) );
  INV_X1 U22105 ( .A(n20064), .ZN(n20066) );
  AOI22_X1 U22106 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20242), .B1(
        n20246), .B2(n20066), .ZN(n20031) );
  OAI211_X1 U22107 ( .C1(n20069), .C2(n20344), .A(n20032), .B(n20031), .ZN(
        P2_U3172) );
  INV_X1 U22108 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20035) );
  AOI22_X1 U22109 ( .A1(n20066), .A2(n20254), .B1(n20065), .B2(n20245), .ZN(
        n20034) );
  INV_X1 U22110 ( .A(n20069), .ZN(n20061) );
  AOI22_X1 U22111 ( .A1(n20029), .A2(n20247), .B1(n20246), .B2(n20061), .ZN(
        n20033) );
  OAI211_X1 U22112 ( .C1(n20035), .C2(n20250), .A(n20034), .B(n20033), .ZN(
        P2_U3164) );
  AOI22_X1 U22113 ( .A1(n20253), .A2(n20029), .B1(n20065), .B2(n20252), .ZN(
        n20037) );
  AOI22_X1 U22114 ( .A1(n20061), .A2(n20254), .B1(n20255), .B2(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n20036) );
  OAI211_X1 U22115 ( .C1(n20064), .C2(n20258), .A(n20037), .B(n20036), .ZN(
        P2_U3156) );
  AOI22_X1 U22116 ( .A1(n20260), .A2(n20029), .B1(n20065), .B2(n20259), .ZN(
        n20039) );
  AOI22_X1 U22117 ( .A1(n20262), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n20261), .B2(n20061), .ZN(n20038) );
  OAI211_X1 U22118 ( .C1(n20064), .C2(n20270), .A(n20039), .B(n20038), .ZN(
        P2_U3148) );
  AOI22_X1 U22119 ( .A1(n20266), .A2(n20029), .B1(n20065), .B2(n20265), .ZN(
        n20042) );
  AOI22_X1 U22120 ( .A1(n20040), .A2(n20061), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n20267), .ZN(n20041) );
  OAI211_X1 U22121 ( .C1(n20064), .C2(n20193), .A(n20042), .B(n20041), .ZN(
        P2_U3140) );
  AOI22_X1 U22122 ( .A1(n20190), .A2(n20066), .B1(n20065), .B2(n20271), .ZN(
        n20044) );
  AOI22_X1 U22123 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20274), .B1(
        n20029), .B2(n20273), .ZN(n20043) );
  OAI211_X1 U22124 ( .C1(n20069), .C2(n20193), .A(n20044), .B(n20043), .ZN(
        P2_U3132) );
  AOI22_X1 U22125 ( .A1(n20066), .A2(n20284), .B1(n20065), .B2(n20277), .ZN(
        n20046) );
  AOI22_X1 U22126 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20279), .B1(
        n20029), .B2(n20278), .ZN(n20045) );
  OAI211_X1 U22127 ( .C1(n20069), .C2(n20282), .A(n20046), .B(n20045), .ZN(
        P2_U3124) );
  AOI22_X1 U22128 ( .A1(n20061), .A2(n20284), .B1(n20065), .B2(n20283), .ZN(
        n20048) );
  AOI22_X1 U22129 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20286), .B1(
        n20029), .B2(n20285), .ZN(n20047) );
  OAI211_X1 U22130 ( .C1(n20064), .C2(n20294), .A(n20048), .B(n20047), .ZN(
        P2_U3116) );
  AOI22_X1 U22131 ( .A1(n20290), .A2(n20029), .B1(n20289), .B2(n20065), .ZN(
        n20050) );
  AOI22_X1 U22132 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20291), .B1(
        n20297), .B2(n20066), .ZN(n20049) );
  OAI211_X1 U22133 ( .C1(n20069), .C2(n20294), .A(n20050), .B(n20049), .ZN(
        P2_U3108) );
  AOI22_X1 U22134 ( .A1(n20296), .A2(n20029), .B1(n20065), .B2(n20295), .ZN(
        n20052) );
  AOI22_X1 U22135 ( .A1(n20298), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n20297), .B2(n20061), .ZN(n20051) );
  OAI211_X1 U22136 ( .C1(n20064), .C2(n20306), .A(n20052), .B(n20051), .ZN(
        P2_U3100) );
  AOI22_X1 U22137 ( .A1(n20308), .A2(n20066), .B1(n20065), .B2(n20301), .ZN(
        n20054) );
  AOI22_X1 U22138 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20303), .B1(
        n20029), .B2(n20302), .ZN(n20053) );
  OAI211_X1 U22139 ( .C1(n20069), .C2(n20306), .A(n20054), .B(n20053), .ZN(
        P2_U3092) );
  AOI22_X1 U22140 ( .A1(n20308), .A2(n20061), .B1(n20065), .B2(n20307), .ZN(
        n20056) );
  AOI22_X1 U22141 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20310), .B1(
        n20029), .B2(n20309), .ZN(n20055) );
  OAI211_X1 U22142 ( .C1(n20064), .C2(n20313), .A(n20056), .B(n20055), .ZN(
        P2_U3084) );
  AOI22_X1 U22143 ( .A1(n20315), .A2(n20061), .B1(n20314), .B2(n20065), .ZN(
        n20058) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20317), .B1(
        n20029), .B2(n20316), .ZN(n20057) );
  OAI211_X1 U22145 ( .C1(n20064), .C2(n20326), .A(n20058), .B(n20057), .ZN(
        P2_U3076) );
  AOI22_X1 U22146 ( .A1(n20321), .A2(n20029), .B1(n20065), .B2(n20320), .ZN(
        n20060) );
  AOI22_X1 U22147 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20323), .B1(
        n20330), .B2(n20066), .ZN(n20059) );
  OAI211_X1 U22148 ( .C1(n20069), .C2(n20326), .A(n20060), .B(n20059), .ZN(
        P2_U3068) );
  AOI22_X1 U22149 ( .A1(n20329), .A2(n20029), .B1(n20065), .B2(n20328), .ZN(
        n20063) );
  AOI22_X1 U22150 ( .A1(n20331), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n20330), .B2(n20061), .ZN(n20062) );
  OAI211_X1 U22151 ( .C1(n20064), .C2(n20334), .A(n20063), .B(n20062), .ZN(
        P2_U3060) );
  AOI22_X1 U22152 ( .A1(n20066), .A2(n20215), .B1(n20065), .B2(n20335), .ZN(
        n20068) );
  AOI22_X1 U22153 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n20029), .ZN(n20067) );
  OAI211_X1 U22154 ( .C1(n20069), .C2(n20334), .A(n20068), .B(n20067), .ZN(
        P2_U3052) );
  AOI22_X1 U22155 ( .A1(n20070), .A2(n20169), .B1(n20221), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n20076) );
  AOI21_X1 U22156 ( .B1(n20073), .B2(n20072), .A(n20071), .ZN(n20074) );
  OR2_X1 U22157 ( .A1(n20074), .A2(n20228), .ZN(n20075) );
  OAI211_X1 U22158 ( .C1(n20077), .C2(n20176), .A(n20076), .B(n20075), .ZN(
        P2_U2916) );
  AOI22_X1 U22159 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n20241), .B1(
        BUF1_REG_19__SCAN_IN), .B2(n20240), .ZN(n20112) );
  NOR2_X2 U22160 ( .A1(n20079), .A2(n20236), .ZN(n20115) );
  AOI22_X1 U22161 ( .A1(n20239), .A2(n20078), .B1(n20238), .B2(n20115), .ZN(
        n20083) );
  INV_X1 U22162 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n21252) );
  OAI22_X1 U22163 ( .A1(n20617), .A2(n20081), .B1(n21252), .B2(n20080), .ZN(
        n20109) );
  AOI22_X1 U22164 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20242), .B1(
        n20246), .B2(n20109), .ZN(n20082) );
  OAI211_X1 U22165 ( .C1(n20112), .C2(n20344), .A(n20083), .B(n20082), .ZN(
        P2_U3171) );
  INV_X1 U22166 ( .A(n20112), .ZN(n20116) );
  AOI22_X1 U22167 ( .A1(n20246), .A2(n20116), .B1(n20115), .B2(n20245), .ZN(
        n20085) );
  AOI22_X1 U22168 ( .A1(n20078), .A2(n20247), .B1(n20254), .B2(n20109), .ZN(
        n20084) );
  OAI211_X1 U22169 ( .C1(n20086), .C2(n20250), .A(n20085), .B(n20084), .ZN(
        P2_U3163) );
  AOI22_X1 U22170 ( .A1(n20253), .A2(n20078), .B1(n20115), .B2(n20252), .ZN(
        n20088) );
  AOI22_X1 U22171 ( .A1(n20255), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n20254), .B2(n20116), .ZN(n20087) );
  OAI211_X1 U22172 ( .C1(n20119), .C2(n20258), .A(n20088), .B(n20087), .ZN(
        P2_U3155) );
  AOI22_X1 U22173 ( .A1(n20260), .A2(n20078), .B1(n20115), .B2(n20259), .ZN(
        n20090) );
  AOI22_X1 U22174 ( .A1(n20262), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n20261), .B2(n20116), .ZN(n20089) );
  OAI211_X1 U22175 ( .C1(n20119), .C2(n20270), .A(n20090), .B(n20089), .ZN(
        P2_U3147) );
  AOI22_X1 U22176 ( .A1(n20266), .A2(n20078), .B1(n20115), .B2(n20265), .ZN(
        n20092) );
  AOI22_X1 U22177 ( .A1(n20272), .A2(n20109), .B1(n20267), .B2(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n20091) );
  OAI211_X1 U22178 ( .C1(n20112), .C2(n20270), .A(n20092), .B(n20091), .ZN(
        P2_U3139) );
  AOI22_X1 U22179 ( .A1(n20190), .A2(n20109), .B1(n20115), .B2(n20271), .ZN(
        n20094) );
  AOI22_X1 U22180 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20274), .B1(
        n20078), .B2(n20273), .ZN(n20093) );
  OAI211_X1 U22181 ( .C1(n20112), .C2(n20193), .A(n20094), .B(n20093), .ZN(
        P2_U3131) );
  AOI22_X1 U22182 ( .A1(n20284), .A2(n20109), .B1(n20115), .B2(n20277), .ZN(
        n20096) );
  AOI22_X1 U22183 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20279), .B1(
        n20078), .B2(n20278), .ZN(n20095) );
  OAI211_X1 U22184 ( .C1(n20112), .C2(n20282), .A(n20096), .B(n20095), .ZN(
        P2_U3123) );
  AOI22_X1 U22185 ( .A1(n20284), .A2(n20116), .B1(n20115), .B2(n20283), .ZN(
        n20098) );
  AOI22_X1 U22186 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20286), .B1(
        n20078), .B2(n20285), .ZN(n20097) );
  OAI211_X1 U22187 ( .C1(n20119), .C2(n20294), .A(n20098), .B(n20097), .ZN(
        P2_U3115) );
  AOI22_X1 U22188 ( .A1(n20290), .A2(n20078), .B1(n20289), .B2(n20115), .ZN(
        n20100) );
  AOI22_X1 U22189 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20291), .B1(
        n20297), .B2(n20109), .ZN(n20099) );
  OAI211_X1 U22190 ( .C1(n20112), .C2(n20294), .A(n20100), .B(n20099), .ZN(
        P2_U3107) );
  AOI22_X1 U22191 ( .A1(n20296), .A2(n20078), .B1(n20115), .B2(n20295), .ZN(
        n20102) );
  AOI22_X1 U22192 ( .A1(n20298), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n20297), .B2(n20116), .ZN(n20101) );
  OAI211_X1 U22193 ( .C1(n20119), .C2(n20306), .A(n20102), .B(n20101), .ZN(
        P2_U3099) );
  AOI22_X1 U22194 ( .A1(n20308), .A2(n20109), .B1(n20115), .B2(n20301), .ZN(
        n20104) );
  AOI22_X1 U22195 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20303), .B1(
        n20078), .B2(n20302), .ZN(n20103) );
  OAI211_X1 U22196 ( .C1(n20112), .C2(n20306), .A(n20104), .B(n20103), .ZN(
        P2_U3091) );
  AOI22_X1 U22197 ( .A1(n20308), .A2(n20116), .B1(n20115), .B2(n20307), .ZN(
        n20106) );
  AOI22_X1 U22198 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20310), .B1(
        n20078), .B2(n20309), .ZN(n20105) );
  OAI211_X1 U22199 ( .C1(n20119), .C2(n20313), .A(n20106), .B(n20105), .ZN(
        P2_U3083) );
  AOI22_X1 U22200 ( .A1(n20315), .A2(n20116), .B1(n20314), .B2(n20115), .ZN(
        n20108) );
  AOI22_X1 U22201 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20317), .B1(
        n20078), .B2(n20316), .ZN(n20107) );
  OAI211_X1 U22202 ( .C1(n20119), .C2(n20326), .A(n20108), .B(n20107), .ZN(
        P2_U3075) );
  AOI22_X1 U22203 ( .A1(n20321), .A2(n20078), .B1(n20115), .B2(n20320), .ZN(
        n20111) );
  AOI22_X1 U22204 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20323), .B1(
        n20330), .B2(n20109), .ZN(n20110) );
  OAI211_X1 U22205 ( .C1(n20112), .C2(n20326), .A(n20111), .B(n20110), .ZN(
        P2_U3067) );
  AOI22_X1 U22206 ( .A1(n20329), .A2(n20078), .B1(n20115), .B2(n20328), .ZN(
        n20114) );
  AOI22_X1 U22207 ( .A1(n20331), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n20330), .B2(n20116), .ZN(n20113) );
  OAI211_X1 U22208 ( .C1(n20119), .C2(n20334), .A(n20114), .B(n20113), .ZN(
        P2_U3059) );
  AOI22_X1 U22209 ( .A1(n20338), .A2(n20116), .B1(n20115), .B2(n20335), .ZN(
        n20118) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n20078), .ZN(n20117) );
  OAI211_X1 U22211 ( .C1(n20119), .C2(n20344), .A(n20118), .B(n20117), .ZN(
        P2_U3051) );
  AOI22_X1 U22212 ( .A1(n20223), .A2(n20120), .B1(n20221), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n20127) );
  AOI22_X1 U22213 ( .A1(n20225), .A2(BUF2_REG_18__SCAN_IN), .B1(n20224), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n20126) );
  INV_X1 U22214 ( .A(n20121), .ZN(n20122) );
  AOI22_X1 U22215 ( .A1(n20124), .A2(n20123), .B1(n20169), .B2(n20122), .ZN(
        n20125) );
  NAND3_X1 U22216 ( .A1(n20127), .A2(n20126), .A3(n20125), .ZN(P2_U2901) );
  AOI22_X1 U22217 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20240), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20241), .ZN(n20167) );
  NOR2_X2 U22218 ( .A1(n20128), .A2(n20234), .ZN(n20164) );
  NOR2_X2 U22219 ( .A1(n14257), .A2(n20236), .ZN(n20162) );
  AOI22_X1 U22220 ( .A1(n20239), .A2(n20164), .B1(n20238), .B2(n20162), .ZN(
        n20130) );
  AOI22_X1 U22221 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20240), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20241), .ZN(n20161) );
  INV_X1 U22222 ( .A(n20161), .ZN(n20163) );
  AOI22_X1 U22223 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20242), .B1(
        n20246), .B2(n20163), .ZN(n20129) );
  OAI211_X1 U22224 ( .C1(n20167), .C2(n20344), .A(n20130), .B(n20129), .ZN(
        P2_U3170) );
  INV_X1 U22225 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20133) );
  AOI22_X1 U22226 ( .A1(n20163), .A2(n20254), .B1(n20162), .B2(n20245), .ZN(
        n20132) );
  INV_X1 U22227 ( .A(n20167), .ZN(n20158) );
  AOI22_X1 U22228 ( .A1(n20164), .A2(n20247), .B1(n20246), .B2(n20158), .ZN(
        n20131) );
  OAI211_X1 U22229 ( .C1(n20133), .C2(n20250), .A(n20132), .B(n20131), .ZN(
        P2_U3162) );
  AOI22_X1 U22230 ( .A1(n20253), .A2(n20164), .B1(n20162), .B2(n20252), .ZN(
        n20135) );
  AOI22_X1 U22231 ( .A1(n20158), .A2(n20254), .B1(n20255), .B2(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20134) );
  OAI211_X1 U22232 ( .C1(n20161), .C2(n20258), .A(n20135), .B(n20134), .ZN(
        P2_U3154) );
  AOI22_X1 U22233 ( .A1(n20260), .A2(n20164), .B1(n20162), .B2(n20259), .ZN(
        n20137) );
  AOI22_X1 U22234 ( .A1(n20262), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n20261), .B2(n20158), .ZN(n20136) );
  OAI211_X1 U22235 ( .C1(n20161), .C2(n20270), .A(n20137), .B(n20136), .ZN(
        P2_U3146) );
  AOI22_X1 U22236 ( .A1(n20266), .A2(n20164), .B1(n20162), .B2(n20265), .ZN(
        n20139) );
  AOI22_X1 U22237 ( .A1(n20163), .A2(n20272), .B1(n20267), .B2(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20138) );
  OAI211_X1 U22238 ( .C1(n20167), .C2(n20270), .A(n20139), .B(n20138), .ZN(
        P2_U3138) );
  AOI22_X1 U22239 ( .A1(n20190), .A2(n20163), .B1(n20162), .B2(n20271), .ZN(
        n20141) );
  AOI22_X1 U22240 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20274), .B1(
        n20164), .B2(n20273), .ZN(n20140) );
  OAI211_X1 U22241 ( .C1(n20167), .C2(n20193), .A(n20141), .B(n20140), .ZN(
        P2_U3130) );
  AOI22_X1 U22242 ( .A1(n20163), .A2(n20284), .B1(n20162), .B2(n20277), .ZN(
        n20143) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20279), .B1(
        n20164), .B2(n20278), .ZN(n20142) );
  OAI211_X1 U22244 ( .C1(n20167), .C2(n20282), .A(n20143), .B(n20142), .ZN(
        P2_U3122) );
  AOI22_X1 U22245 ( .A1(n20158), .A2(n20284), .B1(n20162), .B2(n20283), .ZN(
        n20145) );
  AOI22_X1 U22246 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20286), .B1(
        n20164), .B2(n20285), .ZN(n20144) );
  OAI211_X1 U22247 ( .C1(n20161), .C2(n20294), .A(n20145), .B(n20144), .ZN(
        P2_U3114) );
  AOI22_X1 U22248 ( .A1(n20290), .A2(n20164), .B1(n20289), .B2(n20162), .ZN(
        n20147) );
  AOI22_X1 U22249 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20291), .B1(
        n20297), .B2(n20163), .ZN(n20146) );
  OAI211_X1 U22250 ( .C1(n20167), .C2(n20294), .A(n20147), .B(n20146), .ZN(
        P2_U3106) );
  AOI22_X1 U22251 ( .A1(n20296), .A2(n20164), .B1(n20162), .B2(n20295), .ZN(
        n20149) );
  AOI22_X1 U22252 ( .A1(n20298), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n20297), .B2(n20158), .ZN(n20148) );
  OAI211_X1 U22253 ( .C1(n20161), .C2(n20306), .A(n20149), .B(n20148), .ZN(
        P2_U3098) );
  AOI22_X1 U22254 ( .A1(n20308), .A2(n20163), .B1(n20162), .B2(n20301), .ZN(
        n20151) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20303), .B1(
        n20164), .B2(n20302), .ZN(n20150) );
  OAI211_X1 U22256 ( .C1(n20167), .C2(n20306), .A(n20151), .B(n20150), .ZN(
        P2_U3090) );
  AOI22_X1 U22257 ( .A1(n20308), .A2(n20158), .B1(n20162), .B2(n20307), .ZN(
        n20153) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20310), .B1(
        n20164), .B2(n20309), .ZN(n20152) );
  OAI211_X1 U22259 ( .C1(n20161), .C2(n20313), .A(n20153), .B(n20152), .ZN(
        P2_U3082) );
  AOI22_X1 U22260 ( .A1(n20315), .A2(n20158), .B1(n20314), .B2(n20162), .ZN(
        n20155) );
  AOI22_X1 U22261 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20317), .B1(
        n20164), .B2(n20316), .ZN(n20154) );
  OAI211_X1 U22262 ( .C1(n20161), .C2(n20326), .A(n20155), .B(n20154), .ZN(
        P2_U3074) );
  AOI22_X1 U22263 ( .A1(n20321), .A2(n20164), .B1(n20162), .B2(n20320), .ZN(
        n20157) );
  AOI22_X1 U22264 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20323), .B1(
        n20330), .B2(n20163), .ZN(n20156) );
  OAI211_X1 U22265 ( .C1(n20167), .C2(n20326), .A(n20157), .B(n20156), .ZN(
        P2_U3066) );
  AOI22_X1 U22266 ( .A1(n20329), .A2(n20164), .B1(n20162), .B2(n20328), .ZN(
        n20160) );
  AOI22_X1 U22267 ( .A1(n20331), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n20330), .B2(n20158), .ZN(n20159) );
  OAI211_X1 U22268 ( .C1(n20161), .C2(n20334), .A(n20160), .B(n20159), .ZN(
        P2_U3058) );
  AOI22_X1 U22269 ( .A1(n20163), .A2(n20215), .B1(n20162), .B2(n20335), .ZN(
        n20166) );
  AOI22_X1 U22270 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n20164), .ZN(n20165) );
  OAI211_X1 U22271 ( .C1(n20167), .C2(n20334), .A(n20166), .B(n20165), .ZN(
        P2_U3050) );
  AOI22_X1 U22272 ( .A1(n20169), .A2(n20168), .B1(n20221), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n20175) );
  AOI21_X1 U22273 ( .B1(n20172), .B2(n20171), .A(n20170), .ZN(n20173) );
  OR2_X1 U22274 ( .A1(n20173), .A2(n20228), .ZN(n20174) );
  OAI211_X1 U22275 ( .C1(n20177), .C2(n20176), .A(n20175), .B(n20174), .ZN(
        P2_U2918) );
  AOI22_X1 U22276 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n20241), .B1(
        BUF1_REG_17__SCAN_IN), .B2(n20240), .ZN(n20220) );
  NOR2_X2 U22277 ( .A1(n20177), .A2(n20234), .ZN(n20217) );
  NOR2_X2 U22278 ( .A1(n13109), .A2(n20236), .ZN(n20214) );
  AOI22_X1 U22279 ( .A1(n20239), .A2(n20217), .B1(n20238), .B2(n20214), .ZN(
        n20180) );
  AOI22_X1 U22280 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20240), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20241), .ZN(n20213) );
  INV_X1 U22281 ( .A(n20213), .ZN(n20216) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20242), .B1(
        n20246), .B2(n20216), .ZN(n20179) );
  OAI211_X1 U22283 ( .C1(n20220), .C2(n20344), .A(n20180), .B(n20179), .ZN(
        P2_U3169) );
  INV_X1 U22284 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n20183) );
  AOI22_X1 U22285 ( .A1(n20216), .A2(n20254), .B1(n20214), .B2(n20245), .ZN(
        n20182) );
  INV_X1 U22286 ( .A(n20220), .ZN(n20210) );
  AOI22_X1 U22287 ( .A1(n20217), .A2(n20247), .B1(n20246), .B2(n20210), .ZN(
        n20181) );
  OAI211_X1 U22288 ( .C1(n20183), .C2(n20250), .A(n20182), .B(n20181), .ZN(
        P2_U3161) );
  AOI22_X1 U22289 ( .A1(n20253), .A2(n20217), .B1(n20214), .B2(n20252), .ZN(
        n20185) );
  AOI22_X1 U22290 ( .A1(n20210), .A2(n20254), .B1(n20255), .B2(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n20184) );
  OAI211_X1 U22291 ( .C1(n20213), .C2(n20258), .A(n20185), .B(n20184), .ZN(
        P2_U3153) );
  AOI22_X1 U22292 ( .A1(n20260), .A2(n20217), .B1(n20214), .B2(n20259), .ZN(
        n20187) );
  AOI22_X1 U22293 ( .A1(n20262), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n20261), .B2(n20210), .ZN(n20186) );
  OAI211_X1 U22294 ( .C1(n20213), .C2(n20270), .A(n20187), .B(n20186), .ZN(
        P2_U3145) );
  AOI22_X1 U22295 ( .A1(n20266), .A2(n20217), .B1(n20214), .B2(n20265), .ZN(
        n20189) );
  AOI22_X1 U22296 ( .A1(n20216), .A2(n20272), .B1(n20267), .B2(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n20188) );
  OAI211_X1 U22297 ( .C1(n20220), .C2(n20270), .A(n20189), .B(n20188), .ZN(
        P2_U3137) );
  AOI22_X1 U22298 ( .A1(n20190), .A2(n20216), .B1(n20214), .B2(n20271), .ZN(
        n20192) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20274), .B1(
        n20217), .B2(n20273), .ZN(n20191) );
  OAI211_X1 U22300 ( .C1(n20220), .C2(n20193), .A(n20192), .B(n20191), .ZN(
        P2_U3129) );
  AOI22_X1 U22301 ( .A1(n20216), .A2(n20284), .B1(n20214), .B2(n20277), .ZN(
        n20195) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20279), .B1(
        n20217), .B2(n20278), .ZN(n20194) );
  OAI211_X1 U22303 ( .C1(n20220), .C2(n20282), .A(n20195), .B(n20194), .ZN(
        P2_U3121) );
  AOI22_X1 U22304 ( .A1(n20210), .A2(n20284), .B1(n20214), .B2(n20283), .ZN(
        n20197) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20286), .B1(
        n20217), .B2(n20285), .ZN(n20196) );
  OAI211_X1 U22306 ( .C1(n20213), .C2(n20294), .A(n20197), .B(n20196), .ZN(
        P2_U3113) );
  AOI22_X1 U22307 ( .A1(n20290), .A2(n20217), .B1(n20289), .B2(n20214), .ZN(
        n20199) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20291), .B1(
        n20297), .B2(n20216), .ZN(n20198) );
  OAI211_X1 U22309 ( .C1(n20220), .C2(n20294), .A(n20199), .B(n20198), .ZN(
        P2_U3105) );
  AOI22_X1 U22310 ( .A1(n20296), .A2(n20217), .B1(n20214), .B2(n20295), .ZN(
        n20201) );
  AOI22_X1 U22311 ( .A1(n20298), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n20297), .B2(n20210), .ZN(n20200) );
  OAI211_X1 U22312 ( .C1(n20213), .C2(n20306), .A(n20201), .B(n20200), .ZN(
        P2_U3097) );
  AOI22_X1 U22313 ( .A1(n20308), .A2(n20216), .B1(n20214), .B2(n20301), .ZN(
        n20203) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20303), .B1(
        n20217), .B2(n20302), .ZN(n20202) );
  OAI211_X1 U22315 ( .C1(n20220), .C2(n20306), .A(n20203), .B(n20202), .ZN(
        P2_U3089) );
  AOI22_X1 U22316 ( .A1(n20308), .A2(n20210), .B1(n20214), .B2(n20307), .ZN(
        n20205) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20310), .B1(
        n20217), .B2(n20309), .ZN(n20204) );
  OAI211_X1 U22318 ( .C1(n20213), .C2(n20313), .A(n20205), .B(n20204), .ZN(
        P2_U3081) );
  AOI22_X1 U22319 ( .A1(n20315), .A2(n20210), .B1(n20314), .B2(n20214), .ZN(
        n20207) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20317), .B1(
        n20217), .B2(n20316), .ZN(n20206) );
  OAI211_X1 U22321 ( .C1(n20213), .C2(n20326), .A(n20207), .B(n20206), .ZN(
        P2_U3073) );
  AOI22_X1 U22322 ( .A1(n20321), .A2(n20217), .B1(n20214), .B2(n20320), .ZN(
        n20209) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20323), .B1(
        n20330), .B2(n20216), .ZN(n20208) );
  OAI211_X1 U22324 ( .C1(n20220), .C2(n20326), .A(n20209), .B(n20208), .ZN(
        P2_U3065) );
  AOI22_X1 U22325 ( .A1(n20329), .A2(n20217), .B1(n20214), .B2(n20328), .ZN(
        n20212) );
  AOI22_X1 U22326 ( .A1(n20331), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n20330), .B2(n20210), .ZN(n20211) );
  OAI211_X1 U22327 ( .C1(n20213), .C2(n20334), .A(n20212), .B(n20211), .ZN(
        P2_U3057) );
  AOI22_X1 U22328 ( .A1(n20216), .A2(n20215), .B1(n20214), .B2(n20335), .ZN(
        n20219) );
  AOI22_X1 U22329 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n20217), .ZN(n20218) );
  OAI211_X1 U22330 ( .C1(n20220), .C2(n20334), .A(n20219), .B(n20218), .ZN(
        P2_U3049) );
  INV_X1 U22331 ( .A(n20235), .ZN(n20222) );
  AOI22_X1 U22332 ( .A1(n20223), .A2(n20222), .B1(n20221), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n20233) );
  AOI22_X1 U22333 ( .A1(n20225), .A2(BUF2_REG_16__SCAN_IN), .B1(n20224), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n20232) );
  OAI22_X1 U22334 ( .A1(n20229), .A2(n20228), .B1(n20227), .B2(n20226), .ZN(
        n20230) );
  INV_X1 U22335 ( .A(n20230), .ZN(n20231) );
  NAND3_X1 U22336 ( .A1(n20233), .A2(n20232), .A3(n20231), .ZN(P2_U2903) );
  AOI22_X1 U22337 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n20241), .B1(
        BUF1_REG_16__SCAN_IN), .B2(n20240), .ZN(n20327) );
  NOR2_X2 U22338 ( .A1(n20235), .A2(n20234), .ZN(n20339) );
  NOR2_X2 U22339 ( .A1(n20237), .A2(n20236), .ZN(n20336) );
  AOI22_X1 U22340 ( .A1(n20239), .A2(n20339), .B1(n20238), .B2(n20336), .ZN(
        n20244) );
  AOI22_X1 U22341 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n20241), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n20240), .ZN(n20345) );
  INV_X1 U22342 ( .A(n20345), .ZN(n20322) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20242), .B1(
        n20246), .B2(n20322), .ZN(n20243) );
  OAI211_X1 U22344 ( .C1(n20327), .C2(n20344), .A(n20244), .B(n20243), .ZN(
        P2_U3168) );
  INV_X1 U22345 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n20251) );
  AOI22_X1 U22346 ( .A1(n20322), .A2(n20254), .B1(n20336), .B2(n20245), .ZN(
        n20249) );
  AOI22_X1 U22347 ( .A1(n20339), .A2(n20247), .B1(n20246), .B2(n20337), .ZN(
        n20248) );
  OAI211_X1 U22348 ( .C1(n20251), .C2(n20250), .A(n20249), .B(n20248), .ZN(
        P2_U3160) );
  AOI22_X1 U22349 ( .A1(n20253), .A2(n20339), .B1(n20336), .B2(n20252), .ZN(
        n20257) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20255), .B1(
        n20337), .B2(n20254), .ZN(n20256) );
  OAI211_X1 U22351 ( .C1(n20345), .C2(n20258), .A(n20257), .B(n20256), .ZN(
        P2_U3152) );
  AOI22_X1 U22352 ( .A1(n20260), .A2(n20339), .B1(n20336), .B2(n20259), .ZN(
        n20264) );
  AOI22_X1 U22353 ( .A1(n20262), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n20261), .B2(n20337), .ZN(n20263) );
  OAI211_X1 U22354 ( .C1(n20345), .C2(n20270), .A(n20264), .B(n20263), .ZN(
        P2_U3144) );
  AOI22_X1 U22355 ( .A1(n20266), .A2(n20339), .B1(n20336), .B2(n20265), .ZN(
        n20269) );
  AOI22_X1 U22356 ( .A1(n20322), .A2(n20272), .B1(
        P2_INSTQUEUE_REG_11__0__SCAN_IN), .B2(n20267), .ZN(n20268) );
  OAI211_X1 U22357 ( .C1(n20327), .C2(n20270), .A(n20269), .B(n20268), .ZN(
        P2_U3136) );
  AOI22_X1 U22358 ( .A1(n20337), .A2(n20272), .B1(n20336), .B2(n20271), .ZN(
        n20276) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20274), .B1(
        n20339), .B2(n20273), .ZN(n20275) );
  OAI211_X1 U22360 ( .C1(n20345), .C2(n20282), .A(n20276), .B(n20275), .ZN(
        P2_U3128) );
  AOI22_X1 U22361 ( .A1(n20322), .A2(n20284), .B1(n20336), .B2(n20277), .ZN(
        n20281) );
  AOI22_X1 U22362 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20279), .B1(
        n20339), .B2(n20278), .ZN(n20280) );
  OAI211_X1 U22363 ( .C1(n20327), .C2(n20282), .A(n20281), .B(n20280), .ZN(
        P2_U3120) );
  AOI22_X1 U22364 ( .A1(n20337), .A2(n20284), .B1(n20336), .B2(n20283), .ZN(
        n20288) );
  AOI22_X1 U22365 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20286), .B1(
        n20339), .B2(n20285), .ZN(n20287) );
  OAI211_X1 U22366 ( .C1(n20345), .C2(n20294), .A(n20288), .B(n20287), .ZN(
        P2_U3112) );
  AOI22_X1 U22367 ( .A1(n20290), .A2(n20339), .B1(n20289), .B2(n20336), .ZN(
        n20293) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20291), .B1(
        n20297), .B2(n20322), .ZN(n20292) );
  OAI211_X1 U22369 ( .C1(n20327), .C2(n20294), .A(n20293), .B(n20292), .ZN(
        P2_U3104) );
  AOI22_X1 U22370 ( .A1(n20296), .A2(n20339), .B1(n20336), .B2(n20295), .ZN(
        n20300) );
  AOI22_X1 U22371 ( .A1(n20298), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n20297), .B2(n20337), .ZN(n20299) );
  OAI211_X1 U22372 ( .C1(n20345), .C2(n20306), .A(n20300), .B(n20299), .ZN(
        P2_U3096) );
  AOI22_X1 U22373 ( .A1(n20308), .A2(n20322), .B1(n20336), .B2(n20301), .ZN(
        n20305) );
  AOI22_X1 U22374 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20303), .B1(
        n20339), .B2(n20302), .ZN(n20304) );
  OAI211_X1 U22375 ( .C1(n20327), .C2(n20306), .A(n20305), .B(n20304), .ZN(
        P2_U3088) );
  AOI22_X1 U22376 ( .A1(n20308), .A2(n20337), .B1(n20336), .B2(n20307), .ZN(
        n20312) );
  AOI22_X1 U22377 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20310), .B1(
        n20339), .B2(n20309), .ZN(n20311) );
  OAI211_X1 U22378 ( .C1(n20345), .C2(n20313), .A(n20312), .B(n20311), .ZN(
        P2_U3080) );
  AOI22_X1 U22379 ( .A1(n20315), .A2(n20337), .B1(n20314), .B2(n20336), .ZN(
        n20319) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20317), .B1(
        n20339), .B2(n20316), .ZN(n20318) );
  OAI211_X1 U22381 ( .C1(n20345), .C2(n20326), .A(n20319), .B(n20318), .ZN(
        P2_U3072) );
  AOI22_X1 U22382 ( .A1(n20321), .A2(n20339), .B1(n20336), .B2(n20320), .ZN(
        n20325) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20323), .B1(
        n20330), .B2(n20322), .ZN(n20324) );
  OAI211_X1 U22384 ( .C1(n20327), .C2(n20326), .A(n20325), .B(n20324), .ZN(
        P2_U3064) );
  AOI22_X1 U22385 ( .A1(n20329), .A2(n20339), .B1(n20336), .B2(n20328), .ZN(
        n20333) );
  AOI22_X1 U22386 ( .A1(n20331), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n20330), .B2(n20337), .ZN(n20332) );
  OAI211_X1 U22387 ( .C1(n20345), .C2(n20334), .A(n20333), .B(n20332), .ZN(
        P2_U3056) );
  AOI22_X1 U22388 ( .A1(n20338), .A2(n20337), .B1(n20336), .B2(n20335), .ZN(
        n20343) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n20339), .ZN(n20342) );
  OAI211_X1 U22390 ( .C1(n20345), .C2(n20344), .A(n20343), .B(n20342), .ZN(
        P2_U3048) );
  INV_X1 U22391 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20624) );
  INV_X1 U22392 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20346) );
  AOI222_X1 U22393 ( .A1(n20624), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20627), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n20346), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20347) );
  INV_X1 U22394 ( .A(n20372), .ZN(n20371) );
  OAI22_X1 U22395 ( .A1(n20372), .A2(P3_ADDRESS_REG_0__SCAN_IN), .B1(
        P2_ADDRESS_REG_0__SCAN_IN), .B2(n20371), .ZN(n20348) );
  INV_X1 U22396 ( .A(n20348), .ZN(U376) );
  OAI22_X1 U22397 ( .A1(n20372), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n20371), .ZN(n20349) );
  INV_X1 U22398 ( .A(n20349), .ZN(U365) );
  OAI22_X1 U22399 ( .A1(n20372), .A2(P3_ADDRESS_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n20371), .ZN(n20350) );
  INV_X1 U22400 ( .A(n20350), .ZN(U354) );
  OAI22_X1 U22401 ( .A1(n20372), .A2(P3_ADDRESS_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n20371), .ZN(n20351) );
  INV_X1 U22402 ( .A(n20351), .ZN(U353) );
  OAI22_X1 U22403 ( .A1(n20372), .A2(P3_ADDRESS_REG_4__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n20371), .ZN(n20352) );
  INV_X1 U22404 ( .A(n20352), .ZN(U352) );
  OAI22_X1 U22405 ( .A1(n20372), .A2(P3_ADDRESS_REG_5__SCAN_IN), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(n20371), .ZN(n20353) );
  INV_X1 U22406 ( .A(n20353), .ZN(U351) );
  OAI22_X1 U22407 ( .A1(n20372), .A2(P3_ADDRESS_REG_6__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n20371), .ZN(n20354) );
  INV_X1 U22408 ( .A(n20354), .ZN(U350) );
  OAI22_X1 U22409 ( .A1(n20372), .A2(P3_ADDRESS_REG_7__SCAN_IN), .B1(
        P2_ADDRESS_REG_7__SCAN_IN), .B2(n20371), .ZN(n20355) );
  INV_X1 U22410 ( .A(n20355), .ZN(U349) );
  OAI22_X1 U22411 ( .A1(n20372), .A2(P3_ADDRESS_REG_8__SCAN_IN), .B1(
        P2_ADDRESS_REG_8__SCAN_IN), .B2(n20371), .ZN(n20356) );
  INV_X1 U22412 ( .A(n20356), .ZN(U348) );
  OAI22_X1 U22413 ( .A1(n20372), .A2(P3_ADDRESS_REG_9__SCAN_IN), .B1(
        P2_ADDRESS_REG_9__SCAN_IN), .B2(n20371), .ZN(n20357) );
  INV_X1 U22414 ( .A(n20357), .ZN(U347) );
  OAI22_X1 U22415 ( .A1(n20372), .A2(P3_ADDRESS_REG_10__SCAN_IN), .B1(
        P2_ADDRESS_REG_10__SCAN_IN), .B2(n20371), .ZN(n20358) );
  INV_X1 U22416 ( .A(n20358), .ZN(U375) );
  OAI22_X1 U22417 ( .A1(n20372), .A2(P3_ADDRESS_REG_11__SCAN_IN), .B1(
        P2_ADDRESS_REG_11__SCAN_IN), .B2(n20371), .ZN(n20359) );
  INV_X1 U22418 ( .A(n20359), .ZN(U374) );
  INV_X1 U22419 ( .A(n20372), .ZN(n20379) );
  OAI22_X1 U22420 ( .A1(n20372), .A2(P3_ADDRESS_REG_12__SCAN_IN), .B1(
        P2_ADDRESS_REG_12__SCAN_IN), .B2(n20379), .ZN(n20360) );
  INV_X1 U22421 ( .A(n20360), .ZN(U373) );
  OAI22_X1 U22422 ( .A1(n20372), .A2(P3_ADDRESS_REG_13__SCAN_IN), .B1(
        P2_ADDRESS_REG_13__SCAN_IN), .B2(n20371), .ZN(n20361) );
  INV_X1 U22423 ( .A(n20361), .ZN(U372) );
  OAI22_X1 U22424 ( .A1(n20372), .A2(P3_ADDRESS_REG_14__SCAN_IN), .B1(
        P2_ADDRESS_REG_14__SCAN_IN), .B2(n20371), .ZN(n20362) );
  INV_X1 U22425 ( .A(n20362), .ZN(U371) );
  OAI22_X1 U22426 ( .A1(n20372), .A2(P3_ADDRESS_REG_15__SCAN_IN), .B1(
        P2_ADDRESS_REG_15__SCAN_IN), .B2(n20371), .ZN(n20363) );
  INV_X1 U22427 ( .A(n20363), .ZN(U370) );
  OAI22_X1 U22428 ( .A1(n20372), .A2(P3_ADDRESS_REG_16__SCAN_IN), .B1(
        P2_ADDRESS_REG_16__SCAN_IN), .B2(n20379), .ZN(n20364) );
  INV_X1 U22429 ( .A(n20364), .ZN(U369) );
  OAI22_X1 U22430 ( .A1(n20372), .A2(P3_ADDRESS_REG_17__SCAN_IN), .B1(
        P2_ADDRESS_REG_17__SCAN_IN), .B2(n20371), .ZN(n20365) );
  INV_X1 U22431 ( .A(n20365), .ZN(U368) );
  OAI22_X1 U22432 ( .A1(n20372), .A2(P3_ADDRESS_REG_18__SCAN_IN), .B1(
        P2_ADDRESS_REG_18__SCAN_IN), .B2(n20371), .ZN(n20366) );
  INV_X1 U22433 ( .A(n20366), .ZN(U367) );
  OAI22_X1 U22434 ( .A1(n20372), .A2(P3_ADDRESS_REG_19__SCAN_IN), .B1(
        P2_ADDRESS_REG_19__SCAN_IN), .B2(n20371), .ZN(n20367) );
  INV_X1 U22435 ( .A(n20367), .ZN(U366) );
  OAI22_X1 U22436 ( .A1(n20372), .A2(P3_ADDRESS_REG_20__SCAN_IN), .B1(
        P2_ADDRESS_REG_20__SCAN_IN), .B2(n20371), .ZN(n20368) );
  INV_X1 U22437 ( .A(n20368), .ZN(U364) );
  OAI22_X1 U22438 ( .A1(n20372), .A2(P3_ADDRESS_REG_21__SCAN_IN), .B1(
        P2_ADDRESS_REG_21__SCAN_IN), .B2(n20371), .ZN(n20369) );
  INV_X1 U22439 ( .A(n20369), .ZN(U363) );
  OAI22_X1 U22440 ( .A1(n20372), .A2(P3_ADDRESS_REG_22__SCAN_IN), .B1(
        P2_ADDRESS_REG_22__SCAN_IN), .B2(n20371), .ZN(n20370) );
  INV_X1 U22441 ( .A(n20370), .ZN(U362) );
  OAI22_X1 U22442 ( .A1(n20372), .A2(P3_ADDRESS_REG_23__SCAN_IN), .B1(
        P2_ADDRESS_REG_23__SCAN_IN), .B2(n20371), .ZN(n20373) );
  INV_X1 U22443 ( .A(n20373), .ZN(U361) );
  OAI22_X1 U22444 ( .A1(n20372), .A2(P3_ADDRESS_REG_24__SCAN_IN), .B1(
        P2_ADDRESS_REG_24__SCAN_IN), .B2(n20379), .ZN(n20374) );
  INV_X1 U22445 ( .A(n20374), .ZN(U360) );
  OAI22_X1 U22446 ( .A1(n20372), .A2(P3_ADDRESS_REG_25__SCAN_IN), .B1(
        P2_ADDRESS_REG_25__SCAN_IN), .B2(n20379), .ZN(n20375) );
  INV_X1 U22447 ( .A(n20375), .ZN(U359) );
  OAI22_X1 U22448 ( .A1(n20372), .A2(P3_ADDRESS_REG_26__SCAN_IN), .B1(
        P2_ADDRESS_REG_26__SCAN_IN), .B2(n20379), .ZN(n20376) );
  INV_X1 U22449 ( .A(n20376), .ZN(U358) );
  OAI22_X1 U22450 ( .A1(n20372), .A2(P3_ADDRESS_REG_27__SCAN_IN), .B1(
        P2_ADDRESS_REG_27__SCAN_IN), .B2(n20379), .ZN(n20377) );
  INV_X1 U22451 ( .A(n20377), .ZN(U357) );
  OAI22_X1 U22452 ( .A1(n20372), .A2(P3_ADDRESS_REG_28__SCAN_IN), .B1(
        P2_ADDRESS_REG_28__SCAN_IN), .B2(n20379), .ZN(n20378) );
  INV_X1 U22453 ( .A(n20378), .ZN(U356) );
  OAI22_X1 U22454 ( .A1(n20372), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n20379), .ZN(n20380) );
  INV_X1 U22455 ( .A(n20380), .ZN(U355) );
  AOI22_X1 U22456 ( .A1(n21862), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20393), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20382) );
  OAI21_X1 U22457 ( .B1(n22314), .B2(n20401), .A(n20382), .ZN(P1_U2936) );
  INV_X1 U22458 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n22321) );
  AOI22_X1 U22459 ( .A1(n20390), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20383) );
  OAI21_X1 U22460 ( .B1(n22321), .B2(n20401), .A(n20383), .ZN(P1_U2935) );
  INV_X1 U22461 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n22327) );
  AOI22_X1 U22462 ( .A1(n20390), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20393), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20384) );
  OAI21_X1 U22463 ( .B1(n22327), .B2(n20401), .A(n20384), .ZN(P1_U2934) );
  AOI22_X1 U22464 ( .A1(n20390), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20385) );
  OAI21_X1 U22465 ( .B1(n22333), .B2(n20401), .A(n20385), .ZN(P1_U2933) );
  AOI22_X1 U22466 ( .A1(n20390), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20393), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20386) );
  OAI21_X1 U22467 ( .B1(n22340), .B2(n20401), .A(n20386), .ZN(P1_U2932) );
  AOI22_X1 U22468 ( .A1(n20390), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20387) );
  OAI21_X1 U22469 ( .B1(n12160), .B2(n20401), .A(n20387), .ZN(P1_U2931) );
  AOI22_X1 U22470 ( .A1(n20390), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20393), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20388) );
  OAI21_X1 U22471 ( .B1(n22351), .B2(n20401), .A(n20388), .ZN(P1_U2930) );
  AOI22_X1 U22472 ( .A1(n21862), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20393), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20389) );
  OAI21_X1 U22473 ( .B1(n12149), .B2(n20401), .A(n20389), .ZN(P1_U2929) );
  INV_X1 U22474 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n22361) );
  AOI22_X1 U22475 ( .A1(n20390), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20393), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20391) );
  OAI21_X1 U22476 ( .B1(n22361), .B2(n20401), .A(n20391), .ZN(P1_U2928) );
  INV_X1 U22477 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n22367) );
  AOI22_X1 U22478 ( .A1(n21862), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20393), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20392) );
  OAI21_X1 U22479 ( .B1(n22367), .B2(n20401), .A(n20392), .ZN(P1_U2927) );
  INV_X1 U22480 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n22374) );
  AOI22_X1 U22481 ( .A1(n21862), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20393), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20394) );
  OAI21_X1 U22482 ( .B1(n22374), .B2(n20401), .A(n20394), .ZN(P1_U2926) );
  INV_X1 U22483 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n22381) );
  AOI22_X1 U22484 ( .A1(n21862), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20395) );
  OAI21_X1 U22485 ( .B1(n22381), .B2(n20401), .A(n20395), .ZN(P1_U2925) );
  INV_X1 U22486 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n22389) );
  AOI22_X1 U22487 ( .A1(n21862), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20396) );
  OAI21_X1 U22488 ( .B1(n22389), .B2(n20401), .A(n20396), .ZN(P1_U2924) );
  INV_X1 U22489 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n22396) );
  AOI22_X1 U22490 ( .A1(n21862), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20397) );
  OAI21_X1 U22491 ( .B1(n22396), .B2(n20401), .A(n20397), .ZN(P1_U2923) );
  INV_X1 U22492 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n22406) );
  AOI22_X1 U22493 ( .A1(n21862), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20398) );
  OAI21_X1 U22494 ( .B1(n22406), .B2(n20401), .A(n20398), .ZN(P1_U2922) );
  AOI22_X1 U22495 ( .A1(n21862), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20399), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20400) );
  OAI21_X1 U22496 ( .B1(n20402), .B2(n20401), .A(n20400), .ZN(P1_U2921) );
  OR2_X1 U22497 ( .A1(n20562), .A2(n22806), .ZN(n20426) );
  OR2_X1 U22498 ( .A1(n22806), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20428) );
  OAI222_X1 U22499 ( .A1(n20426), .A2(n22031), .B1(n20403), .B2(n22805), .C1(
        n22032), .C2(n20428), .ZN(P1_U3197) );
  AOI222_X1 U22500 ( .A1(n11169), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n22806), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n11168), .ZN(n20404) );
  INV_X1 U22501 ( .A(n20404), .ZN(P1_U3198) );
  INV_X1 U22502 ( .A(n22805), .ZN(n20434) );
  AOI222_X1 U22503 ( .A1(n11169), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n11168), .ZN(n20405) );
  INV_X1 U22504 ( .A(n20405), .ZN(P1_U3199) );
  AOI222_X1 U22505 ( .A1(n11168), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n11169), .ZN(n20406) );
  INV_X1 U22506 ( .A(n20406), .ZN(P1_U3200) );
  AOI222_X1 U22507 ( .A1(n11169), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n11168), .ZN(n20407) );
  INV_X1 U22508 ( .A(n20407), .ZN(P1_U3201) );
  AOI222_X1 U22509 ( .A1(n11169), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n11168), .ZN(n20408) );
  INV_X1 U22510 ( .A(n20408), .ZN(P1_U3202) );
  AOI222_X1 U22511 ( .A1(n11169), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n11168), .ZN(n20409) );
  INV_X1 U22512 ( .A(n20409), .ZN(P1_U3203) );
  AOI222_X1 U22513 ( .A1(n11168), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n11169), .ZN(n20410) );
  INV_X1 U22514 ( .A(n20410), .ZN(P1_U3204) );
  AOI222_X1 U22515 ( .A1(n11168), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n11169), .ZN(n20411) );
  INV_X1 U22516 ( .A(n20411), .ZN(P1_U3205) );
  AOI222_X1 U22517 ( .A1(n11169), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n11168), .ZN(n20412) );
  INV_X1 U22518 ( .A(n20412), .ZN(P1_U3206) );
  AOI222_X1 U22519 ( .A1(n11168), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n11169), .ZN(n20413) );
  INV_X1 U22520 ( .A(n20413), .ZN(P1_U3207) );
  AOI222_X1 U22521 ( .A1(n11169), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n11168), .ZN(n20414) );
  INV_X1 U22522 ( .A(n20414), .ZN(P1_U3208) );
  AOI222_X1 U22523 ( .A1(n11169), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n11168), .ZN(n20415) );
  INV_X1 U22524 ( .A(n20415), .ZN(P1_U3209) );
  AOI222_X1 U22525 ( .A1(n11169), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n11168), .ZN(n20416) );
  INV_X1 U22526 ( .A(n20416), .ZN(P1_U3210) );
  AOI222_X1 U22527 ( .A1(n11169), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n11168), .ZN(n20417) );
  INV_X1 U22528 ( .A(n20417), .ZN(P1_U3211) );
  AOI222_X1 U22529 ( .A1(n11169), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n11168), .ZN(n20418) );
  INV_X1 U22530 ( .A(n20418), .ZN(P1_U3212) );
  AOI222_X1 U22531 ( .A1(n11169), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n11168), .ZN(n20419) );
  INV_X1 U22532 ( .A(n20419), .ZN(P1_U3213) );
  AOI222_X1 U22533 ( .A1(n11169), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n11168), .ZN(n20420) );
  INV_X1 U22534 ( .A(n20420), .ZN(P1_U3214) );
  AOI222_X1 U22535 ( .A1(n11169), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n11168), .ZN(n20421) );
  INV_X1 U22536 ( .A(n20421), .ZN(P1_U3215) );
  AOI222_X1 U22537 ( .A1(n11168), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n11169), .ZN(n20422) );
  INV_X1 U22538 ( .A(n20422), .ZN(P1_U3216) );
  AOI222_X1 U22539 ( .A1(n11169), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n11168), .ZN(n20423) );
  INV_X1 U22540 ( .A(n20423), .ZN(P1_U3217) );
  AOI222_X1 U22541 ( .A1(n11169), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n11168), .ZN(n20424) );
  INV_X1 U22542 ( .A(n20424), .ZN(P1_U3218) );
  AOI22_X1 U22543 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n11168), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n22806), .ZN(n20425) );
  OAI21_X1 U22544 ( .B1(n22191), .B2(n20426), .A(n20425), .ZN(P1_U3219) );
  AOI22_X1 U22545 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n11169), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n22806), .ZN(n20427) );
  OAI21_X1 U22546 ( .B1(n20429), .B2(n20428), .A(n20427), .ZN(P1_U3220) );
  AOI222_X1 U22547 ( .A1(n11169), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n11168), .ZN(n20430) );
  INV_X1 U22548 ( .A(n20430), .ZN(P1_U3221) );
  AOI222_X1 U22549 ( .A1(n11169), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n11168), .ZN(n20431) );
  INV_X1 U22550 ( .A(n20431), .ZN(P1_U3222) );
  AOI222_X1 U22551 ( .A1(n11169), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n11168), .ZN(n20432) );
  INV_X1 U22552 ( .A(n20432), .ZN(P1_U3223) );
  AOI222_X1 U22553 ( .A1(n11169), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n11168), .ZN(n20433) );
  INV_X1 U22554 ( .A(n20433), .ZN(P1_U3224) );
  AOI222_X1 U22555 ( .A1(n11169), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20434), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n11168), .ZN(n20435) );
  INV_X1 U22556 ( .A(n20435), .ZN(P1_U3225) );
  AOI222_X1 U22557 ( .A1(n11169), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n22806), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n11168), .ZN(n20436) );
  INV_X1 U22558 ( .A(n20436), .ZN(P1_U3226) );
  OAI22_X1 U22559 ( .A1(n22806), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22805), .ZN(n20437) );
  INV_X1 U22560 ( .A(n20437), .ZN(P1_U3458) );
  AOI221_X1 U22561 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20448) );
  NOR4_X1 U22562 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20441) );
  NOR4_X1 U22563 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20440) );
  NOR4_X1 U22564 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20439) );
  NOR4_X1 U22565 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20438) );
  NAND4_X1 U22566 ( .A1(n20441), .A2(n20440), .A3(n20439), .A4(n20438), .ZN(
        n20447) );
  NOR4_X1 U22567 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20445) );
  AOI211_X1 U22568 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20444) );
  NOR4_X1 U22569 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20443) );
  NOR4_X1 U22570 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20442) );
  NAND4_X1 U22571 ( .A1(n20445), .A2(n20444), .A3(n20443), .A4(n20442), .ZN(
        n20446) );
  NOR2_X1 U22572 ( .A1(n20447), .A2(n20446), .ZN(n20460) );
  MUX2_X1 U22573 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n20448), .S(n20460), 
        .Z(P1_U2808) );
  OAI22_X1 U22574 ( .A1(n22806), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22805), .ZN(n20449) );
  INV_X1 U22575 ( .A(n20449), .ZN(P1_U3459) );
  AOI21_X1 U22576 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20450) );
  OAI221_X1 U22577 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20450), .C1(n22031), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20460), .ZN(n20451) );
  OAI21_X1 U22578 ( .B1(n20460), .B2(n20452), .A(n20451), .ZN(P1_U3481) );
  OAI22_X1 U22579 ( .A1(n22806), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22805), .ZN(n20453) );
  INV_X1 U22580 ( .A(n20453), .ZN(P1_U3460) );
  INV_X1 U22581 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20456) );
  NOR3_X1 U22582 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20454) );
  OAI21_X1 U22583 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20454), .A(n20460), .ZN(
        n20455) );
  OAI21_X1 U22584 ( .B1(n20460), .B2(n20456), .A(n20455), .ZN(P1_U2807) );
  OAI22_X1 U22585 ( .A1(n22806), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22805), .ZN(n20457) );
  INV_X1 U22586 ( .A(n20457), .ZN(P1_U3461) );
  OAI21_X1 U22587 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20460), .ZN(n20458) );
  OAI21_X1 U22588 ( .B1(n20460), .B2(n20459), .A(n20458), .ZN(P1_U3482) );
  AOI22_X1 U22589 ( .A1(n20462), .A2(n20489), .B1(n20488), .B2(n20461), .ZN(
        n20463) );
  OAI21_X1 U22590 ( .B1(n20493), .B2(n11742), .A(n20463), .ZN(P1_U2871) );
  AOI22_X1 U22591 ( .A1(n22026), .A2(n20489), .B1(n20488), .B2(n22019), .ZN(
        n20464) );
  OAI21_X1 U22592 ( .B1(n20493), .B2(n20465), .A(n20464), .ZN(P1_U2870) );
  OAI21_X1 U22593 ( .B1(n20467), .B2(n20466), .A(n16580), .ZN(n20468) );
  INV_X1 U22594 ( .A(n20468), .ZN(n22145) );
  AOI22_X1 U22595 ( .A1(n22146), .A2(n20489), .B1(n22145), .B2(n20488), .ZN(
        n20469) );
  OAI21_X1 U22596 ( .B1(n20493), .B2(n22142), .A(n20469), .ZN(P1_U2856) );
  AOI22_X1 U22597 ( .A1(n22173), .A2(n20489), .B1(n20488), .B2(n22164), .ZN(
        n20470) );
  OAI21_X1 U22598 ( .B1(n20493), .B2(n20471), .A(n20470), .ZN(P1_U2854) );
  INV_X1 U22599 ( .A(n20472), .ZN(n22127) );
  AOI22_X1 U22600 ( .A1(n22127), .A2(n20489), .B1(n20488), .B2(n22125), .ZN(
        n20473) );
  OAI21_X1 U22601 ( .B1(n20493), .B2(n22122), .A(n20473), .ZN(P1_U2858) );
  AOI22_X1 U22602 ( .A1(n20547), .A2(n20489), .B1(n21937), .B2(n20488), .ZN(
        n20474) );
  OAI21_X1 U22603 ( .B1(n20493), .B2(n20475), .A(n20474), .ZN(P1_U2850) );
  INV_X1 U22604 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n22202) );
  NAND2_X1 U22605 ( .A1(n20477), .A2(n20476), .ZN(n20478) );
  NAND2_X1 U22606 ( .A1(n20479), .A2(n20478), .ZN(n22207) );
  OAI22_X1 U22607 ( .A1(n22210), .A2(n20483), .B1(n22207), .B2(n20480), .ZN(
        n20481) );
  INV_X1 U22608 ( .A(n20481), .ZN(n20482) );
  OAI21_X1 U22609 ( .B1(n20493), .B2(n22202), .A(n20482), .ZN(P1_U2848) );
  OAI22_X1 U22610 ( .A1(n20539), .A2(n20483), .B1(n21924), .B2(n20480), .ZN(
        n20484) );
  INV_X1 U22611 ( .A(n20484), .ZN(n20485) );
  OAI21_X1 U22612 ( .B1(n20493), .B2(n20486), .A(n20485), .ZN(P1_U2852) );
  AOI22_X1 U22613 ( .A1(n20490), .A2(n20489), .B1(n20488), .B2(n20487), .ZN(
        n20491) );
  OAI21_X1 U22614 ( .B1(n20493), .B2(n20492), .A(n20491), .ZN(P1_U2864) );
  INV_X1 U22615 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20499) );
  INV_X1 U22616 ( .A(n22075), .ZN(n20494) );
  AOI222_X1 U22617 ( .A1(n20495), .A2(n20556), .B1(n20494), .B2(n20520), .C1(
        n20557), .C2(n22070), .ZN(n20498) );
  INV_X1 U22618 ( .A(n20496), .ZN(n20497) );
  OAI211_X1 U22619 ( .C1(n20506), .C2(n20499), .A(n20498), .B(n20497), .ZN(
        P1_U2994) );
  INV_X1 U22620 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20505) );
  INV_X1 U22621 ( .A(n22091), .ZN(n20501) );
  AOI222_X1 U22622 ( .A1(n20502), .A2(n20556), .B1(n20501), .B2(n20520), .C1(
        n20557), .C2(n20500), .ZN(n20504) );
  OAI211_X1 U22623 ( .C1(n20506), .C2(n20505), .A(n20504), .B(n20503), .ZN(
        P1_U2992) );
  AOI22_X1 U22624 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20551), .B1(
        n21999), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n20511) );
  INV_X1 U22625 ( .A(n20507), .ZN(n20508) );
  AOI22_X1 U22626 ( .A1(n20509), .A2(n20557), .B1(n20520), .B2(n20508), .ZN(
        n20510) );
  OAI211_X1 U22627 ( .C1(n22216), .C2(n20512), .A(n20511), .B(n20510), .ZN(
        P1_U2989) );
  AOI22_X1 U22628 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20551), .B1(
        n21999), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n20519) );
  OAI21_X1 U22629 ( .B1(n20517), .B2(n20516), .A(n20515), .ZN(n21887) );
  AOI22_X1 U22630 ( .A1(n20556), .A2(n21887), .B1(n20520), .B2(n22117), .ZN(
        n20518) );
  OAI211_X1 U22631 ( .C1(n20538), .C2(n22120), .A(n20519), .B(n20518), .ZN(
        P1_U2987) );
  AOI22_X1 U22632 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20551), .B1(
        n21999), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n20522) );
  AOI22_X1 U22633 ( .A1(n22127), .A2(n20557), .B1(n20520), .B2(n22126), .ZN(
        n20521) );
  OAI211_X1 U22634 ( .C1(n20523), .C2(n22216), .A(n20522), .B(n20521), .ZN(
        P1_U2985) );
  AOI22_X1 U22635 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n20551), .B1(
        n21999), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n20532) );
  NOR2_X1 U22636 ( .A1(n11861), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n20524) );
  OAI22_X1 U22637 ( .A1(n20525), .A2(n20524), .B1(n20552), .B2(n21901), .ZN(
        n20530) );
  INV_X1 U22638 ( .A(n20526), .ZN(n20527) );
  NOR2_X1 U22639 ( .A1(n20528), .A2(n20527), .ZN(n20529) );
  XNOR2_X1 U22640 ( .A(n20530), .B(n20529), .ZN(n21906) );
  AOI22_X1 U22641 ( .A1(n21906), .A2(n20556), .B1(n20557), .B2(n22146), .ZN(
        n20531) );
  OAI211_X1 U22642 ( .C1(n20561), .C2(n22143), .A(n20532), .B(n20531), .ZN(
        P1_U2983) );
  AOI22_X1 U22643 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20551), .B1(
        n21999), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n20542) );
  NAND2_X1 U22644 ( .A1(n20533), .A2(n21932), .ZN(n20536) );
  NAND2_X1 U22645 ( .A1(n20534), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n20535) );
  NAND2_X1 U22646 ( .A1(n20536), .A2(n20535), .ZN(n20537) );
  XNOR2_X1 U22647 ( .A(n20537), .B(n16725), .ZN(n21923) );
  OAI22_X1 U22648 ( .A1(n20539), .A2(n20538), .B1(n22216), .B2(n21923), .ZN(
        n20540) );
  INV_X1 U22649 ( .A(n20540), .ZN(n20541) );
  OAI211_X1 U22650 ( .C1(n20561), .C2(n20543), .A(n20542), .B(n20541), .ZN(
        P1_U2979) );
  AOI22_X1 U22651 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20551), .B1(
        n21999), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n20549) );
  NAND2_X1 U22652 ( .A1(n20545), .A2(n20544), .ZN(n20546) );
  XNOR2_X1 U22653 ( .A(n20546), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n21938) );
  AOI22_X1 U22654 ( .A1(n20547), .A2(n20557), .B1(n20556), .B2(n21938), .ZN(
        n20548) );
  OAI211_X1 U22655 ( .C1(n20561), .C2(n20550), .A(n20549), .B(n20548), .ZN(
        P1_U2977) );
  AOI22_X1 U22656 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20551), .B1(
        n21999), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n20560) );
  INV_X1 U22657 ( .A(n22210), .ZN(n20558) );
  INV_X1 U22658 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n22003) );
  NAND2_X1 U22659 ( .A1(n11861), .A2(n22003), .ZN(n20554) );
  NAND3_X1 U22660 ( .A1(n16680), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n20552), .ZN(n20553) );
  OAI21_X1 U22661 ( .B1(n16680), .B2(n20554), .A(n20553), .ZN(n20555) );
  XNOR2_X1 U22662 ( .A(n20555), .B(n21960), .ZN(n21958) );
  AOI22_X1 U22663 ( .A1(n20558), .A2(n20557), .B1(n20556), .B2(n21958), .ZN(
        n20559) );
  OAI211_X1 U22664 ( .C1(n20561), .C2(n22204), .A(n20560), .B(n20559), .ZN(
        P1_U2975) );
  OAI21_X1 U22665 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20562), .A(n22259), 
        .ZN(n20563) );
  AOI22_X1 U22666 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n22805), .B1(n20564), 
        .B2(n20563), .ZN(P1_U2804) );
  INV_X1 U22667 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20567) );
  AOI22_X1 U22668 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n20608), .ZN(n20566) );
  OAI21_X1 U22669 ( .B1(n20567), .B2(n20626), .A(n20566), .ZN(U247) );
  AOI22_X1 U22670 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n20608), .ZN(n20568) );
  OAI21_X1 U22671 ( .B1(n20569), .B2(n20626), .A(n20568), .ZN(U246) );
  AOI22_X1 U22672 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n20608), .ZN(n20570) );
  OAI21_X1 U22673 ( .B1(n20571), .B2(n20626), .A(n20570), .ZN(U245) );
  INV_X1 U22674 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20573) );
  AOI22_X1 U22675 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n20608), .ZN(n20572) );
  OAI21_X1 U22676 ( .B1(n20573), .B2(n20626), .A(n20572), .ZN(U244) );
  INV_X1 U22677 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20575) );
  AOI22_X1 U22678 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n20608), .ZN(n20574) );
  OAI21_X1 U22679 ( .B1(n20575), .B2(n20626), .A(n20574), .ZN(U243) );
  INV_X1 U22680 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20577) );
  AOI22_X1 U22681 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n20608), .ZN(n20576) );
  OAI21_X1 U22682 ( .B1(n20577), .B2(n20626), .A(n20576), .ZN(U242) );
  AOI22_X1 U22683 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n20608), .ZN(n20578) );
  OAI21_X1 U22684 ( .B1(n20579), .B2(n20626), .A(n20578), .ZN(U241) );
  INV_X1 U22685 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20581) );
  AOI22_X1 U22686 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n20608), .ZN(n20580) );
  OAI21_X1 U22687 ( .B1(n20581), .B2(n20626), .A(n20580), .ZN(U240) );
  INV_X1 U22688 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20583) );
  AOI22_X1 U22689 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n20608), .ZN(n20582) );
  OAI21_X1 U22690 ( .B1(n20583), .B2(n20626), .A(n20582), .ZN(U239) );
  AOI22_X1 U22691 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n20608), .ZN(n20584) );
  OAI21_X1 U22692 ( .B1(n14610), .B2(n20626), .A(n20584), .ZN(U238) );
  AOI22_X1 U22693 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n20608), .ZN(n20585) );
  OAI21_X1 U22694 ( .B1(n20586), .B2(n20626), .A(n20585), .ZN(U237) );
  INV_X1 U22695 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20588) );
  AOI22_X1 U22696 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n20608), .ZN(n20587) );
  OAI21_X1 U22697 ( .B1(n20588), .B2(n20626), .A(n20587), .ZN(U236) );
  INV_X1 U22698 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20590) );
  AOI22_X1 U22699 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n20608), .ZN(n20589) );
  OAI21_X1 U22700 ( .B1(n20590), .B2(n20626), .A(n20589), .ZN(U235) );
  INV_X1 U22701 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20592) );
  AOI22_X1 U22702 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n20608), .ZN(n20591) );
  OAI21_X1 U22703 ( .B1(n20592), .B2(n20626), .A(n20591), .ZN(U234) );
  INV_X1 U22704 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20594) );
  INV_X1 U22705 ( .A(U212), .ZN(n20621) );
  AOI22_X1 U22706 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n20621), .ZN(n20593) );
  OAI21_X1 U22707 ( .B1(n20594), .B2(n20626), .A(n20593), .ZN(U233) );
  INV_X1 U22708 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20596) );
  AOI22_X1 U22709 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n20608), .ZN(n20595) );
  OAI21_X1 U22710 ( .B1(n20596), .B2(n20626), .A(n20595), .ZN(U232) );
  INV_X1 U22711 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n22421) );
  AOI22_X1 U22712 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n20621), .ZN(n20597) );
  OAI21_X1 U22713 ( .B1(n22421), .B2(n20626), .A(n20597), .ZN(U231) );
  AOI22_X1 U22714 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n20608), .ZN(n20598) );
  OAI21_X1 U22715 ( .B1(n20599), .B2(n20626), .A(n20598), .ZN(U230) );
  INV_X1 U22716 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n22557) );
  AOI22_X1 U22717 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n20608), .ZN(n20600) );
  OAI21_X1 U22718 ( .B1(n22557), .B2(n20626), .A(n20600), .ZN(U229) );
  AOI22_X1 U22719 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n20621), .ZN(n20601) );
  OAI21_X1 U22720 ( .B1(n20602), .B2(n20626), .A(n20601), .ZN(U228) );
  INV_X1 U22721 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n22631) );
  AOI22_X1 U22722 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n20608), .ZN(n20603) );
  OAI21_X1 U22723 ( .B1(n22631), .B2(n20626), .A(n20603), .ZN(U227) );
  AOI22_X1 U22724 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n20621), .ZN(n20604) );
  OAI21_X1 U22725 ( .B1(n20605), .B2(n20626), .A(n20604), .ZN(U226) );
  AOI22_X1 U22726 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n20608), .ZN(n20606) );
  OAI21_X1 U22727 ( .B1(n20607), .B2(n20626), .A(n20606), .ZN(U225) );
  AOI22_X1 U22728 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n20608), .ZN(n20609) );
  OAI21_X1 U22729 ( .B1(n20610), .B2(n20626), .A(n20609), .ZN(U224) );
  INV_X1 U22730 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n22412) );
  AOI22_X1 U22731 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n20621), .ZN(n20611) );
  OAI21_X1 U22732 ( .B1(n22412), .B2(n20626), .A(n20611), .ZN(U223) );
  AOI22_X1 U22733 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n20621), .ZN(n20612) );
  OAI21_X1 U22734 ( .B1(n20613), .B2(n20626), .A(n20612), .ZN(U222) );
  AOI22_X1 U22735 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n20621), .ZN(n20614) );
  OAI21_X1 U22736 ( .B1(n17075), .B2(n20626), .A(n20614), .ZN(U221) );
  AOI22_X1 U22737 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n20621), .ZN(n20616) );
  OAI21_X1 U22738 ( .B1(n20617), .B2(n20626), .A(n20616), .ZN(U220) );
  INV_X1 U22739 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n22628) );
  AOI22_X1 U22740 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n20621), .ZN(n20618) );
  OAI21_X1 U22741 ( .B1(n22628), .B2(n20626), .A(n20618), .ZN(U219) );
  AOI22_X1 U22742 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n20621), .ZN(n20619) );
  OAI21_X1 U22743 ( .B1(n20620), .B2(n20626), .A(n20619), .ZN(U218) );
  AOI22_X1 U22744 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20615), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n20621), .ZN(n20622) );
  OAI21_X1 U22745 ( .B1(n20623), .B2(n20626), .A(n20622), .ZN(U217) );
  OAI222_X1 U22746 ( .A1(U212), .A2(n20627), .B1(n20626), .B2(n20625), .C1(
        U214), .C2(n20624), .ZN(U216) );
  AOI22_X1 U22747 ( .A1(n22805), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20628), 
        .B2(n22806), .ZN(P1_U3483) );
  OAI21_X1 U22748 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n21370), .A(n21371), 
        .ZN(n20630) );
  INV_X1 U22749 ( .A(n22297), .ZN(n22290) );
  AOI211_X1 U22750 ( .C1(n20631), .C2(n20630), .A(n22290), .B(n20629), .ZN(
        n20632) );
  OAI21_X1 U22751 ( .B1(n20632), .B2(n21841), .A(n21843), .ZN(n20637) );
  AOI22_X1 U22752 ( .A1(n21785), .A2(n22297), .B1(n20633), .B2(n21847), .ZN(
        n20635) );
  INV_X1 U22753 ( .A(n20682), .ZN(n20634) );
  NAND2_X1 U22754 ( .A1(n20635), .A2(n20634), .ZN(n20636) );
  MUX2_X1 U22755 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .B(n20637), .S(n20636), 
        .Z(P3_U3296) );
  NAND2_X1 U22756 ( .A1(n20638), .A2(n21118), .ZN(n20672) );
  OR2_X1 U22757 ( .A1(n21827), .A2(n20639), .ZN(n20680) );
  AOI22_X1 U22758 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20677), .ZN(n20640) );
  OAI21_X1 U22759 ( .B1(n21274), .B2(n20672), .A(n20640), .ZN(P3_U2768) );
  AOI22_X1 U22760 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20678), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20677), .ZN(n20641) );
  OAI21_X1 U22761 ( .B1(n21205), .B2(n20680), .A(n20641), .ZN(P3_U2769) );
  AOI22_X1 U22762 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20677), .ZN(n20642) );
  OAI21_X1 U22763 ( .B1(n21211), .B2(n20672), .A(n20642), .ZN(P3_U2770) );
  AOI22_X1 U22764 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20677), .ZN(n20643) );
  OAI21_X1 U22765 ( .B1(n21168), .B2(n20672), .A(n20643), .ZN(P3_U2771) );
  AOI22_X1 U22766 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20669), .ZN(n20644) );
  OAI21_X1 U22767 ( .B1(n21191), .B2(n20672), .A(n20644), .ZN(P3_U2772) );
  AOI22_X1 U22768 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20669), .ZN(n20645) );
  OAI21_X1 U22769 ( .B1(n21159), .B2(n20672), .A(n20645), .ZN(P3_U2773) );
  AOI22_X1 U22770 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20669), .ZN(n20646) );
  OAI21_X1 U22771 ( .B1(n21199), .B2(n20672), .A(n20646), .ZN(P3_U2774) );
  AOI22_X1 U22772 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20669), .ZN(n20647) );
  OAI21_X1 U22773 ( .B1(n21150), .B2(n20672), .A(n20647), .ZN(P3_U2775) );
  AOI22_X1 U22774 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20678), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20677), .ZN(n20648) );
  OAI21_X1 U22775 ( .B1(n21255), .B2(n20680), .A(n20648), .ZN(P3_U2776) );
  INV_X1 U22776 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21146) );
  AOI22_X1 U22777 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20669), .ZN(n20649) );
  OAI21_X1 U22778 ( .B1(n21146), .B2(n20672), .A(n20649), .ZN(P3_U2777) );
  INV_X1 U22779 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n20667) );
  AOI22_X1 U22780 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20669), .ZN(n20650) );
  OAI21_X1 U22781 ( .B1(n20667), .B2(n20672), .A(n20650), .ZN(P3_U2778) );
  INV_X1 U22782 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n21135) );
  AOI22_X1 U22783 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20669), .ZN(n20651) );
  OAI21_X1 U22784 ( .B1(n21135), .B2(n20672), .A(n20651), .ZN(P3_U2779) );
  INV_X1 U22785 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21129) );
  AOI22_X1 U22786 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n20670), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20677), .ZN(n20652) );
  OAI21_X1 U22787 ( .B1(n21129), .B2(n20672), .A(n20652), .ZN(P3_U2780) );
  AOI22_X1 U22788 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20678), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20677), .ZN(n20653) );
  OAI21_X1 U22789 ( .B1(n20654), .B2(n20680), .A(n20653), .ZN(P3_U2781) );
  AOI22_X1 U22790 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20678), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20677), .ZN(n20655) );
  OAI21_X1 U22791 ( .B1(n21236), .B2(n20680), .A(n20655), .ZN(P3_U2782) );
  AOI22_X1 U22792 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20677), .ZN(n20656) );
  OAI21_X1 U22793 ( .B1(n21274), .B2(n20672), .A(n20656), .ZN(P3_U2783) );
  AOI22_X1 U22794 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20678), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20677), .ZN(n20657) );
  OAI21_X1 U22795 ( .B1(n21296), .B2(n20680), .A(n20657), .ZN(P3_U2784) );
  AOI22_X1 U22796 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20677), .ZN(n20658) );
  OAI21_X1 U22797 ( .B1(n21211), .B2(n20672), .A(n20658), .ZN(P3_U2785) );
  AOI22_X1 U22798 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20677), .ZN(n20659) );
  OAI21_X1 U22799 ( .B1(n21168), .B2(n20672), .A(n20659), .ZN(P3_U2786) );
  AOI22_X1 U22800 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20677), .ZN(n20660) );
  OAI21_X1 U22801 ( .B1(n21191), .B2(n20672), .A(n20660), .ZN(P3_U2787) );
  AOI22_X1 U22802 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20677), .ZN(n20661) );
  OAI21_X1 U22803 ( .B1(n21159), .B2(n20672), .A(n20661), .ZN(P3_U2788) );
  AOI22_X1 U22804 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20677), .ZN(n20662) );
  OAI21_X1 U22805 ( .B1(n21199), .B2(n20672), .A(n20662), .ZN(P3_U2789) );
  AOI22_X1 U22806 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20677), .ZN(n20663) );
  OAI21_X1 U22807 ( .B1(n21150), .B2(n20672), .A(n20663), .ZN(P3_U2790) );
  AOI22_X1 U22808 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20678), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20677), .ZN(n20664) );
  OAI21_X1 U22809 ( .B1(n21287), .B2(n20680), .A(n20664), .ZN(P3_U2791) );
  AOI22_X1 U22810 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20669), .ZN(n20665) );
  OAI21_X1 U22811 ( .B1(n21146), .B2(n20672), .A(n20665), .ZN(P3_U2792) );
  AOI22_X1 U22812 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20669), .ZN(n20666) );
  OAI21_X1 U22813 ( .B1(n20667), .B2(n20672), .A(n20666), .ZN(P3_U2793) );
  AOI22_X1 U22814 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20669), .ZN(n20668) );
  OAI21_X1 U22815 ( .B1(n21135), .B2(n20672), .A(n20668), .ZN(P3_U2794) );
  AOI22_X1 U22816 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n20670), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20669), .ZN(n20671) );
  OAI21_X1 U22817 ( .B1(n21129), .B2(n20672), .A(n20671), .ZN(P3_U2795) );
  AOI22_X1 U22818 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20678), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20677), .ZN(n20673) );
  OAI21_X1 U22819 ( .B1(n20674), .B2(n20680), .A(n20673), .ZN(P3_U2796) );
  AOI22_X1 U22820 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20678), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20677), .ZN(n20675) );
  OAI21_X1 U22821 ( .B1(n20676), .B2(n20680), .A(n20675), .ZN(P3_U2797) );
  AOI22_X1 U22822 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20678), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20677), .ZN(n20679) );
  OAI21_X1 U22823 ( .B1(n21282), .B2(n20680), .A(n20679), .ZN(P3_U2798) );
  INV_X1 U22824 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20873) );
  NOR4_X4 U22825 ( .A1(n21314), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .A4(P3_STATEBS16_REG_SCAN_IN), .ZN(n21056)
         );
  OAI21_X1 U22826 ( .B1(n21080), .B2(n20873), .A(n21056), .ZN(n20849) );
  INV_X1 U22827 ( .A(n21056), .ZN(n21833) );
  NOR2_X1 U22828 ( .A1(n21080), .A2(n21833), .ZN(n20846) );
  NOR2_X1 U22829 ( .A1(n21830), .A2(n20681), .ZN(n21837) );
  NOR2_X2 U22830 ( .A1(n21836), .A2(n11157), .ZN(n21023) );
  AOI21_X1 U22831 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20846), .A(
        n21023), .ZN(n20692) );
  OAI211_X1 U22832 ( .C1(n21371), .C2(n21370), .A(n22297), .B(n22243), .ZN(
        n21828) );
  INV_X1 U22833 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n21095) );
  INV_X1 U22834 ( .A(n20686), .ZN(n20683) );
  OAI211_X2 U22835 ( .C1(n21095), .C2(n20684), .A(n21828), .B(n20683), .ZN(
        n21107) );
  OAI22_X1 U22836 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20996), .B1(n21107), 
        .B2(n20694), .ZN(n20690) );
  NAND2_X1 U22837 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n21370), .ZN(n20685) );
  AOI211_X4 U22838 ( .C1(n22297), .C2(n22243), .A(n20686), .B(n20685), .ZN(
        n21072) );
  NAND2_X1 U22839 ( .A1(n20687), .A2(n21344), .ZN(n21313) );
  OAI22_X1 U22840 ( .A1(n21106), .A2(n20688), .B1(n21313), .B2(n21113), .ZN(
        n20689) );
  AOI211_X1 U22841 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n11157), .A(n20690), .B(
        n20689), .ZN(n20691) );
  OAI221_X1 U22842 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20849), .C1(
        n20693), .C2(n20692), .A(n20691), .ZN(P3_U2670) );
  NAND2_X1 U22843 ( .A1(n20695), .A2(n20694), .ZN(n20696) );
  NOR3_X1 U22844 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20715) );
  AOI211_X1 U22845 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20696), .A(n20715), .B(
        n21106), .ZN(n20701) );
  NAND2_X1 U22846 ( .A1(n21056), .A2(n21080), .ZN(n20788) );
  AOI21_X1 U22847 ( .B1(n21342), .B2(n21344), .A(n20710), .ZN(n21330) );
  AOI22_X1 U22848 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n11157), .B1(n21330), 
        .B2(n20721), .ZN(n20698) );
  NAND2_X1 U22849 ( .A1(n20873), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20776) );
  INV_X1 U22850 ( .A(n20776), .ZN(n20834) );
  OAI221_X1 U22851 ( .B1(n20834), .B2(n20699), .C1(n20776), .C2(n18798), .A(
        n20846), .ZN(n20697) );
  OAI211_X1 U22852 ( .C1(n20788), .C2(n20699), .A(n20698), .B(n20697), .ZN(
        n20700) );
  AOI211_X1 U22853 ( .C1(n21023), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n20701), .B(n20700), .ZN(n20703) );
  NAND2_X1 U22854 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20706) );
  OAI211_X1 U22855 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20980), .B(n20706), .ZN(n20702) );
  OAI211_X1 U22856 ( .C1(n20704), .C2(n21107), .A(n20703), .B(n20702), .ZN(
        P3_U2669) );
  NOR2_X1 U22857 ( .A1(n20705), .A2(n20706), .ZN(n20735) );
  INV_X1 U22858 ( .A(n11157), .ZN(n21110) );
  OAI21_X1 U22859 ( .B1(n20735), .B2(n20996), .A(n21110), .ZN(n20731) );
  OAI21_X1 U22860 ( .B1(n20996), .B2(n20706), .A(n20705), .ZN(n20713) );
  OAI21_X1 U22861 ( .B1(n18798), .B2(n20776), .A(n21054), .ZN(n20708) );
  OAI21_X1 U22862 ( .B1(n20709), .B2(n20708), .A(n21056), .ZN(n20707) );
  AOI21_X1 U22863 ( .B1(n20709), .B2(n20708), .A(n20707), .ZN(n20712) );
  NOR2_X1 U22864 ( .A1(n20710), .A2(n21361), .ZN(n21352) );
  NOR2_X1 U22865 ( .A1(n18321), .A2(n21352), .ZN(n21336) );
  OAI22_X1 U22866 ( .A1(n21336), .A2(n21113), .B1(n21107), .B2(n20714), .ZN(
        n20711) );
  AOI211_X1 U22867 ( .C1(n20731), .C2(n20713), .A(n20712), .B(n20711), .ZN(
        n20717) );
  NAND2_X1 U22868 ( .A1(n20715), .A2(n20714), .ZN(n20723) );
  OAI211_X1 U22869 ( .C1(n20715), .C2(n20714), .A(n21072), .B(n20723), .ZN(
        n20716) );
  OAI211_X1 U22870 ( .C1(n21096), .C2(n20718), .A(n20717), .B(n20716), .ZN(
        P3_U2668) );
  AOI21_X1 U22871 ( .B1(n20873), .B2(n20719), .A(n21080), .ZN(n20740) );
  INV_X1 U22872 ( .A(n20740), .ZN(n20738) );
  NOR3_X1 U22873 ( .A1(n20730), .A2(n21833), .A3(n20738), .ZN(n20720) );
  AOI221_X1 U22874 ( .B1(n20722), .B2(n20721), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n20721), .A(n20720), .ZN(
        n20734) );
  NOR2_X1 U22875 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20723), .ZN(n20742) );
  AOI211_X1 U22876 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20723), .A(n20742), .B(
        n21106), .ZN(n20727) );
  NAND2_X1 U22877 ( .A1(n20980), .A2(n20735), .ZN(n20725) );
  OAI22_X1 U22878 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20725), .B1(n20724), 
        .B2(n21096), .ZN(n20726) );
  AOI211_X1 U22879 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n21087), .A(n20727), .B(
        n20726), .ZN(n20733) );
  AOI21_X1 U22880 ( .B1(n20728), .B2(n20788), .A(n20849), .ZN(n20729) );
  AOI22_X1 U22881 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20731), .B1(n20730), 
        .B2(n20729), .ZN(n20732) );
  NAND4_X1 U22882 ( .A1(n20734), .A2(n20733), .A3(n20732), .A4(n11165), .ZN(
        P3_U2667) );
  INV_X1 U22883 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20749) );
  NAND2_X1 U22884 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20735), .ZN(n20737) );
  NOR2_X1 U22885 ( .A1(n20736), .A2(n20737), .ZN(n20765) );
  OAI21_X1 U22886 ( .B1(n20765), .B2(n20996), .A(n21110), .ZN(n20771) );
  OAI21_X1 U22887 ( .B1(n20996), .B2(n20737), .A(n20736), .ZN(n20747) );
  INV_X1 U22888 ( .A(n20739), .ZN(n20741) );
  OAI221_X1 U22889 ( .B1(n20741), .B2(n20740), .C1(n20739), .C2(n20738), .A(
        n21056), .ZN(n20744) );
  NAND2_X1 U22890 ( .A1(n20742), .A2(n20749), .ZN(n20752) );
  OAI211_X1 U22891 ( .C1(n20742), .C2(n20749), .A(n21072), .B(n20752), .ZN(
        n20743) );
  OAI211_X1 U22892 ( .C1(n21096), .C2(n20745), .A(n20744), .B(n20743), .ZN(
        n20746) );
  AOI21_X1 U22893 ( .B1(n20771), .B2(n20747), .A(n20746), .ZN(n20748) );
  OAI211_X1 U22894 ( .C1(n21107), .C2(n20749), .A(n20748), .B(n11165), .ZN(
        P3_U2666) );
  OAI21_X1 U22895 ( .B1(n20750), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21054), .ZN(n20763) );
  NOR3_X1 U22896 ( .A1(n20751), .A2(n21833), .A3(n20763), .ZN(n20754) );
  NOR2_X1 U22897 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20752), .ZN(n20766) );
  AOI211_X1 U22898 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20752), .A(n20766), .B(
        n21106), .ZN(n20753) );
  AOI211_X1 U22899 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n20771), .A(n20754), .B(
        n20753), .ZN(n20762) );
  INV_X1 U22900 ( .A(n20765), .ZN(n20755) );
  NOR3_X1 U22901 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20996), .A3(n20755), .ZN(
        n20772) );
  AOI211_X1 U22902 ( .C1(n20757), .C2(n20788), .A(n20849), .B(n20756), .ZN(
        n20760) );
  AOI22_X1 U22903 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n21023), .B1(
        n21087), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n20758) );
  INV_X1 U22904 ( .A(n20758), .ZN(n20759) );
  NOR4_X1 U22905 ( .A1(n21537), .A2(n20772), .A3(n20760), .A4(n20759), .ZN(
        n20761) );
  NAND2_X1 U22906 ( .A1(n20762), .A2(n20761), .ZN(P3_U2665) );
  XOR2_X1 U22907 ( .A(n20764), .B(n20763), .Z(n20775) );
  NAND2_X1 U22908 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20765), .ZN(n20782) );
  NOR3_X1 U22909 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20996), .A3(n20782), .ZN(
        n20770) );
  NAND2_X1 U22910 ( .A1(n20766), .A2(n20768), .ZN(n20780) );
  OAI211_X1 U22911 ( .C1(n20766), .C2(n20768), .A(n21072), .B(n20780), .ZN(
        n20767) );
  OAI211_X1 U22912 ( .C1(n21107), .C2(n20768), .A(n11165), .B(n20767), .ZN(
        n20769) );
  AOI211_X1 U22913 ( .C1(n21023), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20770), .B(n20769), .ZN(n20774) );
  OAI21_X1 U22914 ( .B1(n20772), .B2(n20771), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n20773) );
  OAI211_X1 U22915 ( .C1(n20775), .C2(n21833), .A(n20774), .B(n20773), .ZN(
        P3_U2664) );
  OAI21_X1 U22916 ( .B1(n20777), .B2(n20776), .A(n21054), .ZN(n20778) );
  XNOR2_X1 U22917 ( .A(n20779), .B(n20778), .ZN(n20787) );
  NOR2_X1 U22918 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20780), .ZN(n20803) );
  OR2_X1 U22919 ( .A1(n21106), .A2(n20803), .ZN(n20801) );
  AOI21_X1 U22920 ( .B1(n20780), .B2(P3_EBX_REG_8__SCAN_IN), .A(n20801), .ZN(
        n20781) );
  AOI21_X1 U22921 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n21087), .A(n20781), .ZN(
        n20786) );
  NOR2_X1 U22922 ( .A1(n21470), .A2(n20782), .ZN(n20783) );
  NAND2_X1 U22923 ( .A1(n20980), .A2(n20783), .ZN(n20791) );
  NAND2_X1 U22924 ( .A1(n20996), .A2(n21110), .ZN(n21108) );
  NAND2_X1 U22925 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n20783), .ZN(n20903) );
  NOR2_X1 U22926 ( .A1(n11157), .A2(n20903), .ZN(n20818) );
  OR2_X1 U22927 ( .A1(n21062), .A2(n20818), .ZN(n20806) );
  AOI21_X1 U22928 ( .B1(n20792), .B2(n20791), .A(n20806), .ZN(n20784) );
  AOI211_X1 U22929 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n21023), .A(
        n21537), .B(n20784), .ZN(n20785) );
  OAI211_X1 U22930 ( .C1(n21833), .C2(n20787), .A(n20786), .B(n20785), .ZN(
        P3_U2663) );
  AOI211_X1 U22931 ( .C1(n20789), .C2(n20788), .A(n20849), .B(n20798), .ZN(
        n20796) );
  AOI21_X1 U22932 ( .B1(n21072), .B2(n20803), .A(n21087), .ZN(n20790) );
  OAI22_X1 U22933 ( .A1(n20811), .A2(n20806), .B1(n20802), .B2(n20790), .ZN(
        n20795) );
  NOR2_X1 U22934 ( .A1(n20792), .A2(n20791), .ZN(n20833) );
  INV_X1 U22935 ( .A(n20833), .ZN(n20891) );
  OAI22_X1 U22936 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20891), .B1(n20793), 
        .B2(n21096), .ZN(n20794) );
  NOR4_X1 U22937 ( .A1(n21537), .A2(n20796), .A3(n20795), .A4(n20794), .ZN(
        n20800) );
  AOI21_X1 U22938 ( .B1(n20797), .B2(n20873), .A(n21080), .ZN(n20809) );
  NAND3_X1 U22939 ( .A1(n21056), .A2(n20809), .A3(n20798), .ZN(n20799) );
  OAI211_X1 U22940 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n20801), .A(n20800), .B(
        n20799), .ZN(P3_U2662) );
  INV_X1 U22941 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20817) );
  NAND2_X1 U22942 ( .A1(n20803), .A2(n20802), .ZN(n20804) );
  NOR2_X1 U22943 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20804), .ZN(n20823) );
  AOI211_X1 U22944 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20804), .A(n20823), .B(
        n21106), .ZN(n20805) );
  AOI211_X1 U22945 ( .C1(n21087), .C2(P3_EBX_REG_10__SCAN_IN), .A(n21780), .B(
        n20805), .ZN(n20816) );
  OAI21_X1 U22946 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n20891), .A(n20806), .ZN(
        n20814) );
  INV_X1 U22947 ( .A(n20808), .ZN(n20810) );
  INV_X1 U22948 ( .A(n20809), .ZN(n20807) );
  AOI221_X1 U22949 ( .B1(n20810), .B2(n20809), .C1(n20808), .C2(n20807), .A(
        n21833), .ZN(n20813) );
  NOR3_X1 U22950 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20811), .A3(n20891), 
        .ZN(n20812) );
  AOI211_X1 U22951 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n20814), .A(n20813), 
        .B(n20812), .ZN(n20815) );
  OAI211_X1 U22952 ( .C1(n20817), .C2(n21096), .A(n20816), .B(n20815), .ZN(
        P3_U2661) );
  INV_X1 U22953 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20830) );
  NAND2_X1 U22954 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n20819) );
  NOR2_X1 U22955 ( .A1(n21503), .A2(n20819), .ZN(n20889) );
  AOI21_X1 U22956 ( .B1(n20889), .B2(n20818), .A(n21062), .ZN(n20862) );
  OAI21_X1 U22957 ( .B1(n20819), .B2(n20891), .A(n21503), .ZN(n20828) );
  AOI21_X1 U22958 ( .B1(n20835), .B2(n20834), .A(n21080), .ZN(n20821) );
  AOI21_X1 U22959 ( .B1(n20822), .B2(n20821), .A(n21833), .ZN(n20820) );
  OAI21_X1 U22960 ( .B1(n20822), .B2(n20821), .A(n20820), .ZN(n20825) );
  NAND2_X1 U22961 ( .A1(n20823), .A2(n20830), .ZN(n20831) );
  OAI211_X1 U22962 ( .C1(n20823), .C2(n20830), .A(n21072), .B(n20831), .ZN(
        n20824) );
  OAI211_X1 U22963 ( .C1(n21096), .C2(n20826), .A(n20825), .B(n20824), .ZN(
        n20827) );
  AOI21_X1 U22964 ( .B1(n20862), .B2(n20828), .A(n20827), .ZN(n20829) );
  OAI211_X1 U22965 ( .C1(n21107), .C2(n20830), .A(n20829), .B(n11165), .ZN(
        P3_U2660) );
  NOR2_X1 U22966 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20831), .ZN(n20851) );
  AOI211_X1 U22967 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20831), .A(n20851), .B(
        n21106), .ZN(n20832) );
  AOI211_X1 U22968 ( .C1(n21087), .C2(P3_EBX_REG_12__SCAN_IN), .A(n21537), .B(
        n20832), .ZN(n20842) );
  NAND2_X1 U22969 ( .A1(n20889), .A2(n20833), .ZN(n20864) );
  INV_X1 U22970 ( .A(n20864), .ZN(n20882) );
  NAND3_X1 U22971 ( .A1(n20835), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n20834), .ZN(n20844) );
  NAND2_X1 U22972 ( .A1(n21054), .A2(n20844), .ZN(n20837) );
  OAI21_X1 U22973 ( .B1(n20838), .B2(n20837), .A(n21056), .ZN(n20836) );
  AOI21_X1 U22974 ( .B1(n20838), .B2(n20837), .A(n20836), .ZN(n20839) );
  AOI221_X1 U22975 ( .B1(n20862), .B2(P3_REIP_REG_12__SCAN_IN), .C1(n20882), 
        .C2(n20840), .A(n20839), .ZN(n20841) );
  OAI211_X1 U22976 ( .C1(n20843), .C2(n21096), .A(n20842), .B(n20841), .ZN(
        P3_U2659) );
  NOR2_X1 U22977 ( .A1(n20845), .A2(n20844), .ZN(n20859) );
  INV_X1 U22978 ( .A(n20846), .ZN(n21092) );
  NOR2_X1 U22979 ( .A1(n20859), .A2(n21092), .ZN(n20847) );
  AOI22_X1 U22980 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n21023), .B1(
        n20847), .B2(n20848), .ZN(n20858) );
  AOI211_X1 U22981 ( .C1(n21054), .C2(n20850), .A(n20849), .B(n20848), .ZN(
        n20855) );
  NAND2_X1 U22982 ( .A1(n20851), .A2(n20853), .ZN(n20867) );
  OAI211_X1 U22983 ( .C1(n20851), .C2(n20853), .A(n21072), .B(n20867), .ZN(
        n20852) );
  OAI21_X1 U22984 ( .B1(n20853), .B2(n21107), .A(n20852), .ZN(n20854) );
  AOI211_X1 U22985 ( .C1(n20862), .C2(P3_REIP_REG_13__SCAN_IN), .A(n20855), 
        .B(n20854), .ZN(n20857) );
  NAND2_X1 U22986 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n20866) );
  OAI211_X1 U22987 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(P3_REIP_REG_12__SCAN_IN), .A(n20882), .B(n20866), .ZN(n20856) );
  NAND4_X1 U22988 ( .A1(n20858), .A2(n20857), .A3(n11165), .A4(n20856), .ZN(
        P3_U2658) );
  NOR2_X1 U22989 ( .A1(n20859), .A2(n21080), .ZN(n20860) );
  XNOR2_X1 U22990 ( .A(n20861), .B(n20860), .ZN(n20872) );
  AOI21_X1 U22991 ( .B1(n21087), .B2(P3_EBX_REG_14__SCAN_IN), .A(n21537), .ZN(
        n20871) );
  NOR2_X1 U22992 ( .A1(n20865), .A2(n20866), .ZN(n20890) );
  INV_X1 U22993 ( .A(n20890), .ZN(n20863) );
  AOI21_X1 U22994 ( .B1(n20980), .B2(n20863), .A(n20862), .ZN(n20893) );
  AOI221_X1 U22995 ( .B1(n20866), .B2(n20865), .C1(n20864), .C2(n20865), .A(
        n20893), .ZN(n20869) );
  NOR2_X1 U22996 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20867), .ZN(n20878) );
  AOI211_X1 U22997 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20867), .A(n20878), .B(
        n21106), .ZN(n20868) );
  AOI211_X1 U22998 ( .C1(n21023), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20869), .B(n20868), .ZN(n20870) );
  OAI211_X1 U22999 ( .C1(n21833), .C2(n20872), .A(n20871), .B(n20870), .ZN(
        P3_U2657) );
  AOI22_X1 U23000 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n21023), .B1(
        n21087), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n20881) );
  AOI21_X1 U23001 ( .B1(n20874), .B2(n20873), .A(n21080), .ZN(n20888) );
  OAI211_X1 U23002 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(n21054), .B(n20876), .ZN(n20875)
         );
  OAI211_X1 U23003 ( .C1(n20876), .C2(n20888), .A(n21056), .B(n20875), .ZN(
        n20880) );
  NAND2_X1 U23004 ( .A1(n20878), .A2(n20877), .ZN(n20885) );
  OAI211_X1 U23005 ( .C1(n20878), .C2(n20877), .A(n21072), .B(n20885), .ZN(
        n20879) );
  AND4_X1 U23006 ( .A1(n20881), .A2(n11165), .A3(n20880), .A4(n20879), .ZN(
        n20883) );
  NAND3_X1 U23007 ( .A1(n20890), .A2(n20882), .A3(n20884), .ZN(n20892) );
  OAI211_X1 U23008 ( .C1(n20893), .C2(n20884), .A(n20883), .B(n20892), .ZN(
        P3_U2656) );
  NOR2_X1 U23009 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20885), .ZN(n20910) );
  AOI211_X1 U23010 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20885), .A(n20910), .B(
        n21106), .ZN(n20886) );
  AOI211_X1 U23011 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n21023), .A(
        n21780), .B(n20886), .ZN(n20898) );
  XNOR2_X1 U23012 ( .A(n20888), .B(n20887), .ZN(n20896) );
  NAND3_X1 U23013 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n20890), .A3(n20889), 
        .ZN(n20902) );
  NOR3_X1 U23014 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n20902), .A3(n20891), 
        .ZN(n20895) );
  AOI21_X1 U23015 ( .B1(n20893), .B2(n20892), .A(n21751), .ZN(n20894) );
  AOI211_X1 U23016 ( .C1(n21056), .C2(n20896), .A(n20895), .B(n20894), .ZN(
        n20897) );
  OAI211_X1 U23017 ( .C1(n21107), .C2(n20899), .A(n20898), .B(n20897), .ZN(
        P3_U2655) );
  OAI21_X1 U23018 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20914), .A(
        n21054), .ZN(n20900) );
  XNOR2_X1 U23019 ( .A(n20901), .B(n20900), .ZN(n20909) );
  NOR3_X1 U23020 ( .A1(n21751), .A2(n20903), .A3(n20902), .ZN(n20905) );
  NAND2_X1 U23021 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n20905), .ZN(n20938) );
  AOI21_X1 U23022 ( .B1(n20980), .B2(n20938), .A(n11157), .ZN(n20922) );
  AND2_X1 U23023 ( .A1(n20938), .A2(n20980), .ZN(n20904) );
  AOI22_X1 U23024 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n21023), .B1(
        n20905), .B2(n20904), .ZN(n20906) );
  OAI211_X1 U23025 ( .C1(n20922), .C2(n20907), .A(n20906), .B(n11165), .ZN(
        n20908) );
  AOI21_X1 U23026 ( .B1(n21056), .B2(n20909), .A(n20908), .ZN(n20912) );
  NAND2_X1 U23027 ( .A1(n20910), .A2(n20913), .ZN(n20916) );
  OAI211_X1 U23028 ( .C1(n20910), .C2(n20913), .A(n21072), .B(n20916), .ZN(
        n20911) );
  OAI211_X1 U23029 ( .C1(n20913), .C2(n21107), .A(n20912), .B(n20911), .ZN(
        P3_U2654) );
  NOR3_X1 U23030 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n11638), .A3(
        n20914), .ZN(n20923) );
  NOR2_X1 U23031 ( .A1(n20923), .A2(n21080), .ZN(n20915) );
  XOR2_X1 U23032 ( .A(n20924), .B(n20915), .Z(n20921) );
  NOR2_X1 U23033 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20916), .ZN(n20933) );
  AOI211_X1 U23034 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20916), .A(n20933), .B(
        n21106), .ZN(n20919) );
  NOR2_X1 U23035 ( .A1(n20996), .A2(n20938), .ZN(n20934) );
  AOI22_X1 U23036 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n21023), .B1(
        n20934), .B2(n21735), .ZN(n20917) );
  OAI211_X1 U23037 ( .C1(n20922), .C2(n21735), .A(n20917), .B(n11165), .ZN(
        n20918) );
  AOI211_X1 U23038 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n21087), .A(n20919), .B(
        n20918), .ZN(n20920) );
  OAI21_X1 U23039 ( .B1(n21833), .B2(n20921), .A(n20920), .ZN(P3_U2653) );
  INV_X1 U23040 ( .A(n20922), .ZN(n20931) );
  AND2_X1 U23041 ( .A1(n20924), .A2(n20923), .ZN(n20925) );
  AOI211_X1 U23042 ( .C1(n20927), .C2(n20926), .A(n20941), .B(n21833), .ZN(
        n20930) );
  INV_X1 U23043 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20932) );
  OAI22_X1 U23044 ( .A1(n20928), .A2(n21096), .B1(n21107), .B2(n20932), .ZN(
        n20929) );
  AOI211_X1 U23045 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n20931), .A(n20930), 
        .B(n20929), .ZN(n20937) );
  NAND2_X1 U23046 ( .A1(n20933), .A2(n20932), .ZN(n20940) );
  OAI211_X1 U23047 ( .C1(n20933), .C2(n20932), .A(n21072), .B(n20940), .ZN(
        n20936) );
  NAND2_X1 U23048 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n20939) );
  OAI211_X1 U23049 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(P3_REIP_REG_19__SCAN_IN), .A(n20934), .B(n20939), .ZN(n20935) );
  NAND4_X1 U23050 ( .A1(n20937), .A2(n11165), .A3(n20936), .A4(n20935), .ZN(
        P3_U2652) );
  NOR2_X1 U23051 ( .A1(n20939), .A2(n20938), .ZN(n20947) );
  NAND2_X1 U23052 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20947), .ZN(n20978) );
  AOI21_X1 U23053 ( .B1(n20980), .B2(n20978), .A(n11157), .ZN(n20976) );
  AOI22_X1 U23054 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n21023), .B1(
        n21087), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n20949) );
  NOR2_X1 U23055 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20996), .ZN(n20946) );
  NOR2_X1 U23056 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20940), .ZN(n20962) );
  AOI211_X1 U23057 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20940), .A(n20962), .B(
        n21106), .ZN(n20945) );
  AOI211_X1 U23058 ( .C1(n20943), .C2(n20942), .A(n20951), .B(n21833), .ZN(
        n20944) );
  AOI211_X1 U23059 ( .C1(n20947), .C2(n20946), .A(n20945), .B(n20944), .ZN(
        n20948) );
  OAI211_X1 U23060 ( .C1(n20950), .C2(n20976), .A(n20949), .B(n20948), .ZN(
        P3_U2651) );
  OR2_X1 U23061 ( .A1(n20996), .A2(n20978), .ZN(n20965) );
  INV_X1 U23062 ( .A(n20976), .ZN(n20960) );
  NOR2_X1 U23063 ( .A1(n20951), .A2(n21080), .ZN(n20955) );
  INV_X1 U23064 ( .A(n20955), .ZN(n20953) );
  INV_X1 U23065 ( .A(n20968), .ZN(n20954) );
  AOI211_X1 U23066 ( .C1(n20956), .C2(n20955), .A(n20954), .B(n21833), .ZN(
        n20959) );
  OAI22_X1 U23067 ( .A1(n20957), .A2(n21096), .B1(n21107), .B2(n20961), .ZN(
        n20958) );
  AOI211_X1 U23068 ( .C1(n20960), .C2(P3_REIP_REG_21__SCAN_IN), .A(n20959), 
        .B(n20958), .ZN(n20964) );
  NAND2_X1 U23069 ( .A1(n20962), .A2(n20961), .ZN(n20967) );
  OAI211_X1 U23070 ( .C1(n20962), .C2(n20961), .A(n21072), .B(n20967), .ZN(
        n20963) );
  OAI211_X1 U23071 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n20965), .A(n20964), 
        .B(n20963), .ZN(P3_U2650) );
  AOI22_X1 U23072 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n21023), .B1(
        n21087), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n20975) );
  AOI211_X1 U23073 ( .C1(n20977), .C2(n20966), .A(n20996), .B(n20978), .ZN(
        n20973) );
  NAND2_X1 U23074 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n20979) );
  NOR2_X1 U23075 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n20967), .ZN(n20990) );
  AOI211_X1 U23076 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20967), .A(n20990), .B(
        n21106), .ZN(n20972) );
  NOR2_X1 U23077 ( .A1(n20970), .A2(n20969), .ZN(n20983) );
  AOI211_X1 U23078 ( .C1(n20970), .C2(n20969), .A(n20983), .B(n21833), .ZN(
        n20971) );
  AOI211_X1 U23079 ( .C1(n20973), .C2(n20979), .A(n20972), .B(n20971), .ZN(
        n20974) );
  OAI211_X1 U23080 ( .C1(n20977), .C2(n20976), .A(n20975), .B(n20974), .ZN(
        P3_U2649) );
  NOR2_X1 U23081 ( .A1(n20979), .A2(n20978), .ZN(n20981) );
  NAND2_X1 U23082 ( .A1(n20980), .A2(n20981), .ZN(n20993) );
  NAND2_X1 U23083 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n20981), .ZN(n20995) );
  NOR2_X1 U23084 ( .A1(n11157), .A2(n20995), .ZN(n21014) );
  NOR2_X1 U23085 ( .A1(n21062), .A2(n21014), .ZN(n20994) );
  NOR2_X1 U23086 ( .A1(n20983), .A2(n21080), .ZN(n20984) );
  NOR2_X1 U23087 ( .A1(n20985), .A2(n20984), .ZN(n20998) );
  AOI211_X1 U23088 ( .C1(n20985), .C2(n20984), .A(n20998), .B(n21833), .ZN(
        n20988) );
  OAI22_X1 U23089 ( .A1(n20986), .A2(n21096), .B1(n21107), .B2(n20989), .ZN(
        n20987) );
  AOI211_X1 U23090 ( .C1(n20994), .C2(P3_REIP_REG_23__SCAN_IN), .A(n20988), 
        .B(n20987), .ZN(n20992) );
  NAND2_X1 U23091 ( .A1(n20990), .A2(n20989), .ZN(n20997) );
  OAI211_X1 U23092 ( .C1(n20990), .C2(n20989), .A(n21072), .B(n20997), .ZN(
        n20991) );
  OAI211_X1 U23093 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n20993), .A(n20992), 
        .B(n20991), .ZN(P3_U2648) );
  INV_X1 U23094 ( .A(n20994), .ZN(n21005) );
  AOI22_X1 U23095 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n21023), .B1(
        n21087), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n21004) );
  NOR2_X1 U23096 ( .A1(n20996), .A2(n20995), .ZN(n21007) );
  NOR2_X1 U23097 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n20997), .ZN(n21013) );
  AOI211_X1 U23098 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n20997), .A(n21013), .B(
        n21106), .ZN(n21002) );
  NOR2_X1 U23099 ( .A1(n20998), .A2(n21080), .ZN(n20999) );
  NOR2_X1 U23100 ( .A1(n21000), .A2(n20999), .ZN(n21008) );
  AOI211_X1 U23101 ( .C1(n21000), .C2(n20999), .A(n21008), .B(n21833), .ZN(
        n21001) );
  AOI211_X1 U23102 ( .C1(n21007), .C2(n21006), .A(n21002), .B(n21001), .ZN(
        n21003) );
  OAI211_X1 U23103 ( .C1(n21006), .C2(n21005), .A(n21004), .B(n21003), .ZN(
        P3_U2647) );
  AOI22_X1 U23104 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n21023), .B1(
        n21087), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n21018) );
  AND2_X1 U23105 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21007), .ZN(n21019) );
  NOR2_X1 U23106 ( .A1(n21008), .A2(n21080), .ZN(n21009) );
  NOR2_X1 U23107 ( .A1(n21010), .A2(n21009), .ZN(n21027) );
  AOI211_X1 U23108 ( .C1(n21010), .C2(n21009), .A(n21027), .B(n21833), .ZN(
        n21011) );
  AOI21_X1 U23109 ( .B1(n21019), .B2(n21021), .A(n21011), .ZN(n21017) );
  NAND2_X1 U23110 ( .A1(n21013), .A2(n21012), .ZN(n21022) );
  OAI211_X1 U23111 ( .C1(n21013), .C2(n21012), .A(n21072), .B(n21022), .ZN(
        n21016) );
  NAND2_X1 U23112 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21014), .ZN(n21020) );
  NAND3_X1 U23113 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n21108), .A3(n21020), 
        .ZN(n21015) );
  NAND4_X1 U23114 ( .A1(n21018), .A2(n21017), .A3(n21016), .A4(n21015), .ZN(
        P3_U2646) );
  NAND2_X1 U23115 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n21019), .ZN(n21032) );
  NOR3_X1 U23116 ( .A1(n21021), .A2(n21033), .A3(n21020), .ZN(n21049) );
  NOR2_X1 U23117 ( .A1(n21062), .A2(n21049), .ZN(n21036) );
  NOR2_X1 U23118 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n21022), .ZN(n21038) );
  AOI211_X1 U23119 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n21022), .A(n21038), .B(
        n21106), .ZN(n21026) );
  AOI22_X1 U23120 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n21023), .B1(
        n21087), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n21024) );
  INV_X1 U23121 ( .A(n21024), .ZN(n21025) );
  AOI211_X1 U23122 ( .C1(n21036), .C2(P3_REIP_REG_26__SCAN_IN), .A(n21026), 
        .B(n21025), .ZN(n21031) );
  INV_X1 U23123 ( .A(n21029), .ZN(n21040) );
  NOR2_X1 U23124 ( .A1(n21027), .A2(n21080), .ZN(n21039) );
  INV_X1 U23125 ( .A(n21039), .ZN(n21028) );
  OAI221_X1 U23126 ( .B1(n21040), .B2(n21039), .C1(n21029), .C2(n21028), .A(
        n21056), .ZN(n21030) );
  OAI211_X1 U23127 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n21032), .A(n21031), 
        .B(n21030), .ZN(P3_U2645) );
  NOR2_X1 U23128 ( .A1(n21033), .A2(n21032), .ZN(n21047) );
  INV_X1 U23129 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n21037) );
  OAI22_X1 U23130 ( .A1(n11647), .A2(n21096), .B1(n21107), .B2(n21037), .ZN(
        n21034) );
  AOI221_X1 U23131 ( .B1(n21036), .B2(P3_REIP_REG_27__SCAN_IN), .C1(n21047), 
        .C2(n21035), .A(n21034), .ZN(n21046) );
  NAND2_X1 U23132 ( .A1(n21038), .A2(n21037), .ZN(n21048) );
  OAI211_X1 U23133 ( .C1(n21038), .C2(n21037), .A(n21072), .B(n21048), .ZN(
        n21045) );
  AOI21_X1 U23134 ( .B1(n21040), .B2(n21054), .A(n21039), .ZN(n21043) );
  INV_X1 U23135 ( .A(n21041), .ZN(n21042) );
  OAI211_X1 U23136 ( .C1(n21043), .C2(n21042), .A(n21056), .B(n21055), .ZN(
        n21044) );
  NAND3_X1 U23137 ( .A1(n21046), .A2(n21045), .A3(n21044), .ZN(P3_U2644) );
  NAND2_X1 U23138 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n21047), .ZN(n21064) );
  NOR2_X1 U23139 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n21048), .ZN(n21071) );
  AOI211_X1 U23140 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n21048), .A(n21071), .B(
        n21106), .ZN(n21053) );
  NAND2_X1 U23141 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n21049), .ZN(n21061) );
  NAND2_X1 U23142 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n21061), .ZN(n21051) );
  OAI22_X1 U23143 ( .A1(n21062), .A2(n21051), .B1(n21050), .B2(n21096), .ZN(
        n21052) );
  AOI211_X1 U23144 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n21087), .A(n21053), .B(
        n21052), .ZN(n21060) );
  NAND2_X1 U23145 ( .A1(n21055), .A2(n21054), .ZN(n21067) );
  INV_X1 U23146 ( .A(n21067), .ZN(n21057) );
  OAI221_X1 U23147 ( .B1(n21058), .B2(n21057), .C1(n21066), .C2(n21067), .A(
        n21056), .ZN(n21059) );
  OAI211_X1 U23148 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n21064), .A(n21060), 
        .B(n21059), .ZN(P3_U2643) );
  NOR2_X1 U23149 ( .A1(n21065), .A2(n21061), .ZN(n21063) );
  AOI21_X1 U23150 ( .B1(n21063), .B2(P3_REIP_REG_29__SCAN_IN), .A(n21062), 
        .ZN(n21101) );
  AOI22_X1 U23151 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n21101), .B1(n21087), 
        .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n21078) );
  NOR2_X1 U23152 ( .A1(n21065), .A2(n21064), .ZN(n21082) );
  NOR2_X1 U23153 ( .A1(n21068), .A2(n21069), .ZN(n21081) );
  AOI211_X1 U23154 ( .C1(n21069), .C2(n21068), .A(n21081), .B(n21833), .ZN(
        n21075) );
  INV_X1 U23155 ( .A(n21071), .ZN(n21073) );
  NAND2_X1 U23156 ( .A1(n21071), .A2(n21070), .ZN(n21086) );
  NAND2_X1 U23157 ( .A1(n21072), .A2(n21086), .ZN(n21084) );
  AOI21_X1 U23158 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n21073), .A(n21084), .ZN(
        n21074) );
  OAI211_X1 U23159 ( .C1(n21079), .C2(n21096), .A(n21078), .B(n21077), .ZN(
        P3_U2642) );
  XNOR2_X1 U23160 ( .A(n21094), .B(n21093), .ZN(n21090) );
  NAND2_X1 U23161 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n21082), .ZN(n21105) );
  NOR2_X1 U23162 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n21105), .ZN(n21102) );
  OAI22_X1 U23163 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n21084), .B1(n21083), 
        .B2(n21096), .ZN(n21085) );
  AOI211_X1 U23164 ( .C1(P3_REIP_REG_30__SCAN_IN), .C2(n21101), .A(n21102), 
        .B(n21085), .ZN(n21089) );
  NOR2_X1 U23165 ( .A1(n21106), .A2(n21086), .ZN(n21100) );
  OAI21_X1 U23166 ( .B1(n21087), .B2(n21100), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n21088) );
  OAI211_X1 U23167 ( .C1(n21833), .C2(n21090), .A(n21089), .B(n21088), .ZN(
        P3_U2641) );
  NAND2_X1 U23168 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n21091), .ZN(n21104) );
  OAI22_X1 U23169 ( .A1(n21097), .A2(n21096), .B1(n21095), .B2(n21107), .ZN(
        n21098) );
  OAI21_X1 U23170 ( .B1(n21102), .B2(n21101), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n21103) );
  NAND2_X1 U23171 ( .A1(n21107), .A2(n21106), .ZN(n21109) );
  AOI22_X1 U23172 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n21109), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n21108), .ZN(n21112) );
  NAND3_X1 U23173 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21110), .A3(
        n21308), .ZN(n21111) );
  OAI211_X1 U23174 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n21113), .A(
        n21112), .B(n21111), .ZN(P3_U2671) );
  NOR3_X1 U23175 ( .A1(n21370), .A2(n21115), .A3(n21114), .ZN(n21116) );
  NAND4_X1 U23176 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n21119) );
  NOR3_X1 U23177 ( .A1(n21148), .A2(n21170), .A3(n21119), .ZN(n21176) );
  AND3_X1 U23178 ( .A1(n21219), .A2(n21294), .A3(n21176), .ZN(n21288) );
  NAND2_X1 U23179 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21288), .ZN(n21140) );
  NOR2_X1 U23180 ( .A1(n21141), .A2(n21140), .ZN(n21145) );
  NAND2_X1 U23181 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n21145), .ZN(n21137) );
  NOR2_X1 U23182 ( .A1(n21130), .A2(n21137), .ZN(n21134) );
  NAND2_X1 U23183 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n21134), .ZN(n21126) );
  NAND2_X1 U23184 ( .A1(n21126), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n21125) );
  NOR2_X1 U23185 ( .A1(n21120), .A2(n21121), .ZN(n21303) );
  AOI22_X1 U23186 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21303), .B1(n21302), .B2(
        n21123), .ZN(n21124) );
  OAI221_X1 U23187 ( .B1(n21126), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n21125), 
        .C2(n21295), .A(n21124), .ZN(P3_U2722) );
  INV_X1 U23188 ( .A(n21126), .ZN(n21276) );
  AOI21_X1 U23189 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n21290), .A(n21134), .ZN(
        n21128) );
  OAI222_X1 U23190 ( .A1(n21175), .A2(n21129), .B1(n21276), .B2(n21128), .C1(
        n21300), .C2(n21127), .ZN(P3_U2723) );
  OAI21_X1 U23191 ( .B1(n21130), .B2(n21295), .A(n21137), .ZN(n21131) );
  INV_X1 U23192 ( .A(n21131), .ZN(n21133) );
  OAI222_X1 U23193 ( .A1(n21175), .A2(n21135), .B1(n21134), .B2(n21133), .C1(
        n21300), .C2(n21132), .ZN(P3_U2724) );
  AOI22_X1 U23194 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21303), .B1(n21302), .B2(
        n21136), .ZN(n21139) );
  OAI211_X1 U23195 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n21145), .A(n21290), .B(
        n21137), .ZN(n21138) );
  NAND2_X1 U23196 ( .A1(n21139), .A2(n21138), .ZN(P3_U2725) );
  OAI21_X1 U23197 ( .B1(n21141), .B2(n21295), .A(n21140), .ZN(n21142) );
  INV_X1 U23198 ( .A(n21142), .ZN(n21144) );
  OAI222_X1 U23199 ( .A1(n21175), .A2(n21146), .B1(n21145), .B2(n21144), .C1(
        n21300), .C2(n21143), .ZN(P3_U2726) );
  NAND2_X1 U23200 ( .A1(n21219), .A2(n21294), .ZN(n21169) );
  NOR2_X1 U23201 ( .A1(n21170), .A2(n21169), .ZN(n21174) );
  NAND2_X1 U23202 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n21174), .ZN(n21160) );
  NOR2_X1 U23203 ( .A1(n21147), .A2(n21160), .ZN(n21164) );
  NAND2_X1 U23204 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n21164), .ZN(n21151) );
  NOR2_X1 U23205 ( .A1(n21148), .A2(n21151), .ZN(n21155) );
  AOI21_X1 U23206 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n21290), .A(n21155), .ZN(
        n21149) );
  OAI222_X1 U23207 ( .A1(n21175), .A2(n21150), .B1(n21288), .B2(n21149), .C1(
        n21300), .C2(n21655), .ZN(P3_U2728) );
  INV_X1 U23208 ( .A(n21151), .ZN(n21158) );
  AOI21_X1 U23209 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n21290), .A(n21158), .ZN(
        n21154) );
  INV_X1 U23210 ( .A(n21152), .ZN(n21153) );
  OAI222_X1 U23211 ( .A1(n21199), .A2(n21175), .B1(n21155), .B2(n21154), .C1(
        n21300), .C2(n21153), .ZN(P3_U2729) );
  AOI21_X1 U23212 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n21290), .A(n21164), .ZN(
        n21157) );
  OAI222_X1 U23213 ( .A1(n21159), .A2(n21175), .B1(n21158), .B2(n21157), .C1(
        n21300), .C2(n21156), .ZN(P3_U2730) );
  INV_X1 U23214 ( .A(n21160), .ZN(n21167) );
  AOI21_X1 U23215 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n21290), .A(n21167), .ZN(
        n21163) );
  INV_X1 U23216 ( .A(n21161), .ZN(n21162) );
  OAI222_X1 U23217 ( .A1(n21191), .A2(n21175), .B1(n21164), .B2(n21163), .C1(
        n21300), .C2(n21162), .ZN(P3_U2731) );
  AOI21_X1 U23218 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n21290), .A(n21174), .ZN(
        n21166) );
  OAI222_X1 U23219 ( .A1(n21168), .A2(n21175), .B1(n21167), .B2(n21166), .C1(
        n21300), .C2(n21165), .ZN(P3_U2732) );
  OAI21_X1 U23220 ( .B1(n21170), .B2(n21295), .A(n21169), .ZN(n21171) );
  INV_X1 U23221 ( .A(n21171), .ZN(n21173) );
  OAI222_X1 U23222 ( .A1(n21211), .A2(n21175), .B1(n21174), .B2(n21173), .C1(
        n21300), .C2(n21172), .ZN(P3_U2733) );
  NAND4_X1 U23223 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(P3_EAX_REG_13__SCAN_IN), .ZN(n21177)
         );
  NAND4_X1 U23224 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(n21178), .ZN(n21283) );
  NAND2_X1 U23225 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n21218) );
  NAND2_X1 U23226 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n21206), .ZN(n21200) );
  INV_X1 U23227 ( .A(n21200), .ZN(n21188) );
  NAND2_X1 U23228 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n21188), .ZN(n21187) );
  NAND2_X1 U23229 ( .A1(n21290), .A2(n21187), .ZN(n21192) );
  NAND2_X1 U23230 ( .A1(n15979), .A2(n21295), .ZN(n21275) );
  NOR2_X1 U23231 ( .A1(n21290), .A2(n21180), .ZN(n21270) );
  OAI22_X1 U23232 ( .A1(n21182), .A2(n21300), .B1(n21181), .B2(n21253), .ZN(
        n21183) );
  AOI21_X1 U23233 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n21266), .A(n21183), .ZN(
        n21184) );
  OAI221_X1 U23234 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21187), .C1(n21185), 
        .C2(n21192), .A(n21184), .ZN(P3_U2714) );
  AOI22_X1 U23235 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n21270), .B1(n21302), .B2(
        n21186), .ZN(n21190) );
  OAI211_X1 U23236 ( .C1(n21188), .C2(P3_EAX_REG_20__SCAN_IN), .A(n21290), .B(
        n21187), .ZN(n21189) );
  OAI211_X1 U23237 ( .C1(n21275), .C2(n21191), .A(n21190), .B(n21189), .ZN(
        P3_U2715) );
  NAND2_X1 U23238 ( .A1(n21219), .A2(n21305), .ZN(n21306) );
  OAI21_X1 U23239 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21306), .A(n21192), .ZN(
        n21197) );
  NAND2_X1 U23240 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .ZN(n21217) );
  NOR3_X1 U23241 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n21217), .A3(n21200), .ZN(
        n21196) );
  OAI22_X1 U23242 ( .A1(n21194), .A2(n21300), .B1(n21193), .B2(n21253), .ZN(
        n21195) );
  AOI211_X1 U23243 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n21197), .A(n21196), .B(
        n21195), .ZN(n21198) );
  OAI21_X1 U23244 ( .B1(n21199), .B2(n21275), .A(n21198), .ZN(P3_U2713) );
  AOI22_X1 U23245 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21266), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n21270), .ZN(n21202) );
  OAI211_X1 U23246 ( .C1(n21206), .C2(P3_EAX_REG_19__SCAN_IN), .A(n21290), .B(
        n21200), .ZN(n21201) );
  OAI211_X1 U23247 ( .C1(n21203), .C2(n21300), .A(n21202), .B(n21201), .ZN(
        P3_U2716) );
  AOI22_X1 U23248 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n21270), .B1(n21302), .B2(
        n21204), .ZN(n21210) );
  OR2_X1 U23249 ( .A1(n21205), .A2(n21271), .ZN(n21212) );
  AOI211_X1 U23250 ( .C1(n21207), .C2(n21212), .A(n21206), .B(n21295), .ZN(
        n21208) );
  INV_X1 U23251 ( .A(n21208), .ZN(n21209) );
  OAI211_X1 U23252 ( .C1(n21275), .C2(n21211), .A(n21210), .B(n21209), .ZN(
        P3_U2717) );
  AOI22_X1 U23253 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21266), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n21270), .ZN(n21214) );
  OAI211_X1 U23254 ( .C1(n11423), .C2(P3_EAX_REG_17__SCAN_IN), .A(n21290), .B(
        n21212), .ZN(n21213) );
  OAI211_X1 U23255 ( .C1(n21215), .C2(n21300), .A(n21214), .B(n21213), .ZN(
        P3_U2718) );
  AOI22_X1 U23256 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21266), .B1(n21302), .B2(
        n21216), .ZN(n21223) );
  NAND2_X1 U23257 ( .A1(n21219), .A2(n21262), .ZN(n21254) );
  AOI211_X1 U23258 ( .C1(n21220), .C2(n21256), .A(n21225), .B(n21295), .ZN(
        n21221) );
  INV_X1 U23259 ( .A(n21221), .ZN(n21222) );
  OAI211_X1 U23260 ( .C1(n21253), .C2(n21224), .A(n21223), .B(n21222), .ZN(
        P3_U2710) );
  AOI22_X1 U23261 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21266), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n21270), .ZN(n21227) );
  OAI211_X1 U23262 ( .C1(n21225), .C2(P3_EAX_REG_26__SCAN_IN), .A(n21290), .B(
        n21247), .ZN(n21226) );
  OAI211_X1 U23263 ( .C1(n21228), .C2(n21300), .A(n21227), .B(n21226), .ZN(
        P3_U2709) );
  NAND2_X1 U23264 ( .A1(n21239), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n21238) );
  NOR2_X1 U23265 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n21238), .ZN(n21229) );
  OAI22_X1 U23266 ( .A1(n21232), .A2(n21300), .B1(n21231), .B2(n21253), .ZN(
        n21233) );
  AOI21_X1 U23267 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n21266), .A(n21233), .ZN(
        n21234) );
  OAI221_X1 U23268 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n21238), .C1(n21236), 
        .C2(n21235), .A(n21234), .ZN(P3_U2705) );
  AOI22_X1 U23269 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21266), .B1(n21302), .B2(
        n21237), .ZN(n21241) );
  OAI211_X1 U23270 ( .C1(n21239), .C2(P3_EAX_REG_29__SCAN_IN), .A(n21290), .B(
        n21238), .ZN(n21240) );
  OAI211_X1 U23271 ( .C1(n21253), .C2(n17051), .A(n21241), .B(n21240), .ZN(
        P3_U2706) );
  AOI22_X1 U23272 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21266), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n21270), .ZN(n21244) );
  OAI211_X1 U23273 ( .C1(n11265), .C2(P3_EAX_REG_28__SCAN_IN), .A(n21290), .B(
        n21242), .ZN(n21243) );
  OAI211_X1 U23274 ( .C1(n21245), .C2(n21300), .A(n21244), .B(n21243), .ZN(
        P3_U2707) );
  AOI22_X1 U23275 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21266), .B1(n21302), .B2(
        n21246), .ZN(n21251) );
  AOI211_X1 U23276 ( .C1(n21248), .C2(n21247), .A(n11265), .B(n21295), .ZN(
        n21249) );
  INV_X1 U23277 ( .A(n21249), .ZN(n21250) );
  OAI211_X1 U23278 ( .C1(n21253), .C2(n21252), .A(n21251), .B(n21250), .ZN(
        P3_U2708) );
  AOI22_X1 U23279 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21266), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n21270), .ZN(n21259) );
  OAI21_X1 U23280 ( .B1(n21255), .B2(n21295), .A(n21254), .ZN(n21257) );
  NAND2_X1 U23281 ( .A1(n21257), .A2(n21256), .ZN(n21258) );
  OAI211_X1 U23282 ( .C1(n21260), .C2(n21300), .A(n21259), .B(n21258), .ZN(
        P3_U2711) );
  AOI22_X1 U23283 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n21270), .B1(n21302), .B2(
        n21261), .ZN(n21268) );
  AOI211_X1 U23284 ( .C1(n21264), .C2(n21263), .A(n21295), .B(n21262), .ZN(
        n21265) );
  AOI21_X1 U23285 ( .B1(n21266), .B2(BUF2_REG_7__SCAN_IN), .A(n21265), .ZN(
        n21267) );
  NAND2_X1 U23286 ( .A1(n21268), .A2(n21267), .ZN(P3_U2712) );
  AOI22_X1 U23287 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n21270), .B1(n21302), .B2(
        n21269), .ZN(n21273) );
  OAI211_X1 U23288 ( .C1(n21281), .C2(P3_EAX_REG_16__SCAN_IN), .A(n21290), .B(
        n21271), .ZN(n21272) );
  OAI211_X1 U23289 ( .C1(n21275), .C2(n21274), .A(n21273), .B(n21272), .ZN(
        P3_U2719) );
  NAND2_X1 U23290 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n21276), .ZN(n21280) );
  AOI22_X1 U23291 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21303), .B1(n21302), .B2(
        n21277), .ZN(n21279) );
  NAND3_X1 U23292 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n21290), .A3(n21283), 
        .ZN(n21278) );
  OAI211_X1 U23293 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n21280), .A(n21279), .B(
        n21278), .ZN(P3_U2721) );
  AOI211_X1 U23294 ( .C1(n21283), .C2(n21282), .A(n21295), .B(n21281), .ZN(
        n21284) );
  AOI21_X1 U23295 ( .B1(n21303), .B2(BUF2_REG_15__SCAN_IN), .A(n21284), .ZN(
        n21285) );
  OAI21_X1 U23296 ( .B1(n21286), .B2(n21300), .A(n21285), .ZN(P3_U2720) );
  AOI22_X1 U23297 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21303), .B1(n21288), .B2(
        n21287), .ZN(n21292) );
  NAND3_X1 U23298 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21290), .A3(n21289), .ZN(
        n21291) );
  OAI211_X1 U23299 ( .C1(n21293), .C2(n21300), .A(n21292), .B(n21291), .ZN(
        P3_U2727) );
  AOI211_X1 U23300 ( .C1(n21297), .C2(n21296), .A(n21295), .B(n21294), .ZN(
        n21298) );
  AOI21_X1 U23301 ( .B1(n21303), .B2(BUF2_REG_1__SCAN_IN), .A(n21298), .ZN(
        n21299) );
  OAI21_X1 U23302 ( .B1(n21301), .B2(n21300), .A(n21299), .ZN(P3_U2734) );
  AOI22_X1 U23303 ( .A1(n21303), .A2(BUF2_REG_0__SCAN_IN), .B1(n21302), .B2(
        n11540), .ZN(n21304) );
  OAI221_X1 U23304 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n21306), .C1(n11420), 
        .C2(n21305), .A(n21304), .ZN(P3_U2735) );
  NOR2_X1 U23305 ( .A1(n21307), .A2(n21606), .ZN(n21312) );
  AOI22_X1 U23306 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21601), .B1(
        n21312), .B2(n21310), .ZN(n21810) );
  INV_X1 U23307 ( .A(n21308), .ZN(n21356) );
  AOI222_X1 U23308 ( .A1(n21532), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21810), 
        .B2(n21356), .C1(n21310), .C2(n21358), .ZN(n21309) );
  INV_X1 U23309 ( .A(n21362), .ZN(n21359) );
  AOI22_X1 U23310 ( .A1(n21362), .A2(n21310), .B1(n21309), .B2(n21359), .ZN(
        P3_U3290) );
  OAI21_X1 U23311 ( .B1(n21775), .B2(n21310), .A(n21318), .ZN(n21323) );
  OAI21_X1 U23312 ( .B1(n21327), .B2(n21323), .A(n21324), .ZN(n21311) );
  OAI21_X1 U23313 ( .B1(n21312), .B2(n21313), .A(n21311), .ZN(n21808) );
  INV_X1 U23314 ( .A(n21313), .ZN(n21315) );
  INV_X1 U23315 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21416) );
  OAI22_X1 U23316 ( .A1(n21416), .A2(n21646), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21317) );
  NOR2_X1 U23317 ( .A1(n21314), .A2(n21532), .ZN(n21332) );
  AOI222_X1 U23318 ( .A1(n21808), .A2(n21356), .B1(n21315), .B2(n21358), .C1(
        n21317), .C2(n21332), .ZN(n21316) );
  AOI22_X1 U23319 ( .A1(n21362), .A2(n21324), .B1(n21316), .B2(n21359), .ZN(
        P3_U3289) );
  INV_X1 U23320 ( .A(n21317), .ZN(n21331) );
  OAI21_X1 U23321 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21318), .A(
        n21348), .ZN(n21322) );
  OAI22_X1 U23322 ( .A1(n21321), .A2(n21320), .B1(n21337), .B2(n21319), .ZN(
        n21351) );
  OAI211_X1 U23323 ( .C1(n21322), .C2(n21351), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n21344), .ZN(n21329) );
  NAND2_X1 U23324 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21323), .ZN(
        n21354) );
  INV_X1 U23325 ( .A(n21354), .ZN(n21326) );
  NAND2_X1 U23326 ( .A1(n21342), .A2(n21324), .ZN(n21325) );
  OAI211_X1 U23327 ( .C1(n21327), .C2(n21326), .A(n21325), .B(n21341), .ZN(
        n21328) );
  OAI211_X1 U23328 ( .C1(n21330), .C2(n21728), .A(n21329), .B(n21328), .ZN(
        n21805) );
  AOI22_X1 U23329 ( .A1(n21332), .A2(n21331), .B1(n21356), .B2(n21805), .ZN(
        n21335) );
  OR3_X1 U23330 ( .A1(n21344), .A2(n21842), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21334) );
  OAI221_X1 U23331 ( .B1(n21362), .B2(n21358), .C1(n21362), .C2(n21344), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21333) );
  OAI221_X1 U23332 ( .B1(n21362), .B2(n21335), .C1(n21362), .C2(n21334), .A(
        n21333), .ZN(P3_U3288) );
  INV_X1 U23333 ( .A(n21336), .ZN(n21357) );
  INV_X1 U23334 ( .A(n21337), .ZN(n21340) );
  AOI21_X1 U23335 ( .B1(n21340), .B2(n21361), .A(n21341), .ZN(n21338) );
  AOI221_X1 U23336 ( .B1(n21341), .B2(n21361), .C1(n21340), .C2(n21339), .A(
        n21338), .ZN(n21350) );
  NAND2_X1 U23337 ( .A1(n21342), .A2(n21344), .ZN(n21343) );
  AOI22_X1 U23338 ( .A1(n21345), .A2(n21344), .B1(n21361), .B2(n21343), .ZN(
        n21346) );
  OAI22_X1 U23339 ( .A1(n21348), .A2(n21347), .B1(n21346), .B2(n21728), .ZN(
        n21349) );
  AOI211_X1 U23340 ( .C1(n21352), .C2(n21351), .A(n21350), .B(n21349), .ZN(
        n21353) );
  OAI21_X1 U23341 ( .B1(n21355), .B2(n21354), .A(n21353), .ZN(n21804) );
  AOI22_X1 U23342 ( .A1(n21358), .A2(n21357), .B1(n21356), .B2(n21804), .ZN(
        n21360) );
  AOI22_X1 U23343 ( .A1(n21362), .A2(n21361), .B1(n21360), .B2(n21359), .ZN(
        P3_U3285) );
  INV_X1 U23344 ( .A(n21363), .ZN(n21365) );
  OAI21_X1 U23345 ( .B1(n21366), .B2(n21365), .A(n21364), .ZN(n21376) );
  AND3_X1 U23346 ( .A1(n21368), .A2(n21367), .A3(n21794), .ZN(n21375) );
  XNOR2_X1 U23347 ( .A(n21370), .B(n21369), .ZN(n21372) );
  OAI21_X1 U23348 ( .B1(n21372), .B2(n21371), .A(n22297), .ZN(n21796) );
  NOR3_X1 U23349 ( .A1(n21373), .A2(n21797), .A3(n21796), .ZN(n21374) );
  AOI211_X1 U23350 ( .C1(n21790), .C2(n21376), .A(n21375), .B(n21374), .ZN(
        n21377) );
  AOI21_X2 U23351 ( .B1(n21378), .B2(n21377), .A(n21847), .ZN(n21653) );
  OAI22_X1 U23352 ( .A1(n21720), .A2(n21489), .B1(n21675), .B2(n21379), .ZN(
        n21498) );
  INV_X1 U23353 ( .A(n21498), .ZN(n21385) );
  NAND2_X1 U23354 ( .A1(n21382), .A2(n21380), .ZN(n21384) );
  INV_X1 U23355 ( .A(n21381), .ZN(n21497) );
  NAND3_X1 U23356 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21455) );
  NAND2_X1 U23357 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21427) );
  NOR2_X1 U23358 ( .A1(n21455), .A2(n21427), .ZN(n21445) );
  NAND2_X1 U23359 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21445), .ZN(
        n21469) );
  NOR2_X1 U23360 ( .A1(n21497), .A2(n21469), .ZN(n21535) );
  INV_X1 U23361 ( .A(n21535), .ZN(n21765) );
  NOR2_X1 U23362 ( .A1(n21532), .A2(n21765), .ZN(n21774) );
  INV_X1 U23363 ( .A(n21774), .ZN(n21507) );
  NOR2_X1 U23364 ( .A1(n21384), .A2(n21507), .ZN(n21605) );
  INV_X1 U23365 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21465) );
  AOI21_X1 U23366 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21428) );
  OR2_X1 U23367 ( .A1(n21455), .A2(n21428), .ZN(n21446) );
  NOR2_X1 U23368 ( .A1(n21465), .A2(n21446), .ZN(n21467) );
  NAND2_X1 U23369 ( .A1(n21381), .A2(n21467), .ZN(n21716) );
  NOR2_X1 U23370 ( .A1(n21384), .A2(n21716), .ZN(n21566) );
  NAND2_X1 U23371 ( .A1(n21382), .A2(n21535), .ZN(n21725) );
  NOR2_X1 U23372 ( .A1(n21383), .A2(n21725), .ZN(n21603) );
  AOI222_X1 U23373 ( .A1(n21606), .A2(n21605), .B1(n21566), .B2(n21789), .C1(
        n21766), .C2(n21603), .ZN(n21615) );
  OAI21_X1 U23374 ( .B1(n21385), .B2(n21384), .A(n21615), .ZN(n21678) );
  NAND2_X1 U23375 ( .A1(n21653), .A2(n21678), .ZN(n21715) );
  INV_X1 U23376 ( .A(n21566), .ZN(n21588) );
  NAND2_X1 U23377 ( .A1(n21789), .A2(n21588), .ZN(n21386) );
  OAI221_X1 U23378 ( .B1(n21601), .B2(n21603), .C1(n21601), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n21386), .ZN(n21696) );
  OAI22_X1 U23379 ( .A1(n21601), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n21387), .B2(n21728), .ZN(n21391) );
  OAI22_X1 U23380 ( .A1(n21389), .A2(n21675), .B1(n21388), .B2(n21720), .ZN(
        n21390) );
  NOR3_X1 U23381 ( .A1(n21696), .A2(n21391), .A3(n21390), .ZN(n21552) );
  OAI21_X1 U23382 ( .B1(n21775), .B2(n21605), .A(n21653), .ZN(n21697) );
  AOI21_X1 U23383 ( .B1(n21606), .B2(n21392), .A(n21697), .ZN(n21393) );
  AOI211_X1 U23384 ( .C1(n21552), .C2(n21393), .A(n21780), .B(n21554), .ZN(
        n21394) );
  AOI21_X1 U23385 ( .B1(n21779), .B2(n21395), .A(n21394), .ZN(n21397) );
  OAI211_X1 U23386 ( .C1(n21398), .C2(n21715), .A(n21397), .B(n21396), .ZN(
        P3_U2841) );
  NAND2_X1 U23387 ( .A1(n21653), .A2(n21788), .ZN(n21458) );
  NAND2_X1 U23388 ( .A1(n11165), .A2(n21764), .ZN(n21755) );
  NOR2_X1 U23389 ( .A1(n11165), .A2(n21399), .ZN(n21402) );
  NAND2_X1 U23390 ( .A1(n21775), .A2(n21728), .ZN(n21705) );
  INV_X1 U23391 ( .A(n21705), .ZN(n21400) );
  AOI221_X1 U23392 ( .B1(n21400), .B2(n21532), .C1(n21601), .C2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n21764), .ZN(n21401) );
  AOI211_X1 U23393 ( .C1(n21681), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n21402), .B(n21401), .ZN(n21403) );
  OAI221_X1 U23394 ( .B1(n21405), .B2(n21458), .C1(n21404), .C2(n21476), .A(
        n21403), .ZN(P3_U2862) );
  NAND3_X1 U23395 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21532), .A3(
        n21705), .ZN(n21407) );
  OAI211_X1 U23396 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n21766), .A(
        n21416), .B(n21748), .ZN(n21406) );
  OAI211_X1 U23397 ( .C1(n21408), .C2(n21795), .A(n21407), .B(n21406), .ZN(
        n21410) );
  INV_X1 U23398 ( .A(n21458), .ZN(n21577) );
  AOI22_X1 U23399 ( .A1(n21653), .A2(n21410), .B1(n21577), .B2(n21409), .ZN(
        n21412) );
  NAND2_X1 U23400 ( .A1(n21780), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n21411) );
  OAI211_X1 U23401 ( .C1(n21755), .C2(n21416), .A(n21412), .B(n21411), .ZN(
        P3_U2861) );
  NOR2_X1 U23402 ( .A1(n21532), .A2(n21427), .ZN(n21424) );
  OAI21_X1 U23403 ( .B1(n21428), .B2(n21424), .A(n21789), .ZN(n21414) );
  NOR2_X1 U23404 ( .A1(n21775), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21722) );
  NOR2_X1 U23405 ( .A1(n21766), .A2(n21606), .ZN(n21565) );
  INV_X1 U23406 ( .A(n21565), .ZN(n21730) );
  OAI211_X1 U23407 ( .C1(n21722), .C2(n21416), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n21730), .ZN(n21413) );
  OAI211_X1 U23408 ( .C1(n21415), .C2(n21795), .A(n21414), .B(n21413), .ZN(
        n21420) );
  AOI21_X1 U23409 ( .B1(n21606), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n21766), .ZN(n21426) );
  OR3_X1 U23410 ( .A1(n21416), .A2(n21426), .A3(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21417) );
  OAI21_X1 U23411 ( .B1(n21418), .B2(n21675), .A(n21417), .ZN(n21419) );
  OAI21_X1 U23412 ( .B1(n21420), .B2(n21419), .A(n21653), .ZN(n21421) );
  OAI211_X1 U23413 ( .C1(n21755), .C2(n18364), .A(n21422), .B(n21421), .ZN(
        P3_U2860) );
  AND2_X1 U23414 ( .A1(n21789), .A2(n21428), .ZN(n21423) );
  AOI211_X1 U23415 ( .C1(n21766), .C2(n21427), .A(n21423), .B(n21443), .ZN(
        n21425) );
  AOI221_X1 U23416 ( .B1(n21775), .B2(n21425), .C1(n21424), .C2(n21425), .A(
        n21764), .ZN(n21435) );
  OAI22_X1 U23417 ( .A1(n21728), .A2(n21428), .B1(n21427), .B2(n21426), .ZN(
        n21434) );
  OAI22_X1 U23418 ( .A1(n21476), .A2(n21430), .B1(n21458), .B2(n21429), .ZN(
        n21431) );
  AOI221_X1 U23419 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21435), .C1(
        n21434), .C2(n21435), .A(n21431), .ZN(n21433) );
  OAI211_X1 U23420 ( .C1(n21755), .C2(n21443), .A(n21433), .B(n21432), .ZN(
        P3_U2859) );
  INV_X1 U23421 ( .A(n21434), .ZN(n21456) );
  NOR4_X1 U23422 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21456), .A3(
        n21764), .A4(n21443), .ZN(n21439) );
  AOI21_X1 U23423 ( .B1(n21435), .B2(n21748), .A(n21681), .ZN(n21437) );
  OAI22_X1 U23424 ( .A1(n21437), .A2(n21444), .B1(n21458), .B2(n21436), .ZN(
        n21438) );
  NOR2_X1 U23425 ( .A1(n21439), .A2(n21438), .ZN(n21441) );
  NAND2_X1 U23426 ( .A1(n18728), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n21440) );
  OAI211_X1 U23427 ( .C1(n21476), .C2(n21442), .A(n21441), .B(n21440), .ZN(
        P3_U2858) );
  NOR4_X1 U23428 ( .A1(n21456), .A2(n21444), .A3(n21764), .A4(n21443), .ZN(
        n21451) );
  INV_X1 U23429 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21450) );
  INV_X1 U23430 ( .A(n21722), .ZN(n21589) );
  OAI211_X1 U23431 ( .C1(n21445), .C2(n21565), .A(n21653), .B(n21589), .ZN(
        n21447) );
  OAI221_X1 U23432 ( .B1(n21447), .B2(n21789), .C1(n21447), .C2(n21446), .A(
        n11165), .ZN(n21464) );
  OAI22_X1 U23433 ( .A1(n21450), .A2(n21464), .B1(n21458), .B2(n21448), .ZN(
        n21449) );
  AOI21_X1 U23434 ( .B1(n21451), .B2(n21450), .A(n21449), .ZN(n21453) );
  OAI211_X1 U23435 ( .C1(n21454), .C2(n21476), .A(n21453), .B(n21452), .ZN(
        P3_U2857) );
  NOR2_X1 U23436 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21764), .ZN(
        n21461) );
  NOR2_X1 U23437 ( .A1(n21456), .A2(n21455), .ZN(n21466) );
  OAI22_X1 U23438 ( .A1(n21476), .A2(n21459), .B1(n21458), .B2(n21457), .ZN(
        n21460) );
  AOI21_X1 U23439 ( .B1(n21461), .B2(n21466), .A(n21460), .ZN(n21463) );
  NAND2_X1 U23440 ( .A1(n21780), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n21462) );
  OAI211_X1 U23441 ( .C1(n21465), .C2(n21464), .A(n21463), .B(n21462), .ZN(
        P3_U2856) );
  NAND2_X1 U23442 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21466), .ZN(
        n21496) );
  OAI211_X1 U23443 ( .C1(n21467), .C2(n21728), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n21589), .ZN(n21468) );
  AOI21_X1 U23444 ( .B1(n21469), .B2(n21730), .A(n21468), .ZN(n21478) );
  AOI211_X1 U23445 ( .C1(n21479), .C2(n21496), .A(n21478), .B(n21764), .ZN(
        n21472) );
  OAI22_X1 U23446 ( .A1(n11165), .A2(n21470), .B1(n21479), .B2(n21755), .ZN(
        n21471) );
  AOI211_X1 U23447 ( .C1(n21473), .C2(n21577), .A(n21472), .B(n21471), .ZN(
        n21474) );
  OAI21_X1 U23448 ( .B1(n21476), .B2(n21475), .A(n21474), .ZN(P3_U2855) );
  NOR3_X1 U23449 ( .A1(n21628), .A2(n21478), .A3(n21477), .ZN(n21481) );
  NOR3_X1 U23450 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21479), .A3(
        n21496), .ZN(n21480) );
  AOI211_X1 U23451 ( .C1(n21487), .C2(n21673), .A(n21481), .B(n21480), .ZN(
        n21482) );
  OAI21_X1 U23452 ( .B1(n21675), .B2(n21483), .A(n21482), .ZN(n21484) );
  AOI22_X1 U23453 ( .A1(n21653), .A2(n21484), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21681), .ZN(n21486) );
  OAI211_X1 U23454 ( .C1(n21487), .C2(n21741), .A(n21486), .B(n21485), .ZN(
        P3_U2854) );
  OR2_X1 U23455 ( .A1(n21728), .A2(n21488), .ZN(n21511) );
  OAI211_X1 U23456 ( .C1(n21775), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n21653), .B(n21511), .ZN(n21495) );
  NAND2_X1 U23457 ( .A1(n21720), .A2(n21675), .ZN(n21724) );
  AOI21_X1 U23458 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21774), .A(
        n21775), .ZN(n21492) );
  NAND2_X1 U23459 ( .A1(n21673), .A2(n21489), .ZN(n21490) );
  NAND2_X1 U23460 ( .A1(n21789), .A2(n21716), .ZN(n21533) );
  OAI211_X1 U23461 ( .C1(n21491), .C2(n21675), .A(n21490), .B(n21533), .ZN(
        n21777) );
  AOI211_X1 U23462 ( .C1(n21499), .C2(n21724), .A(n21492), .B(n21777), .ZN(
        n21767) );
  OAI221_X1 U23463 ( .B1(n21601), .B2(n21493), .C1(n21601), .C2(n21535), .A(
        n21767), .ZN(n21494) );
  OAI21_X1 U23464 ( .B1(n21495), .B2(n21494), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21504) );
  NOR2_X1 U23465 ( .A1(n21497), .A2(n21496), .ZN(n21540) );
  OAI21_X1 U23466 ( .B1(n21540), .B2(n21498), .A(n21653), .ZN(n21784) );
  NOR3_X1 U23467 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21499), .A3(
        n21784), .ZN(n21500) );
  AOI21_X1 U23468 ( .B1(n21779), .B2(n21501), .A(n21500), .ZN(n21502) );
  OAI221_X1 U23469 ( .B1(n18728), .B2(n21504), .C1(n11165), .C2(n21503), .A(
        n21502), .ZN(P3_U2851) );
  AOI22_X1 U23470 ( .A1(n21780), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n21779), 
        .B2(n21505), .ZN(n21516) );
  INV_X1 U23471 ( .A(n21506), .ZN(n21512) );
  OAI21_X1 U23472 ( .B1(n21508), .B2(n21507), .A(n21606), .ZN(n21510) );
  OAI21_X1 U23473 ( .B1(n21508), .B2(n21765), .A(n21766), .ZN(n21509) );
  NAND4_X1 U23474 ( .A1(n21533), .A2(n21511), .A3(n21510), .A4(n21509), .ZN(
        n21519) );
  AOI21_X1 U23475 ( .B1(n21788), .B2(n21512), .A(n21519), .ZN(n21513) );
  OAI21_X1 U23476 ( .B1(n21514), .B2(n21720), .A(n21513), .ZN(n21752) );
  OAI211_X1 U23477 ( .C1(n21764), .C2(n21752), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n11165), .ZN(n21515) );
  OAI211_X1 U23478 ( .C1(n21784), .C2(n21517), .A(n21516), .B(n21515), .ZN(
        P3_U2850) );
  NAND2_X1 U23479 ( .A1(n21518), .A2(n21540), .ZN(n21524) );
  NOR2_X1 U23480 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21728), .ZN(
        n21753) );
  AOI211_X1 U23481 ( .C1(n21748), .C2(n21754), .A(n21753), .B(n21519), .ZN(
        n21523) );
  AOI22_X1 U23482 ( .A1(n21673), .A2(n21521), .B1(n21788), .B2(n21520), .ZN(
        n21522) );
  OAI221_X1 U23483 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21524), 
        .C1(n21529), .C2(n21523), .A(n21522), .ZN(n21526) );
  AOI22_X1 U23484 ( .A1(n21653), .A2(n21526), .B1(n21779), .B2(n21525), .ZN(
        n21528) );
  OAI211_X1 U23485 ( .C1(n21755), .C2(n21529), .A(n21528), .B(n21527), .ZN(
        P3_U2848) );
  INV_X1 U23486 ( .A(n21768), .ZN(n21555) );
  NOR2_X1 U23487 ( .A1(n21720), .A2(n21530), .ZN(n21543) );
  INV_X1 U23488 ( .A(n21543), .ZN(n21531) );
  OAI211_X1 U23489 ( .C1(n21718), .C2(n21675), .A(n21653), .B(n21531), .ZN(
        n21747) );
  OAI22_X1 U23490 ( .A1(n21606), .A2(n21545), .B1(n21532), .B2(n21725), .ZN(
        n21534) );
  OAI211_X1 U23491 ( .C1(n21601), .C2(n21535), .A(n21534), .B(n21533), .ZN(
        n21541) );
  AOI211_X1 U23492 ( .C1(n21555), .C2(n21539), .A(n21747), .B(n21541), .ZN(
        n21536) );
  NOR2_X1 U23493 ( .A1(n21537), .A2(n21536), .ZN(n21746) );
  AOI22_X1 U23494 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21746), .B1(
        n21779), .B2(n21538), .ZN(n21550) );
  AND3_X1 U23495 ( .A1(n21541), .A2(n21540), .A3(n11527), .ZN(n21544) );
  OAI221_X1 U23496 ( .B1(n21544), .B2(n21543), .C1(n21544), .C2(n21542), .A(
        n21653), .ZN(n21549) );
  NAND3_X1 U23497 ( .A1(n21546), .A2(n21577), .A3(n21545), .ZN(n21548) );
  NAND4_X1 U23498 ( .A1(n21550), .A2(n21549), .A3(n21548), .A4(n21547), .ZN(
        P3_U2847) );
  NOR2_X1 U23499 ( .A1(n21551), .A2(n21715), .ZN(n21689) );
  AOI21_X1 U23500 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n21653), .A(
        n21689), .ZN(n21561) );
  AND3_X1 U23501 ( .A1(n21677), .A2(n21603), .A3(n21589), .ZN(n21564) );
  OAI211_X1 U23502 ( .C1(n21775), .C2(n21564), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n21552), .ZN(n21553) );
  AOI21_X1 U23503 ( .B1(n21555), .B2(n21554), .A(n21553), .ZN(n21560) );
  INV_X1 U23504 ( .A(n21556), .ZN(n21557) );
  AOI22_X1 U23505 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21681), .B1(
        n21779), .B2(n21557), .ZN(n21559) );
  OAI211_X1 U23506 ( .C1(n21561), .C2(n21560), .A(n21559), .B(n21558), .ZN(
        P3_U2840) );
  OAI21_X1 U23507 ( .B1(n21615), .B2(n21563), .A(n21562), .ZN(n21571) );
  NOR2_X1 U23508 ( .A1(n21565), .A2(n21564), .ZN(n21671) );
  OAI221_X1 U23509 ( .B1(n21728), .B2(n21566), .C1(n21728), .C2(n21677), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21686) );
  NOR3_X1 U23510 ( .A1(n21671), .A2(n21694), .A3(n21686), .ZN(n21567) );
  OAI21_X1 U23511 ( .B1(n21628), .B2(n21567), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21580) );
  INV_X1 U23512 ( .A(n21568), .ZN(n21570) );
  AOI222_X1 U23513 ( .A1(n21571), .A2(n21580), .B1(n21788), .B2(n21570), .C1(
        n21673), .C2(n21569), .ZN(n21575) );
  AOI22_X1 U23514 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21681), .B1(
        n21779), .B2(n21572), .ZN(n21574) );
  NAND2_X1 U23515 ( .A1(n18728), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21573) );
  OAI211_X1 U23516 ( .C1(n21575), .C2(n21764), .A(n21574), .B(n21573), .ZN(
        P3_U2837) );
  NAND2_X1 U23517 ( .A1(n21577), .A2(n21576), .ZN(n21592) );
  NOR2_X1 U23518 ( .A1(n21590), .A2(n21720), .ZN(n21579) );
  AOI211_X1 U23519 ( .C1(n21748), .C2(n21580), .A(n21579), .B(n21578), .ZN(
        n21583) );
  AOI21_X1 U23520 ( .B1(n21581), .B2(n21678), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21582) );
  AOI211_X1 U23521 ( .C1(n21592), .C2(n21583), .A(n21582), .B(n21764), .ZN(
        n21584) );
  AOI21_X1 U23522 ( .B1(n21681), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n21584), .ZN(n21586) );
  OAI211_X1 U23523 ( .C1(n21587), .C2(n21741), .A(n21586), .B(n21585), .ZN(
        P3_U2836) );
  NAND2_X1 U23524 ( .A1(n21604), .A2(n21678), .ZN(n21650) );
  INV_X1 U23525 ( .A(n21604), .ZN(n21614) );
  OAI21_X1 U23526 ( .B1(n21588), .B2(n21614), .A(n21789), .ZN(n21623) );
  AND2_X1 U23527 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21623), .ZN(
        n21608) );
  OAI211_X1 U23528 ( .C1(n21590), .C2(n21720), .A(n21608), .B(n21589), .ZN(
        n21591) );
  NAND2_X1 U23529 ( .A1(n21603), .A2(n21604), .ZN(n21657) );
  OAI221_X1 U23530 ( .B1(n21591), .B2(n21657), .C1(n21591), .C2(n21730), .A(
        n21653), .ZN(n21593) );
  AOI22_X1 U23531 ( .A1(n21598), .A2(n21650), .B1(n21593), .B2(n21592), .ZN(
        n21594) );
  AOI211_X1 U23532 ( .C1(n21779), .C2(n21596), .A(n21595), .B(n21594), .ZN(
        n21597) );
  OAI21_X1 U23533 ( .B1(n21598), .B2(n21755), .A(n21597), .ZN(P3_U2835) );
  AOI22_X1 U23534 ( .A1(n21673), .A2(n21600), .B1(n21788), .B2(n21599), .ZN(
        n21622) );
  NOR2_X1 U23535 ( .A1(n21614), .A2(n21613), .ZN(n21602) );
  AOI21_X1 U23536 ( .B1(n21603), .B2(n21602), .A(n21601), .ZN(n21625) );
  NAND3_X1 U23537 ( .A1(n21605), .A2(n21604), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21607) );
  NAND2_X1 U23538 ( .A1(n21607), .A2(n21606), .ZN(n21624) );
  OAI211_X1 U23539 ( .C1(n21608), .C2(n21728), .A(n21653), .B(n21624), .ZN(
        n21609) );
  AOI211_X1 U23540 ( .C1(n21610), .C2(n21705), .A(n21625), .B(n21609), .ZN(
        n21611) );
  AOI21_X1 U23541 ( .B1(n21622), .B2(n21611), .A(n21618), .ZN(n21612) );
  AOI22_X1 U23542 ( .A1(n21780), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n21612), 
        .B2(n11165), .ZN(n21620) );
  INV_X1 U23543 ( .A(n21660), .ZN(n21617) );
  NOR3_X1 U23544 ( .A1(n21615), .A2(n21614), .A3(n21613), .ZN(n21638) );
  AOI21_X1 U23545 ( .B1(n21659), .B2(n21673), .A(n21638), .ZN(n21616) );
  OAI21_X1 U23546 ( .B1(n21675), .B2(n21617), .A(n21616), .ZN(n21633) );
  NAND3_X1 U23547 ( .A1(n21653), .A2(n21618), .A3(n21633), .ZN(n21619) );
  OAI211_X1 U23548 ( .C1(n21621), .C2(n21741), .A(n21620), .B(n21619), .ZN(
        P3_U2833) );
  INV_X1 U23549 ( .A(n21622), .ZN(n21629) );
  NAND2_X1 U23550 ( .A1(n21624), .A2(n21623), .ZN(n21656) );
  NOR3_X1 U23551 ( .A1(n21625), .A2(n21630), .A3(n21656), .ZN(n21626) );
  OAI21_X1 U23552 ( .B1(n21628), .B2(n21627), .A(n21626), .ZN(n21641) );
  OAI22_X1 U23553 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(n21629), .B2(n21641), .ZN(
        n21631) );
  OAI22_X1 U23554 ( .A1(n21764), .A2(n21631), .B1(n21755), .B2(n21630), .ZN(
        n21632) );
  OAI21_X1 U23555 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n21633), .A(
        n21632), .ZN(n21634) );
  OAI211_X1 U23556 ( .C1(n21636), .C2(n21741), .A(n21635), .B(n21634), .ZN(
        P3_U2832) );
  AND2_X1 U23557 ( .A1(n21646), .A2(n21637), .ZN(n21639) );
  NAND3_X1 U23558 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21748), .A3(
        n21641), .ZN(n21642) );
  NAND2_X1 U23559 ( .A1(n21648), .A2(n21647), .ZN(n21654) );
  OAI22_X1 U23560 ( .A1(n21651), .A2(n21650), .B1(n21649), .B2(n21654), .ZN(
        n21652) );
  AOI22_X1 U23561 ( .A1(n21653), .A2(n21652), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n11165), .ZN(n21670) );
  OAI21_X1 U23562 ( .B1(n21655), .B2(n21654), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21663) );
  AOI211_X1 U23563 ( .C1(n21766), .C2(n21657), .A(n21681), .B(n21656), .ZN(
        n21658) );
  OAI21_X1 U23564 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21768), .A(
        n21658), .ZN(n21662) );
  OAI22_X1 U23565 ( .A1(n21660), .A2(n21675), .B1(n21659), .B2(n21720), .ZN(
        n21661) );
  AOI211_X1 U23566 ( .C1(n21664), .C2(n21663), .A(n21662), .B(n21661), .ZN(
        n21669) );
  OR3_X1 U23567 ( .A1(n21666), .A2(n21741), .A3(n21665), .ZN(n21667) );
  OAI211_X1 U23568 ( .C1(n21670), .C2(n21669), .A(n21668), .B(n21667), .ZN(
        P3_U2834) );
  AOI211_X1 U23569 ( .C1(n21673), .C2(n21672), .A(n21681), .B(n21671), .ZN(
        n21674) );
  OAI21_X1 U23570 ( .B1(n21676), .B2(n21675), .A(n21674), .ZN(n21687) );
  NAND2_X1 U23571 ( .A1(n21678), .A2(n21677), .ZN(n21680) );
  OAI21_X1 U23572 ( .B1(n21681), .B2(n21680), .A(n21679), .ZN(n21682) );
  OAI211_X1 U23573 ( .C1(n21686), .C2(n21687), .A(n11165), .B(n21682), .ZN(
        n21684) );
  OAI211_X1 U23574 ( .C1(n21741), .C2(n21685), .A(n21684), .B(n21683), .ZN(
        P3_U2839) );
  OAI221_X1 U23575 ( .B1(n21687), .B2(n21748), .C1(n21687), .C2(n21686), .A(
        n11165), .ZN(n21693) );
  AOI22_X1 U23576 ( .A1(n21779), .A2(n21690), .B1(n21689), .B2(n21688), .ZN(
        n21692) );
  OAI211_X1 U23577 ( .C1(n21694), .C2(n21693), .A(n21692), .B(n21691), .ZN(
        P3_U2838) );
  INV_X1 U23578 ( .A(n21695), .ZN(n21700) );
  AOI211_X1 U23579 ( .C1(n21788), .C2(n21698), .A(n21697), .B(n21696), .ZN(
        n21699) );
  OAI21_X1 U23580 ( .B1(n21720), .B2(n21700), .A(n21699), .ZN(n21701) );
  NAND2_X1 U23581 ( .A1(n21701), .A2(n11165), .ZN(n21709) );
  AOI21_X1 U23582 ( .B1(n21779), .B2(n21703), .A(n21702), .ZN(n21704) );
  OAI221_X1 U23583 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21715), 
        .C1(n21706), .C2(n21709), .A(n21704), .ZN(P3_U2843) );
  NAND3_X1 U23584 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21706), .A3(n21705), 
        .ZN(n21708) );
  AOI21_X1 U23585 ( .B1(n21709), .B2(n21708), .A(n21707), .ZN(n21710) );
  AOI211_X1 U23586 ( .C1(n21712), .C2(n21779), .A(n21711), .B(n21710), .ZN(
        n21713) );
  OAI21_X1 U23587 ( .B1(n21715), .B2(n21714), .A(n21713), .ZN(P3_U2842) );
  NOR3_X1 U23588 ( .A1(n21731), .A2(n21717), .A3(n21716), .ZN(n21729) );
  OAI211_X1 U23589 ( .C1(n21721), .C2(n21720), .A(n21719), .B(n21718), .ZN(
        n21723) );
  AOI211_X1 U23590 ( .C1(n21724), .C2(n21723), .A(n21722), .B(n21764), .ZN(
        n21727) );
  OAI21_X1 U23591 ( .B1(n21725), .B2(n21743), .A(n21730), .ZN(n21726) );
  OAI211_X1 U23592 ( .C1(n21729), .C2(n21728), .A(n21727), .B(n21726), .ZN(
        n21737) );
  OAI221_X1 U23593 ( .B1(n21737), .B2(n21738), .C1(n21737), .C2(n21730), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21736) );
  NOR2_X1 U23594 ( .A1(n21731), .A2(n21784), .ZN(n21744) );
  AOI22_X1 U23595 ( .A1(n21779), .A2(n21733), .B1(n21744), .B2(n21732), .ZN(
        n21734) );
  OAI221_X1 U23596 ( .B1(n18728), .B2(n21736), .C1(n11165), .C2(n21735), .A(
        n21734), .ZN(P3_U2844) );
  OAI221_X1 U23597 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n11165), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18728), .A(n21737), .ZN(
        n21740) );
  NAND3_X1 U23598 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21744), .A3(
        n21738), .ZN(n21739) );
  OAI211_X1 U23599 ( .C1(n21742), .C2(n21741), .A(n21740), .B(n21739), .ZN(
        P3_U2845) );
  AOI22_X1 U23600 ( .A1(n21745), .A2(n21779), .B1(n21744), .B2(n21743), .ZN(
        n21750) );
  OAI211_X1 U23601 ( .C1(n21748), .C2(n21747), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n21746), .ZN(n21749) );
  OAI211_X1 U23602 ( .C1(n21751), .C2(n11165), .A(n21750), .B(n21749), .ZN(
        P3_U2846) );
  NOR2_X1 U23603 ( .A1(n21753), .A2(n21752), .ZN(n21756) );
  AOI21_X1 U23604 ( .B1(n21756), .B2(n21755), .A(n21754), .ZN(n21757) );
  AOI22_X1 U23605 ( .A1(n21758), .A2(n21779), .B1(n21757), .B2(n11165), .ZN(
        n21760) );
  OAI211_X1 U23606 ( .C1(n21784), .C2(n21761), .A(n21760), .B(n21759), .ZN(
        P3_U2849) );
  NAND2_X1 U23607 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21762), .ZN(
        n21772) );
  AOI22_X1 U23608 ( .A1(n21780), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21779), 
        .B2(n21763), .ZN(n21771) );
  AOI21_X1 U23609 ( .B1(n21766), .B2(n21765), .A(n21764), .ZN(n21773) );
  OAI211_X1 U23610 ( .C1(n21768), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n21767), .B(n21773), .ZN(n21769) );
  NAND3_X1 U23611 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n11165), .A3(
        n21769), .ZN(n21770) );
  OAI211_X1 U23612 ( .C1(n21772), .C2(n21784), .A(n21771), .B(n21770), .ZN(
        P3_U2852) );
  OAI21_X1 U23613 ( .B1(n21775), .B2(n21774), .A(n21773), .ZN(n21776) );
  OAI21_X1 U23614 ( .B1(n21777), .B2(n21776), .A(n11165), .ZN(n21782) );
  AOI22_X1 U23615 ( .A1(n21780), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n21779), 
        .B2(n21778), .ZN(n21781) );
  OAI221_X1 U23616 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21784), .C1(
        n21783), .C2(n21782), .A(n21781), .ZN(P3_U2853) );
  NAND2_X1 U23617 ( .A1(n22290), .A2(n21785), .ZN(n21840) );
  INV_X1 U23618 ( .A(n21786), .ZN(n21832) );
  INV_X1 U23619 ( .A(n21787), .ZN(n21825) );
  NOR2_X1 U23620 ( .A1(n21789), .A2(n21788), .ZN(n21791) );
  OAI222_X1 U23621 ( .A1(n21795), .A2(n21794), .B1(n21793), .B2(n21792), .C1(
        n21791), .C2(n21790), .ZN(n21849) );
  INV_X1 U23622 ( .A(n21796), .ZN(n21799) );
  NOR3_X1 U23623 ( .A1(n21799), .A2(n21798), .A3(n21797), .ZN(n21848) );
  OAI21_X1 U23624 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21848), .ZN(n21800) );
  OAI211_X1 U23625 ( .C1(n21803), .C2(n21802), .A(n21801), .B(n21800), .ZN(
        n21824) );
  INV_X1 U23626 ( .A(n21803), .ZN(n21813) );
  AOI22_X1 U23627 ( .A1(n21813), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21804), .B2(n21803), .ZN(n21822) );
  MUX2_X1 U23628 ( .A(n21805), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n21813), .Z(n21817) );
  OR3_X1 U23629 ( .A1(n21810), .A2(n21809), .A3(n21806), .ZN(n21807) );
  AOI22_X1 U23630 ( .A1(n21810), .A2(n21809), .B1(n21808), .B2(n21807), .ZN(
        n21812) );
  OAI21_X1 U23631 ( .B1(n21813), .B2(n21812), .A(n21811), .ZN(n21816) );
  AND2_X1 U23632 ( .A1(n21817), .A2(n21816), .ZN(n21814) );
  OAI221_X1 U23633 ( .B1(n21817), .B2(n21816), .C1(n21815), .C2(n21814), .A(
        n21819), .ZN(n21821) );
  AOI21_X1 U23634 ( .B1(n21819), .B2(n21818), .A(n21817), .ZN(n21820) );
  AOI222_X1 U23635 ( .A1(n21822), .A2(n21821), .B1(n21822), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n21821), .C2(n21820), .ZN(
        n21823) );
  NOR4_X1 U23636 ( .A1(n21825), .A2(n21849), .A3(n21824), .A4(n21823), .ZN(
        n21846) );
  OAI211_X1 U23637 ( .C1(n21828), .C2(n21827), .A(n21826), .B(n21846), .ZN(
        n21835) );
  OAI21_X1 U23638 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n22297), .A(n21835), 
        .ZN(n21838) );
  OR3_X1 U23639 ( .A1(n21830), .A2(n21838), .A3(n21829), .ZN(n21831) );
  NAND4_X1 U23640 ( .A1(n21833), .A2(n21840), .A3(n21832), .A4(n21831), .ZN(
        P3_U2997) );
  OAI221_X1 U23641 ( .B1(n21836), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21836), 
        .C2(n21835), .A(n21834), .ZN(P3_U3282) );
  AOI221_X1 U23642 ( .B1(n21839), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21838), 
        .C2(P3_STATE2_REG_0__SCAN_IN), .A(n21837), .ZN(n21845) );
  OAI211_X1 U23643 ( .C1(n21843), .C2(n21842), .A(n21841), .B(n21840), .ZN(
        n21844) );
  OAI211_X1 U23644 ( .C1(n21846), .C2(n21847), .A(n21845), .B(n21844), .ZN(
        P3_U2996) );
  NOR2_X1 U23645 ( .A1(n21848), .A2(n21847), .ZN(n21853) );
  MUX2_X1 U23646 ( .A(P3_MORE_REG_SCAN_IN), .B(n21849), .S(n21853), .Z(
        P3_U3295) );
  INV_X1 U23647 ( .A(n21850), .ZN(n21851) );
  OAI21_X1 U23648 ( .B1(n21853), .B2(n21852), .A(n21851), .ZN(P3_U2637) );
  AOI211_X1 U23649 ( .C1(n21857), .C2(n21856), .A(n21855), .B(n21854), .ZN(
        n21859) );
  OAI21_X1 U23650 ( .B1(n21859), .B2(n22225), .A(n21858), .ZN(n21864) );
  AOI211_X1 U23651 ( .C1(n21862), .C2(n22253), .A(n21861), .B(n21860), .ZN(
        n21863) );
  MUX2_X1 U23652 ( .A(n21864), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21863), 
        .Z(P1_U3485) );
  AOI22_X1 U23653 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21865), .B1(
        n21999), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n21869) );
  AOI22_X1 U23654 ( .A1(n21867), .A2(n22004), .B1(n16757), .B2(n21866), .ZN(
        n21868) );
  OAI211_X1 U23655 ( .C1(n22009), .C2(n21870), .A(n21869), .B(n21868), .ZN(
        P1_U3018) );
  INV_X1 U23656 ( .A(n21871), .ZN(n21875) );
  OAI22_X1 U23657 ( .A1(n21873), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n21872), .B2(n22010), .ZN(n21874) );
  AOI21_X1 U23658 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21875), .A(
        n21874), .ZN(n21877) );
  NAND2_X1 U23659 ( .A1(n21999), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n21876) );
  OAI211_X1 U23660 ( .C1(n22009), .C2(n22036), .A(n21877), .B(n21876), .ZN(
        P1_U3028) );
  OAI22_X1 U23661 ( .A1(n21879), .A2(n22010), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21878), .ZN(n21880) );
  AOI21_X1 U23662 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21881), .A(
        n21880), .ZN(n21883) );
  NAND2_X1 U23663 ( .A1(n21999), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n21882) );
  OAI211_X1 U23664 ( .C1(n22009), .C2(n21884), .A(n21883), .B(n21882), .ZN(
        P1_U3022) );
  INV_X1 U23665 ( .A(n21885), .ZN(n22111) );
  AOI22_X1 U23666 ( .A1(n21999), .A2(P1_REIP_REG_12__SCAN_IN), .B1(n21993), 
        .B2(n22111), .ZN(n21893) );
  AOI22_X1 U23667 ( .A1(n21887), .A2(n22004), .B1(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21886), .ZN(n21892) );
  NAND3_X1 U23668 ( .A1(n21890), .A2(n21889), .A3(n21888), .ZN(n21891) );
  NAND3_X1 U23669 ( .A1(n21893), .A2(n21892), .A3(n21891), .ZN(P1_U3019) );
  NAND2_X1 U23670 ( .A1(n21999), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n21894) );
  OAI221_X1 U23671 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21915), 
        .C1(n21901), .C2(n21907), .A(n21894), .ZN(n21895) );
  AOI21_X1 U23672 ( .B1(n21896), .B2(n22004), .A(n21895), .ZN(n21897) );
  OAI21_X1 U23673 ( .B1(n22009), .B2(n22134), .A(n21897), .ZN(P1_U3016) );
  OAI21_X1 U23674 ( .B1(n21899), .B2(n22010), .A(n21898), .ZN(n21900) );
  INV_X1 U23675 ( .A(n21900), .ZN(n21905) );
  NOR2_X1 U23676 ( .A1(n21901), .A2(n21915), .ZN(n21912) );
  OAI211_X1 U23677 ( .C1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n21912), .A(
        n21903), .B(n21902), .ZN(n21904) );
  OAI211_X1 U23678 ( .C1(n22009), .C2(n22163), .A(n21905), .B(n21904), .ZN(
        P1_U3014) );
  AOI22_X1 U23679 ( .A1(n21906), .A2(n22004), .B1(n21993), .B2(n22145), .ZN(
        n21914) );
  OAI21_X1 U23680 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21915), .A(
        n21907), .ZN(n21910) );
  NOR2_X1 U23681 ( .A1(n21975), .A2(n21908), .ZN(n21909) );
  AOI221_X1 U23682 ( .B1(n21912), .B2(n21911), .C1(n21910), .C2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n21909), .ZN(n21913) );
  NAND2_X1 U23683 ( .A1(n21914), .A2(n21913), .ZN(P1_U3015) );
  NOR2_X1 U23684 ( .A1(n21916), .A2(n21915), .ZN(n21945) );
  NAND2_X1 U23685 ( .A1(n21945), .A2(n21944), .ZN(n21929) );
  NAND2_X1 U23686 ( .A1(n21918), .A2(n21917), .ZN(n21919) );
  OAI211_X1 U23687 ( .C1(n21922), .C2(n21921), .A(n21920), .B(n21919), .ZN(
        n21939) );
  AOI22_X1 U23688 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21939), .B1(
        n21999), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n21928) );
  INV_X1 U23689 ( .A(n21923), .ZN(n21926) );
  INV_X1 U23690 ( .A(n21924), .ZN(n21925) );
  AOI22_X1 U23691 ( .A1(n21926), .A2(n22004), .B1(n21993), .B2(n21925), .ZN(
        n21927) );
  OAI211_X1 U23692 ( .C1(n21930), .C2(n21929), .A(n21928), .B(n21927), .ZN(
        P1_U3011) );
  AOI22_X1 U23693 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21939), .B1(
        n21999), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n21935) );
  INV_X1 U23694 ( .A(n21931), .ZN(n21933) );
  AOI22_X1 U23695 ( .A1(n21933), .A2(n22004), .B1(n21932), .B2(n21945), .ZN(
        n21934) );
  OAI211_X1 U23696 ( .C1(n22009), .C2(n21936), .A(n21935), .B(n21934), .ZN(
        P1_U3012) );
  AOI22_X1 U23697 ( .A1(n21938), .A2(n22004), .B1(n21993), .B2(n21937), .ZN(
        n21950) );
  NAND2_X1 U23698 ( .A1(n21999), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n21949) );
  INV_X1 U23699 ( .A(n21939), .ZN(n21942) );
  AOI21_X1 U23700 ( .B1(n21942), .B2(n21941), .A(n21940), .ZN(n21953) );
  INV_X1 U23701 ( .A(n21945), .ZN(n21943) );
  NOR3_X1 U23702 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21944), .A3(
        n21943), .ZN(n21951) );
  OAI21_X1 U23703 ( .B1(n21953), .B2(n21951), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21948) );
  NAND3_X1 U23704 ( .A1(n21946), .A2(n21945), .A3(n11778), .ZN(n21947) );
  NAND4_X1 U23705 ( .A1(n21950), .A2(n21949), .A3(n21948), .A4(n21947), .ZN(
        P1_U3009) );
  AOI21_X1 U23706 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n21999), .A(n21951), 
        .ZN(n21956) );
  INV_X1 U23707 ( .A(n21952), .ZN(n21954) );
  AOI22_X1 U23708 ( .A1(n21954), .A2(n22004), .B1(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n21953), .ZN(n21955) );
  OAI211_X1 U23709 ( .C1(n22009), .C2(n22186), .A(n21956), .B(n21955), .ZN(
        P1_U3010) );
  INV_X1 U23710 ( .A(n22207), .ZN(n21957) );
  AOI22_X1 U23711 ( .A1(n21958), .A2(n22004), .B1(n21993), .B2(n21957), .ZN(
        n21964) );
  NAND2_X1 U23712 ( .A1(n21999), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n21963) );
  OAI221_X1 U23713 ( .B1(n22000), .B2(n21959), .C1(n22000), .C2(n22003), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21962) );
  INV_X1 U23714 ( .A(n21970), .ZN(n22002) );
  NAND3_X1 U23715 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21960), .A3(
        n22002), .ZN(n21961) );
  NAND4_X1 U23716 ( .A1(n21964), .A2(n21963), .A3(n21962), .A4(n21961), .ZN(
        P1_U3007) );
  INV_X1 U23717 ( .A(n21965), .ZN(n21968) );
  INV_X1 U23718 ( .A(n21966), .ZN(n21967) );
  AOI22_X1 U23719 ( .A1(n21968), .A2(n22004), .B1(n21993), .B2(n21967), .ZN(
        n21974) );
  NOR3_X1 U23720 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21970), .A3(
        n21969), .ZN(n21989) );
  OAI22_X1 U23721 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21972), .B1(
        n21989), .B2(n21971), .ZN(n21973) );
  OAI211_X1 U23722 ( .C1(n21976), .C2(n21975), .A(n21974), .B(n21973), .ZN(
        P1_U3005) );
  INV_X1 U23723 ( .A(n21977), .ZN(n21983) );
  INV_X1 U23724 ( .A(n21978), .ZN(n21982) );
  NOR3_X1 U23725 ( .A1(n21980), .A2(n12927), .A3(n21979), .ZN(n21981) );
  AOI211_X1 U23726 ( .C1(n21983), .C2(n22004), .A(n21982), .B(n21981), .ZN(
        n21988) );
  INV_X1 U23727 ( .A(n21984), .ZN(n21985) );
  AOI22_X1 U23728 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n21986), .B1(
        n21993), .B2(n21985), .ZN(n21987) );
  NAND2_X1 U23729 ( .A1(n21988), .A2(n21987), .ZN(P1_U3003) );
  AOI21_X1 U23730 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n21999), .A(n21989), 
        .ZN(n21996) );
  INV_X1 U23731 ( .A(n21990), .ZN(n21994) );
  INV_X1 U23732 ( .A(n21991), .ZN(n21992) );
  AOI22_X1 U23733 ( .A1(n21994), .A2(n22004), .B1(n21993), .B2(n21992), .ZN(
        n21995) );
  OAI211_X1 U23734 ( .C1(n21998), .C2(n21997), .A(n21996), .B(n21995), .ZN(
        P1_U3006) );
  AOI22_X1 U23735 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n22000), .B1(
        n21999), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n22007) );
  INV_X1 U23736 ( .A(n22001), .ZN(n22005) );
  AOI22_X1 U23737 ( .A1(n22005), .A2(n22004), .B1(n22003), .B2(n22002), .ZN(
        n22006) );
  OAI211_X1 U23738 ( .C1(n22009), .C2(n22192), .A(n22007), .B(n22006), .ZN(
        P1_U3008) );
  OAI22_X1 U23739 ( .A1(n22011), .A2(n22010), .B1(n22009), .B2(n22008), .ZN(
        n22012) );
  INV_X1 U23740 ( .A(n22012), .ZN(n22018) );
  OAI22_X1 U23741 ( .A1(n22015), .A2(n22014), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n22013), .ZN(n22016) );
  NAND3_X1 U23742 ( .A1(n22018), .A2(n22017), .A3(n22016), .ZN(P1_U3031) );
  AOI21_X1 U23743 ( .B1(n22034), .B2(n22031), .A(n22030), .ZN(n22029) );
  AOI22_X1 U23744 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(n22166), .B1(n22165), .B2(
        n22019), .ZN(n22028) );
  INV_X1 U23745 ( .A(n22020), .ZN(n22021) );
  AOI22_X1 U23746 ( .A1(n22021), .A2(n22187), .B1(n22206), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n22023) );
  NAND3_X1 U23747 ( .A1(n22034), .A2(n22032), .A3(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n22022) );
  OAI211_X1 U23748 ( .C1(n22024), .C2(n22050), .A(n22023), .B(n22022), .ZN(
        n22025) );
  AOI21_X1 U23749 ( .B1(n22026), .B2(n22069), .A(n22025), .ZN(n22027) );
  OAI211_X1 U23750 ( .C1(n22029), .C2(n22032), .A(n22028), .B(n22027), .ZN(
        P1_U2838) );
  AOI221_X1 U23751 ( .B1(n22031), .B2(n22034), .C1(n22032), .C2(n22034), .A(
        n22030), .ZN(n22049) );
  INV_X1 U23752 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n22048) );
  NOR3_X1 U23753 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n22032), .A3(n22031), .ZN(
        n22033) );
  NAND2_X1 U23754 ( .A1(n22034), .A2(n22033), .ZN(n22035) );
  OAI21_X1 U23755 ( .B1(n22208), .B2(n22036), .A(n22035), .ZN(n22040) );
  OAI22_X1 U23756 ( .A1(n22201), .A2(n22038), .B1(n22037), .B2(n22152), .ZN(
        n22039) );
  AOI211_X1 U23757 ( .C1(n22042), .C2(n22041), .A(n22040), .B(n22039), .ZN(
        n22047) );
  INV_X1 U23758 ( .A(n22043), .ZN(n22044) );
  AOI22_X1 U23759 ( .A1(n22045), .A2(n22069), .B1(n22044), .B2(n22187), .ZN(
        n22046) );
  OAI211_X1 U23760 ( .C1(n22049), .C2(n22048), .A(n22047), .B(n22046), .ZN(
        P1_U2837) );
  OAI22_X1 U23761 ( .A1(n22208), .A2(n22052), .B1(n22051), .B2(n22050), .ZN(
        n22053) );
  AOI211_X1 U23762 ( .C1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n22206), .A(
        n22170), .B(n22053), .ZN(n22063) );
  NOR2_X1 U23763 ( .A1(n22189), .A2(n22054), .ZN(n22065) );
  NAND2_X1 U23764 ( .A1(n22056), .A2(n22055), .ZN(n22061) );
  OAI22_X1 U23765 ( .A1(n22059), .A2(n22058), .B1(n22057), .B2(n22203), .ZN(
        n22060) );
  AOI21_X1 U23766 ( .B1(n22065), .B2(n22061), .A(n22060), .ZN(n22062) );
  OAI211_X1 U23767 ( .C1(n22064), .C2(n22201), .A(n22063), .B(n22062), .ZN(
        P1_U2836) );
  AOI22_X1 U23768 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n22166), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n22065), .ZN(n22066) );
  OAI21_X1 U23769 ( .B1(n22208), .B2(n22067), .A(n22066), .ZN(n22068) );
  AOI211_X1 U23770 ( .C1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n22206), .A(
        n22170), .B(n22068), .ZN(n22074) );
  AOI22_X1 U23771 ( .A1(n22072), .A2(n22071), .B1(n22070), .B2(n22069), .ZN(
        n22073) );
  OAI211_X1 U23772 ( .C1(n22075), .C2(n22203), .A(n22074), .B(n22073), .ZN(
        P1_U2835) );
  INV_X1 U23773 ( .A(n22076), .ZN(n22085) );
  NAND2_X1 U23774 ( .A1(n22200), .A2(n22077), .ZN(n22089) );
  OAI22_X1 U23775 ( .A1(n22079), .A2(n22201), .B1(n22208), .B2(n22078), .ZN(
        n22080) );
  AOI211_X1 U23776 ( .C1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n22206), .A(
        n22170), .B(n22080), .ZN(n22081) );
  OAI221_X1 U23777 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n22083), .C1(n22082), 
        .C2(n22089), .A(n22081), .ZN(n22084) );
  AOI21_X1 U23778 ( .B1(n22085), .B2(n22172), .A(n22084), .ZN(n22086) );
  OAI21_X1 U23779 ( .B1(n22087), .B2(n22203), .A(n22086), .ZN(P1_U2834) );
  OAI22_X1 U23780 ( .A1(n22094), .A2(n22089), .B1(n22208), .B2(n22088), .ZN(
        n22090) );
  AOI211_X1 U23781 ( .C1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n22206), .A(
        n22170), .B(n22090), .ZN(n22097) );
  OAI22_X1 U23782 ( .A1(n22092), .A2(n22209), .B1(n22091), .B2(n22203), .ZN(
        n22093) );
  AOI21_X1 U23783 ( .B1(n22095), .B2(n22094), .A(n22093), .ZN(n22096) );
  OAI211_X1 U23784 ( .C1(n22098), .C2(n22201), .A(n22097), .B(n22096), .ZN(
        P1_U2833) );
  AOI22_X1 U23785 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n22166), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n22099), .ZN(n22100) );
  OAI21_X1 U23786 ( .B1(n22208), .B2(n22101), .A(n22100), .ZN(n22102) );
  AOI211_X1 U23787 ( .C1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n22206), .A(
        n22170), .B(n22102), .ZN(n22107) );
  OAI22_X1 U23788 ( .A1(n22104), .A2(n22209), .B1(n22103), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n22105) );
  INV_X1 U23789 ( .A(n22105), .ZN(n22106) );
  OAI211_X1 U23790 ( .C1(n22108), .C2(n22203), .A(n22107), .B(n22106), .ZN(
        P1_U2829) );
  AOI22_X1 U23791 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n22206), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(n22166), .ZN(n22109) );
  INV_X1 U23792 ( .A(n22109), .ZN(n22110) );
  AOI211_X1 U23793 ( .C1(n22165), .C2(n22111), .A(n22170), .B(n22110), .ZN(
        n22119) );
  AOI221_X1 U23794 ( .B1(n22114), .B2(n22113), .C1(n22112), .C2(n22113), .A(
        n22189), .ZN(n22116) );
  AOI22_X1 U23795 ( .A1(n22117), .A2(n22187), .B1(n22116), .B2(n22115), .ZN(
        n22118) );
  OAI211_X1 U23796 ( .C1(n22209), .C2(n22120), .A(n22119), .B(n22118), .ZN(
        P1_U2828) );
  NOR2_X1 U23797 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n22121), .ZN(n22130) );
  NAND2_X1 U23798 ( .A1(n22200), .A2(n22140), .ZN(n22138) );
  OAI22_X1 U23799 ( .A1(n22123), .A2(n22152), .B1(n22122), .B2(n22201), .ZN(
        n22124) );
  AOI211_X1 U23800 ( .C1(n22165), .C2(n22125), .A(n22170), .B(n22124), .ZN(
        n22129) );
  AOI22_X1 U23801 ( .A1(n22127), .A2(n22172), .B1(n22187), .B2(n22126), .ZN(
        n22128) );
  OAI211_X1 U23802 ( .C1(n22130), .C2(n22138), .A(n22129), .B(n22128), .ZN(
        P1_U2826) );
  AOI22_X1 U23803 ( .A1(n22131), .A2(n22187), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n22166), .ZN(n22133) );
  AOI21_X1 U23804 ( .B1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n22206), .A(
        n22170), .ZN(n22132) );
  OAI211_X1 U23805 ( .C1(n22208), .C2(n22134), .A(n22133), .B(n22132), .ZN(
        n22135) );
  AOI21_X1 U23806 ( .B1(n22136), .B2(n22172), .A(n22135), .ZN(n22137) );
  OAI221_X1 U23807 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n22140), .C1(n22139), 
        .C2(n22138), .A(n22137), .ZN(P1_U2825) );
  AOI21_X1 U23808 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n22200), .A(n22141), 
        .ZN(n22149) );
  OAI22_X1 U23809 ( .A1(n22143), .A2(n22203), .B1(n22142), .B2(n22201), .ZN(
        n22144) );
  AOI211_X1 U23810 ( .C1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n22206), .A(
        n22170), .B(n22144), .ZN(n22148) );
  AOI22_X1 U23811 ( .A1(n22146), .A2(n22172), .B1(n22165), .B2(n22145), .ZN(
        n22147) );
  OAI211_X1 U23812 ( .C1(n22150), .C2(n22149), .A(n22148), .B(n22147), .ZN(
        P1_U2824) );
  OAI22_X1 U23813 ( .A1(n22153), .A2(n22152), .B1(n22151), .B2(n22201), .ZN(
        n22154) );
  AOI211_X1 U23814 ( .C1(n22187), .C2(n22155), .A(n22170), .B(n22154), .ZN(
        n22162) );
  INV_X1 U23815 ( .A(n22156), .ZN(n22160) );
  NAND2_X1 U23816 ( .A1(n22158), .A2(n22157), .ZN(n22159) );
  AOI22_X1 U23817 ( .A1(n22160), .A2(n22172), .B1(n22171), .B2(n22159), .ZN(
        n22161) );
  OAI211_X1 U23818 ( .C1(n22208), .C2(n22163), .A(n22162), .B(n22161), .ZN(
        P1_U2823) );
  AOI22_X1 U23819 ( .A1(P1_EBX_REG_18__SCAN_IN), .A2(n22166), .B1(n22165), 
        .B2(n22164), .ZN(n22167) );
  OAI21_X1 U23820 ( .B1(n22168), .B2(n22203), .A(n22167), .ZN(n22169) );
  AOI211_X1 U23821 ( .C1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n22206), .A(
        n22170), .B(n22169), .ZN(n22175) );
  AOI22_X1 U23822 ( .A1(n22173), .A2(n22172), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n22171), .ZN(n22174) );
  OAI211_X1 U23823 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n22176), .A(n22175), 
        .B(n22174), .ZN(P1_U2822) );
  AOI22_X1 U23824 ( .A1(n22178), .A2(n22187), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n22177), .ZN(n22179) );
  OAI21_X1 U23825 ( .B1(n22180), .B2(n22201), .A(n22179), .ZN(n22184) );
  OAI22_X1 U23826 ( .A1(n22182), .A2(n22209), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n22181), .ZN(n22183) );
  AOI211_X1 U23827 ( .C1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n22206), .A(
        n22184), .B(n22183), .ZN(n22185) );
  OAI21_X1 U23828 ( .B1(n22208), .B2(n22186), .A(n22185), .ZN(P1_U2819) );
  AOI22_X1 U23829 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n22206), .B1(
        n22188), .B2(n22187), .ZN(n22197) );
  AOI211_X1 U23830 ( .C1(n22191), .C2(n22190), .A(n22199), .B(n22189), .ZN(
        n22195) );
  OAI22_X1 U23831 ( .A1(n22193), .A2(n22209), .B1(n22208), .B2(n22192), .ZN(
        n22194) );
  NOR2_X1 U23832 ( .A1(n22195), .A2(n22194), .ZN(n22196) );
  OAI211_X1 U23833 ( .C1(n22198), .C2(n22201), .A(n22197), .B(n22196), .ZN(
        P1_U2817) );
  AOI21_X1 U23834 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n22200), .A(n22199), 
        .ZN(n22214) );
  OAI22_X1 U23835 ( .A1(n22204), .A2(n22203), .B1(n22202), .B2(n22201), .ZN(
        n22205) );
  AOI21_X1 U23836 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n22206), .A(
        n22205), .ZN(n22213) );
  OAI22_X1 U23837 ( .A1(n22210), .A2(n22209), .B1(n22208), .B2(n22207), .ZN(
        n22211) );
  INV_X1 U23838 ( .A(n22211), .ZN(n22212) );
  OAI211_X1 U23839 ( .C1(n22215), .C2(n22214), .A(n22213), .B(n22212), .ZN(
        P1_U2816) );
  OAI21_X1 U23840 ( .B1(n22218), .B2(n22217), .A(n22216), .ZN(P1_U2806) );
  AOI21_X1 U23841 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n22226), .A(n21855), 
        .ZN(n22219) );
  INV_X1 U23842 ( .A(n22219), .ZN(n22221) );
  OAI211_X1 U23843 ( .C1(n22223), .C2(n22222), .A(n22221), .B(n22220), .ZN(
        P1_U3163) );
  OAI22_X1 U23844 ( .A1(n22226), .A2(n22464), .B1(n22225), .B2(n22224), .ZN(
        P1_U3466) );
  AOI21_X1 U23845 ( .B1(n22229), .B2(n22228), .A(n22227), .ZN(n22230) );
  OAI22_X1 U23846 ( .A1(n22232), .A2(n22231), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n22230), .ZN(n22233) );
  OAI21_X1 U23847 ( .B1(n22235), .B2(n22234), .A(n22233), .ZN(P1_U3161) );
  AOI21_X1 U23848 ( .B1(n17710), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n22237), 
        .ZN(n22236) );
  INV_X1 U23849 ( .A(n22236), .ZN(P1_U2805) );
  AOI21_X1 U23850 ( .B1(n17710), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n22237), 
        .ZN(n22238) );
  INV_X1 U23851 ( .A(n22238), .ZN(P1_U3465) );
  OAI21_X1 U23852 ( .B1(n22242), .B2(n22239), .A(n22240), .ZN(P2_U2818) );
  OAI21_X1 U23853 ( .B1(n22242), .B2(n22241), .A(n22240), .ZN(P2_U3592) );
  OAI21_X1 U23854 ( .B1(n22246), .B2(n22243), .A(n22244), .ZN(P3_U2636) );
  INV_X1 U23855 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22245) );
  OAI21_X1 U23856 ( .B1(n22246), .B2(n22245), .A(n22244), .ZN(P3_U3281) );
  INV_X1 U23857 ( .A(HOLD), .ZN(n22299) );
  OAI21_X1 U23858 ( .B1(n22299), .B2(n22247), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22248) );
  INV_X1 U23859 ( .A(n22248), .ZN(n22251) );
  AOI21_X1 U23860 ( .B1(n22290), .B2(P3_STATE_REG_1__SCAN_IN), .A(n22249), 
        .ZN(n22307) );
  AOI21_X1 U23861 ( .B1(n22250), .B2(NA), .A(n22300), .ZN(n22305) );
  OAI22_X1 U23862 ( .A1(n22252), .A2(n22251), .B1(n22307), .B2(n22305), .ZN(
        P3_U3029) );
  AOI221_X1 U23863 ( .B1(NA), .B2(P1_STATE_REG_1__SCAN_IN), .C1(n22253), .C2(
        P1_STATE_REG_1__SCAN_IN), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n22257) );
  NAND2_X1 U23864 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n22254), .ZN(n22264) );
  NOR3_X1 U23865 ( .A1(NA), .A2(n22255), .A3(n22264), .ZN(n22256) );
  AOI221_X1 U23866 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n22257), 
        .C2(HOLD), .A(n22256), .ZN(n22260) );
  NAND2_X1 U23867 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n22264), .ZN(n22267) );
  OAI211_X1 U23868 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n22302), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n22267), .ZN(n22258) );
  OAI21_X1 U23869 ( .B1(n22260), .B2(n22259), .A(n22258), .ZN(P1_U3196) );
  NAND2_X1 U23870 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22268) );
  INV_X1 U23871 ( .A(n22268), .ZN(n22263) );
  NAND2_X1 U23872 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n22262) );
  AOI21_X1 U23873 ( .B1(n22263), .B2(n22262), .A(n22261), .ZN(n22265) );
  OAI211_X1 U23874 ( .C1(n22299), .C2(n22266), .A(n22265), .B(n22264), .ZN(
        P1_U3195) );
  INV_X1 U23875 ( .A(n22267), .ZN(n22272) );
  NAND2_X1 U23876 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(n22302), .ZN(
        n22269) );
  AOI22_X1 U23877 ( .A1(HOLD), .A2(n22270), .B1(n22269), .B2(n22268), .ZN(
        n22271) );
  OAI22_X1 U23878 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22272), .B1(n22805), 
        .B2(n22271), .ZN(P1_U3194) );
  OAI22_X1 U23879 ( .A1(n22299), .A2(n22273), .B1(n22302), .B2(
        P2_STATE_REG_0__SCAN_IN), .ZN(n22277) );
  NAND2_X1 U23880 ( .A1(n22274), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n22285) );
  NAND2_X1 U23881 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n22285), .ZN(n22284) );
  INV_X1 U23882 ( .A(n22284), .ZN(n22275) );
  OAI21_X1 U23883 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n22275), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22276) );
  AOI22_X1 U23884 ( .A1(n22278), .A2(n22277), .B1(n17900), .B2(n22276), .ZN(
        n22279) );
  INV_X1 U23885 ( .A(n22279), .ZN(P2_U3209) );
  NAND2_X1 U23886 ( .A1(n22280), .A2(HOLD), .ZN(n22282) );
  OAI211_X1 U23887 ( .C1(n22289), .C2(n22299), .A(P2_STATE_REG_0__SCAN_IN), 
        .B(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22281) );
  NAND4_X1 U23888 ( .A1(n22283), .A2(n22282), .A3(n22285), .A4(n22281), .ZN(
        P2_U3210) );
  OAI22_X1 U23889 ( .A1(HOLD), .A2(n22284), .B1(P2_STATE_REG_0__SCAN_IN), .B2(
        n22302), .ZN(n22288) );
  OAI22_X1 U23890 ( .A1(NA), .A2(n22285), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22286) );
  OAI211_X1 U23891 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n22286), .ZN(n22287) );
  OAI211_X1 U23892 ( .C1(n22289), .C2(n22288), .A(n17900), .B(n22287), .ZN(
        P2_U3211) );
  NOR2_X1 U23893 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22309)
         );
  OAI21_X1 U23894 ( .B1(n22299), .B2(n22300), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n22291) );
  NAND2_X1 U23895 ( .A1(n22290), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n22301) );
  OAI21_X1 U23896 ( .B1(n22309), .B2(n22291), .A(n22301), .ZN(n22294) );
  OAI211_X1 U23897 ( .C1(n22299), .C2(n22300), .A(P3_STATE_REG_0__SCAN_IN), 
        .B(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22292) );
  AOI21_X1 U23898 ( .B1(n22292), .B2(n22295), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n22293) );
  AOI21_X1 U23899 ( .B1(n22295), .B2(n22294), .A(n22293), .ZN(n22296) );
  OAI221_X1 U23900 ( .B1(n22298), .B2(P3_STATE_REG_2__SCAN_IN), .C1(n22298), 
        .C2(n22297), .A(n22296), .ZN(P3_U3030) );
  OAI22_X1 U23901 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n22300), .B2(n22299), .ZN(n22304)
         );
  INV_X1 U23902 ( .A(n22301), .ZN(n22303) );
  OAI221_X1 U23903 ( .B1(n22304), .B2(n22303), .C1(n22304), .C2(n22302), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n22308) );
  INV_X1 U23904 ( .A(n22305), .ZN(n22306) );
  OAI22_X1 U23905 ( .A1(n22309), .A2(n22308), .B1(n22307), .B2(n22306), .ZN(
        P3_U3031) );
  NOR2_X1 U23906 ( .A1(n22399), .A2(n22410), .ZN(n22312) );
  AOI21_X1 U23907 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n22400), .A(n22312), 
        .ZN(n22310) );
  OAI21_X1 U23908 ( .B1(n22311), .B2(n22405), .A(n22310), .ZN(P1_U2937) );
  AOI21_X1 U23909 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(n22400), .A(n22312), 
        .ZN(n22313) );
  OAI21_X1 U23910 ( .B1(n22314), .B2(n22405), .A(n22313), .ZN(P1_U2952) );
  INV_X1 U23911 ( .A(n22315), .ZN(n22316) );
  NOR2_X1 U23912 ( .A1(n22399), .A2(n22316), .ZN(n22319) );
  AOI21_X1 U23913 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n22400), .A(n22319), 
        .ZN(n22317) );
  OAI21_X1 U23914 ( .B1(n22318), .B2(n22405), .A(n22317), .ZN(P1_U2938) );
  AOI21_X1 U23915 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n22400), .A(n22319), 
        .ZN(n22320) );
  OAI21_X1 U23916 ( .B1(n22321), .B2(n22405), .A(n22320), .ZN(P1_U2953) );
  INV_X1 U23917 ( .A(n22555), .ZN(n22322) );
  NOR2_X1 U23918 ( .A1(n22399), .A2(n22322), .ZN(n22325) );
  AOI21_X1 U23919 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n22400), .A(n22325), 
        .ZN(n22323) );
  OAI21_X1 U23920 ( .B1(n22324), .B2(n22405), .A(n22323), .ZN(P1_U2939) );
  AOI21_X1 U23921 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n22400), .A(n22325), 
        .ZN(n22326) );
  OAI21_X1 U23922 ( .B1(n22327), .B2(n22405), .A(n22326), .ZN(P1_U2954) );
  NOR2_X1 U23923 ( .A1(n22399), .A2(n22328), .ZN(n22331) );
  AOI21_X1 U23924 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n22400), .A(n22331), 
        .ZN(n22329) );
  OAI21_X1 U23925 ( .B1(n22330), .B2(n22405), .A(n22329), .ZN(P1_U2940) );
  AOI21_X1 U23926 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n22400), .A(n22331), 
        .ZN(n22332) );
  OAI21_X1 U23927 ( .B1(n22333), .B2(n22405), .A(n22332), .ZN(P1_U2955) );
  NOR2_X1 U23928 ( .A1(n22399), .A2(n22334), .ZN(n22338) );
  AOI21_X1 U23929 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n22400), .A(n22338), 
        .ZN(n22335) );
  OAI21_X1 U23930 ( .B1(n22336), .B2(n22405), .A(n22335), .ZN(P1_U2941) );
  AOI21_X1 U23931 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n22387), .A(n22338), 
        .ZN(n22339) );
  OAI21_X1 U23932 ( .B1(n22340), .B2(n22405), .A(n22339), .ZN(P1_U2956) );
  NOR2_X1 U23933 ( .A1(n22399), .A2(n22341), .ZN(n22344) );
  AOI21_X1 U23934 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n22387), .A(n22344), 
        .ZN(n22342) );
  OAI21_X1 U23935 ( .B1(n22343), .B2(n22405), .A(n22342), .ZN(P1_U2942) );
  AOI21_X1 U23936 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n22387), .A(n22344), 
        .ZN(n22345) );
  OAI21_X1 U23937 ( .B1(n12160), .B2(n22405), .A(n22345), .ZN(P1_U2957) );
  NOR2_X1 U23938 ( .A1(n22399), .A2(n22346), .ZN(n22349) );
  AOI21_X1 U23939 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n22387), .A(n22349), 
        .ZN(n22347) );
  OAI21_X1 U23940 ( .B1(n22348), .B2(n22405), .A(n22347), .ZN(P1_U2943) );
  AOI21_X1 U23941 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n22400), .A(n22349), 
        .ZN(n22350) );
  OAI21_X1 U23942 ( .B1(n22351), .B2(n22405), .A(n22350), .ZN(P1_U2958) );
  NOR2_X1 U23943 ( .A1(n22399), .A2(n22352), .ZN(n22355) );
  AOI21_X1 U23944 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n22400), .A(n22355), 
        .ZN(n22353) );
  OAI21_X1 U23945 ( .B1(n22354), .B2(n22405), .A(n22353), .ZN(P1_U2944) );
  AOI21_X1 U23946 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n22400), .A(n22355), 
        .ZN(n22356) );
  OAI21_X1 U23947 ( .B1(n12149), .B2(n22405), .A(n22356), .ZN(P1_U2959) );
  NOR2_X1 U23948 ( .A1(n22399), .A2(n22357), .ZN(n22359) );
  AOI21_X1 U23949 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n22400), .A(n22359), 
        .ZN(n22358) );
  OAI21_X1 U23950 ( .B1(n16619), .B2(n22405), .A(n22358), .ZN(P1_U2945) );
  AOI21_X1 U23951 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n22400), .A(n22359), 
        .ZN(n22360) );
  OAI21_X1 U23952 ( .B1(n22361), .B2(n22405), .A(n22360), .ZN(P1_U2960) );
  NOR2_X1 U23953 ( .A1(n22399), .A2(n22362), .ZN(n22365) );
  AOI21_X1 U23954 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n22400), .A(n22365), 
        .ZN(n22363) );
  OAI21_X1 U23955 ( .B1(n22364), .B2(n22405), .A(n22363), .ZN(P1_U2946) );
  AOI21_X1 U23956 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n22400), .A(n22365), 
        .ZN(n22366) );
  OAI21_X1 U23957 ( .B1(n22367), .B2(n22405), .A(n22366), .ZN(P1_U2961) );
  INV_X1 U23958 ( .A(n22368), .ZN(n22369) );
  NOR2_X1 U23959 ( .A1(n22399), .A2(n22369), .ZN(n22372) );
  AOI21_X1 U23960 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n22387), .A(n22372), 
        .ZN(n22370) );
  OAI21_X1 U23961 ( .B1(n22371), .B2(n22405), .A(n22370), .ZN(P1_U2947) );
  AOI21_X1 U23962 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n22387), .A(n22372), 
        .ZN(n22373) );
  OAI21_X1 U23963 ( .B1(n22374), .B2(n22405), .A(n22373), .ZN(P1_U2962) );
  INV_X1 U23964 ( .A(n22375), .ZN(n22376) );
  NOR2_X1 U23965 ( .A1(n22399), .A2(n22376), .ZN(n22379) );
  AOI21_X1 U23966 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n22387), .A(n22379), 
        .ZN(n22377) );
  OAI21_X1 U23967 ( .B1(n22378), .B2(n22405), .A(n22377), .ZN(P1_U2948) );
  AOI21_X1 U23968 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n22387), .A(n22379), 
        .ZN(n22380) );
  OAI21_X1 U23969 ( .B1(n22381), .B2(n22405), .A(n22380), .ZN(P1_U2963) );
  INV_X1 U23970 ( .A(n22382), .ZN(n22383) );
  NOR2_X1 U23971 ( .A1(n22399), .A2(n22383), .ZN(n22386) );
  AOI21_X1 U23972 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n22387), .A(n22386), 
        .ZN(n22384) );
  OAI21_X1 U23973 ( .B1(n22385), .B2(n22405), .A(n22384), .ZN(P1_U2949) );
  AOI21_X1 U23974 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n22387), .A(n22386), 
        .ZN(n22388) );
  OAI21_X1 U23975 ( .B1(n22389), .B2(n22405), .A(n22388), .ZN(P1_U2964) );
  INV_X1 U23976 ( .A(n22390), .ZN(n22391) );
  NOR2_X1 U23977 ( .A1(n22399), .A2(n22391), .ZN(n22394) );
  AOI21_X1 U23978 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n22400), .A(n22394), 
        .ZN(n22392) );
  OAI21_X1 U23979 ( .B1(n22393), .B2(n22405), .A(n22392), .ZN(P1_U2950) );
  AOI21_X1 U23980 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n22400), .A(n22394), 
        .ZN(n22395) );
  OAI21_X1 U23981 ( .B1(n22396), .B2(n22405), .A(n22395), .ZN(P1_U2965) );
  INV_X1 U23982 ( .A(n22397), .ZN(n22398) );
  NOR2_X1 U23983 ( .A1(n22399), .A2(n22398), .ZN(n22403) );
  AOI21_X1 U23984 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n22400), .A(n22403), 
        .ZN(n22401) );
  OAI21_X1 U23985 ( .B1(n22402), .B2(n22405), .A(n22401), .ZN(P1_U2951) );
  AOI21_X1 U23986 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n22400), .A(n22403), 
        .ZN(n22404) );
  OAI21_X1 U23987 ( .B1(n22406), .B2(n22405), .A(n22404), .ZN(P1_U2966) );
  NOR3_X1 U23988 ( .A1(n22737), .A2(n22800), .A3(n22497), .ZN(n22407) );
  NOR2_X1 U23989 ( .A1(n22497), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22498) );
  NOR2_X1 U23990 ( .A1(n22407), .A2(n22498), .ZN(n22420) );
  INV_X1 U23991 ( .A(n22420), .ZN(n22409) );
  NOR2_X1 U23992 ( .A1(n22431), .A2(n22500), .ZN(n22419) );
  INV_X1 U23993 ( .A(n22417), .ZN(n22408) );
  INV_X1 U23994 ( .A(n22522), .ZN(n22514) );
  NOR2_X2 U23995 ( .A1(n22629), .A2(n22414), .ZN(n22521) );
  NOR2_X1 U23996 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22415), .ZN(
        n22736) );
  AOI22_X1 U23997 ( .A1(n22800), .A2(n22517), .B1(n22521), .B2(n22736), .ZN(
        n22424) );
  INV_X1 U23998 ( .A(n22736), .ZN(n22416) );
  AOI22_X1 U23999 ( .A1(n22417), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n22416), .ZN(n22418) );
  OAI211_X1 U24000 ( .C1(n22420), .C2(n22419), .A(n22490), .B(n22418), .ZN(
        n22738) );
  AOI22_X1 U24001 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22738), .B1(
        n22737), .B2(n22523), .ZN(n22423) );
  OAI211_X1 U24002 ( .C1(n22741), .C2(n22514), .A(n22424), .B(n22423), .ZN(
        P1_U3033) );
  INV_X1 U24003 ( .A(n22523), .ZN(n22520) );
  AOI22_X1 U24004 ( .A1(n22522), .A2(n22689), .B1(n22521), .B2(n22688), .ZN(
        n22426) );
  AOI22_X1 U24005 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22690), .B1(
        n22737), .B2(n22517), .ZN(n22425) );
  OAI211_X1 U24006 ( .C1(n22520), .C2(n22693), .A(n22426), .B(n22425), .ZN(
        P1_U3041) );
  NOR3_X1 U24007 ( .A1(n22749), .A2(n22743), .A3(n22497), .ZN(n22429) );
  NOR2_X1 U24008 ( .A1(n22429), .A2(n22498), .ZN(n22437) );
  INV_X1 U24009 ( .A(n22437), .ZN(n22433) );
  NOR2_X1 U24010 ( .A1(n22431), .A2(n22430), .ZN(n22436) );
  NOR2_X1 U24011 ( .A1(n22432), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22461) );
  AOI22_X1 U24012 ( .A1(n22433), .A2(n22436), .B1(n22481), .B2(n22461), .ZN(
        n22747) );
  NAND3_X1 U24013 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n12668), .A3(
        n12665), .ZN(n22449) );
  NOR2_X1 U24014 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22449), .ZN(
        n22742) );
  AOI22_X1 U24015 ( .A1(n22743), .A2(n22517), .B1(n22521), .B2(n22742), .ZN(
        n22439) );
  INV_X1 U24016 ( .A(n22742), .ZN(n22434) );
  NOR2_X1 U24017 ( .A1(n22461), .A2(n21855), .ZN(n22465) );
  AOI21_X1 U24018 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22434), .A(n22465), 
        .ZN(n22435) );
  OAI211_X1 U24019 ( .C1(n22437), .C2(n22436), .A(n22490), .B(n22435), .ZN(
        n22744) );
  AOI22_X1 U24020 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22744), .B1(
        n22749), .B2(n22523), .ZN(n22438) );
  OAI211_X1 U24021 ( .C1(n22747), .C2(n22514), .A(n22439), .B(n22438), .ZN(
        P1_U3049) );
  OAI21_X1 U24022 ( .B1(n22442), .B2(n22441), .A(n22440), .ZN(n22452) );
  NOR2_X1 U24023 ( .A1(n22485), .A2(n22449), .ZN(n22748) );
  AOI21_X1 U24024 ( .B1(n22444), .B2(n22443), .A(n22748), .ZN(n22446) );
  OAI22_X1 U24025 ( .A1(n21855), .A2(n22449), .B1(n22452), .B2(n22446), .ZN(
        n22445) );
  AOI22_X1 U24026 ( .A1(n22749), .A2(n22517), .B1(n22521), .B2(n22748), .ZN(
        n22454) );
  INV_X1 U24027 ( .A(n22446), .ZN(n22451) );
  INV_X1 U24028 ( .A(n22447), .ZN(n22448) );
  AOI21_X1 U24029 ( .B1(n22497), .B2(n22449), .A(n22448), .ZN(n22450) );
  OAI21_X1 U24030 ( .B1(n22452), .B2(n22451), .A(n22450), .ZN(n22751) );
  AOI22_X1 U24031 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22751), .B1(
        n22750), .B2(n22523), .ZN(n22453) );
  OAI211_X1 U24032 ( .C1(n22754), .C2(n22514), .A(n22454), .B(n22453), .ZN(
        P1_U3057) );
  AOI22_X1 U24033 ( .A1(n22522), .A2(n22699), .B1(n22521), .B2(n22698), .ZN(
        n22456) );
  AOI22_X1 U24034 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n22700), .B1(
        n22750), .B2(n22517), .ZN(n22455) );
  OAI211_X1 U24035 ( .C1(n22520), .C2(n22760), .A(n22456), .B(n22455), .ZN(
        P1_U3065) );
  INV_X1 U24036 ( .A(n22517), .ZN(n22526) );
  AOI22_X1 U24037 ( .A1(n22522), .A2(n22756), .B1(n22521), .B2(n22755), .ZN(
        n22458) );
  AOI22_X1 U24038 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n22757), .B1(
        n22762), .B2(n22523), .ZN(n22457) );
  OAI211_X1 U24039 ( .C1(n22526), .C2(n22760), .A(n22458), .B(n22457), .ZN(
        P1_U3073) );
  NOR3_X1 U24040 ( .A1(n22762), .A2(n22761), .A3(n22497), .ZN(n22459) );
  NOR2_X1 U24041 ( .A1(n22459), .A2(n22498), .ZN(n22468) );
  INV_X1 U24042 ( .A(n22468), .ZN(n22462) );
  AND2_X1 U24043 ( .A1(n22460), .A2(n22500), .ZN(n22467) );
  AOI22_X1 U24044 ( .A1(n22462), .A2(n22467), .B1(n22503), .B2(n22461), .ZN(
        n22766) );
  AOI22_X1 U24045 ( .A1(n22762), .A2(n22517), .B1(n22521), .B2(n11343), .ZN(
        n22470) );
  AOI21_X1 U24046 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n11221), .A(n22465), 
        .ZN(n22466) );
  OAI211_X1 U24047 ( .C1(n22468), .C2(n22467), .A(n22509), .B(n22466), .ZN(
        n22763) );
  AOI22_X1 U24048 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n22763), .B1(
        n22761), .B2(n22523), .ZN(n22469) );
  OAI211_X1 U24049 ( .C1(n22766), .C2(n22514), .A(n22470), .B(n22469), .ZN(
        P1_U3081) );
  AOI22_X1 U24050 ( .A1(n22522), .A2(n22706), .B1(n22705), .B2(n22521), .ZN(
        n22472) );
  AOI22_X1 U24051 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n22707), .B1(
        n22761), .B2(n22517), .ZN(n22471) );
  OAI211_X1 U24052 ( .C1(n22520), .C2(n22710), .A(n22472), .B(n22471), .ZN(
        P1_U3089) );
  INV_X1 U24053 ( .A(n22473), .ZN(n22712) );
  AOI22_X1 U24054 ( .A1(n22522), .A2(n22712), .B1(n22521), .B2(n22711), .ZN(
        n22475) );
  AOI22_X1 U24055 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n22714), .B1(
        n22713), .B2(n22517), .ZN(n22474) );
  OAI211_X1 U24056 ( .C1(n22520), .C2(n22772), .A(n22475), .B(n22474), .ZN(
        P1_U3097) );
  AOI22_X1 U24057 ( .A1(n22522), .A2(n22768), .B1(n22521), .B2(n22767), .ZN(
        n22477) );
  AOI22_X1 U24058 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22769), .B1(
        n22774), .B2(n22523), .ZN(n22476) );
  OAI211_X1 U24059 ( .C1(n22526), .C2(n22772), .A(n22477), .B(n22476), .ZN(
        P1_U3105) );
  NOR3_X1 U24060 ( .A1(n22774), .A2(n22775), .A3(n22497), .ZN(n22478) );
  NOR2_X1 U24061 ( .A1(n22478), .A2(n22498), .ZN(n22492) );
  INV_X1 U24062 ( .A(n22492), .ZN(n22483) );
  AND2_X1 U24063 ( .A1(n22479), .A2(n22500), .ZN(n22491) );
  INV_X1 U24064 ( .A(n22480), .ZN(n22482) );
  NAND2_X1 U24065 ( .A1(n22485), .A2(n22484), .ZN(n22488) );
  INV_X1 U24066 ( .A(n22488), .ZN(n22773) );
  AOI22_X1 U24067 ( .A1(n22775), .A2(n22523), .B1(n22521), .B2(n22773), .ZN(
        n22494) );
  INV_X1 U24068 ( .A(n22486), .ZN(n22487) );
  AOI21_X1 U24069 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22488), .A(n22487), 
        .ZN(n22489) );
  OAI211_X1 U24070 ( .C1(n22492), .C2(n22491), .A(n22490), .B(n22489), .ZN(
        n22776) );
  AOI22_X1 U24071 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22776), .B1(
        n22774), .B2(n22517), .ZN(n22493) );
  OAI211_X1 U24072 ( .C1(n22779), .C2(n22514), .A(n22494), .B(n22493), .ZN(
        P1_U3113) );
  INV_X1 U24073 ( .A(n22783), .ZN(n22724) );
  AOI22_X1 U24074 ( .A1(n22522), .A2(n22720), .B1(n22521), .B2(n22719), .ZN(
        n22496) );
  AOI22_X1 U24075 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n22721), .B1(
        n22775), .B2(n22517), .ZN(n22495) );
  OAI211_X1 U24076 ( .C1(n22520), .C2(n22724), .A(n22496), .B(n22495), .ZN(
        P1_U3121) );
  NOR3_X1 U24077 ( .A1(n22783), .A2(n22781), .A3(n22497), .ZN(n22499) );
  NOR2_X1 U24078 ( .A1(n22499), .A2(n22498), .ZN(n22511) );
  INV_X1 U24079 ( .A(n22511), .ZN(n22504) );
  NOR2_X1 U24080 ( .A1(n22501), .A2(n22500), .ZN(n22510) );
  AOI22_X1 U24081 ( .A1(n22504), .A2(n22510), .B1(n22503), .B2(n22502), .ZN(
        n22788) );
  NOR2_X1 U24082 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22505), .ZN(
        n22780) );
  AOI22_X1 U24083 ( .A1(n22781), .A2(n22523), .B1(n22521), .B2(n22780), .ZN(
        n22513) );
  INV_X1 U24084 ( .A(n22780), .ZN(n22506) );
  AOI22_X1 U24085 ( .A1(n22507), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n22506), .ZN(n22508) );
  OAI211_X1 U24086 ( .C1(n22511), .C2(n22510), .A(n22509), .B(n22508), .ZN(
        n22784) );
  AOI22_X1 U24087 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n22784), .B1(
        n22783), .B2(n22517), .ZN(n22512) );
  OAI211_X1 U24088 ( .C1(n22788), .C2(n22514), .A(n22513), .B(n22512), .ZN(
        P1_U3129) );
  AOI22_X1 U24089 ( .A1(n22522), .A2(n22790), .B1(n22521), .B2(n22789), .ZN(
        n22516) );
  AOI22_X1 U24090 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22792), .B1(
        n22791), .B2(n22523), .ZN(n22515) );
  OAI211_X1 U24091 ( .C1(n22526), .C2(n22795), .A(n22516), .B(n22515), .ZN(
        P1_U3137) );
  AOI22_X1 U24092 ( .A1(n22522), .A2(n22731), .B1(n22521), .B2(n22729), .ZN(
        n22519) );
  AOI22_X1 U24093 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22733), .B1(
        n22791), .B2(n22517), .ZN(n22518) );
  OAI211_X1 U24094 ( .C1(n22520), .C2(n22804), .A(n22519), .B(n22518), .ZN(
        P1_U3145) );
  AOI22_X1 U24095 ( .A1(n22522), .A2(n22798), .B1(n22796), .B2(n22521), .ZN(
        n22525) );
  AOI22_X1 U24096 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n22801), .B1(
        n22800), .B2(n22523), .ZN(n22524) );
  OAI211_X1 U24097 ( .C1(n22526), .C2(n22804), .A(n22525), .B(n22524), .ZN(
        P1_U3153) );
  AOI22_X1 U24098 ( .A1(n22800), .A2(n15390), .B1(n22551), .B2(n22736), .ZN(
        n22528) );
  AOI22_X1 U24099 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22738), .B1(
        n22737), .B2(n11342), .ZN(n22527) );
  OAI211_X1 U24100 ( .C1(n22741), .C2(n22550), .A(n22528), .B(n22527), .ZN(
        P1_U3034) );
  AOI22_X1 U24101 ( .A1(n22552), .A2(n22689), .B1(n22551), .B2(n22688), .ZN(
        n22530) );
  AOI22_X1 U24102 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n22737), .B2(n15390), .ZN(n22529) );
  OAI211_X1 U24103 ( .C1(n11341), .C2(n22693), .A(n22530), .B(n22529), .ZN(
        P1_U3042) );
  AOI22_X1 U24104 ( .A1(n22749), .A2(n11342), .B1(n22551), .B2(n22742), .ZN(
        n22532) );
  AOI22_X1 U24105 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n22743), .B2(n15390), .ZN(n22531) );
  OAI211_X1 U24106 ( .C1(n22747), .C2(n22550), .A(n22532), .B(n22531), .ZN(
        P1_U3050) );
  AOI22_X1 U24107 ( .A1(n22750), .A2(n11342), .B1(n22551), .B2(n22748), .ZN(
        n22534) );
  AOI22_X1 U24108 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n22749), .B2(n15390), .ZN(n22533) );
  OAI211_X1 U24109 ( .C1(n22754), .C2(n22550), .A(n22534), .B(n22533), .ZN(
        P1_U3058) );
  AOI22_X1 U24110 ( .A1(n22552), .A2(n22699), .B1(n22551), .B2(n22698), .ZN(
        n22536) );
  AOI22_X1 U24111 ( .A1(n22700), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n22750), .B2(n15390), .ZN(n22535) );
  OAI211_X1 U24112 ( .C1(n11341), .C2(n22760), .A(n22536), .B(n22535), .ZN(
        P1_U3066) );
  AOI22_X1 U24113 ( .A1(n22762), .A2(n15390), .B1(n11343), .B2(n22551), .ZN(
        n22538) );
  AOI22_X1 U24114 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n22763), .B1(
        n22761), .B2(n11342), .ZN(n22537) );
  OAI211_X1 U24115 ( .C1(n22766), .C2(n22550), .A(n22538), .B(n22537), .ZN(
        P1_U3082) );
  AOI22_X1 U24116 ( .A1(n22552), .A2(n22706), .B1(n22551), .B2(n22705), .ZN(
        n22540) );
  AOI22_X1 U24117 ( .A1(n22707), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n22761), .B2(n15390), .ZN(n22539) );
  OAI211_X1 U24118 ( .C1(n11341), .C2(n22710), .A(n22540), .B(n22539), .ZN(
        P1_U3090) );
  AOI22_X1 U24119 ( .A1(n22712), .A2(n22552), .B1(n22551), .B2(n22711), .ZN(
        n22542) );
  AOI22_X1 U24120 ( .A1(n22714), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n22713), .B2(n15390), .ZN(n22541) );
  OAI211_X1 U24121 ( .C1(n11341), .C2(n22772), .A(n22542), .B(n22541), .ZN(
        P1_U3098) );
  AOI22_X1 U24122 ( .A1(n22775), .A2(n11342), .B1(n22551), .B2(n22773), .ZN(
        n22544) );
  AOI22_X1 U24123 ( .A1(n22776), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n22774), .B2(n15390), .ZN(n22543) );
  OAI211_X1 U24124 ( .C1(n22779), .C2(n22550), .A(n22544), .B(n22543), .ZN(
        P1_U3114) );
  AOI22_X1 U24125 ( .A1(n22552), .A2(n22720), .B1(n22551), .B2(n22719), .ZN(
        n22546) );
  AOI22_X1 U24126 ( .A1(n22721), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n22775), .B2(n15390), .ZN(n22545) );
  OAI211_X1 U24127 ( .C1(n11341), .C2(n22724), .A(n22546), .B(n22545), .ZN(
        P1_U3122) );
  AOI22_X1 U24128 ( .A1(n22781), .A2(n11342), .B1(n22551), .B2(n22780), .ZN(
        n22549) );
  AOI22_X1 U24129 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n22783), .B2(n15390), .ZN(n22548) );
  OAI211_X1 U24130 ( .C1(n22788), .C2(n22550), .A(n22549), .B(n22548), .ZN(
        P1_U3130) );
  AOI22_X1 U24131 ( .A1(n22552), .A2(n22731), .B1(n22551), .B2(n22729), .ZN(
        n22554) );
  AOI22_X1 U24132 ( .A1(n22733), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n22791), .B2(n15390), .ZN(n22553) );
  OAI211_X1 U24133 ( .C1(n11341), .C2(n22804), .A(n22554), .B(n22553), .ZN(
        P1_U3146) );
  NAND2_X1 U24134 ( .A1(n22626), .A2(n22555), .ZN(n22585) );
  INV_X1 U24135 ( .A(DATAI_26_), .ZN(n22556) );
  OAI22_X1 U24136 ( .A1(n22556), .A2(n22632), .B1(n17075), .B2(n22630), .ZN(
        n22588) );
  NOR2_X2 U24137 ( .A1(n22629), .A2(n14540), .ZN(n22592) );
  AOI22_X1 U24138 ( .A1(n22800), .A2(n11347), .B1(n22592), .B2(n22736), .ZN(
        n22560) );
  AOI22_X1 U24139 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22738), .B1(
        n22737), .B2(n22594), .ZN(n22559) );
  OAI211_X1 U24140 ( .C1(n22741), .C2(n22585), .A(n22560), .B(n22559), .ZN(
        P1_U3035) );
  INV_X1 U24141 ( .A(n22594), .ZN(n22591) );
  AOI22_X1 U24142 ( .A1(n22593), .A2(n22689), .B1(n22592), .B2(n22688), .ZN(
        n22562) );
  AOI22_X1 U24143 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22690), .B1(
        n22737), .B2(n11347), .ZN(n22561) );
  OAI211_X1 U24144 ( .C1(n22591), .C2(n22693), .A(n22562), .B(n22561), .ZN(
        P1_U3043) );
  AOI22_X1 U24145 ( .A1(n22749), .A2(n22594), .B1(n22592), .B2(n22742), .ZN(
        n22564) );
  AOI22_X1 U24146 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22744), .B1(
        n22743), .B2(n11347), .ZN(n22563) );
  OAI211_X1 U24147 ( .C1(n22747), .C2(n22585), .A(n22564), .B(n22563), .ZN(
        P1_U3051) );
  AOI22_X1 U24148 ( .A1(n22749), .A2(n11347), .B1(n22592), .B2(n22748), .ZN(
        n22566) );
  AOI22_X1 U24149 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22751), .B1(
        n22750), .B2(n22594), .ZN(n22565) );
  OAI211_X1 U24150 ( .C1(n22754), .C2(n22585), .A(n22566), .B(n22565), .ZN(
        P1_U3059) );
  AOI22_X1 U24151 ( .A1(n22593), .A2(n22699), .B1(n22592), .B2(n22698), .ZN(
        n22568) );
  AOI22_X1 U24152 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n22700), .B1(
        n22750), .B2(n11347), .ZN(n22567) );
  OAI211_X1 U24153 ( .C1(n22591), .C2(n22760), .A(n22568), .B(n22567), .ZN(
        P1_U3067) );
  AOI22_X1 U24154 ( .A1(n22593), .A2(n22756), .B1(n22592), .B2(n22755), .ZN(
        n22570) );
  AOI22_X1 U24155 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n22757), .B1(
        n22762), .B2(n22594), .ZN(n22569) );
  OAI211_X1 U24156 ( .C1(n11346), .C2(n22760), .A(n22570), .B(n22569), .ZN(
        P1_U3075) );
  AOI22_X1 U24157 ( .A1(n22761), .A2(n22594), .B1(n22592), .B2(n11343), .ZN(
        n22572) );
  AOI22_X1 U24158 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n22763), .B1(
        n22762), .B2(n11347), .ZN(n22571) );
  OAI211_X1 U24159 ( .C1(n22766), .C2(n22585), .A(n22572), .B(n22571), .ZN(
        P1_U3083) );
  AOI22_X1 U24160 ( .A1(n22593), .A2(n22706), .B1(n22592), .B2(n22705), .ZN(
        n22574) );
  AOI22_X1 U24161 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n22707), .B1(
        n22761), .B2(n11347), .ZN(n22573) );
  OAI211_X1 U24162 ( .C1(n22591), .C2(n22710), .A(n22574), .B(n22573), .ZN(
        P1_U3091) );
  AOI22_X1 U24163 ( .A1(n22712), .A2(n22593), .B1(n22592), .B2(n22711), .ZN(
        n22576) );
  AOI22_X1 U24164 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n22714), .B1(
        n22713), .B2(n11347), .ZN(n22575) );
  OAI211_X1 U24165 ( .C1(n22591), .C2(n22772), .A(n22576), .B(n22575), .ZN(
        P1_U3099) );
  AOI22_X1 U24166 ( .A1(n22593), .A2(n22768), .B1(n22592), .B2(n22767), .ZN(
        n22578) );
  AOI22_X1 U24167 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22769), .B1(
        n22774), .B2(n22594), .ZN(n22577) );
  OAI211_X1 U24168 ( .C1(n11346), .C2(n22772), .A(n22578), .B(n22577), .ZN(
        P1_U3107) );
  AOI22_X1 U24169 ( .A1(n22775), .A2(n22594), .B1(n22592), .B2(n22773), .ZN(
        n22580) );
  AOI22_X1 U24170 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22776), .B1(
        n22774), .B2(n11347), .ZN(n22579) );
  OAI211_X1 U24171 ( .C1(n22779), .C2(n22585), .A(n22580), .B(n22579), .ZN(
        P1_U3115) );
  AOI22_X1 U24172 ( .A1(n22593), .A2(n22720), .B1(n22592), .B2(n22719), .ZN(
        n22582) );
  AOI22_X1 U24173 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n22721), .B1(
        n22775), .B2(n11347), .ZN(n22581) );
  OAI211_X1 U24174 ( .C1(n22591), .C2(n22724), .A(n22582), .B(n22581), .ZN(
        P1_U3123) );
  AOI22_X1 U24175 ( .A1(n22781), .A2(n22594), .B1(n22592), .B2(n22780), .ZN(
        n22584) );
  AOI22_X1 U24176 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n22784), .B1(
        n22783), .B2(n11347), .ZN(n22583) );
  OAI211_X1 U24177 ( .C1(n22788), .C2(n22585), .A(n22584), .B(n22583), .ZN(
        P1_U3131) );
  AOI22_X1 U24178 ( .A1(n22593), .A2(n22790), .B1(n22592), .B2(n22789), .ZN(
        n22587) );
  AOI22_X1 U24179 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22792), .B1(
        n22791), .B2(n22594), .ZN(n22586) );
  OAI211_X1 U24180 ( .C1(n11346), .C2(n22795), .A(n22587), .B(n22586), .ZN(
        P1_U3139) );
  AOI22_X1 U24181 ( .A1(n22593), .A2(n22731), .B1(n22592), .B2(n22729), .ZN(
        n22590) );
  AOI22_X1 U24182 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22733), .B1(
        n22791), .B2(n11347), .ZN(n22589) );
  OAI211_X1 U24183 ( .C1(n22591), .C2(n22804), .A(n22590), .B(n22589), .ZN(
        P1_U3147) );
  AOI22_X1 U24184 ( .A1(n22593), .A2(n22798), .B1(n22592), .B2(n22796), .ZN(
        n22596) );
  AOI22_X1 U24185 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n22801), .B1(
        n22800), .B2(n22594), .ZN(n22595) );
  OAI211_X1 U24186 ( .C1(n11346), .C2(n22804), .A(n22596), .B(n22595), .ZN(
        P1_U3155) );
  AOI22_X1 U24187 ( .A1(n22800), .A2(n15382), .B1(n22621), .B2(n22736), .ZN(
        n22598) );
  AOI22_X1 U24188 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22738), .B1(
        n22737), .B2(n11340), .ZN(n22597) );
  OAI211_X1 U24189 ( .C1(n22741), .C2(n22620), .A(n22598), .B(n22597), .ZN(
        P1_U3036) );
  AOI22_X1 U24190 ( .A1(n22622), .A2(n22689), .B1(n22621), .B2(n22688), .ZN(
        n22600) );
  AOI22_X1 U24191 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n22737), .B2(n15382), .ZN(n22599) );
  OAI211_X1 U24192 ( .C1(n11339), .C2(n22693), .A(n22600), .B(n22599), .ZN(
        P1_U3044) );
  AOI22_X1 U24193 ( .A1(n22743), .A2(n15382), .B1(n22742), .B2(n22621), .ZN(
        n22602) );
  AOI22_X1 U24194 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22744), .B1(
        n22749), .B2(n11340), .ZN(n22601) );
  OAI211_X1 U24195 ( .C1(n22747), .C2(n22620), .A(n22602), .B(n22601), .ZN(
        P1_U3052) );
  AOI22_X1 U24196 ( .A1(n22750), .A2(n11340), .B1(n22621), .B2(n22748), .ZN(
        n22604) );
  AOI22_X1 U24197 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n22749), .B2(n15382), .ZN(n22603) );
  OAI211_X1 U24198 ( .C1(n22754), .C2(n22620), .A(n22604), .B(n22603), .ZN(
        P1_U3060) );
  AOI22_X1 U24199 ( .A1(n22622), .A2(n22699), .B1(n22621), .B2(n22698), .ZN(
        n22606) );
  AOI22_X1 U24200 ( .A1(n22700), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n22750), .B2(n15382), .ZN(n22605) );
  OAI211_X1 U24201 ( .C1(n11339), .C2(n22760), .A(n22606), .B(n22605), .ZN(
        P1_U3068) );
  AOI22_X1 U24202 ( .A1(n22762), .A2(n15382), .B1(n11343), .B2(n22621), .ZN(
        n22608) );
  AOI22_X1 U24203 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n22763), .B1(
        n22761), .B2(n11340), .ZN(n22607) );
  OAI211_X1 U24204 ( .C1(n22766), .C2(n22620), .A(n22608), .B(n22607), .ZN(
        P1_U3084) );
  AOI22_X1 U24205 ( .A1(n22622), .A2(n22706), .B1(n22621), .B2(n22705), .ZN(
        n22610) );
  AOI22_X1 U24206 ( .A1(n22707), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n22761), .B2(n15382), .ZN(n22609) );
  OAI211_X1 U24207 ( .C1(n11339), .C2(n22710), .A(n22610), .B(n22609), .ZN(
        P1_U3092) );
  AOI22_X1 U24208 ( .A1(n22712), .A2(n22622), .B1(n22621), .B2(n22711), .ZN(
        n22612) );
  AOI22_X1 U24209 ( .A1(n22714), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n22713), .B2(n15382), .ZN(n22611) );
  OAI211_X1 U24210 ( .C1(n11339), .C2(n22772), .A(n22612), .B(n22611), .ZN(
        P1_U3100) );
  AOI22_X1 U24211 ( .A1(n22775), .A2(n11340), .B1(n22621), .B2(n22773), .ZN(
        n22614) );
  AOI22_X1 U24212 ( .A1(n22776), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n22774), .B2(n15382), .ZN(n22613) );
  OAI211_X1 U24213 ( .C1(n22779), .C2(n22620), .A(n22614), .B(n22613), .ZN(
        P1_U3116) );
  AOI22_X1 U24214 ( .A1(n22622), .A2(n22720), .B1(n22621), .B2(n22719), .ZN(
        n22616) );
  AOI22_X1 U24215 ( .A1(n22721), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n22775), .B2(n15382), .ZN(n22615) );
  OAI211_X1 U24216 ( .C1(n11339), .C2(n22724), .A(n22616), .B(n22615), .ZN(
        P1_U3124) );
  AOI22_X1 U24217 ( .A1(n22781), .A2(n11340), .B1(n22621), .B2(n22780), .ZN(
        n22619) );
  AOI22_X1 U24218 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22783), .B2(n15382), .ZN(n22618) );
  OAI211_X1 U24219 ( .C1(n22788), .C2(n22620), .A(n22619), .B(n22618), .ZN(
        P1_U3132) );
  AOI22_X1 U24220 ( .A1(n22622), .A2(n22731), .B1(n22621), .B2(n22729), .ZN(
        n22624) );
  AOI22_X1 U24221 ( .A1(n22733), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n22791), .B2(n15382), .ZN(n22623) );
  OAI211_X1 U24222 ( .C1(n11339), .C2(n22804), .A(n22624), .B(n22623), .ZN(
        P1_U3148) );
  NAND2_X1 U24223 ( .A1(n22626), .A2(n22625), .ZN(n22660) );
  INV_X1 U24224 ( .A(DATAI_28_), .ZN(n22627) );
  OAI22_X1 U24225 ( .A1(n22628), .A2(n22630), .B1(n22627), .B2(n22632), .ZN(
        n22663) );
  NOR2_X2 U24226 ( .A1(n22629), .A2(n14550), .ZN(n22666) );
  AOI22_X1 U24227 ( .A1(n22800), .A2(n11349), .B1(n22666), .B2(n22736), .ZN(
        n22635) );
  OAI22_X1 U24228 ( .A1(n22633), .A2(n22632), .B1(n22631), .B2(n22630), .ZN(
        n22668) );
  AOI22_X1 U24229 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22738), .B1(
        n22737), .B2(n11336), .ZN(n22634) );
  OAI211_X1 U24230 ( .C1(n22741), .C2(n22660), .A(n22635), .B(n22634), .ZN(
        P1_U3037) );
  AOI22_X1 U24231 ( .A1(n22667), .A2(n22689), .B1(n22666), .B2(n22688), .ZN(
        n22637) );
  AOI22_X1 U24232 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22690), .B1(
        n22737), .B2(n11349), .ZN(n22636) );
  OAI211_X1 U24233 ( .C1(n11335), .C2(n22693), .A(n22637), .B(n22636), .ZN(
        P1_U3045) );
  AOI22_X1 U24234 ( .A1(n22743), .A2(n11349), .B1(n22666), .B2(n22742), .ZN(
        n22639) );
  AOI22_X1 U24235 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22744), .B1(
        n22749), .B2(n11336), .ZN(n22638) );
  OAI211_X1 U24236 ( .C1(n22747), .C2(n22660), .A(n22639), .B(n22638), .ZN(
        P1_U3053) );
  AOI22_X1 U24237 ( .A1(n22750), .A2(n11336), .B1(n22666), .B2(n22748), .ZN(
        n22641) );
  AOI22_X1 U24238 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n22751), .B1(
        n22749), .B2(n11349), .ZN(n22640) );
  OAI211_X1 U24239 ( .C1(n22754), .C2(n22660), .A(n22641), .B(n22640), .ZN(
        P1_U3061) );
  AOI22_X1 U24240 ( .A1(n22667), .A2(n22699), .B1(n22666), .B2(n22698), .ZN(
        n22643) );
  AOI22_X1 U24241 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n22700), .B1(
        n22750), .B2(n11349), .ZN(n22642) );
  OAI211_X1 U24242 ( .C1(n11335), .C2(n22760), .A(n22643), .B(n22642), .ZN(
        P1_U3069) );
  AOI22_X1 U24243 ( .A1(n22667), .A2(n22756), .B1(n22666), .B2(n22755), .ZN(
        n22645) );
  AOI22_X1 U24244 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n22757), .B1(
        n22762), .B2(n11336), .ZN(n22644) );
  OAI211_X1 U24245 ( .C1(n11348), .C2(n22760), .A(n22645), .B(n22644), .ZN(
        P1_U3077) );
  AOI22_X1 U24246 ( .A1(n22761), .A2(n11336), .B1(n22666), .B2(n11343), .ZN(
        n22647) );
  AOI22_X1 U24247 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n22763), .B1(
        n22762), .B2(n11349), .ZN(n22646) );
  OAI211_X1 U24248 ( .C1(n22766), .C2(n22660), .A(n22647), .B(n22646), .ZN(
        P1_U3085) );
  AOI22_X1 U24249 ( .A1(n22667), .A2(n22706), .B1(n22666), .B2(n22705), .ZN(
        n22649) );
  AOI22_X1 U24250 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n22707), .B1(
        n22761), .B2(n11349), .ZN(n22648) );
  OAI211_X1 U24251 ( .C1(n11335), .C2(n22710), .A(n22649), .B(n22648), .ZN(
        P1_U3093) );
  AOI22_X1 U24252 ( .A1(n22712), .A2(n22667), .B1(n22666), .B2(n22711), .ZN(
        n22651) );
  AOI22_X1 U24253 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n22714), .B1(
        n22713), .B2(n11349), .ZN(n22650) );
  OAI211_X1 U24254 ( .C1(n11335), .C2(n22772), .A(n22651), .B(n22650), .ZN(
        P1_U3101) );
  AOI22_X1 U24255 ( .A1(n22667), .A2(n22768), .B1(n22666), .B2(n22767), .ZN(
        n22653) );
  AOI22_X1 U24256 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22769), .B1(
        n22774), .B2(n11336), .ZN(n22652) );
  OAI211_X1 U24257 ( .C1(n11348), .C2(n22772), .A(n22653), .B(n22652), .ZN(
        P1_U3109) );
  AOI22_X1 U24258 ( .A1(n22774), .A2(n11349), .B1(n22666), .B2(n22773), .ZN(
        n22655) );
  AOI22_X1 U24259 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22776), .B1(
        n22775), .B2(n11336), .ZN(n22654) );
  OAI211_X1 U24260 ( .C1(n22779), .C2(n22660), .A(n22655), .B(n22654), .ZN(
        P1_U3117) );
  AOI22_X1 U24261 ( .A1(n22667), .A2(n22720), .B1(n22666), .B2(n22719), .ZN(
        n22657) );
  AOI22_X1 U24262 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n22721), .B1(
        n22775), .B2(n11349), .ZN(n22656) );
  OAI211_X1 U24263 ( .C1(n11335), .C2(n22724), .A(n22657), .B(n22656), .ZN(
        P1_U3125) );
  AOI22_X1 U24264 ( .A1(n22781), .A2(n11336), .B1(n22666), .B2(n22780), .ZN(
        n22659) );
  AOI22_X1 U24265 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n22784), .B1(
        n22783), .B2(n11349), .ZN(n22658) );
  OAI211_X1 U24266 ( .C1(n22788), .C2(n22660), .A(n22659), .B(n22658), .ZN(
        P1_U3133) );
  AOI22_X1 U24267 ( .A1(n22667), .A2(n22790), .B1(n22666), .B2(n22789), .ZN(
        n22662) );
  AOI22_X1 U24268 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22792), .B1(
        n22791), .B2(n11336), .ZN(n22661) );
  OAI211_X1 U24269 ( .C1(n11348), .C2(n22795), .A(n22662), .B(n22661), .ZN(
        P1_U3141) );
  AOI22_X1 U24270 ( .A1(n22667), .A2(n22731), .B1(n22666), .B2(n22729), .ZN(
        n22665) );
  AOI22_X1 U24271 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22733), .B1(
        n22791), .B2(n11349), .ZN(n22664) );
  OAI211_X1 U24272 ( .C1(n11335), .C2(n22804), .A(n22665), .B(n22664), .ZN(
        P1_U3149) );
  AOI22_X1 U24273 ( .A1(n22667), .A2(n22798), .B1(n22666), .B2(n22796), .ZN(
        n22670) );
  AOI22_X1 U24274 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n22801), .B1(
        n22800), .B2(n11336), .ZN(n22669) );
  OAI211_X1 U24275 ( .C1(n11348), .C2(n22804), .A(n22670), .B(n22669), .ZN(
        P1_U3157) );
  AOI22_X1 U24276 ( .A1(n22800), .A2(n22682), .B1(n22681), .B2(n22736), .ZN(
        n22672) );
  AOI22_X1 U24277 ( .A1(n22738), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n22737), .B2(n15591), .ZN(n22671) );
  OAI211_X1 U24278 ( .C1(n22741), .C2(n22685), .A(n22672), .B(n22671), .ZN(
        P1_U3038) );
  AOI22_X1 U24279 ( .A1(n22743), .A2(n22682), .B1(n22742), .B2(n22681), .ZN(
        n22674) );
  AOI22_X1 U24280 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n22749), .B2(n15591), .ZN(n22673) );
  OAI211_X1 U24281 ( .C1(n22747), .C2(n22685), .A(n22674), .B(n22673), .ZN(
        P1_U3054) );
  AOI22_X1 U24282 ( .A1(n22749), .A2(n22682), .B1(n22748), .B2(n22681), .ZN(
        n22676) );
  AOI22_X1 U24283 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n22750), .B2(n15591), .ZN(n22675) );
  OAI211_X1 U24284 ( .C1(n22754), .C2(n22685), .A(n22676), .B(n22675), .ZN(
        P1_U3062) );
  AOI22_X1 U24285 ( .A1(n22761), .A2(n15591), .B1(n11343), .B2(n22681), .ZN(
        n22678) );
  AOI22_X1 U24286 ( .A1(n22763), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22762), .B2(n22682), .ZN(n22677) );
  OAI211_X1 U24287 ( .C1(n22766), .C2(n22685), .A(n22678), .B(n22677), .ZN(
        P1_U3086) );
  AOI22_X1 U24288 ( .A1(n22774), .A2(n22682), .B1(n22773), .B2(n22681), .ZN(
        n22680) );
  AOI22_X1 U24289 ( .A1(n22776), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n22775), .B2(n15591), .ZN(n22679) );
  OAI211_X1 U24290 ( .C1(n22779), .C2(n22685), .A(n22680), .B(n22679), .ZN(
        P1_U3118) );
  AOI22_X1 U24291 ( .A1(n22781), .A2(n15591), .B1(n22780), .B2(n22681), .ZN(
        n22684) );
  AOI22_X1 U24292 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n22783), .B2(n22682), .ZN(n22683) );
  OAI211_X1 U24293 ( .C1(n22788), .C2(n22685), .A(n22684), .B(n22683), .ZN(
        P1_U3134) );
  AOI22_X1 U24294 ( .A1(n22800), .A2(n15528), .B1(n22730), .B2(n22736), .ZN(
        n22687) );
  AOI22_X1 U24295 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22738), .B1(
        n22737), .B2(n11338), .ZN(n22686) );
  OAI211_X1 U24296 ( .C1(n22741), .C2(n22728), .A(n22687), .B(n22686), .ZN(
        P1_U3039) );
  AOI22_X1 U24297 ( .A1(n22732), .A2(n22689), .B1(n22730), .B2(n22688), .ZN(
        n22692) );
  AOI22_X1 U24298 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n22737), .B2(n15528), .ZN(n22691) );
  OAI211_X1 U24299 ( .C1(n11337), .C2(n22693), .A(n22692), .B(n22691), .ZN(
        P1_U3047) );
  AOI22_X1 U24300 ( .A1(n22743), .A2(n15528), .B1(n22742), .B2(n22730), .ZN(
        n22695) );
  AOI22_X1 U24301 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22744), .B1(
        n22749), .B2(n11338), .ZN(n22694) );
  OAI211_X1 U24302 ( .C1(n22747), .C2(n22728), .A(n22695), .B(n22694), .ZN(
        P1_U3055) );
  AOI22_X1 U24303 ( .A1(n22750), .A2(n11338), .B1(n22730), .B2(n22748), .ZN(
        n22697) );
  AOI22_X1 U24304 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22749), .B2(n15528), .ZN(n22696) );
  OAI211_X1 U24305 ( .C1(n22754), .C2(n22728), .A(n22697), .B(n22696), .ZN(
        P1_U3063) );
  AOI22_X1 U24306 ( .A1(n22732), .A2(n22699), .B1(n22730), .B2(n22698), .ZN(
        n22702) );
  AOI22_X1 U24307 ( .A1(n22700), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n22750), .B2(n15528), .ZN(n22701) );
  OAI211_X1 U24308 ( .C1(n11337), .C2(n22760), .A(n22702), .B(n22701), .ZN(
        P1_U3071) );
  AOI22_X1 U24309 ( .A1(n22762), .A2(n15528), .B1(n11343), .B2(n22730), .ZN(
        n22704) );
  AOI22_X1 U24310 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n22763), .B1(
        n22761), .B2(n11338), .ZN(n22703) );
  OAI211_X1 U24311 ( .C1(n22766), .C2(n22728), .A(n22704), .B(n22703), .ZN(
        P1_U3087) );
  AOI22_X1 U24312 ( .A1(n22732), .A2(n22706), .B1(n22730), .B2(n22705), .ZN(
        n22709) );
  AOI22_X1 U24313 ( .A1(n22707), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n22761), .B2(n15528), .ZN(n22708) );
  OAI211_X1 U24314 ( .C1(n11337), .C2(n22710), .A(n22709), .B(n22708), .ZN(
        P1_U3095) );
  AOI22_X1 U24315 ( .A1(n22712), .A2(n22732), .B1(n22730), .B2(n22711), .ZN(
        n22716) );
  AOI22_X1 U24316 ( .A1(n22714), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n22713), .B2(n15528), .ZN(n22715) );
  OAI211_X1 U24317 ( .C1(n11337), .C2(n22772), .A(n22716), .B(n22715), .ZN(
        P1_U3103) );
  AOI22_X1 U24318 ( .A1(n22775), .A2(n11338), .B1(n22730), .B2(n22773), .ZN(
        n22718) );
  AOI22_X1 U24319 ( .A1(n22776), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n22774), .B2(n15528), .ZN(n22717) );
  OAI211_X1 U24320 ( .C1(n22779), .C2(n22728), .A(n22718), .B(n22717), .ZN(
        P1_U3119) );
  AOI22_X1 U24321 ( .A1(n22732), .A2(n22720), .B1(n22730), .B2(n22719), .ZN(
        n22723) );
  AOI22_X1 U24322 ( .A1(n22721), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n22775), .B2(n15528), .ZN(n22722) );
  OAI211_X1 U24323 ( .C1(n11337), .C2(n22724), .A(n22723), .B(n22722), .ZN(
        P1_U3127) );
  AOI22_X1 U24324 ( .A1(n22781), .A2(n11338), .B1(n22730), .B2(n22780), .ZN(
        n22727) );
  AOI22_X1 U24325 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22783), .B2(n15528), .ZN(n22726) );
  OAI211_X1 U24326 ( .C1(n22788), .C2(n22728), .A(n22727), .B(n22726), .ZN(
        P1_U3135) );
  AOI22_X1 U24327 ( .A1(n22732), .A2(n22731), .B1(n22730), .B2(n22729), .ZN(
        n22735) );
  AOI22_X1 U24328 ( .A1(n22733), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n22791), .B2(n15528), .ZN(n22734) );
  OAI211_X1 U24329 ( .C1(n11337), .C2(n22804), .A(n22735), .B(n22734), .ZN(
        P1_U3151) );
  AOI22_X1 U24330 ( .A1(n22800), .A2(n11345), .B1(n22797), .B2(n22736), .ZN(
        n22740) );
  AOI22_X1 U24331 ( .A1(n22738), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n22737), .B2(n15142), .ZN(n22739) );
  OAI211_X1 U24332 ( .C1(n22741), .C2(n22787), .A(n22740), .B(n22739), .ZN(
        P1_U3040) );
  AOI22_X1 U24333 ( .A1(n22743), .A2(n11345), .B1(n22797), .B2(n22742), .ZN(
        n22746) );
  AOI22_X1 U24334 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n22749), .B2(n15142), .ZN(n22745) );
  OAI211_X1 U24335 ( .C1(n22747), .C2(n22787), .A(n22746), .B(n22745), .ZN(
        P1_U3056) );
  AOI22_X1 U24336 ( .A1(n22749), .A2(n11345), .B1(n22797), .B2(n22748), .ZN(
        n22753) );
  AOI22_X1 U24337 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n22750), .B2(n15142), .ZN(n22752) );
  OAI211_X1 U24338 ( .C1(n22754), .C2(n22787), .A(n22753), .B(n22752), .ZN(
        P1_U3064) );
  AOI22_X1 U24339 ( .A1(n22799), .A2(n22756), .B1(n22797), .B2(n22755), .ZN(
        n22759) );
  AOI22_X1 U24340 ( .A1(n22757), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n22762), .B2(n15142), .ZN(n22758) );
  OAI211_X1 U24341 ( .C1(n11344), .C2(n22760), .A(n22759), .B(n22758), .ZN(
        P1_U3080) );
  AOI22_X1 U24342 ( .A1(n22761), .A2(n15142), .B1(n11343), .B2(n22797), .ZN(
        n22765) );
  AOI22_X1 U24343 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n22763), .B1(
        n22762), .B2(n11345), .ZN(n22764) );
  OAI211_X1 U24344 ( .C1(n22766), .C2(n22787), .A(n22765), .B(n22764), .ZN(
        P1_U3088) );
  AOI22_X1 U24345 ( .A1(n22799), .A2(n22768), .B1(n22797), .B2(n22767), .ZN(
        n22771) );
  AOI22_X1 U24346 ( .A1(n22769), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n22774), .B2(n15142), .ZN(n22770) );
  OAI211_X1 U24347 ( .C1(n11344), .C2(n22772), .A(n22771), .B(n22770), .ZN(
        P1_U3112) );
  AOI22_X1 U24348 ( .A1(n22774), .A2(n11345), .B1(n22797), .B2(n22773), .ZN(
        n22778) );
  AOI22_X1 U24349 ( .A1(n22776), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n22775), .B2(n15142), .ZN(n22777) );
  OAI211_X1 U24350 ( .C1(n22779), .C2(n22787), .A(n22778), .B(n22777), .ZN(
        P1_U3120) );
  AOI22_X1 U24351 ( .A1(n22781), .A2(n15142), .B1(n22780), .B2(n22797), .ZN(
        n22786) );
  AOI22_X1 U24352 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22784), .B1(
        n22783), .B2(n11345), .ZN(n22785) );
  OAI211_X1 U24353 ( .C1(n22788), .C2(n22787), .A(n22786), .B(n22785), .ZN(
        P1_U3136) );
  AOI22_X1 U24354 ( .A1(n22799), .A2(n22790), .B1(n22797), .B2(n22789), .ZN(
        n22794) );
  AOI22_X1 U24355 ( .A1(n22792), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n22791), .B2(n15142), .ZN(n22793) );
  OAI211_X1 U24356 ( .C1(n11344), .C2(n22795), .A(n22794), .B(n22793), .ZN(
        P1_U3144) );
  AOI22_X1 U24357 ( .A1(n22799), .A2(n22798), .B1(n22797), .B2(n22796), .ZN(
        n22803) );
  AOI22_X1 U24358 ( .A1(n22801), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n22800), .B2(n15142), .ZN(n22802) );
  OAI211_X1 U24359 ( .C1(n11344), .C2(n22804), .A(n22803), .B(n22802), .ZN(
        P1_U3160) );
  OAI22_X1 U24360 ( .A1(n22806), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n22805), .ZN(n22807) );
  INV_X1 U24361 ( .A(n22807), .ZN(P1_U3486) );
  NAND3_X1 U24362 ( .A1(n22810), .A2(n22809), .A3(n22808), .ZN(n22811) );
  NAND2_X1 U24363 ( .A1(n22811), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22812)
         );
  NAND3_X1 U24364 ( .A1(n22814), .A2(n22813), .A3(n22812), .ZN(P1_U2801) );
  INV_X2 U11407 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15200) );
  CLKBUF_X2 U14960 ( .A(n13320), .Z(n16397) );
  CLKBUF_X3 U11404 ( .A(n18122), .Z(n11164) );
  AND2_X1 U14957 ( .A1(n11162), .A2(n15200), .ZN(n16232) );
  OR2_X1 U13488 ( .A1(n12001), .A2(n12000), .ZN(n12059) );
  AND4_X1 U11351 ( .A1(n14119), .A2(n14124), .A3(n14123), .A4(n14125), .ZN(
        n11483) );
  CLKBUF_X1 U11312 ( .A(n12037), .Z(n12638) );
  NAND2_X1 U11315 ( .A1(n12029), .A2(n12028), .ZN(n12163) );
  XNOR2_X1 U11327 ( .A(n14203), .B(n14204), .ZN(n14312) );
  CLKBUF_X1 U11330 ( .A(n11921), .Z(n14580) );
  CLKBUF_X1 U11368 ( .A(n13104), .Z(n16136) );
  CLKBUF_X1 U11644 ( .A(n13109), .Z(n20178) );
  CLKBUF_X1 U11645 ( .A(n12179), .Z(n15412) );
  CLKBUF_X1 U12108 ( .A(n17836), .Z(n17850) );
  CLKBUF_X1 U12358 ( .A(n20669), .Z(n20677) );
endmodule

