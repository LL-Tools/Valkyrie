

module b21_C_SARLock_k_64_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4264, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10017;

  OAI21_X1 U4770 ( .B1(n4452), .B2(n8197), .A(n8196), .ZN(n9191) );
  NAND2_X1 U4771 ( .A1(n8361), .A2(n8362), .ZN(n8435) );
  INV_X1 U4772 ( .A(n5050), .ZN(n5628) );
  NAND2_X2 U4773 ( .A1(n5561), .A2(n5585), .ZN(n5650) );
  NAND2_X1 U4774 ( .A1(n6456), .A2(n7244), .ZN(n6499) );
  XNOR2_X1 U4775 ( .A(n4861), .B(SI_5_), .ZN(n5095) );
  INV_X1 U4776 ( .A(n10017), .ZN(n4264) );
  INV_X2 U4777 ( .A(n4264), .ZN(P2_U3152) );
  INV_X1 U4778 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n10017) );
  AND2_X1 U4779 ( .A1(n4638), .A2(n7017), .ZN(n5829) );
  AND2_X1 U4780 ( .A1(n5427), .A2(n5426), .ZN(n8367) );
  AND2_X1 U4781 ( .A1(n5009), .A2(n8262), .ZN(n5051) );
  OR2_X1 U4782 ( .A1(n5856), .A2(n4831), .ZN(n5857) );
  NOR2_X2 U4783 ( .A1(n9268), .A2(n9442), .ZN(n9260) );
  AND2_X1 U4784 ( .A1(n4623), .A2(n5095), .ZN(n4627) );
  AND2_X1 U4785 ( .A1(n5411), .A2(n4827), .ZN(n5427) );
  NAND2_X1 U4786 ( .A1(n8311), .A2(n4654), .ZN(n8393) );
  INV_X1 U4787 ( .A(n5012), .ZN(n5629) );
  NOR2_X1 U4788 ( .A1(n8703), .A2(n8853), .ZN(n8687) );
  NAND2_X1 U4789 ( .A1(n7303), .A2(n7302), .ZN(n7751) );
  INV_X2 U4791 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5528) );
  INV_X1 U4792 ( .A(n6452), .ZN(n6387) );
  INV_X1 U4793 ( .A(n4446), .ZN(n7939) );
  INV_X1 U4794 ( .A(n6025), .ZN(n7942) );
  OAI21_X1 U4795 ( .B1(n6067), .B2(n6583), .A(n4447), .ZN(n9730) );
  XNOR2_X1 U4796 ( .A(n5427), .B(n5416), .ZN(n8287) );
  NAND2_X1 U4797 ( .A1(n8342), .A2(n8341), .ZN(n8447) );
  NAND2_X1 U4798 ( .A1(n8401), .A2(n8402), .ZN(n8400) );
  AND4_X1 U4799 ( .A1(n5090), .A2(n5089), .A3(n5088), .A4(n4833), .ZN(n7224)
         );
  NAND2_X1 U4800 ( .A1(n4684), .A2(n4322), .ZN(n7722) );
  NAND2_X1 U4801 ( .A1(n5850), .A2(n5893), .ZN(n9624) );
  XNOR2_X1 U4802 ( .A(n4989), .B(n4988), .ZN(n5562) );
  INV_X1 U4803 ( .A(n4266), .ZN(n4267) );
  OAI211_X2 U4804 ( .C1(n6067), .C2(n6591), .A(n5987), .B(n5986), .ZN(n7107)
         );
  OAI21_X2 U4805 ( .B1(n9191), .B2(n4329), .A(n4783), .ZN(n4782) );
  OAI222_X1 U4806 ( .A1(n9524), .A2(n6598), .B1(n9522), .B2(n6032), .C1(
        P1_U3084), .C2(n6597), .ZN(P1_U3347) );
  OAI222_X1 U4807 ( .A1(n6913), .A2(P2_U3152), .B1(n8920), .B2(n6032), .C1(
        n6580), .C2(n8259), .ZN(P2_U3352) );
  NOR3_X2 U4808 ( .A1(n6884), .A2(n6883), .A3(n6971), .ZN(n6972) );
  INV_X1 U4809 ( .A(n8250), .ZN(n4266) );
  AOI21_X2 U4810 ( .B1(n6266), .B2(n6265), .A(n8969), .ZN(n9007) );
  OAI21_X2 U4811 ( .B1(n5805), .B2(n7605), .A(n5673), .ZN(n7015) );
  NOR2_X2 U4812 ( .A1(n9378), .A2(n9470), .ZN(n9379) );
  XNOR2_X2 U4813 ( .A(n5005), .B(n5004), .ZN(n8262) );
  NAND2_X2 U4814 ( .A1(n5140), .A2(n5139), .ZN(n9904) );
  NAND2_X1 U4815 ( .A1(n4990), .A2(n7262), .ZN(n4268) );
  NAND2_X1 U4816 ( .A1(n4990), .A2(n7262), .ZN(n4269) );
  NAND2_X1 U4817 ( .A1(n4990), .A2(n7262), .ZN(n5049) );
  OAI21_X1 U4818 ( .B1(n5776), .B2(n4503), .A(n4501), .ZN(n4505) );
  AND3_X1 U4819 ( .A1(n5774), .A2(n5773), .A3(n5772), .ZN(n5776) );
  OAI21_X1 U4820 ( .B1(n8631), .B2(n4271), .A(n4272), .ZN(n8604) );
  NAND2_X1 U4821 ( .A1(n5653), .A2(n4274), .ZN(n4273) );
  AND2_X1 U4822 ( .A1(n7214), .A2(n7220), .ZN(n7312) );
  INV_X2 U4823 ( .A(n8387), .ZN(n7215) );
  NOR2_X1 U4824 ( .A1(n7606), .A2(n5496), .ZN(n5036) );
  INV_X1 U4826 ( .A(n8301), .ZN(n7492) );
  AND2_X1 U4827 ( .A1(n5914), .A2(n5880), .ZN(n6456) );
  NAND2_X1 U4828 ( .A1(n5914), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5915) );
  INV_X4 U4829 ( .A(n5650), .ZN(n5496) );
  NAND2_X1 U4830 ( .A1(n5879), .A2(n5878), .ZN(n5914) );
  AND4_X1 U4831 ( .A1(n5984), .A2(n5983), .A3(n5982), .A4(n5981), .ZN(n7192)
         );
  CLKBUF_X3 U4832 ( .A(n5051), .Z(n4284) );
  INV_X4 U4833 ( .A(n5790), .ZN(n4270) );
  NAND2_X2 U4834 ( .A1(n8245), .A2(n5900), .ZN(n5989) );
  NOR2_X1 U4835 ( .A1(n5007), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U4836 ( .A1(n5022), .A2(n4549), .ZN(n6978) );
  OAI21_X1 U4837 ( .B1(n5651), .B2(n4822), .A(n4520), .ZN(n4477) );
  NOR2_X1 U4838 ( .A1(n4633), .A2(n8816), .ZN(n8819) );
  NAND2_X1 U4839 ( .A1(n4395), .A2(n4649), .ZN(n8448) );
  AND2_X1 U4840 ( .A1(n9389), .A2(n9113), .ZN(n8170) );
  AND2_X1 U4841 ( .A1(n5792), .A2(n5782), .ZN(n5823) );
  AOI21_X1 U4842 ( .B1(n8239), .B2(n9725), .A(n8238), .ZN(n9398) );
  NAND2_X1 U4843 ( .A1(n4392), .A2(n4310), .ZN(n6380) );
  AOI21_X1 U4844 ( .B1(n7935), .B2(n5489), .A(n5645), .ZN(n8810) );
  NAND2_X1 U4845 ( .A1(n8604), .A2(n8610), .ZN(n8603) );
  XNOR2_X1 U4846 ( .A(n5643), .B(n5642), .ZN(n7935) );
  NAND2_X1 U4847 ( .A1(n8631), .A2(n8562), .ZN(n8618) );
  NAND2_X1 U4848 ( .A1(n4407), .A2(n8317), .ZN(n8320) );
  NAND2_X1 U4849 ( .A1(n8667), .A2(n8556), .ZN(n8666) );
  NAND2_X1 U4850 ( .A1(n4590), .A2(n4589), .ZN(n9215) );
  AND2_X1 U4851 ( .A1(n4273), .A2(n8564), .ZN(n4272) );
  NAND2_X1 U4852 ( .A1(n4332), .A2(n8127), .ZN(n4589) );
  AOI21_X1 U4853 ( .B1(n4749), .B2(n4747), .A(n4830), .ZN(n8667) );
  NAND2_X1 U4854 ( .A1(n4604), .A2(n4603), .ZN(n8747) );
  NAND2_X1 U4855 ( .A1(n8714), .A2(n4339), .ZN(n4749) );
  AOI22_X1 U4856 ( .A1(n8732), .A2(n8550), .B1(n8750), .B2(n8737), .ZN(n8714)
         );
  INV_X1 U4857 ( .A(n5653), .ZN(n4271) );
  NOR2_X1 U4858 ( .A1(n4320), .A2(n4376), .ZN(n4375) );
  INV_X1 U4859 ( .A(n8562), .ZN(n4274) );
  AND2_X1 U4860 ( .A1(n8554), .A2(n4748), .ZN(n4747) );
  NAND2_X1 U4861 ( .A1(n8775), .A2(n4341), .ZN(n4754) );
  NAND2_X1 U4862 ( .A1(n4690), .A2(n4688), .ZN(n7529) );
  NAND2_X1 U4863 ( .A1(n6383), .A2(n6382), .ZN(n9415) );
  NAND2_X1 U4864 ( .A1(n7828), .A2(n7829), .ZN(n7827) );
  NAND2_X1 U4865 ( .A1(n8777), .A2(n8776), .ZN(n8775) );
  NAND2_X1 U4866 ( .A1(n4462), .A2(n5399), .ZN(n8853) );
  AOI22_X1 U4867 ( .A1(n8791), .A2(n8797), .B1(n8796), .B2(n8546), .ZN(n8777)
         );
  AOI21_X1 U4868 ( .B1(n9348), .B2(n8189), .A(n8188), .ZN(n9333) );
  AOI21_X1 U4869 ( .B1(n4608), .B2(n4610), .A(n4607), .ZN(n4606) );
  AND2_X1 U4870 ( .A1(n5387), .A2(n5386), .ZN(n8706) );
  OR2_X1 U4871 ( .A1(n8778), .A2(n8880), .ZN(n8766) );
  NAND2_X1 U4872 ( .A1(n4277), .A2(n4275), .ZN(n4276) );
  AND2_X1 U4873 ( .A1(n4277), .A2(n7769), .ZN(n7772) );
  NAND2_X1 U4874 ( .A1(n6284), .A2(n6283), .ZN(n9446) );
  OR2_X1 U4875 ( .A1(n6182), .A2(n6181), .ZN(n7873) );
  OR2_X1 U4876 ( .A1(n7562), .A2(n7561), .ZN(n4277) );
  AND2_X1 U4877 ( .A1(n4337), .A2(n7769), .ZN(n4275) );
  NAND2_X1 U4878 ( .A1(n6205), .A2(n6206), .ZN(n7871) );
  NAND2_X1 U4879 ( .A1(n9797), .A2(n7557), .ZN(n7575) );
  NAND2_X1 U4880 ( .A1(n7555), .A2(n4761), .ZN(n9797) );
  NAND2_X1 U4881 ( .A1(n6168), .A2(n6167), .ZN(n9470) );
  NAND2_X1 U4882 ( .A1(n5250), .A2(n5249), .ZN(n8894) );
  NAND2_X1 U4883 ( .A1(n7751), .A2(n4762), .ZN(n7555) );
  NAND2_X1 U4884 ( .A1(n8427), .A2(n8482), .ZN(n7769) );
  NAND2_X1 U4885 ( .A1(n6187), .A2(n6186), .ZN(n9597) );
  NAND2_X1 U4886 ( .A1(n6136), .A2(n6135), .ZN(n9479) );
  XNOR2_X1 U4887 ( .A(n5246), .B(n4836), .ZN(n6790) );
  OAI21_X1 U4888 ( .B1(n5209), .B2(n4887), .A(n4886), .ZN(n5226) );
  NAND2_X1 U4889 ( .A1(n5198), .A2(n5197), .ZN(n9928) );
  NAND2_X2 U4890 ( .A1(n7270), .A2(n8678), .ZN(n9829) );
  AND2_X1 U4891 ( .A1(n5684), .A2(n5685), .ZN(n7290) );
  NAND2_X1 U4892 ( .A1(n4279), .A2(n7045), .ZN(n7293) );
  INV_X4 U4893 ( .A(n9740), .ZN(n9743) );
  XNOR2_X1 U4894 ( .A(n5192), .B(n4832), .ZN(n6732) );
  INV_X1 U4895 ( .A(n7444), .ZN(n9766) );
  INV_X1 U4896 ( .A(n7754), .ZN(n9900) );
  NAND2_X1 U4897 ( .A1(n4476), .A2(n4877), .ZN(n5192) );
  NAND2_X1 U4898 ( .A1(n4683), .A2(n4319), .ZN(n7444) );
  NAND2_X1 U4899 ( .A1(n4628), .A2(n4824), .ZN(n7754) );
  INV_X1 U4900 ( .A(n5805), .ZN(n7010) );
  NAND2_X1 U4901 ( .A1(n4714), .A2(n4717), .ZN(n5134) );
  NAND2_X1 U4902 ( .A1(n5673), .A2(n5674), .ZN(n5805) );
  NAND2_X1 U4903 ( .A1(n8491), .A2(n4266), .ZN(n5674) );
  NAND2_X1 U4904 ( .A1(n5659), .A2(n9874), .ZN(n9877) );
  CLKBUF_X1 U4905 ( .A(n6456), .Z(n8172) );
  NAND4_X1 U4906 ( .A1(n5105), .A2(n5104), .A3(n5103), .A4(n5102), .ZN(n8488)
         );
  NAND3_X1 U4907 ( .A1(n4842), .A2(n5026), .A3(n5025), .ZN(n8492) );
  NOR2_X1 U4908 ( .A1(n9730), .A2(n9731), .ZN(n9729) );
  INV_X1 U4909 ( .A(n4528), .ZN(n4527) );
  AND4_X1 U4910 ( .A1(n5076), .A2(n5075), .A3(n5074), .A4(n5073), .ZN(n7607)
         );
  OAI211_X1 U4911 ( .C1(n6877), .C2(n6991), .A(n5048), .B(n5047), .ZN(n8250)
         );
  AOI21_X1 U4912 ( .B1(n4381), .B2(n4383), .A(n4379), .ZN(n4378) );
  NAND4_X1 U4913 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n6544)
         );
  NAND2_X1 U4914 ( .A1(n4602), .A2(n4854), .ZN(n5069) );
  OAI21_X1 U4915 ( .B1(n6877), .B2(n6978), .A(n4488), .ZN(n7272) );
  CLKBUF_X1 U4916 ( .A(n4284), .Z(n5577) );
  NAND2_X1 U4917 ( .A1(n5877), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5879) );
  OR2_X1 U4918 ( .A1(n5097), .A2(n4479), .ZN(n5047) );
  AND2_X2 U4919 ( .A1(n6539), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NOR2_X1 U4920 ( .A1(n4718), .A2(n4716), .ZN(n4715) );
  AND2_X2 U4921 ( .A1(n5011), .A2(n5009), .ZN(n5072) );
  INV_X1 U4922 ( .A(n5876), .ZN(n5881) );
  AND2_X1 U4923 ( .A1(n5562), .A2(n7139), .ZN(n5585) );
  NOR2_X1 U4924 ( .A1(n5565), .A2(n5652), .ZN(n5790) );
  OR2_X1 U4925 ( .A1(n5565), .A2(n5662), .ZN(n4638) );
  AND2_X1 U4926 ( .A1(n8916), .A2(n5010), .ZN(n5009) );
  NAND2_X1 U4927 ( .A1(n4973), .A2(n4278), .ZN(n5832) );
  XNOR2_X1 U4928 ( .A(n5533), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U4929 ( .A1(n4987), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4989) );
  MUX2_X1 U4930 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5008), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5010) );
  OR2_X1 U4931 ( .A1(n4971), .A2(n4966), .ZN(n4973) );
  INV_X1 U4932 ( .A(n5662), .ZN(n7362) );
  AND2_X1 U4933 ( .A1(n4972), .A2(n4311), .ZN(n4278) );
  OR2_X1 U4934 ( .A1(n5006), .A2(n5528), .ZN(n5005) );
  NAND2_X1 U4935 ( .A1(n5527), .A2(n4490), .ZN(n4972) );
  INV_X8 U4936 ( .A(n4282), .ZN(n6581) );
  NAND2_X1 U4937 ( .A1(n4282), .A2(n4847), .ZN(n5029) );
  XNOR2_X1 U4938 ( .A(n4986), .B(n4985), .ZN(n7139) );
  NAND2_X1 U4939 ( .A1(P1_U3084), .A2(n4282), .ZN(n9524) );
  XNOR2_X1 U4940 ( .A(n4984), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5662) );
  OR2_X1 U4941 ( .A1(n4982), .A2(n5528), .ZN(n4986) );
  AND2_X1 U4942 ( .A1(n5263), .A2(n4962), .ZN(n5527) );
  NOR2_X1 U4943 ( .A1(n5860), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6120) );
  AND2_X1 U4944 ( .A1(n5263), .A2(n4976), .ZN(n5304) );
  AND3_X1 U4945 ( .A1(n4564), .A2(n4334), .A3(n4563), .ZN(n5888) );
  NAND3_X1 U4946 ( .A1(n4564), .A2(n4334), .A3(n4562), .ZN(n6475) );
  AND3_X1 U4947 ( .A1(n4568), .A2(n4567), .A3(n5845), .ZN(n4563) );
  NOR2_X1 U4948 ( .A1(n5997), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6013) );
  INV_X4 U4949 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U4950 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4951) );
  NOR2_X1 U4951 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4950) );
  NOR2_X1 U4952 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4952) );
  INV_X1 U4953 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4844) );
  INV_X1 U4954 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6633) );
  NOR2_X2 U4955 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5021) );
  INV_X1 U4956 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5535) );
  INV_X1 U4957 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5284) );
  INV_X1 U4958 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U4959 ( .A1(n8618), .A2(n5653), .ZN(n8617) );
  INV_X1 U4960 ( .A(n4277), .ZN(n7770) );
  NAND2_X1 U4961 ( .A1(n4276), .A2(n4765), .ZN(n9579) );
  NAND2_X1 U4962 ( .A1(n4280), .A2(n4279), .ZN(n7489) );
  NAND2_X1 U4963 ( .A1(n7011), .A2(n7014), .ZN(n4279) );
  OR2_X1 U4964 ( .A1(n7011), .A2(n7014), .ZN(n4280) );
  NAND2_X1 U4965 ( .A1(n9577), .A2(n8545), .ZN(n8791) );
  INV_X1 U4966 ( .A(n4846), .ZN(n4281) );
  INV_X4 U4967 ( .A(n4281), .ZN(n4282) );
  NAND2_X1 U4968 ( .A1(n4601), .A2(n4598), .ZN(n4846) );
  BUF_X4 U4969 ( .A(n6012), .Z(n6408) );
  CLKBUF_X1 U4970 ( .A(n5051), .Z(n4283) );
  OR2_X2 U4971 ( .A1(n9283), .A2(n9446), .ZN(n9268) );
  NAND2_X1 U4972 ( .A1(n6877), .A2(n6581), .ZN(n4285) );
  AOI21_X1 U4973 ( .B1(n4729), .B2(n4887), .A(n4728), .ZN(n4726) );
  INV_X1 U4974 ( .A(n4892), .ZN(n4728) );
  OR2_X1 U4975 ( .A1(n8853), .A2(n8671), .ZN(n5751) );
  NOR2_X1 U4976 ( .A1(n9796), .A2(n4763), .ZN(n4761) );
  INV_X1 U4977 ( .A(n7554), .ZN(n4763) );
  NAND2_X1 U4978 ( .A1(n9182), .A2(n9044), .ZN(n4795) );
  NAND2_X1 U4979 ( .A1(n5369), .A2(n5368), .ZN(n4742) );
  OAI21_X1 U4980 ( .B1(n5350), .B2(n5349), .A(n4928), .ZN(n5369) );
  AOI21_X1 U4981 ( .B1(n4466), .B2(n4302), .A(n4465), .ZN(n4464) );
  NAND2_X1 U4982 ( .A1(n5898), .A2(n5899), .ZN(n6025) );
  NAND2_X1 U4983 ( .A1(n4525), .A2(n4524), .ZN(n4523) );
  AND2_X1 U4984 ( .A1(n5755), .A2(n5757), .ZN(n4524) );
  NAND2_X1 U4985 ( .A1(n4744), .A2(n4743), .ZN(n5755) );
  NAND2_X1 U4986 ( .A1(n4910), .A2(n4909), .ZN(n4913) );
  NAND2_X1 U4987 ( .A1(n4766), .A2(n4770), .ZN(n4767) );
  NAND2_X1 U4988 ( .A1(n7319), .A2(n7754), .ZN(n5683) );
  OR2_X1 U4989 ( .A1(n6220), .A2(n6221), .ZN(n6240) );
  XNOR2_X1 U4990 ( .A(n4679), .B(n6368), .ZN(n6053) );
  NAND2_X1 U4991 ( .A1(n4682), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U4992 ( .A1(n6343), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U4993 ( .A1(n7444), .A2(n6388), .ZN(n4682) );
  NAND2_X1 U4994 ( .A1(n8226), .A2(n4577), .ZN(n4575) );
  OR2_X1 U4995 ( .A1(n9462), .A2(n9329), .ZN(n8215) );
  NOR2_X1 U4996 ( .A1(n9465), .A2(n9354), .ZN(n8190) );
  OAI21_X1 U4997 ( .B1(n8208), .B2(n8207), .A(n8206), .ZN(n9369) );
  NAND2_X1 U4998 ( .A1(n6547), .A2(n6546), .ZN(n7994) );
  NAND2_X1 U4999 ( .A1(n6551), .A2(n9716), .ZN(n6547) );
  NAND2_X1 U5000 ( .A1(n6544), .A2(n9730), .ZN(n6553) );
  AND2_X1 U5001 ( .A1(n4568), .A2(n4567), .ZN(n4562) );
  NOR2_X1 U5002 ( .A1(n5847), .A2(n4820), .ZN(n4819) );
  NAND2_X1 U5003 ( .A1(n4821), .A2(n5890), .ZN(n4820) );
  INV_X1 U5004 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4821) );
  NAND2_X1 U5005 ( .A1(n5612), .A2(n5611), .ZN(n5622) );
  NAND2_X1 U5006 ( .A1(n5608), .A2(n5607), .ZN(n5612) );
  OAI21_X1 U5007 ( .B1(n5457), .B2(n5456), .A(n5455), .ZN(n5481) );
  NOR2_X1 U5008 ( .A1(n4565), .A2(n5997), .ZN(n4564) );
  INV_X1 U5009 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4566) );
  INV_X1 U5010 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5839) );
  INV_X1 U5011 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4804) );
  AND2_X1 U5012 ( .A1(n4933), .A2(n4932), .ZN(n5368) );
  NAND2_X1 U5013 ( .A1(n4923), .A2(n4922), .ZN(n5350) );
  NAND2_X1 U5014 ( .A1(n4719), .A2(n4723), .ZN(n4898) );
  AOI21_X1 U5015 ( .B1(n4726), .B2(n4727), .A(n4724), .ZN(n4723) );
  INV_X1 U5016 ( .A(n4836), .ZN(n4724) );
  AND2_X1 U5017 ( .A1(n8263), .A2(n4647), .ZN(n4646) );
  NAND2_X1 U5018 ( .A1(n8446), .A2(n5479), .ZN(n4647) );
  AND3_X1 U5019 ( .A1(n5392), .A2(n5391), .A3(n5390), .ZN(n8552) );
  INV_X1 U5020 ( .A(n5072), .ZN(n5467) );
  AND4_X1 U5021 ( .A1(n5301), .A2(n5300), .A3(n5299), .A4(n5298), .ZN(n8546)
         );
  INV_X1 U5022 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U5023 ( .A1(n5779), .A2(n5778), .ZN(n8575) );
  AND2_X1 U5024 ( .A1(n5521), .A2(n5520), .ZN(n8579) );
  AND2_X1 U5025 ( .A1(n8558), .A2(n5655), .ZN(n4636) );
  AOI21_X1 U5026 ( .B1(n4619), .B2(n4480), .A(n4617), .ZN(n4616) );
  INV_X1 U5027 ( .A(n4619), .ZN(n4618) );
  INV_X1 U5028 ( .A(n5751), .ZN(n4617) );
  OR2_X1 U5029 ( .A1(n8863), .A2(n8551), .ZN(n5744) );
  NAND2_X1 U5030 ( .A1(n4754), .A2(n4752), .ZN(n8732) );
  OR2_X1 U5031 ( .A1(n8547), .A2(n4753), .ZN(n4752) );
  AND2_X1 U5032 ( .A1(n8548), .A2(n4757), .ZN(n4753) );
  NAND2_X1 U5033 ( .A1(n8772), .A2(n8749), .ZN(n4757) );
  INV_X1 U5034 ( .A(n5097), .ZN(n5352) );
  NOR2_X1 U5035 ( .A1(n7307), .A2(n4764), .ZN(n4762) );
  INV_X1 U5036 ( .A(n7304), .ZN(n4764) );
  NAND2_X1 U5037 ( .A1(n6877), .A2(n6581), .ZN(n5097) );
  NAND2_X2 U5038 ( .A1(n5576), .A2(n5832), .ZN(n6877) );
  INV_X1 U5039 ( .A(n9029), .ZN(n4698) );
  NOR2_X1 U5040 ( .A1(n5934), .A2(n5933), .ZN(n6806) );
  AND2_X1 U5041 ( .A1(n9719), .A2(n6452), .ZN(n5933) );
  AND2_X1 U5042 ( .A1(n6497), .A2(n6496), .ZN(n9131) );
  NAND2_X1 U5043 ( .A1(n5941), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5945) );
  OR2_X1 U5044 ( .A1(n9141), .A2(n6491), .ZN(n6447) );
  NAND2_X1 U5045 ( .A1(n4786), .A2(n4794), .ZN(n4785) );
  INV_X1 U5046 ( .A(n4789), .ZN(n4786) );
  AOI21_X1 U5047 ( .B1(n4791), .B2(n4790), .A(n4323), .ZN(n4789) );
  NAND2_X1 U5048 ( .A1(n4791), .A2(n4794), .ZN(n4787) );
  OR2_X1 U5049 ( .A1(n9442), .A2(n9245), .ZN(n8220) );
  AOI22_X1 U5050 ( .A1(n9306), .A2(n8218), .B1(n8217), .B2(n8216), .ZN(n9274)
         );
  NOR2_X1 U5051 ( .A1(n9719), .A2(n6841), .ZN(n9716) );
  NAND2_X1 U5052 ( .A1(n6473), .A2(n5892), .ZN(n6513) );
  NOR2_X1 U5053 ( .A1(n7850), .A2(n7782), .ZN(n5892) );
  OR2_X1 U5054 ( .A1(n5895), .A2(n9517), .ZN(n5894) );
  OAI21_X1 U5055 ( .B1(n4282), .B2(n4445), .A(n4526), .ZN(n5018) );
  NAND2_X1 U5056 ( .A1(n4282), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4526) );
  INV_X1 U5057 ( .A(n7272), .ZN(n9885) );
  AOI21_X1 U5058 ( .B1(n4704), .B2(n4293), .A(n4360), .ZN(n4700) );
  NAND2_X1 U5059 ( .A1(n4704), .A2(n4703), .ZN(n4702) );
  OAI21_X1 U5060 ( .B1(n9109), .B2(n9108), .A(n4531), .ZN(n4530) );
  AOI21_X1 U5061 ( .B1(n9110), .B2(n9712), .A(n9704), .ZN(n4531) );
  NAND2_X1 U5062 ( .A1(n5669), .A2(n5668), .ZN(n4514) );
  AND2_X1 U5063 ( .A1(n5759), .A2(n4270), .ZN(n4521) );
  AND2_X1 U5064 ( .A1(n5819), .A2(n5758), .ZN(n4522) );
  NAND2_X1 U5065 ( .A1(n5778), .A2(n8473), .ZN(n4504) );
  NOR2_X1 U5066 ( .A1(n4428), .A2(n9332), .ZN(n4427) );
  NAND2_X1 U5067 ( .A1(n9307), .A2(n4429), .ZN(n4428) );
  NOR2_X1 U5068 ( .A1(n9315), .A2(n9349), .ZN(n4429) );
  INV_X1 U5069 ( .A(n9904), .ZN(n7552) );
  INV_X1 U5070 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5532) );
  OAI21_X1 U5071 ( .B1(n5622), .B2(n5621), .A(n5620), .ZN(n5638) );
  INV_X1 U5072 ( .A(n4834), .ZN(n4379) );
  NOR2_X1 U5073 ( .A1(n5150), .A2(n4385), .ZN(n4384) );
  INV_X1 U5074 ( .A(n4867), .ZN(n4385) );
  NAND2_X1 U5075 ( .A1(n5148), .A2(n5149), .ZN(n4406) );
  AND2_X1 U5076 ( .A1(n4663), .A2(n4301), .ZN(n4658) );
  INV_X1 U5077 ( .A(n5049), .ZN(n5444) );
  AND2_X1 U5078 ( .A1(n5795), .A2(n4739), .ZN(n4737) );
  NOR2_X1 U5079 ( .A1(n5824), .A2(n5790), .ZN(n4740) );
  NOR2_X1 U5080 ( .A1(n5791), .A2(n4270), .ZN(n4738) );
  NOR2_X1 U5081 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4771) );
  NOR2_X1 U5082 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4652) );
  INV_X1 U5083 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5229) );
  INV_X1 U5084 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n4954) );
  OR2_X1 U5085 ( .A1(n8822), .A2(n8579), .ZN(n5773) );
  NOR2_X1 U5086 ( .A1(n5653), .A2(n5761), .ZN(n4629) );
  OR2_X1 U5087 ( .A1(n8842), .A2(n8672), .ZN(n5756) );
  AND2_X1 U5088 ( .A1(n8707), .A2(n5744), .ZN(n4622) );
  NOR2_X1 U5089 ( .A1(n8869), .A2(n8875), .ZN(n4494) );
  INV_X1 U5090 ( .A(n8760), .ZN(n4607) );
  AND2_X1 U5091 ( .A1(n8755), .A2(n8477), .ZN(n5798) );
  NOR2_X1 U5092 ( .A1(n8760), .A2(n4760), .ZN(n4756) );
  NOR2_X1 U5093 ( .A1(n8338), .A2(n8894), .ZN(n4481) );
  OR2_X1 U5094 ( .A1(n5180), .A2(n5179), .ZN(n5200) );
  OR2_X1 U5095 ( .A1(n9928), .A2(n7691), .ZN(n5697) );
  NAND2_X1 U5096 ( .A1(n5565), .A2(n9823), .ZN(n7017) );
  AND2_X1 U5097 ( .A1(n5551), .A2(n9833), .ZN(n7259) );
  OAI21_X1 U5098 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n5541), .A(n9867), .ZN(n7255)
         );
  INV_X1 U5099 ( .A(n7722), .ZN(n4376) );
  NAND2_X1 U5100 ( .A1(n8225), .A2(n4422), .ZN(n4421) );
  NOR2_X1 U5101 ( .A1(n9216), .A2(n4423), .ZN(n4422) );
  INV_X1 U5102 ( .A(n9255), .ZN(n4424) );
  MUX2_X1 U5103 ( .A(n8163), .B(n8059), .S(n8158), .Z(n8165) );
  NAND2_X1 U5104 ( .A1(n4440), .A2(n8201), .ZN(n4439) );
  OR2_X1 U5105 ( .A1(n9396), .A2(n9131), .ZN(n8159) );
  NOR2_X1 U5106 ( .A1(n9153), .A2(n8230), .ZN(n9127) );
  OR2_X1 U5107 ( .A1(n9401), .A2(n9152), .ZN(n8152) );
  OAI21_X1 U5108 ( .B1(n4785), .B2(n4570), .A(n4287), .ZN(n4784) );
  OR2_X1 U5109 ( .A1(n9405), .A2(n9130), .ZN(n8149) );
  NAND2_X1 U5110 ( .A1(n9410), .A2(n9186), .ZN(n4794) );
  NAND2_X1 U5111 ( .A1(n4597), .A2(n8222), .ZN(n4596) );
  NOR2_X1 U5112 ( .A1(n9242), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U5113 ( .A1(n8221), .A2(n8220), .ZN(n4592) );
  NOR2_X1 U5114 ( .A1(n9242), .A2(n4594), .ZN(n4593) );
  INV_X1 U5115 ( .A(n8220), .ZN(n4594) );
  OR2_X1 U5116 ( .A1(n9437), .A2(n9259), .ZN(n8123) );
  NOR2_X1 U5117 ( .A1(n9359), .A2(n9465), .ZN(n4450) );
  INV_X1 U5118 ( .A(n8209), .ZN(n4586) );
  AOI21_X1 U5119 ( .B1(n9368), .B2(n4585), .A(n4583), .ZN(n4582) );
  INV_X1 U5120 ( .A(n8210), .ZN(n4583) );
  NAND2_X1 U5121 ( .A1(n4313), .A2(n7730), .ZN(n4781) );
  NAND2_X1 U5122 ( .A1(n7733), .A2(n8078), .ZN(n8208) );
  NAND2_X1 U5123 ( .A1(n7405), .A2(n9047), .ZN(n8071) );
  AND2_X1 U5124 ( .A1(n7244), .A2(n9204), .ZN(n6483) );
  NAND2_X1 U5125 ( .A1(n9718), .A2(n4837), .ZN(n9717) );
  NAND2_X1 U5126 ( .A1(n4282), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n4390) );
  XNOR2_X1 U5127 ( .A(n5638), .B(n5637), .ZN(n5635) );
  NAND2_X1 U5128 ( .A1(n5507), .A2(n5506), .ZN(n5608) );
  NAND2_X1 U5129 ( .A1(n5505), .A2(n5504), .ZN(n5507) );
  OAI21_X1 U5130 ( .B1(n5316), .B2(n4919), .A(n4918), .ZN(n5333) );
  INV_X1 U5131 ( .A(n4902), .ZN(n4468) );
  INV_X1 U5132 ( .A(n4467), .ZN(n4466) );
  OAI21_X1 U5133 ( .B1(n4470), .B2(n4302), .A(n4907), .ZN(n4467) );
  NAND2_X1 U5134 ( .A1(n4894), .A2(n4893), .ZN(n4897) );
  INV_X1 U5135 ( .A(n4726), .ZN(n4725) );
  INV_X1 U5136 ( .A(n4886), .ZN(n4730) );
  AOI21_X1 U5137 ( .B1(n5133), .B2(n4384), .A(n4382), .ZN(n4381) );
  INV_X1 U5138 ( .A(n4872), .ZN(n4382) );
  INV_X1 U5139 ( .A(n4384), .ZN(n4383) );
  INV_X1 U5140 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U5141 ( .A1(n4599), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4598) );
  INV_X1 U5142 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4600) );
  OAI21_X1 U5143 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n4844), .ZN(n4601) );
  AND2_X1 U5144 ( .A1(n5503), .A2(n5501), .ZN(n8263) );
  NOR2_X1 U5145 ( .A1(n5502), .A2(n5454), .ZN(n4648) );
  NOR2_X1 U5146 ( .A1(n7245), .A2(n4405), .ZN(n4404) );
  INV_X1 U5147 ( .A(n5132), .ZN(n4405) );
  INV_X1 U5148 ( .A(n4409), .ZN(n4408) );
  OAI21_X1 U5149 ( .B1(n4655), .B2(n4288), .A(n8422), .ZN(n4409) );
  NOR2_X1 U5150 ( .A1(n8380), .A2(n4664), .ZN(n4663) );
  INV_X1 U5151 ( .A(n5081), .ZN(n4664) );
  NAND2_X1 U5152 ( .A1(n5001), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U5153 ( .A1(n7232), .A2(n4400), .ZN(n4399) );
  NOR2_X1 U5154 ( .A1(n4401), .A2(n4403), .ZN(n4400) );
  INV_X1 U5155 ( .A(n7233), .ZN(n4401) );
  AND2_X1 U5156 ( .A1(n5382), .A2(n5367), .ZN(n4654) );
  INV_X1 U5157 ( .A(n8396), .ZN(n5382) );
  OR2_X1 U5158 ( .A1(n5200), .A2(n5199), .ZN(n5214) );
  INV_X1 U5159 ( .A(n5191), .ZN(n4657) );
  AOI21_X1 U5160 ( .B1(n4655), .B2(n7686), .A(n4288), .ZN(n4411) );
  OR2_X1 U5161 ( .A1(n6032), .A2(n5046), .ZN(n4628) );
  OAI21_X1 U5162 ( .B1(n5647), .B2(n4456), .A(n5823), .ZN(n5648) );
  AOI21_X1 U5163 ( .B1(n5616), .B2(n4454), .A(n4362), .ZN(n4456) );
  AND4_X1 U5164 ( .A1(n5147), .A2(n5146), .A3(n5145), .A4(n5144), .ZN(n7553)
         );
  XNOR2_X1 U5165 ( .A(n6978), .B(n4548), .ZN(n6967) );
  AOI21_X1 U5166 ( .B1(n6988), .B2(n6960), .A(n6959), .ZN(n6958) );
  NOR2_X1 U5167 ( .A1(n7122), .A2(n4547), .ZN(n7125) );
  AND2_X1 U5168 ( .A1(n7128), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4547) );
  NOR2_X1 U5169 ( .A1(n7888), .A2(n7887), .ZN(n7910) );
  NOR2_X1 U5170 ( .A1(n8511), .A2(n4538), .ZN(n8521) );
  AND2_X1 U5171 ( .A1(n7924), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4538) );
  NAND2_X1 U5172 ( .A1(n5615), .A2(n5614), .ZN(n8818) );
  AOI21_X1 U5173 ( .B1(n8607), .B2(n5072), .A(n5495), .ZN(n8588) );
  XNOR2_X1 U5174 ( .A(n8828), .B(n8588), .ZN(n8610) );
  AND2_X1 U5175 ( .A1(n5452), .A2(n5451), .ZN(n8659) );
  NOR2_X1 U5176 ( .A1(n8554), .A2(n4621), .ZN(n4619) );
  NAND2_X1 U5177 ( .A1(n8723), .A2(n4622), .ZN(n4620) );
  INV_X1 U5178 ( .A(n8554), .ZN(n8693) );
  INV_X1 U5179 ( .A(n5722), .ZN(n4612) );
  AND2_X1 U5180 ( .A1(n5729), .A2(n5732), .ZN(n8760) );
  NAND2_X1 U5181 ( .A1(n8775), .A2(n4756), .ZN(n4758) );
  INV_X1 U5182 ( .A(n8797), .ZN(n4614) );
  INV_X1 U5183 ( .A(n8798), .ZN(n4615) );
  NOR2_X1 U5184 ( .A1(n9578), .A2(n5714), .ZN(n4630) );
  NAND2_X1 U5185 ( .A1(n4767), .A2(n4769), .ZN(n4765) );
  INV_X1 U5186 ( .A(n4767), .ZN(n4768) );
  NAND2_X1 U5187 ( .A1(n7772), .A2(n7771), .ZN(n7822) );
  AND2_X1 U5188 ( .A1(n6873), .A2(n5576), .ZN(n8801) );
  INV_X1 U5189 ( .A(n8801), .ZN(n8765) );
  INV_X1 U5190 ( .A(n8817), .ZN(n4635) );
  NAND2_X1 U5191 ( .A1(n8818), .A2(n9929), .ZN(n4634) );
  NAND2_X1 U5192 ( .A1(n5443), .A2(n5442), .ZN(n8838) );
  INV_X1 U5193 ( .A(n8755), .ZN(n8875) );
  OAI21_X1 U5194 ( .B1(n6877), .B2(n6898), .A(n5098), .ZN(n4528) );
  NAND2_X1 U5195 ( .A1(n9799), .A2(n9931), .ZN(n9947) );
  NOR2_X1 U5196 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4967) );
  AND2_X1 U5197 ( .A1(n4772), .A2(n4966), .ZN(n4490) );
  NAND2_X1 U5198 ( .A1(n4981), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5533) );
  AND2_X1 U5199 ( .A1(n4958), .A2(n4668), .ZN(n4667) );
  NAND2_X1 U5200 ( .A1(n5304), .A2(n4977), .ZN(n5283) );
  NAND2_X1 U5201 ( .A1(n5528), .A2(n4552), .ZN(n4551) );
  INV_X1 U5202 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4552) );
  NAND2_X1 U5203 ( .A1(n6223), .A2(n6224), .ZN(n7854) );
  NAND2_X1 U5204 ( .A1(n7529), .A2(n6130), .ZN(n6217) );
  NAND2_X1 U5205 ( .A1(n6435), .A2(n4677), .ZN(n4676) );
  INV_X1 U5206 ( .A(n6413), .ZN(n4677) );
  XNOR2_X1 U5207 ( .A(n6200), .B(n6368), .ZN(n6205) );
  NAND2_X1 U5208 ( .A1(n4689), .A2(n4691), .ZN(n4688) );
  INV_X1 U5209 ( .A(n7494), .ZN(n4689) );
  INV_X1 U5210 ( .A(n6130), .ZN(n4687) );
  NOR2_X1 U5211 ( .A1(n4687), .A2(n6111), .ZN(n4685) );
  OR2_X1 U5212 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  AND2_X1 U5213 ( .A1(n6405), .A2(n6404), .ZN(n8198) );
  OR2_X1 U5214 ( .A1(n9020), .A2(n6491), .ZN(n6405) );
  NOR2_X1 U5215 ( .A1(n9655), .A2(n4511), .ZN(n4510) );
  AND2_X1 U5216 ( .A1(n9638), .A2(n4299), .ZN(n4511) );
  OR2_X1 U5217 ( .A1(n6780), .A2(n6779), .ZN(n4500) );
  NAND2_X1 U5218 ( .A1(n4500), .A2(n4499), .ZN(n9676) );
  OR2_X1 U5219 ( .A1(n6786), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4499) );
  NOR2_X1 U5220 ( .A1(n6857), .A2(n4349), .ZN(n9691) );
  OR2_X1 U5221 ( .A1(n9691), .A2(n9690), .ZN(n4498) );
  NOR2_X1 U5222 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5861) );
  OR2_X1 U5223 ( .A1(n9069), .A2(n9068), .ZN(n4518) );
  INV_X1 U5224 ( .A(n4438), .ZN(n4434) );
  NOR2_X1 U5225 ( .A1(n9118), .A2(n4439), .ZN(n4438) );
  NAND2_X1 U5226 ( .A1(n8159), .A2(n8160), .ZN(n8232) );
  NAND2_X1 U5227 ( .A1(n4572), .A2(n4574), .ZN(n4571) );
  AOI21_X1 U5228 ( .B1(n4574), .B2(n8227), .A(n7950), .ZN(n4573) );
  AND2_X1 U5229 ( .A1(n4571), .A2(n4569), .ZN(n9153) );
  AND2_X1 U5230 ( .A1(n4573), .A2(n4570), .ZN(n4569) );
  AND2_X1 U5231 ( .A1(n4795), .A2(n4796), .ZN(n4792) );
  NAND2_X1 U5232 ( .A1(n4796), .A2(n4309), .ZN(n4793) );
  NAND2_X1 U5233 ( .A1(n9192), .A2(n8957), .ZN(n4796) );
  OR2_X1 U5234 ( .A1(n9256), .A2(n8221), .ZN(n4595) );
  AOI21_X1 U5235 ( .B1(n9316), .B2(n8215), .A(n8214), .ZN(n9306) );
  NAND2_X1 U5236 ( .A1(n9462), .A2(n9308), .ZN(n4816) );
  INV_X1 U5237 ( .A(n9294), .ZN(n9320) );
  NAND2_X1 U5238 ( .A1(n4806), .A2(n4805), .ZN(n9314) );
  INV_X1 U5239 ( .A(n4808), .ZN(n4805) );
  OR2_X1 U5240 ( .A1(n4815), .A2(n8190), .ZN(n4806) );
  AOI21_X1 U5241 ( .B1(n7731), .B2(n4778), .A(n4774), .ZN(n4773) );
  NAND2_X1 U5242 ( .A1(n4775), .A2(n8185), .ZN(n4774) );
  INV_X1 U5243 ( .A(n7786), .ZN(n4780) );
  INV_X1 U5244 ( .A(n4781), .ZN(n4777) );
  INV_X1 U5245 ( .A(n4799), .ZN(n4798) );
  OAI21_X1 U5246 ( .B1(n4306), .B2(n4801), .A(n4800), .ZN(n4799) );
  OR2_X1 U5247 ( .A1(n9486), .A2(n9546), .ZN(n4800) );
  NAND2_X1 U5248 ( .A1(n4441), .A2(n7405), .ZN(n7401) );
  INV_X1 U5249 ( .A(n7442), .ZN(n4441) );
  AND2_X1 U5250 ( .A1(n7378), .A2(n7377), .ZN(n7439) );
  NAND2_X1 U5251 ( .A1(n7160), .A2(n7999), .ZN(n7371) );
  NAND2_X1 U5252 ( .A1(n4554), .A2(n4553), .ZN(n7160) );
  AND4_X1 U5253 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n7101)
         );
  AND2_X1 U5254 ( .A1(n4282), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4443) );
  OR2_X1 U5255 ( .A1(n6544), .A2(n9730), .ZN(n6545) );
  INV_X1 U5256 ( .A(n9328), .ZN(n9721) );
  NAND2_X1 U5257 ( .A1(n6485), .A2(n9515), .ZN(n6834) );
  NAND2_X1 U5258 ( .A1(n6461), .A2(n6473), .ZN(n6734) );
  XNOR2_X1 U5259 ( .A(n6476), .B(n6701), .ZN(n6512) );
  INV_X1 U5260 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4817) );
  XNOR2_X1 U5261 ( .A(n5883), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U5262 ( .A1(n5887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U5263 ( .A1(n4937), .A2(n4936), .ZN(n5398) );
  XNOR2_X1 U5264 ( .A(n5398), .B(n5397), .ZN(n7462) );
  NAND2_X1 U5265 ( .A1(n4469), .A2(n4902), .ZN(n5303) );
  NAND2_X1 U5266 ( .A1(n4898), .A2(n4470), .ZN(n4469) );
  AOI21_X1 U5267 ( .B1(n5112), .B2(n4294), .A(n4330), .ZN(n4717) );
  NAND2_X1 U5268 ( .A1(n4624), .A2(n4459), .ZN(n4623) );
  INV_X1 U5269 ( .A(n4857), .ZN(n4461) );
  NAND2_X1 U5270 ( .A1(n4670), .A2(n4857), .ZN(n5084) );
  NAND2_X1 U5271 ( .A1(n5415), .A2(n5414), .ZN(n8848) );
  AOI21_X1 U5272 ( .B1(n4642), .B2(n4645), .A(n4354), .ZN(n4640) );
  AND4_X1 U5273 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n8335)
         );
  AND4_X1 U5274 ( .A1(n5256), .A2(n5255), .A3(n5254), .A4(n5253), .ZN(n8480)
         );
  NAND2_X1 U5275 ( .A1(n5288), .A2(n5287), .ZN(n8884) );
  AND4_X1 U5276 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n8763)
         );
  INV_X1 U5277 ( .A(n8469), .ZN(n8458) );
  AND2_X1 U5278 ( .A1(n5473), .A2(n5472), .ZN(n8563) );
  OR2_X1 U5279 ( .A1(n8626), .A2(n5467), .ZN(n5473) );
  INV_X1 U5280 ( .A(n8659), .ZN(n8561) );
  AND3_X1 U5281 ( .A1(n5377), .A2(n5376), .A3(n5375), .ZN(n8551) );
  AND4_X1 U5282 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n8749)
         );
  NAND2_X1 U5283 ( .A1(n4300), .A2(n5126), .ZN(n8487) );
  NAND2_X1 U5284 ( .A1(n6936), .A2(n6935), .ZN(n6934) );
  NAND2_X1 U5285 ( .A1(n8494), .A2(n4539), .ZN(n8513) );
  NAND2_X1 U5286 ( .A1(n4541), .A2(n4540), .ZN(n4539) );
  INV_X1 U5287 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n4540) );
  INV_X1 U5288 ( .A(n8503), .ZN(n4541) );
  NAND2_X1 U5289 ( .A1(n6893), .A2(n6892), .ZN(n9788) );
  AND2_X1 U5290 ( .A1(n6893), .A2(n5576), .ZN(n8529) );
  NAND2_X1 U5291 ( .A1(n4631), .A2(n8581), .ZN(n8816) );
  NAND2_X1 U5292 ( .A1(n4632), .A2(n9803), .ZN(n4631) );
  NAND2_X1 U5293 ( .A1(n6877), .A2(n4489), .ZN(n4488) );
  OAI21_X1 U5294 ( .B1(n6583), .B2(n6581), .A(n4331), .ZN(n4489) );
  NAND2_X1 U5295 ( .A1(n6413), .A2(n9018), .ZN(n4367) );
  OAI21_X1 U5296 ( .B1(n8922), .B2(n4355), .A(n8928), .ZN(n4370) );
  OAI21_X1 U5297 ( .B1(n9007), .B2(n4707), .A(n4699), .ZN(n8937) );
  INV_X1 U5298 ( .A(n4701), .ZN(n4699) );
  NAND2_X1 U5299 ( .A1(n4675), .A2(n4676), .ZN(n8924) );
  NAND2_X1 U5300 ( .A1(n4697), .A2(n4841), .ZN(n4695) );
  NAND2_X1 U5301 ( .A1(n5871), .A2(n5870), .ZN(n9455) );
  NAND2_X1 U5302 ( .A1(n6301), .A2(n6300), .ZN(n9442) );
  OR2_X1 U5303 ( .A1(n6032), .A2(n6067), .ZN(n4683) );
  NAND2_X1 U5304 ( .A1(n4415), .A2(n4414), .ZN(n4413) );
  AOI21_X1 U5305 ( .B1(n8057), .B2(n4417), .A(n4416), .ZN(n4415) );
  OR2_X1 U5306 ( .A1(n8169), .A2(n9204), .ZN(n4414) );
  NAND2_X1 U5307 ( .A1(n8176), .A2(n7244), .ZN(n4412) );
  INV_X1 U5308 ( .A(n9329), .ZN(n9308) );
  INV_X1 U5309 ( .A(n7373), .ZN(n9046) );
  NAND4_X1 U5310 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(n9719)
         );
  OR2_X1 U5311 ( .A1(n6025), .A2(n5928), .ZN(n5931) );
  NOR2_X1 U5312 ( .A1(n9678), .A2(n6524), .ZN(n6857) );
  AND2_X1 U5313 ( .A1(n6123), .A2(n6133), .ZN(n9695) );
  AND2_X1 U5314 ( .A1(n6537), .A2(n6536), .ZN(n9712) );
  NOR2_X1 U5315 ( .A1(n9112), .A2(n4844), .ZN(n4533) );
  AND2_X1 U5316 ( .A1(n6393), .A2(n6392), .ZN(n9167) );
  OR2_X1 U5317 ( .A1(n9767), .A2(n6568), .ZN(n9142) );
  INV_X1 U5318 ( .A(n4746), .ZN(n5660) );
  NAND2_X1 U5319 ( .A1(n5656), .A2(n5790), .ZN(n4515) );
  NAND2_X1 U5320 ( .A1(n7312), .A2(n4270), .ZN(n4516) );
  NAND2_X1 U5321 ( .A1(n5756), .A2(n4745), .ZN(n4744) );
  AOI21_X1 U5322 ( .B1(n8675), .B2(n8695), .A(n4270), .ZN(n4745) );
  NAND2_X1 U5323 ( .A1(n5655), .A2(n4270), .ZN(n4743) );
  AOI21_X1 U5324 ( .B1(n4523), .B2(n4522), .A(n4521), .ZN(n5764) );
  OR2_X1 U5325 ( .A1(n5646), .A2(n8536), .ZN(n5792) );
  INV_X1 U5326 ( .A(n4502), .ZN(n4501) );
  OAI21_X1 U5327 ( .B1(n4503), .B2(n5778), .A(n4270), .ZN(n4502) );
  NAND2_X1 U5328 ( .A1(n5779), .A2(n4504), .ZN(n4503) );
  INV_X1 U5329 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U5330 ( .A1(n8487), .A2(n9900), .ZN(n5678) );
  NAND2_X1 U5331 ( .A1(n7874), .A2(n7871), .ZN(n4394) );
  INV_X1 U5332 ( .A(n7873), .ZN(n6210) );
  INV_X1 U5333 ( .A(n8997), .ZN(n4393) );
  NOR2_X1 U5334 ( .A1(n9242), .A2(n4327), .ZN(n4425) );
  OAI21_X1 U5335 ( .B1(n4282), .B2(n4389), .A(n4388), .ZN(n5637) );
  NAND2_X1 U5336 ( .A1(n4282), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n4388) );
  INV_X1 U5337 ( .A(n4942), .ZN(n4712) );
  INV_X1 U5338 ( .A(n5281), .ZN(n4465) );
  NOR2_X1 U5339 ( .A1(n4725), .A2(n4721), .ZN(n4720) );
  INV_X1 U5340 ( .A(n4882), .ZN(n4721) );
  NOR2_X1 U5341 ( .A1(n5789), .A2(n4455), .ZN(n4454) );
  INV_X1 U5342 ( .A(n5779), .ZN(n4455) );
  NAND2_X1 U5343 ( .A1(n7890), .A2(n4536), .ZN(n7920) );
  OR2_X1 U5344 ( .A1(n7891), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4536) );
  NAND2_X1 U5345 ( .A1(n8818), .A2(n8587), .ZN(n5778) );
  OR2_X1 U5346 ( .A1(n8818), .A2(n8587), .ZN(n5779) );
  AND2_X1 U5347 ( .A1(n4485), .A2(n4486), .ZN(n4484) );
  NOR2_X1 U5348 ( .A1(n8838), .A2(n8842), .ZN(n4486) );
  INV_X1 U5349 ( .A(n4622), .ZN(n4480) );
  NAND2_X1 U5350 ( .A1(n8720), .A2(n4494), .ZN(n4493) );
  INV_X1 U5351 ( .A(n8547), .ZN(n4755) );
  OR2_X1 U5352 ( .A1(n5295), .A2(n5294), .ZN(n5297) );
  NAND2_X1 U5353 ( .A1(n8894), .A2(n8544), .ZN(n4769) );
  NOR2_X1 U5354 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4772) );
  NAND2_X1 U5355 ( .A1(n5534), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5556) );
  AND2_X1 U5356 ( .A1(n4977), .A2(n4669), .ZN(n4668) );
  INV_X1 U5357 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4669) );
  AND2_X1 U5358 ( .A1(n4771), .A2(n5066), .ZN(n4653) );
  AND2_X1 U5359 ( .A1(n6371), .A2(n6370), .ZN(n6373) );
  NAND2_X1 U5360 ( .A1(n6499), .A2(n6513), .ZN(n5935) );
  NOR2_X1 U5361 ( .A1(n7352), .A2(n4672), .ZN(n4671) );
  INV_X1 U5362 ( .A(n6056), .ZN(n4672) );
  INV_X1 U5363 ( .A(n5935), .ZN(n5919) );
  NAND2_X1 U5364 ( .A1(n9735), .A2(n6513), .ZN(n6012) );
  INV_X1 U5365 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5846) );
  OR2_X1 U5366 ( .A1(n5852), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5847) );
  NOR2_X1 U5367 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5862) );
  AND2_X1 U5368 ( .A1(n4507), .A2(n4506), .ZN(n7618) );
  NAND2_X1 U5369 ( .A1(n7283), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4506) );
  INV_X1 U5370 ( .A(n4792), .ZN(n4790) );
  OR2_X1 U5371 ( .A1(n9421), .A2(n8957), .ZN(n8137) );
  NOR2_X1 U5372 ( .A1(n9430), .A2(n9437), .ZN(n4453) );
  AND2_X1 U5373 ( .A1(n9446), .A2(n9258), .ZN(n8019) );
  INV_X1 U5374 ( .A(n8190), .ZN(n4810) );
  NOR2_X1 U5375 ( .A1(n4814), .A2(n8191), .ZN(n4813) );
  NOR2_X1 U5376 ( .A1(n9342), .A2(n9319), .ZN(n4808) );
  NAND2_X1 U5377 ( .A1(n5906), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6232) );
  AND2_X1 U5378 ( .A1(n8183), .A2(n4779), .ZN(n4778) );
  NAND2_X1 U5379 ( .A1(n4781), .A2(n7786), .ZN(n4779) );
  NAND2_X1 U5380 ( .A1(n4778), .A2(n4780), .ZN(n4775) );
  NAND2_X1 U5381 ( .A1(n4588), .A2(n4587), .ZN(n9371) );
  INV_X1 U5382 ( .A(n9369), .ZN(n4588) );
  OR2_X1 U5383 ( .A1(n7728), .A2(n4802), .ZN(n4801) );
  INV_X1 U5384 ( .A(n7501), .ZN(n4802) );
  NAND2_X1 U5385 ( .A1(n4561), .A2(n4560), .ZN(n7372) );
  AOI21_X1 U5386 ( .B1(n8000), .B2(n7395), .A(n8069), .ZN(n4560) );
  NOR2_X1 U5387 ( .A1(n7163), .A2(n7199), .ZN(n7164) );
  NOR2_X1 U5388 ( .A1(n8075), .A2(n8076), .ZN(n4559) );
  AND2_X1 U5389 ( .A1(n5506), .A2(n5488), .ZN(n5504) );
  AND2_X1 U5390 ( .A1(n5482), .A2(n5461), .ZN(n5480) );
  OAI21_X1 U5391 ( .B1(n5437), .B2(n5436), .A(n5435), .ZN(n5457) );
  AND2_X1 U5392 ( .A1(n5844), .A2(n5842), .ZN(n4567) );
  AND2_X1 U5393 ( .A1(n5841), .A2(n5843), .ZN(n4568) );
  OAI21_X1 U5394 ( .B1(n5398), .B2(n4709), .A(n4710), .ZN(n5437) );
  AOI21_X1 U5395 ( .B1(n5413), .B2(n4712), .A(n4711), .ZN(n4710) );
  NAND2_X1 U5396 ( .A1(n5413), .A2(n4713), .ZN(n4709) );
  INV_X1 U5397 ( .A(n4948), .ZN(n4711) );
  NOR2_X1 U5398 ( .A1(n4899), .A2(n4471), .ZN(n4470) );
  INV_X1 U5399 ( .A(n4897), .ZN(n4471) );
  NAND2_X1 U5400 ( .A1(n4380), .A2(n4378), .ZN(n4476) );
  AND2_X1 U5401 ( .A1(n4882), .A2(n4881), .ZN(n4832) );
  INV_X1 U5402 ( .A(n5112), .ZN(n4718) );
  INV_X1 U5403 ( .A(n5095), .ZN(n4716) );
  INV_X1 U5404 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5837) );
  AND2_X1 U5405 ( .A1(n5837), .A2(n5838), .ZN(n4803) );
  INV_X1 U5406 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5838) );
  INV_X1 U5407 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4432) );
  INV_X1 U5408 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4430) );
  OAI21_X1 U5409 ( .B1(n4282), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n4387), .ZN(
        n4855) );
  NAND2_X1 U5410 ( .A1(n4282), .A2(n6577), .ZN(n4387) );
  AOI21_X1 U5411 ( .B1(n4646), .B2(n4644), .A(n4643), .ZN(n4642) );
  INV_X1 U5412 ( .A(n5503), .ZN(n4643) );
  INV_X1 U5413 ( .A(n4648), .ZN(n4644) );
  INV_X1 U5414 ( .A(n4646), .ZN(n4645) );
  INV_X1 U5415 ( .A(n4406), .ZN(n4403) );
  OR2_X1 U5416 ( .A1(n5428), .A2(n8475), .ZN(n5425) );
  NOR2_X1 U5417 ( .A1(n5308), .A2(n4666), .ZN(n4665) );
  INV_X1 U5418 ( .A(n5280), .ZN(n4666) );
  NAND2_X1 U5419 ( .A1(n8400), .A2(n5276), .ZN(n8281) );
  NAND2_X1 U5420 ( .A1(n5000), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5419) );
  INV_X1 U5421 ( .A(n5417), .ZN(n5000) );
  NAND2_X1 U5422 ( .A1(n8298), .A2(n5081), .ZN(n8381) );
  NAND2_X1 U5423 ( .A1(n4397), .A2(n4406), .ZN(n4396) );
  NAND2_X1 U5424 ( .A1(n5190), .A2(n5189), .ZN(n7684) );
  NAND2_X1 U5425 ( .A1(n4999), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5388) );
  OR2_X1 U5426 ( .A1(n5388), .A2(n8324), .ZN(n5400) );
  OR2_X1 U5427 ( .A1(n5400), .A2(n8415), .ZN(n5417) );
  NAND2_X1 U5428 ( .A1(n4994), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5235) );
  INV_X1 U5429 ( .A(n5214), .ZN(n4994) );
  INV_X1 U5430 ( .A(n8247), .ZN(n5061) );
  NAND2_X1 U5431 ( .A1(n4661), .A2(n4301), .ZN(n4660) );
  NAND2_X1 U5432 ( .A1(n5110), .A2(n8379), .ZN(n4661) );
  NAND2_X1 U5433 ( .A1(n7232), .A2(n7233), .ZN(n7231) );
  NAND2_X1 U5434 ( .A1(n8281), .A2(n5280), .ZN(n8350) );
  INV_X1 U5435 ( .A(n7017), .ZN(n5826) );
  AND4_X1 U5436 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n7830)
         );
  NAND2_X1 U5437 ( .A1(n5052), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5053) );
  NOR2_X1 U5438 ( .A1(n6953), .A2(n4543), .ZN(n6942) );
  AND2_X1 U5439 ( .A1(n6887), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4543) );
  NOR2_X1 U5440 ( .A1(n6942), .A2(n6941), .ZN(n6940) );
  NOR2_X1 U5441 ( .A1(n7125), .A2(n7124), .ZN(n7340) );
  NOR2_X1 U5442 ( .A1(n7340), .A2(n4546), .ZN(n7344) );
  AND2_X1 U5443 ( .A1(n7341), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4546) );
  NOR2_X1 U5444 ( .A1(n7344), .A2(n7343), .ZN(n7472) );
  NAND2_X1 U5445 ( .A1(n7811), .A2(n4537), .ZN(n7815) );
  OR2_X1 U5446 ( .A1(n7812), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4537) );
  NAND2_X1 U5447 ( .A1(n7815), .A2(n7814), .ZN(n7890) );
  AND3_X1 U5448 ( .A1(n4952), .A2(n4950), .A3(n4652), .ZN(n4651) );
  AND2_X1 U5449 ( .A1(n4951), .A2(n5021), .ZN(n4650) );
  XNOR2_X1 U5450 ( .A(n7920), .B(n7921), .ZN(n7892) );
  AOI21_X1 U5451 ( .B1(n8521), .B2(n8522), .A(n7925), .ZN(n7926) );
  AND2_X1 U5452 ( .A1(n8570), .A2(n8595), .ZN(n8568) );
  AND2_X1 U5453 ( .A1(n8606), .A2(n8599), .ZN(n8595) );
  INV_X1 U5454 ( .A(n4473), .ZN(n4472) );
  AND2_X1 U5455 ( .A1(n8677), .A2(n4482), .ZN(n8606) );
  NOR2_X1 U5456 ( .A1(n8828), .A2(n4483), .ZN(n4482) );
  INV_X1 U5457 ( .A(n4484), .ZN(n4483) );
  OR2_X1 U5458 ( .A1(n8838), .A2(n8561), .ZN(n8562) );
  NAND2_X1 U5459 ( .A1(n8677), .A2(n4486), .ZN(n8634) );
  NAND2_X1 U5460 ( .A1(n8677), .A2(n8655), .ZN(n8649) );
  AND2_X1 U5461 ( .A1(n5017), .A2(n5016), .ZN(n8672) );
  AND2_X1 U5462 ( .A1(n5407), .A2(n5406), .ZN(n8671) );
  AND2_X1 U5463 ( .A1(n8687), .A2(n8675), .ZN(n8677) );
  INV_X1 U5464 ( .A(n4750), .ZN(n4748) );
  OAI21_X1 U5465 ( .B1(n4751), .B2(n4829), .A(n4326), .ZN(n4750) );
  INV_X1 U5466 ( .A(n8553), .ZN(n4751) );
  NOR2_X1 U5467 ( .A1(n8766), .A2(n4492), .ZN(n8733) );
  INV_X1 U5468 ( .A(n4494), .ZN(n4492) );
  AND2_X1 U5469 ( .A1(n5740), .A2(n8722), .ZN(n8739) );
  NAND2_X1 U5470 ( .A1(n4998), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5356) );
  INV_X1 U5471 ( .A(n5338), .ZN(n4998) );
  AOI21_X1 U5472 ( .B1(n4606), .B2(n4609), .A(n5730), .ZN(n4603) );
  NAND2_X1 U5473 ( .A1(n4997), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5321) );
  INV_X1 U5474 ( .A(n5297), .ZN(n4997) );
  OR2_X1 U5475 ( .A1(n5321), .A2(n8363), .ZN(n5338) );
  AND2_X1 U5476 ( .A1(n7773), .A2(n4296), .ZN(n8792) );
  OR2_X1 U5477 ( .A1(n5251), .A2(n7706), .ZN(n5269) );
  NAND2_X1 U5478 ( .A1(n4996), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5295) );
  INV_X1 U5479 ( .A(n5269), .ZN(n4996) );
  NAND2_X1 U5480 ( .A1(n7773), .A2(n9942), .ZN(n7825) );
  AND2_X1 U5481 ( .A1(n7677), .A2(n9938), .ZN(n7773) );
  INV_X1 U5482 ( .A(n7563), .ZN(n7561) );
  OR2_X1 U5483 ( .A1(n9809), .A2(n7690), .ZN(n7678) );
  NOR2_X1 U5484 ( .A1(n7678), .A2(n9928), .ZN(n7677) );
  AND4_X1 U5485 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n7670)
         );
  AND2_X1 U5486 ( .A1(n7555), .A2(n7554), .ZN(n9798) );
  NAND2_X1 U5487 ( .A1(n5598), .A2(n4637), .ZN(n7321) );
  AND4_X1 U5488 ( .A1(n5165), .A2(n5164), .A3(n5163), .A4(n5162), .ZN(n7318)
         );
  NOR2_X1 U5489 ( .A1(n9890), .A2(n8301), .ZN(n7050) );
  AND2_X1 U5490 ( .A1(n9885), .A2(n9873), .ZN(n7271) );
  NAND2_X1 U5491 ( .A1(n5624), .A2(n5623), .ZN(n8811) );
  NAND2_X1 U5492 ( .A1(n5510), .A2(n5509), .ZN(n8822) );
  INV_X1 U5493 ( .A(n8706), .ZN(n8859) );
  NAND2_X1 U5494 ( .A1(n5320), .A2(n5319), .ZN(n8880) );
  INV_X1 U5495 ( .A(n9905), .ZN(n9943) );
  AND2_X1 U5496 ( .A1(n5561), .A2(n5562), .ZN(n9905) );
  INV_X1 U5497 ( .A(n9929), .ZN(n9941) );
  INV_X1 U5498 ( .A(n7024), .ZN(n7256) );
  AND2_X1 U5499 ( .A1(n5540), .A2(n5539), .ZN(n9833) );
  NAND2_X1 U5500 ( .A1(n5556), .A2(n6633), .ZN(n5558) );
  INV_X1 U5501 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4985) );
  INV_X1 U5502 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4955) );
  AND2_X1 U5503 ( .A1(n5176), .A2(n5175), .ZN(n7128) );
  AND2_X1 U5504 ( .A1(n5118), .A2(n5135), .ZN(n6921) );
  AND2_X1 U5505 ( .A1(n5021), .A2(n4949), .ZN(n5066) );
  INV_X1 U5506 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4949) );
  INV_X1 U5507 ( .A(n6380), .ZN(n6377) );
  NAND2_X1 U5508 ( .A1(n6994), .A2(n5978), .ZN(n7084) );
  NOR2_X1 U5509 ( .A1(n9005), .A2(n4708), .ZN(n4707) );
  NOR2_X1 U5510 ( .A1(n9004), .A2(n6281), .ZN(n4701) );
  INV_X1 U5511 ( .A(n4707), .ZN(n4703) );
  INV_X1 U5512 ( .A(n4705), .ZN(n4704) );
  OAI21_X1 U5513 ( .B1(n8938), .B2(n4303), .A(n4706), .ZN(n4705) );
  INV_X1 U5514 ( .A(n8986), .ZN(n4706) );
  INV_X1 U5515 ( .A(n8963), .ZN(n4696) );
  INV_X1 U5516 ( .A(n8970), .ZN(n4697) );
  OR2_X1 U5517 ( .A1(n6360), .A2(n6359), .ZN(n6398) );
  NAND2_X1 U5518 ( .A1(n6182), .A2(n6181), .ZN(n7874) );
  NAND2_X1 U5519 ( .A1(n6334), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6351) );
  INV_X1 U5520 ( .A(n6336), .ZN(n6334) );
  OR2_X1 U5521 ( .A1(n6250), .A2(n5908), .ZN(n6273) );
  NAND2_X1 U5522 ( .A1(n6271), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6287) );
  INV_X1 U5523 ( .A(n6273), .ZN(n6271) );
  INV_X1 U5524 ( .A(n9036), .ZN(n9021) );
  AND2_X1 U5525 ( .A1(n6501), .A2(n6753), .ZN(n9033) );
  INV_X1 U5526 ( .A(n6242), .ZN(n4372) );
  OAI21_X1 U5527 ( .B1(n4307), .B2(n4375), .A(n4374), .ZN(n4373) );
  INV_X1 U5528 ( .A(n7856), .ZN(n4374) );
  OAI21_X1 U5529 ( .B1(n7853), .B2(n7856), .A(n7854), .ZN(n6243) );
  NOR4_X1 U5530 ( .A1(n8170), .A2(n8037), .A3(n8232), .A4(n8036), .ZN(n8039)
         );
  NOR2_X1 U5531 ( .A1(n4421), .A2(n9184), .ZN(n8035) );
  NAND2_X1 U5532 ( .A1(n8174), .A2(n8175), .ZN(n4416) );
  NOR2_X1 U5533 ( .A1(n8056), .A2(n9736), .ZN(n4417) );
  INV_X1 U5534 ( .A(n5848), .ZN(n5856) );
  INV_X1 U5535 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U5536 ( .A1(n5888), .A2(n4818), .ZN(n5848) );
  NOR2_X1 U5537 ( .A1(n5847), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4818) );
  AND4_X1 U5538 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n7373)
         );
  AND4_X1 U5539 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n7380)
         );
  OR2_X1 U5540 ( .A1(n6026), .A2(n6027), .ZN(n6028) );
  OR2_X1 U5541 ( .A1(n9639), .A2(n9638), .ZN(n4513) );
  NAND2_X1 U5542 ( .A1(n9695), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4497) );
  OR2_X1 U5543 ( .A1(n7069), .A2(n7068), .ZN(n4507) );
  XNOR2_X1 U5544 ( .A(n7618), .B(n7617), .ZN(n7285) );
  AND2_X1 U5545 ( .A1(n4518), .A2(n4517), .ZN(n9092) );
  NAND2_X1 U5546 ( .A1(n9089), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4517) );
  NOR2_X1 U5547 ( .A1(n9092), .A2(n9091), .ZN(n9097) );
  INV_X1 U5548 ( .A(n9624), .ZN(n6753) );
  INV_X1 U5549 ( .A(n4439), .ZN(n4437) );
  INV_X1 U5550 ( .A(n4782), .ZN(n9125) );
  INV_X1 U5551 ( .A(n4784), .ZN(n4783) );
  AND2_X1 U5552 ( .A1(n6440), .A2(n6417), .ZN(n9149) );
  OR2_X1 U5553 ( .A1(n9415), .A2(n9044), .ZN(n9168) );
  NOR2_X1 U5554 ( .A1(n9193), .A2(n8227), .ZN(n9170) );
  NAND2_X1 U5555 ( .A1(n9260), .A2(n4451), .ZN(n9201) );
  AND2_X1 U5556 ( .A1(n4291), .A2(n9192), .ZN(n4451) );
  NOR2_X1 U5557 ( .A1(n9201), .A2(n9415), .ZN(n9179) );
  NAND2_X1 U5558 ( .A1(n9256), .A2(n4314), .ZN(n4590) );
  NAND2_X1 U5559 ( .A1(n9260), .A2(n4291), .ZN(n9210) );
  AND2_X1 U5560 ( .A1(n9260), .A2(n9251), .ZN(n9246) );
  NAND2_X1 U5561 ( .A1(n9260), .A2(n4453), .ZN(n9224) );
  OR2_X1 U5562 ( .A1(n6318), .A2(n6317), .ZN(n6336) );
  OR2_X1 U5563 ( .A1(n9264), .A2(n9245), .ZN(n4828) );
  OR2_X1 U5564 ( .A1(n9442), .A2(n9276), .ZN(n8193) );
  OR2_X1 U5565 ( .A1(n6303), .A2(n6302), .ZN(n6318) );
  AND4_X1 U5566 ( .A1(n6325), .A2(n6324), .A3(n6323), .A4(n6322), .ZN(n9259)
         );
  NAND2_X1 U5567 ( .A1(n4809), .A2(n4807), .ZN(n9282) );
  AOI21_X1 U5568 ( .B1(n4813), .B2(n4808), .A(n4812), .ZN(n4807) );
  NAND2_X1 U5569 ( .A1(n9333), .A2(n4315), .ZN(n4809) );
  OAI22_X1 U5570 ( .A1(n8191), .A2(n4816), .B1(n9320), .B2(n9305), .ZN(n4812)
         );
  AND2_X1 U5571 ( .A1(n9379), .A2(n4448), .ZN(n9301) );
  AND2_X1 U5572 ( .A1(n4292), .A2(n9305), .ZN(n4448) );
  AND2_X1 U5573 ( .A1(n9379), .A2(n4292), .ZN(n9321) );
  NAND2_X1 U5574 ( .A1(n5907), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6250) );
  INV_X1 U5575 ( .A(n6248), .ZN(n5907) );
  NOR2_X1 U5576 ( .A1(n4584), .A2(n8021), .ZN(n4581) );
  OAI21_X1 U5577 ( .B1(n4582), .B2(n8021), .A(n4580), .ZN(n4579) );
  NAND2_X1 U5578 ( .A1(n9379), .A2(n4450), .ZN(n9337) );
  OR2_X1 U5579 ( .A1(n8211), .A2(n8021), .ZN(n9332) );
  NAND2_X1 U5580 ( .A1(n4578), .A2(n4582), .ZN(n9327) );
  NAND2_X1 U5581 ( .A1(n9369), .A2(n4585), .ZN(n4578) );
  NAND2_X1 U5582 ( .A1(n9379), .A2(n9592), .ZN(n9357) );
  NAND2_X1 U5583 ( .A1(n9371), .A2(n8209), .ZN(n9351) );
  OR2_X1 U5584 ( .A1(n6191), .A2(n6169), .ZN(n6171) );
  NAND2_X1 U5585 ( .A1(n5904), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6189) );
  INV_X1 U5586 ( .A(n6138), .ZN(n5904) );
  OR2_X1 U5587 ( .A1(n7797), .A2(n9597), .ZN(n9378) );
  OR2_X1 U5588 ( .A1(n9553), .A2(n9479), .ZN(n7797) );
  AND4_X1 U5589 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n7788)
         );
  OR2_X1 U5590 ( .A1(n6094), .A2(n6093), .ZN(n6112) );
  OR2_X1 U5591 ( .A1(n6112), .A2(n7530), .ZN(n6138) );
  AND2_X1 U5592 ( .A1(n7509), .A2(n7514), .ZN(n9555) );
  NAND2_X1 U5593 ( .A1(n7505), .A2(n8073), .ZN(n7732) );
  NOR2_X1 U5594 ( .A1(n7401), .A2(n7598), .ZN(n7509) );
  NAND2_X1 U5595 ( .A1(n7440), .A2(n9766), .ZN(n7442) );
  AND2_X1 U5596 ( .A1(n7540), .A2(n7164), .ZN(n7440) );
  INV_X1 U5597 ( .A(n7995), .ZN(n4556) );
  INV_X1 U5598 ( .A(n7989), .ZN(n4557) );
  INV_X1 U5599 ( .A(n8024), .ZN(n4558) );
  AND4_X1 U5600 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n7145)
         );
  OR2_X1 U5601 ( .A1(n5989), .A2(n5990), .ZN(n5995) );
  NAND2_X1 U5602 ( .A1(n7102), .A2(n7989), .ZN(n7158) );
  INV_X1 U5603 ( .A(n6499), .ZN(n9735) );
  INV_X1 U5604 ( .A(n9167), .ZN(n9410) );
  NAND2_X1 U5605 ( .A1(n6270), .A2(n6269), .ZN(n9450) );
  INV_X1 U5606 ( .A(n9552), .ZN(n9565) );
  AND2_X1 U5607 ( .A1(n6458), .A2(n6457), .ZN(n9487) );
  INV_X1 U5608 ( .A(n9767), .ZN(n9554) );
  NOR2_X1 U5609 ( .A1(n6834), .A2(n6567), .ZN(n6844) );
  OAI21_X1 U5610 ( .B1(n4282), .B2(n4391), .A(n4390), .ZN(n5641) );
  XNOR2_X1 U5611 ( .A(n5622), .B(n5613), .ZN(n7947) );
  XNOR2_X1 U5612 ( .A(n5608), .B(n5607), .ZN(n7903) );
  XNOR2_X1 U5613 ( .A(n5505), .B(n5504), .ZN(n7884) );
  INV_X1 U5614 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U5615 ( .A1(n5885), .A2(n5884), .ZN(n5887) );
  XNOR2_X1 U5616 ( .A(n5437), .B(n5432), .ZN(n7780) );
  NAND2_X1 U5617 ( .A1(n4742), .A2(n4933), .ZN(n5385) );
  NOR2_X1 U5618 ( .A1(n6225), .A2(n5874), .ZN(n5916) );
  OAI21_X1 U5619 ( .B1(n4898), .B2(n4302), .A(n4466), .ZN(n5282) );
  NAND2_X1 U5620 ( .A1(n6147), .A2(n5864), .ZN(n6225) );
  INV_X1 U5621 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U5622 ( .A1(n4898), .A2(n4897), .ZN(n5262) );
  INV_X1 U5623 ( .A(n4722), .ZN(n5246) );
  AOI21_X1 U5624 ( .B1(n5209), .B2(n4729), .A(n4725), .ZN(n4722) );
  AND2_X1 U5625 ( .A1(n6185), .A2(n6184), .ZN(n7065) );
  NAND2_X1 U5626 ( .A1(n4377), .A2(n4381), .ZN(n5171) );
  OR2_X1 U5627 ( .A1(n5134), .A2(n4383), .ZN(n4377) );
  NAND2_X1 U5628 ( .A1(n5019), .A2(n5018), .ZN(n4851) );
  AOI21_X1 U5629 ( .B1(n5966), .B2(P1_IR_REG_2__SCAN_IN), .A(n4534), .ZN(n6527) );
  NAND2_X1 U5630 ( .A1(n5967), .A2(n4535), .ZN(n4534) );
  NAND2_X1 U5631 ( .A1(n9517), .A2(n4797), .ZN(n4535) );
  OR3_X1 U5632 ( .A1(n7785), .A2(n7870), .A3(n7849), .ZN(n6870) );
  NAND2_X1 U5633 ( .A1(n7231), .A2(n5132), .ZN(n7246) );
  NAND2_X1 U5634 ( .A1(n4641), .A2(n4646), .ZN(n8266) );
  NAND2_X1 U5635 ( .A1(n7684), .A2(n5191), .ZN(n7712) );
  NAND2_X1 U5636 ( .A1(n5354), .A2(n5353), .ZN(n8869) );
  OAI21_X1 U5637 ( .B1(n8447), .B2(n4645), .A(n4642), .ZN(n5574) );
  INV_X1 U5638 ( .A(n9806), .ZN(n9914) );
  INV_X1 U5639 ( .A(n4402), .ZN(n7364) );
  AOI21_X1 U5640 ( .B1(n7231), .B2(n4404), .A(n4403), .ZN(n4402) );
  NAND2_X1 U5641 ( .A1(n8393), .A2(n5383), .ZN(n4407) );
  NAND2_X1 U5642 ( .A1(n5224), .A2(n5223), .ZN(n8331) );
  NAND2_X1 U5643 ( .A1(n8298), .A2(n4663), .ZN(n4662) );
  AND4_X1 U5644 ( .A1(n5205), .A2(n5204), .A3(n5203), .A4(n5202), .ZN(n7691)
         );
  NAND2_X1 U5645 ( .A1(n8311), .A2(n5367), .ZN(n8395) );
  NAND2_X1 U5646 ( .A1(n5371), .A2(n5370), .ZN(n8863) );
  NAND2_X1 U5647 ( .A1(n7462), .A2(n5489), .ZN(n4462) );
  OAI21_X1 U5648 ( .B1(n5190), .B2(n4656), .A(n4411), .ZN(n8421) );
  NAND2_X1 U5649 ( .A1(n7073), .A2(n5039), .ZN(n8248) );
  NAND2_X1 U5650 ( .A1(n5575), .A2(n5566), .ZN(n8445) );
  INV_X1 U5651 ( .A(n8454), .ZN(n8464) );
  NAND2_X1 U5652 ( .A1(n8447), .A2(n5478), .ZN(n4395) );
  NAND2_X1 U5653 ( .A1(n5563), .A2(n8678), .ZN(n8469) );
  INV_X2 U5654 ( .A(P2_U3966), .ZN(n8493) );
  NOR2_X1 U5655 ( .A1(n6940), .A2(n4542), .ZN(n6881) );
  AND2_X1 U5656 ( .A1(n6888), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4542) );
  NOR2_X1 U5657 ( .A1(n6881), .A2(n6880), .ZN(n6899) );
  OR2_X1 U5658 ( .A1(n6945), .A2(n6946), .ZN(n6889) );
  NOR2_X1 U5659 ( .A1(n6915), .A2(n4545), .ZN(n6932) );
  AND2_X1 U5660 ( .A1(n6921), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4545) );
  NOR2_X1 U5661 ( .A1(n6932), .A2(n6931), .ZN(n6930) );
  NOR2_X1 U5662 ( .A1(n6930), .A2(n4544), .ZN(n6918) );
  AND2_X1 U5663 ( .A1(n6920), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4544) );
  NOR2_X1 U5664 ( .A1(n6918), .A2(n6917), .ZN(n7029) );
  NAND2_X1 U5665 ( .A1(n6934), .A2(n4321), .ZN(n6927) );
  OAI21_X1 U5666 ( .B1(n7039), .B2(n6925), .A(n7038), .ZN(n7040) );
  AOI21_X1 U5667 ( .B1(n7468), .B2(n7336), .A(n7467), .ZN(n7471) );
  AOI21_X1 U5668 ( .B1(n7805), .B2(n7804), .A(n7803), .ZN(n7810) );
  NOR2_X1 U5669 ( .A1(n7913), .A2(n7912), .ZN(n8502) );
  NOR2_X1 U5670 ( .A1(n8513), .A2(n8512), .ZN(n8511) );
  NAND2_X1 U5671 ( .A1(n4365), .A2(n4364), .ZN(n8520) );
  NAND2_X1 U5672 ( .A1(n7916), .A2(n8530), .ZN(n4364) );
  INV_X1 U5673 ( .A(n7917), .ZN(n4365) );
  INV_X1 U5674 ( .A(n8822), .ZN(n8599) );
  NAND2_X1 U5675 ( .A1(n8620), .A2(n4475), .ZN(n8611) );
  NAND2_X1 U5676 ( .A1(n8643), .A2(n5760), .ZN(n8622) );
  NAND2_X1 U5677 ( .A1(n8670), .A2(n5655), .ZN(n8657) );
  NAND2_X1 U5678 ( .A1(n8666), .A2(n8557), .ZN(n8648) );
  NAND2_X1 U5679 ( .A1(n4620), .A2(n4619), .ZN(n8692) );
  NAND2_X1 U5680 ( .A1(n8713), .A2(n4829), .ZN(n8702) );
  AND2_X1 U5681 ( .A1(n5336), .A2(n5335), .ZN(n8755) );
  AND2_X1 U5682 ( .A1(n4758), .A2(n4757), .ZN(n8745) );
  NAND2_X1 U5683 ( .A1(n4605), .A2(n4608), .ZN(n8761) );
  NAND2_X1 U5684 ( .A1(n8798), .A2(n4611), .ZN(n4605) );
  NAND2_X1 U5685 ( .A1(n8775), .A2(n4759), .ZN(n8759) );
  NAND2_X1 U5686 ( .A1(n4613), .A2(n5722), .ZN(n8785) );
  NAND2_X1 U5687 ( .A1(n4615), .A2(n4614), .ZN(n4613) );
  NAND2_X1 U5688 ( .A1(n7827), .A2(n5711), .ZN(n9571) );
  NAND2_X1 U5689 ( .A1(n7822), .A2(n4770), .ZN(n7823) );
  NAND2_X1 U5690 ( .A1(n7751), .A2(n7304), .ZN(n7306) );
  INV_X1 U5691 ( .A(n5138), .ZN(n5139) );
  OAI21_X1 U5692 ( .B1(n5097), .B2(n6595), .A(n5137), .ZN(n5138) );
  NAND2_X1 U5693 ( .A1(n9829), .A2(n9819), .ZN(n8795) );
  INV_X1 U5694 ( .A(n8808), .ZN(n9581) );
  INV_X1 U5695 ( .A(n8795), .ZN(n9805) );
  NOR2_X1 U5696 ( .A1(n8539), .A2(n9943), .ZN(n8806) );
  AND2_X2 U5697 ( .A1(n7025), .A2(n7024), .ZN(n9967) );
  NAND2_X1 U5698 ( .A1(n4635), .A2(n4634), .ZN(n4633) );
  NOR2_X1 U5699 ( .A1(n4964), .A2(n5528), .ZN(n4965) );
  INV_X1 U5700 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7783) );
  XNOR2_X1 U5701 ( .A(n5536), .B(n5535), .ZN(n7785) );
  NAND2_X1 U5702 ( .A1(n5558), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5536) );
  AND2_X1 U5703 ( .A1(P2_U3152), .A2(n4282), .ZN(n7592) );
  INV_X1 U5704 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7464) );
  INV_X1 U5705 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7360) );
  INV_X1 U5706 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7252) );
  INV_X1 U5707 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7138) );
  INV_X1 U5708 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6993) );
  AND2_X1 U5709 ( .A1(n5317), .A2(n5286), .ZN(n8503) );
  NOR2_X1 U5710 ( .A1(n4282), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8918) );
  INV_X1 U5711 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6829) );
  INV_X1 U5712 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6797) );
  INV_X1 U5713 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6792) );
  INV_X1 U5714 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6747) );
  INV_X1 U5715 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6743) );
  INV_X1 U5716 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6730) );
  INV_X1 U5717 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6599) );
  INV_X1 U5718 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6580) );
  INV_X1 U5719 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6579) );
  INV_X1 U5720 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6578) );
  INV_X1 U5721 ( .A(n4550), .ZN(n4549) );
  OAI21_X1 U5722 ( .B1(n5020), .B2(n4552), .A(n4551), .ZN(n4550) );
  NAND2_X1 U5723 ( .A1(n4282), .A2(SI_0_), .ZN(n5028) );
  NOR2_X1 U5724 ( .A1(n6513), .A2(n7572), .ZN(n6539) );
  NAND2_X1 U5725 ( .A1(n7428), .A2(n6056), .ZN(n7355) );
  NAND2_X1 U5726 ( .A1(n6804), .A2(n5940), .ZN(n6815) );
  NOR2_X1 U5727 ( .A1(n8962), .A2(n8963), .ZN(n8961) );
  NAND2_X1 U5728 ( .A1(n4694), .A2(n9028), .ZN(n8962) );
  NAND2_X1 U5729 ( .A1(n6092), .A2(n7410), .ZN(n7493) );
  AOI21_X1 U5730 ( .B1(n8937), .B2(n8938), .A(n4303), .ZN(n8988) );
  INV_X1 U5731 ( .A(n9373), .ZN(n9331) );
  NAND2_X1 U5732 ( .A1(n6345), .A2(n6346), .ZN(n8995) );
  OR2_X1 U5733 ( .A1(n6345), .A2(n6346), .ZN(n8994) );
  AND4_X1 U5734 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n7734)
         );
  OR2_X1 U5735 ( .A1(n4688), .A2(n4687), .ZN(n4686) );
  NAND2_X1 U5736 ( .A1(n6810), .A2(n6484), .ZN(n9027) );
  NAND2_X1 U5737 ( .A1(n6490), .A2(n6810), .ZN(n9031) );
  NAND2_X1 U5738 ( .A1(n9016), .A2(n9015), .ZN(n9019) );
  NAND2_X1 U5739 ( .A1(n8952), .A2(n6413), .ZN(n9017) );
  AND4_X1 U5740 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n9329)
         );
  NAND2_X1 U5741 ( .A1(n6230), .A2(n6229), .ZN(n9465) );
  INV_X1 U5742 ( .A(n9259), .ZN(n9235) );
  INV_X1 U5743 ( .A(n7788), .ZN(n9374) );
  INV_X1 U5744 ( .A(n7380), .ZN(n9047) );
  NAND4_X1 U5745 ( .A1(n6011), .A2(n6010), .A3(n6009), .A4(n6008), .ZN(n9048)
         );
  INV_X1 U5746 ( .A(n7145), .ZN(n9049) );
  INV_X1 U5747 ( .A(n7192), .ZN(n9050) );
  OR2_X1 U5748 ( .A1(n6025), .A2(n9742), .ZN(n5943) );
  NAND2_X1 U5749 ( .A1(n6798), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5942) );
  AND2_X1 U5750 ( .A1(n4513), .A2(n4299), .ZN(n9656) );
  AND2_X1 U5751 ( .A1(n4512), .A2(n4308), .ZN(n6774) );
  INV_X1 U5752 ( .A(n4500), .ZN(n6778) );
  INV_X1 U5753 ( .A(n9676), .ZN(n6522) );
  INV_X1 U5754 ( .A(n4498), .ZN(n9689) );
  NOR2_X1 U5755 ( .A1(n7064), .A2(n4508), .ZN(n7069) );
  AND2_X1 U5756 ( .A1(n7065), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4508) );
  INV_X1 U5757 ( .A(n4507), .ZN(n7282) );
  NOR2_X1 U5758 ( .A1(n9065), .A2(n9066), .ZN(n9069) );
  INV_X1 U5759 ( .A(n4518), .ZN(n9088) );
  AND2_X1 U5760 ( .A1(n9673), .A2(n9624), .ZN(n9704) );
  OR2_X1 U5761 ( .A1(n9147), .A2(n8015), .ZN(n4436) );
  NAND2_X1 U5762 ( .A1(n4434), .A2(n9389), .ZN(n4433) );
  NAND2_X1 U5763 ( .A1(n9147), .A2(n4317), .ZN(n4435) );
  NAND2_X1 U5764 ( .A1(n9147), .A2(n4438), .ZN(n9390) );
  NAND2_X1 U5765 ( .A1(n8237), .A2(n8236), .ZN(n8238) );
  NOR2_X1 U5766 ( .A1(n9133), .A2(n9132), .ZN(n9134) );
  AOI211_X1 U5767 ( .C1(n9720), .C2(n9186), .A(n9157), .B(n9156), .ZN(n9408)
         );
  OAI21_X1 U5768 ( .B1(n9191), .B2(n4787), .A(n4785), .ZN(n9146) );
  NAND2_X1 U5769 ( .A1(n4788), .A2(n4791), .ZN(n9162) );
  NAND2_X1 U5770 ( .A1(n9191), .A2(n4792), .ZN(n4788) );
  NAND2_X1 U5771 ( .A1(n4595), .A2(n8220), .ZN(n9241) );
  INV_X1 U5772 ( .A(n9450), .ZN(n9288) );
  AOI21_X1 U5773 ( .B1(n9314), .B2(n9315), .A(n4811), .ZN(n9300) );
  INV_X1 U5774 ( .A(n4816), .ZN(n4811) );
  INV_X1 U5775 ( .A(n9465), .ZN(n9342) );
  INV_X1 U5776 ( .A(n4776), .ZN(n8184) );
  AOI21_X1 U5777 ( .B1(n7731), .B2(n4777), .A(n4780), .ZN(n4776) );
  NAND2_X1 U5778 ( .A1(n7502), .A2(n7501), .ZN(n7729) );
  NOR2_X1 U5779 ( .A1(n4316), .A2(n4290), .ZN(n4419) );
  NAND2_X1 U5780 ( .A1(n6065), .A2(n6082), .ZN(n4420) );
  INV_X1 U5781 ( .A(n6543), .ZN(n9755) );
  NAND2_X1 U5782 ( .A1(n9740), .A2(n9727), .ZN(n9341) );
  AND2_X1 U5783 ( .A1(n4442), .A2(n4444), .ZN(n4447) );
  NAND2_X1 U5784 ( .A1(n6511), .A2(n4443), .ZN(n4442) );
  XNOR2_X1 U5785 ( .A(n6551), .B(n9716), .ZN(n9726) );
  INV_X1 U5786 ( .A(n9341), .ZN(n9551) );
  AND2_X1 U5787 ( .A1(n9740), .A2(n6571), .ZN(n9346) );
  AND2_X2 U5788 ( .A1(n6843), .A2(n6835), .ZN(n9782) );
  AND2_X2 U5789 ( .A1(n6844), .A2(n6843), .ZN(n9774) );
  MUX2_X1 U5790 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5896), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5897) );
  INV_X1 U5791 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7781) );
  XNOR2_X1 U5792 ( .A(n5891), .B(n5890), .ZN(n7782) );
  XNOR2_X1 U5793 ( .A(n5412), .B(n5413), .ZN(n7593) );
  INV_X1 U5794 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7463) );
  INV_X1 U5795 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7333) );
  INV_X1 U5796 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7243) );
  INV_X1 U5797 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7141) );
  AND2_X1 U5798 ( .A1(n5869), .A2(n6267), .ZN(n9104) );
  INV_X1 U5799 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6828) );
  INV_X1 U5800 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6795) );
  INV_X1 U5801 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6791) );
  INV_X1 U5802 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6749) );
  INV_X1 U5803 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6741) );
  INV_X1 U5804 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U5805 ( .A1(n4386), .A2(n4867), .ZN(n5151) );
  NAND2_X1 U5806 ( .A1(n5134), .A2(n4865), .ZN(n4386) );
  INV_X1 U5807 ( .A(n6065), .ZN(n6596) );
  INV_X1 U5808 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U5809 ( .A1(n4626), .A2(n4625), .ZN(n5111) );
  AOI21_X1 U5810 ( .B1(n4627), .B2(n4286), .A(n4294), .ZN(n4626) );
  XNOR2_X1 U5811 ( .A(n5096), .B(n5095), .ZN(n6585) );
  OAI21_X1 U5812 ( .B1(n4282), .B2(n5924), .A(n5923), .ZN(n5926) );
  NOR2_X1 U5813 ( .A1(n7656), .A2(n10001), .ZN(n9996) );
  AOI21_X1 U5814 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9994), .ZN(n9993) );
  NOR2_X1 U5815 ( .A1(n9993), .A2(n9992), .ZN(n9991) );
  NAND2_X1 U5816 ( .A1(n4477), .A2(n5831), .ZN(n4519) );
  NAND2_X1 U5817 ( .A1(n4369), .A2(n4368), .ZN(P1_U3212) );
  NAND2_X1 U5818 ( .A1(n8952), .A2(n4366), .ZN(n4368) );
  NOR2_X1 U5819 ( .A1(n8922), .A2(n4367), .ZN(n4366) );
  NOR4_X1 U5820 ( .A1(n4674), .A2(n6480), .A3(n6481), .A4(n4371), .ZN(n4673)
         );
  NAND2_X1 U5821 ( .A1(n4413), .A2(n4412), .ZN(n8182) );
  OAI211_X1 U5822 ( .C1(n9111), .C2(n9736), .A(n4532), .B(n4529), .ZN(P1_U3260) );
  NOR2_X1 U5823 ( .A1(n4533), .A2(n4363), .ZN(n4532) );
  NAND2_X1 U5824 ( .A1(n4530), .A2(n9736), .ZN(n4529) );
  INV_X1 U5825 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9517) );
  AND2_X1 U5826 ( .A1(n4859), .A2(SI_4_), .ZN(n4286) );
  XNOR2_X1 U5827 ( .A(n8834), .B(n8563), .ZN(n5653) );
  OR2_X1 U5828 ( .A1(n9405), .A2(n9173), .ZN(n4287) );
  NAND2_X1 U5829 ( .A1(n5267), .A2(n5266), .ZN(n9576) );
  NAND2_X1 U5830 ( .A1(n6877), .A2(n4282), .ZN(n5046) );
  AND2_X1 U5831 ( .A1(n5888), .A2(n4340), .ZN(n5895) );
  AND2_X1 U5832 ( .A1(n4576), .A2(n4575), .ZN(n4574) );
  AND2_X1 U5833 ( .A1(n5207), .A2(n5206), .ZN(n4288) );
  AND2_X1 U5834 ( .A1(n4481), .A2(n9586), .ZN(n4289) );
  AND2_X1 U5835 ( .A1(n6282), .A2(n6786), .ZN(n4290) );
  XNOR2_X1 U5836 ( .A(n5894), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5898) );
  XNOR2_X1 U5837 ( .A(n4858), .B(SI_4_), .ZN(n5083) );
  INV_X1 U5838 ( .A(n5083), .ZN(n4459) );
  AND2_X1 U5839 ( .A1(n4453), .A2(n4452), .ZN(n4291) );
  OR2_X1 U5840 ( .A1(n9430), .A2(n9244), .ZN(n8127) );
  AND2_X1 U5841 ( .A1(n4450), .A2(n4449), .ZN(n4292) );
  INV_X1 U5842 ( .A(n9232), .ZN(n4597) );
  OR2_X1 U5843 ( .A1(n4303), .A2(n4701), .ZN(n4293) );
  INV_X1 U5844 ( .A(n4609), .ZN(n4608) );
  OAI21_X1 U5845 ( .B1(n4614), .B2(n4610), .A(n5725), .ZN(n4609) );
  OR2_X1 U5846 ( .A1(n8838), .A2(n8659), .ZN(n5760) );
  INV_X1 U5847 ( .A(n9430), .ZN(n9230) );
  NAND2_X1 U5848 ( .A1(n6333), .A2(n6332), .ZN(n9430) );
  AND2_X1 U5849 ( .A1(n4862), .A2(SI_5_), .ZN(n4294) );
  INV_X1 U5850 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U5851 ( .A1(n4333), .A2(n4795), .ZN(n4791) );
  AND2_X1 U5852 ( .A1(n4393), .A2(n6346), .ZN(n4295) );
  INV_X1 U5853 ( .A(n9405), .ZN(n9151) );
  NAND2_X1 U5854 ( .A1(n6415), .A2(n6414), .ZN(n9405) );
  AND2_X1 U5855 ( .A1(n4289), .A2(n8796), .ZN(n4296) );
  NAND2_X1 U5856 ( .A1(n7773), .A2(n4289), .ZN(n4297) );
  AND4_X1 U5857 ( .A1(n4952), .A2(n4950), .A3(n5114), .A4(n4951), .ZN(n4298)
         );
  NAND2_X1 U5858 ( .A1(n7392), .A2(n4306), .ZN(n7502) );
  INV_X1 U5860 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5114) );
  OR2_X1 U5861 ( .A1(n6526), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4299) );
  INV_X1 U5862 ( .A(n4446), .ZN(n6033) );
  NAND2_X1 U5863 ( .A1(n6511), .A2(n4282), .ZN(n4446) );
  AND3_X1 U5864 ( .A1(n5125), .A2(n5124), .A3(n5123), .ZN(n4300) );
  NAND2_X1 U5865 ( .A1(n5109), .A2(n5108), .ZN(n4301) );
  NAND2_X1 U5866 ( .A1(n6013), .A2(n4334), .ZN(n5860) );
  NAND2_X1 U5867 ( .A1(n9885), .A2(n8492), .ZN(n4746) );
  OR2_X1 U5868 ( .A1(n5302), .A2(n4468), .ZN(n4302) );
  AND2_X1 U5869 ( .A1(n6299), .A2(n6298), .ZN(n4303) );
  NAND2_X1 U5870 ( .A1(n5947), .A2(n4797), .ZN(n5967) );
  INV_X2 U5871 ( .A(n6026), .ZN(n5941) );
  NAND2_X1 U5872 ( .A1(n9118), .A2(n8051), .ZN(n4304) );
  NOR2_X1 U5873 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5947) );
  INV_X1 U5874 ( .A(n5791), .ZN(n4739) );
  NAND2_X1 U5875 ( .A1(n6013), .A2(n4803), .ZN(n6036) );
  INV_X1 U5876 ( .A(n8227), .ZN(n4577) );
  NAND2_X1 U5877 ( .A1(n8859), .A2(n8552), .ZN(n4305) );
  AND2_X1 U5878 ( .A1(n7382), .A2(n7381), .ZN(n4306) );
  NOR2_X1 U5879 ( .A1(n6212), .A2(n6239), .ZN(n4307) );
  AND4_X1 U5880 ( .A1(n5056), .A2(n5055), .A3(n5054), .A4(n5053), .ZN(n4835)
         );
  OR2_X1 U5881 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9653), .ZN(n4308) );
  NOR2_X1 U5882 ( .A1(n9192), .A2(n8957), .ZN(n4309) );
  NAND2_X1 U5883 ( .A1(n7937), .A2(n7936), .ZN(n8015) );
  NAND2_X1 U5884 ( .A1(n6511), .A2(n6581), .ZN(n6067) );
  OR2_X1 U5885 ( .A1(n4393), .A2(n6346), .ZN(n4310) );
  NAND2_X1 U5886 ( .A1(n4975), .A2(n4974), .ZN(n8842) );
  INV_X1 U5887 ( .A(n9155), .ZN(n4570) );
  INV_X1 U5888 ( .A(n6877), .ZN(n5351) );
  INV_X1 U5889 ( .A(n9004), .ZN(n4708) );
  AND2_X1 U5890 ( .A1(n6013), .A2(n5837), .ZN(n6034) );
  OR2_X1 U5891 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4311) );
  AND2_X1 U5892 ( .A1(n4595), .A2(n4593), .ZN(n4312) );
  NAND4_X1 U5893 ( .A1(n4797), .A2(n4432), .A3(n4431), .A4(n4430), .ZN(n5997)
         );
  NAND2_X1 U5894 ( .A1(n6152), .A2(n6151), .ZN(n9359) );
  OR2_X1 U5895 ( .A1(n9479), .A2(n9545), .ZN(n4313) );
  AND2_X1 U5896 ( .A1(n4620), .A2(n4305), .ZN(n8691) );
  INV_X1 U5897 ( .A(n4729), .ZN(n4727) );
  NOR2_X1 U5898 ( .A1(n5225), .A2(n4730), .ZN(n4729) );
  AND4_X1 U5899 ( .A1(n6031), .A2(n6030), .A3(n6029), .A4(n6028), .ZN(n7537)
         );
  INV_X1 U5900 ( .A(n7537), .ZN(n4681) );
  AND2_X1 U5901 ( .A1(n4593), .A2(n8127), .ZN(n4314) );
  AND2_X1 U5902 ( .A1(n4813), .A2(n4810), .ZN(n4315) );
  AND2_X1 U5903 ( .A1(n7939), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4316) );
  AND2_X1 U5904 ( .A1(n8015), .A2(n4438), .ZN(n4317) );
  INV_X1 U5905 ( .A(n8828), .ZN(n8609) );
  NAND2_X1 U5906 ( .A1(n5491), .A2(n5490), .ZN(n8828) );
  NAND2_X1 U5907 ( .A1(n6316), .A2(n6315), .ZN(n9437) );
  INV_X1 U5908 ( .A(n7405), .ZN(n7454) );
  AND2_X1 U5909 ( .A1(n4420), .A2(n4419), .ZN(n7405) );
  INV_X1 U5910 ( .A(n8957), .ZN(n9218) );
  AND2_X1 U5911 ( .A1(n6367), .A2(n6366), .ZN(n8957) );
  AND2_X1 U5912 ( .A1(n4498), .A2(n4497), .ZN(n4318) );
  NAND2_X1 U5913 ( .A1(n8677), .A2(n4484), .ZN(n4487) );
  NAND2_X1 U5914 ( .A1(n5483), .A2(n5482), .ZN(n5505) );
  OR2_X1 U5915 ( .A1(n9425), .A2(n8197), .ZN(n8224) );
  NAND2_X1 U5916 ( .A1(n7941), .A2(n7940), .ZN(n9118) );
  AND2_X1 U5917 ( .A1(n6040), .A2(n6039), .ZN(n4319) );
  NAND2_X1 U5918 ( .A1(n7721), .A2(n6240), .ZN(n4320) );
  OR2_X1 U5919 ( .A1(n6939), .A2(n6924), .ZN(n4321) );
  AND2_X1 U5920 ( .A1(n5689), .A2(n5688), .ZN(n9796) );
  INV_X1 U5921 ( .A(n4760), .ZN(n4759) );
  AND2_X1 U5922 ( .A1(n4686), .A2(n6215), .ZN(n4322) );
  INV_X1 U5923 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4797) );
  INV_X1 U5924 ( .A(n8211), .ZN(n4580) );
  AND2_X1 U5925 ( .A1(n9167), .A2(n8198), .ZN(n4323) );
  AND2_X1 U5926 ( .A1(n5839), .A2(n4804), .ZN(n4324) );
  NAND2_X1 U5927 ( .A1(n8620), .A2(n5769), .ZN(n4325) );
  OR2_X1 U5928 ( .A1(n8880), .A2(n8749), .ZN(n5729) );
  OR2_X1 U5929 ( .A1(n8706), .A2(n8552), .ZN(n4326) );
  OR2_X1 U5930 ( .A1(n8034), .A2(n4426), .ZN(n4327) );
  INV_X1 U5931 ( .A(n6111), .ZN(n4691) );
  INV_X1 U5932 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5890) );
  INV_X1 U5933 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U5934 ( .A1(n7579), .A2(n7558), .ZN(n4328) );
  INV_X1 U5935 ( .A(n4305), .ZN(n4621) );
  OR2_X1 U5936 ( .A1(n4787), .A2(n4570), .ZN(n4329) );
  AND2_X1 U5937 ( .A1(n4864), .A2(SI_6_), .ZN(n4330) );
  NAND2_X1 U5938 ( .A1(n6581), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4331) );
  INV_X1 U5939 ( .A(n4474), .ZN(n4475) );
  NAND2_X1 U5940 ( .A1(n5770), .A2(n5769), .ZN(n4474) );
  OR2_X1 U5941 ( .A1(n4596), .A2(n4591), .ZN(n4332) );
  NAND2_X1 U5942 ( .A1(n9184), .A2(n4793), .ZN(n4333) );
  AND2_X1 U5943 ( .A1(n4803), .A2(n4324), .ZN(n4334) );
  AND2_X1 U5944 ( .A1(n8723), .A2(n5744), .ZN(n4335) );
  AND2_X1 U5945 ( .A1(n4749), .A2(n4748), .ZN(n4336) );
  AND2_X1 U5946 ( .A1(n5712), .A2(n5711), .ZN(n7829) );
  INV_X1 U5947 ( .A(n7829), .ZN(n4766) );
  AND2_X1 U5948 ( .A1(n7771), .A2(n4769), .ZN(n4337) );
  AND3_X1 U5949 ( .A1(n4958), .A2(n4668), .A3(n4979), .ZN(n4338) );
  INV_X1 U5950 ( .A(n8229), .ZN(n4576) );
  AND2_X1 U5951 ( .A1(n8553), .A2(n8726), .ZN(n4339) );
  INV_X1 U5952 ( .A(n9192), .ZN(n9421) );
  AND2_X1 U5953 ( .A1(n6358), .A2(n6357), .ZN(n9192) );
  AND2_X1 U5954 ( .A1(n4819), .A2(n4817), .ZN(n4340) );
  INV_X1 U5955 ( .A(n4286), .ZN(n4624) );
  INV_X1 U5956 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4964) );
  AND2_X1 U5957 ( .A1(n4755), .A2(n4756), .ZN(n4341) );
  AND2_X1 U5958 ( .A1(n8656), .A2(n8557), .ZN(n4342) );
  INV_X1 U5959 ( .A(n8558), .ZN(n8656) );
  AND2_X1 U5960 ( .A1(n5756), .A2(n5757), .ZN(n8558) );
  AND2_X1 U5961 ( .A1(n5786), .A2(n4738), .ZN(n4343) );
  AND2_X1 U5962 ( .A1(n4696), .A2(n4697), .ZN(n4344) );
  AND2_X1 U5963 ( .A1(n5229), .A2(n4954), .ZN(n4345) );
  AND2_X1 U5964 ( .A1(n4966), .A2(n4964), .ZN(n4346) );
  INV_X1 U5965 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U5966 ( .A1(n6348), .A2(n6347), .ZN(n9425) );
  INV_X1 U5967 ( .A(n9425), .ZN(n4452) );
  AND2_X1 U5968 ( .A1(n4298), .A2(n5066), .ZN(n5174) );
  INV_X1 U5969 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4479) );
  NAND2_X1 U5970 ( .A1(n5463), .A2(n5462), .ZN(n8834) );
  INV_X1 U5971 ( .A(n8834), .ZN(n4485) );
  AND2_X1 U5972 ( .A1(n7773), .A2(n4481), .ZN(n4347) );
  NAND2_X1 U5973 ( .A1(n7836), .A2(n7835), .ZN(n4348) );
  AND2_X1 U5974 ( .A1(n6858), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4349) );
  AND4_X1 U5975 ( .A1(n4771), .A2(n4651), .A3(n4345), .A4(n4650), .ZN(n5263)
         );
  AND2_X1 U5976 ( .A1(n6120), .A2(n5863), .ZN(n6147) );
  OR2_X1 U5977 ( .A1(n6036), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n4350) );
  NAND2_X1 U5978 ( .A1(n8714), .A2(n8726), .ZN(n8713) );
  NAND2_X1 U5979 ( .A1(n7949), .A2(n7948), .ZN(n9396) );
  INV_X1 U5980 ( .A(n9396), .ZN(n4440) );
  NOR3_X1 U5981 ( .A1(n8766), .A2(n4493), .A3(n8859), .ZN(n4495) );
  NAND2_X1 U5982 ( .A1(n4653), .A2(n4298), .ZN(n5227) );
  AND4_X1 U5983 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n8479)
         );
  NOR2_X1 U5984 ( .A1(n8961), .A2(n4841), .ZN(n4351) );
  INV_X1 U5985 ( .A(n4585), .ZN(n4584) );
  NOR2_X1 U5986 ( .A1(n9349), .A2(n4586), .ZN(n4585) );
  NAND2_X1 U5987 ( .A1(n6437), .A2(n6436), .ZN(n9401) );
  INV_X1 U5988 ( .A(n4611), .ZN(n4610) );
  NOR2_X1 U5989 ( .A1(n5602), .A2(n4612), .ZN(n4611) );
  NAND2_X1 U5990 ( .A1(n5307), .A2(n5306), .ZN(n8888) );
  NOR2_X1 U5991 ( .A1(n8766), .A2(n8875), .ZN(n4496) );
  AND2_X1 U5992 ( .A1(n5425), .A2(n8288), .ZN(n4352) );
  AND2_X1 U5993 ( .A1(n6423), .A2(n6422), .ZN(n9130) );
  INV_X1 U5994 ( .A(n9130), .ZN(n9173) );
  AND2_X1 U5995 ( .A1(n7822), .A2(n4768), .ZN(n4353) );
  INV_X1 U5996 ( .A(n4491), .ZN(n8715) );
  NOR2_X1 U5997 ( .A1(n8766), .A2(n4493), .ZN(n4491) );
  INV_X1 U5998 ( .A(n8446), .ZN(n4649) );
  NOR2_X1 U5999 ( .A1(n5570), .A2(n5569), .ZN(n4354) );
  OR2_X1 U6000 ( .A1(n8923), .A2(n4371), .ZN(n4355) );
  AND2_X1 U6001 ( .A1(n4948), .A2(n4947), .ZN(n5413) );
  AND2_X1 U6002 ( .A1(n5384), .A2(n4933), .ZN(n4356) );
  OR2_X1 U6003 ( .A1(n5283), .A2(n4978), .ZN(n4357) );
  OR2_X1 U6004 ( .A1(n8369), .A2(n8372), .ZN(n4358) );
  INV_X1 U6005 ( .A(n4638), .ZN(n5561) );
  NAND2_X1 U6006 ( .A1(n5527), .A2(n4963), .ZN(n5524) );
  NOR2_X1 U6007 ( .A1(n7770), .A2(n7565), .ZN(n4359) );
  INV_X1 U6008 ( .A(n9368), .ZN(n4587) );
  NAND2_X1 U6009 ( .A1(n6246), .A2(n6245), .ZN(n9462) );
  INV_X1 U6010 ( .A(n9462), .ZN(n4449) );
  AOI21_X1 U6011 ( .B1(n8024), .B2(n4557), .A(n4556), .ZN(n4555) );
  AND2_X1 U6012 ( .A1(n6314), .A2(n6313), .ZN(n4360) );
  INV_X1 U6013 ( .A(n9018), .ZN(n4371) );
  AND2_X1 U6014 ( .A1(n9765), .A2(n6479), .ZN(n9018) );
  NAND2_X1 U6015 ( .A1(n6052), .A2(n6051), .ZN(n7428) );
  INV_X1 U6016 ( .A(n4656), .ZN(n4655) );
  OR2_X1 U6017 ( .A1(n7711), .A2(n4657), .ZN(n4656) );
  AND2_X1 U6018 ( .A1(n7392), .A2(n7381), .ZN(n4361) );
  INV_X1 U6019 ( .A(n5397), .ZN(n4713) );
  XNOR2_X1 U6020 ( .A(n5918), .B(n5875), .ZN(n9204) );
  OAI21_X1 U6021 ( .B1(n7009), .B2(n9885), .A(n7008), .ZN(n7610) );
  INV_X1 U6022 ( .A(n7101), .ZN(n6818) );
  NOR2_X1 U6023 ( .A1(n6744), .A2(n7362), .ZN(n4362) );
  AND2_X1 U6024 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n4363) );
  XNOR2_X1 U6025 ( .A(n5881), .B(n5882), .ZN(n7244) );
  INV_X1 U6026 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4431) );
  INV_X1 U6027 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4445) );
  INV_X1 U6028 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n4389) );
  INV_X1 U6029 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n4391) );
  INV_X1 U6030 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n4548) );
  INV_X1 U6031 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7661) );
  AOI21_X1 U6032 ( .B1(n8924), .B2(n9018), .A(n4370), .ZN(n4369) );
  NAND3_X1 U6033 ( .A1(n7854), .A2(n4373), .A3(n4372), .ZN(n4692) );
  NAND2_X1 U6034 ( .A1(n5134), .A2(n4381), .ZN(n4380) );
  OR2_X2 U6035 ( .A1(n6345), .A2(n4295), .ZN(n4392) );
  NAND2_X1 U6036 ( .A1(n4394), .A2(n7873), .ZN(n6221) );
  NAND3_X1 U6037 ( .A1(n5431), .A2(n5430), .A3(n4358), .ZN(n8342) );
  AND2_X1 U6038 ( .A1(n7363), .A2(n4396), .ZN(n4398) );
  INV_X1 U6039 ( .A(n4404), .ZN(n4397) );
  NAND2_X1 U6040 ( .A1(n4399), .A2(n4398), .ZN(n5170) );
  NAND2_X1 U6042 ( .A1(n5190), .A2(n4411), .ZN(n4410) );
  NAND2_X1 U6043 ( .A1(n4410), .A2(n4408), .ZN(n5224) );
  NAND3_X1 U6044 ( .A1(n5263), .A2(n4962), .A3(n4772), .ZN(n5523) );
  NAND4_X1 U6045 ( .A1(n5263), .A2(n4962), .A3(n4772), .A4(n4346), .ZN(n5007)
         );
  OAI21_X1 U6046 ( .B1(n4282), .B2(P2_DATAO_REG_4__SCAN_IN), .A(n4418), .ZN(
        n4858) );
  NAND2_X1 U6047 ( .A1(n4282), .A2(n6578), .ZN(n4418) );
  NAND3_X1 U6048 ( .A1(n4597), .A2(n4425), .A3(n4424), .ZN(n4423) );
  NAND3_X1 U6049 ( .A1(n9275), .A2(n9292), .A3(n4427), .ZN(n4426) );
  AND2_X1 U6050 ( .A1(n9147), .A2(n4437), .ZN(n9117) );
  NAND2_X1 U6051 ( .A1(n9147), .A2(n8201), .ZN(n9137) );
  NAND3_X1 U6052 ( .A1(n4436), .A2(n4435), .A3(n4433), .ZN(n9387) );
  INV_X1 U6053 ( .A(n6511), .ZN(n6282) );
  NAND2_X2 U6054 ( .A1(n9620), .A2(n9624), .ZN(n6511) );
  NAND3_X1 U6055 ( .A1(n9620), .A2(n9624), .A3(n9608), .ZN(n4444) );
  NAND2_X1 U6056 ( .A1(n5616), .A2(n5779), .ZN(n5634) );
  AOI22_X1 U6057 ( .A1(n4459), .A2(n4624), .B1(n4670), .B2(n4460), .ZN(n4458)
         );
  OAI21_X1 U6058 ( .B1(n4670), .B2(n4459), .A(n4457), .ZN(n5096) );
  AOI21_X1 U6059 ( .B1(n4461), .B2(n5083), .A(n4286), .ZN(n4457) );
  NAND2_X1 U6060 ( .A1(n4715), .A2(n4458), .ZN(n4714) );
  NOR2_X1 U6061 ( .A1(n4286), .A2(n4461), .ZN(n4460) );
  NAND2_X1 U6062 ( .A1(n4898), .A2(n4466), .ZN(n4463) );
  NAND2_X1 U6063 ( .A1(n4463), .A2(n4464), .ZN(n4914) );
  OAI21_X1 U6064 ( .B1(n4474), .B2(n4629), .A(n5768), .ZN(n4473) );
  OAI21_X2 U6065 ( .B1(n4474), .B2(n8643), .A(n4472), .ZN(n8585) );
  NAND2_X2 U6066 ( .A1(n8643), .A2(n4629), .ZN(n8620) );
  NAND2_X1 U6067 ( .A1(n4282), .A2(n4479), .ZN(n4478) );
  OAI21_X1 U6068 ( .B1(n4282), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n4478), .ZN(
        n4852) );
  INV_X1 U6069 ( .A(n4487), .ZN(n8625) );
  INV_X1 U6070 ( .A(n4495), .ZN(n8703) );
  INV_X1 U6071 ( .A(n4496), .ZN(n8751) );
  NAND2_X1 U6072 ( .A1(n4505), .A2(n5775), .ZN(n5788) );
  NAND2_X1 U6073 ( .A1(n9639), .A2(n4299), .ZN(n4509) );
  NAND2_X1 U6074 ( .A1(n4509), .A2(n4510), .ZN(n4512) );
  INV_X1 U6075 ( .A(n4513), .ZN(n9637) );
  INV_X1 U6076 ( .A(n4512), .ZN(n9654) );
  AND2_X1 U6077 ( .A1(n5667), .A2(n4514), .ZN(n5670) );
  NAND2_X1 U6078 ( .A1(n4516), .A2(n4515), .ZN(n5667) );
  NAND2_X1 U6079 ( .A1(n4519), .A2(n5836), .ZN(P2_U3244) );
  NAND2_X1 U6080 ( .A1(n4734), .A2(n4735), .ZN(n4520) );
  NAND3_X1 U6081 ( .A1(n5754), .A2(n5753), .A3(n8555), .ZN(n4525) );
  NAND3_X1 U6082 ( .A1(n4601), .A2(n4598), .A3(n4845), .ZN(n5925) );
  XNOR2_X1 U6083 ( .A(n4849), .B(n4848), .ZN(n5019) );
  NAND2_X1 U6084 ( .A1(n5029), .A2(n5925), .ZN(n4849) );
  OAI21_X2 U6085 ( .B1(n6585), .B2(n5046), .A(n4527), .ZN(n9818) );
  MUX2_X1 U6086 ( .A(n5960), .B(P1_REG2_REG_2__SCAN_IN), .S(n6527), .Z(n6514)
         );
  NAND3_X1 U6087 ( .A1(n8025), .A2(n6551), .A3(n8024), .ZN(n8027) );
  OAI21_X1 U6088 ( .B1(n7102), .B2(n4558), .A(n4555), .ZN(n7189) );
  NAND2_X1 U6089 ( .A1(n7102), .A2(n4555), .ZN(n4553) );
  AOI21_X1 U6090 ( .B1(n4555), .B2(n4558), .A(n7148), .ZN(n4554) );
  NAND2_X1 U6091 ( .A1(n7505), .A2(n4559), .ZN(n9542) );
  NAND2_X1 U6092 ( .A1(n9542), .A2(n8074), .ZN(n7733) );
  NAND2_X1 U6093 ( .A1(n7371), .A2(n7395), .ZN(n4561) );
  NAND2_X1 U6094 ( .A1(n7397), .A2(n7395), .ZN(n8070) );
  OR2_X1 U6095 ( .A1(n7371), .A2(n8000), .ZN(n7397) );
  NAND4_X1 U6096 ( .A1(n5840), .A2(n5862), .A3(n5873), .A4(n4566), .ZN(n4565)
         );
  NOR2_X1 U6097 ( .A1(n9196), .A2(n8226), .ZN(n9193) );
  NAND2_X1 U6098 ( .A1(n4571), .A2(n4573), .ZN(n9154) );
  INV_X1 U6099 ( .A(n9196), .ZN(n4572) );
  AOI21_X1 U6100 ( .B1(n9369), .B2(n4581), .A(n4579), .ZN(n9316) );
  NOR2_X2 U6101 ( .A1(n7756), .A2(n9904), .ZN(n9810) );
  AOI21_X2 U6102 ( .B1(n5858), .B2(P1_IR_REG_27__SCAN_IN), .A(n5857), .ZN(
        n5859) );
  NAND2_X1 U6103 ( .A1(n4600), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4599) );
  NAND2_X1 U6104 ( .A1(n5069), .A2(n5068), .ZN(n4670) );
  NAND2_X1 U6105 ( .A1(n5045), .A2(n5044), .ZN(n4602) );
  NAND2_X1 U6106 ( .A1(n4851), .A2(n4850), .ZN(n5045) );
  NAND2_X1 U6107 ( .A1(n8798), .A2(n4606), .ZN(n4604) );
  OAI21_X1 U6108 ( .B1(n8723), .B2(n4618), .A(n4616), .ZN(n8668) );
  NAND2_X1 U6109 ( .A1(n5084), .A2(n4627), .ZN(n4625) );
  NAND2_X2 U6110 ( .A1(n8639), .A2(n5819), .ZN(n8643) );
  NAND2_X1 U6111 ( .A1(n7827), .A2(n4630), .ZN(n9573) );
  XNOR2_X1 U6112 ( .A(n8576), .B(n8575), .ZN(n4632) );
  NAND2_X1 U6113 ( .A1(n8670), .A2(n4636), .ZN(n8661) );
  NAND2_X2 U6114 ( .A1(n5605), .A2(n8555), .ZN(n8670) );
  AND2_X1 U6115 ( .A1(n7321), .A2(n5685), .ZN(n9794) );
  NAND3_X1 U6116 ( .A1(n4826), .A2(n5597), .A3(n7312), .ZN(n4637) );
  INV_X2 U6117 ( .A(n7139), .ZN(n9823) );
  NAND2_X1 U6118 ( .A1(n8447), .A2(n4642), .ZN(n4639) );
  NAND2_X1 U6119 ( .A1(n4639), .A2(n4640), .ZN(n5571) );
  NAND2_X1 U6120 ( .A1(n8447), .A2(n4648), .ZN(n4641) );
  NAND3_X1 U6121 ( .A1(n5061), .A2(n5039), .A3(n7073), .ZN(n8296) );
  NAND2_X1 U6122 ( .A1(n7074), .A2(n7075), .ZN(n7073) );
  NAND2_X1 U6123 ( .A1(n8298), .A2(n4658), .ZN(n4659) );
  NAND2_X1 U6124 ( .A1(n4659), .A2(n4660), .ZN(n7232) );
  NAND2_X1 U6125 ( .A1(n4662), .A2(n8379), .ZN(n7115) );
  NAND2_X1 U6126 ( .A1(n8281), .A2(n4665), .ZN(n5314) );
  AND2_X1 U6127 ( .A1(n5304), .A2(n4667), .ZN(n4982) );
  NAND2_X1 U6128 ( .A1(n5304), .A2(n4338), .ZN(n4983) );
  NAND2_X1 U6129 ( .A1(n7428), .A2(n4671), .ZN(n6074) );
  NAND2_X1 U6130 ( .A1(n8953), .A2(n8954), .ZN(n8952) );
  NAND2_X1 U6131 ( .A1(n4675), .A2(n4673), .ZN(n6509) );
  INV_X1 U6132 ( .A(n4676), .ZN(n4674) );
  NAND2_X1 U6133 ( .A1(n8953), .A2(n4678), .ZN(n4675) );
  AND2_X1 U6134 ( .A1(n6435), .A2(n8954), .ZN(n4678) );
  NAND3_X1 U6135 ( .A1(n6092), .A2(n4685), .A3(n7410), .ZN(n4684) );
  NAND3_X1 U6136 ( .A1(n6092), .A2(n7410), .A3(n4691), .ZN(n4690) );
  NAND2_X1 U6137 ( .A1(n4692), .A2(n4698), .ZN(n4694) );
  NAND3_X1 U6138 ( .A1(n4694), .A2(n9028), .A3(n4344), .ZN(n4693) );
  NAND2_X1 U6139 ( .A1(n4693), .A2(n4695), .ZN(n8969) );
  OAI21_X1 U6140 ( .B1(n9007), .B2(n4702), .A(n4700), .ZN(n8946) );
  OAI21_X1 U6141 ( .B1(n5398), .B2(n5397), .A(n4942), .ZN(n5412) );
  NAND2_X1 U6142 ( .A1(n4883), .A2(n4882), .ZN(n5209) );
  NAND2_X1 U6143 ( .A1(n4883), .A2(n4720), .ZN(n4719) );
  NAND3_X1 U6144 ( .A1(n4733), .A2(n4731), .A3(n4732), .ZN(n4736) );
  NAND4_X1 U6145 ( .A1(n4733), .A2(n4732), .A3(n4731), .A4(n4741), .ZN(n4735)
         );
  NAND3_X1 U6146 ( .A1(n4737), .A2(n5788), .A3(n5787), .ZN(n4731) );
  AOI21_X1 U6147 ( .B1(n4740), .B2(n5795), .A(n5794), .ZN(n4732) );
  NAND2_X1 U6148 ( .A1(n4343), .A2(n5795), .ZN(n4733) );
  NAND2_X1 U6149 ( .A1(n5828), .A2(n4736), .ZN(n4734) );
  INV_X1 U6150 ( .A(n5829), .ZN(n4741) );
  NAND2_X1 U6151 ( .A1(n4742), .A2(n4356), .ZN(n4937) );
  NAND2_X1 U6152 ( .A1(n5802), .A2(n4746), .ZN(n7009) );
  NAND2_X1 U6153 ( .A1(n5674), .A2(n4746), .ZN(n5665) );
  NAND2_X1 U6154 ( .A1(n5661), .A2(n4746), .ZN(n7605) );
  NAND2_X1 U6155 ( .A1(n8666), .A2(n4342), .ZN(n8560) );
  INV_X1 U6156 ( .A(n4758), .ZN(n8758) );
  NOR2_X1 U6157 ( .A1(n8783), .A2(n8763), .ZN(n4760) );
  OR2_X1 U6158 ( .A1(n8338), .A2(n8481), .ZN(n4770) );
  NAND3_X1 U6159 ( .A1(n4298), .A2(n5066), .A3(n4953), .ZN(n5193) );
  INV_X1 U6160 ( .A(n4773), .ZN(n9367) );
  NAND2_X1 U6161 ( .A1(n7731), .A2(n7730), .ZN(n7787) );
  OAI21_X1 U6162 ( .B1(n9191), .B2(n4309), .A(n4796), .ZN(n9178) );
  OAI21_X1 U6163 ( .B1(n7392), .B2(n4801), .A(n4798), .ZN(n9540) );
  INV_X1 U6164 ( .A(n9315), .ZN(n4814) );
  INV_X1 U6165 ( .A(n9333), .ZN(n4815) );
  NAND2_X1 U6166 ( .A1(n5888), .A2(n5890), .ZN(n5851) );
  NAND2_X1 U6167 ( .A1(n5888), .A2(n4819), .ZN(n5893) );
  INV_X1 U6168 ( .A(n8015), .ZN(n9389) );
  OR2_X1 U6169 ( .A1(n8058), .A2(n4304), .ZN(n8059) );
  NAND2_X1 U6170 ( .A1(n4972), .A2(n4965), .ZN(n4970) );
  AND2_X1 U6171 ( .A1(n7181), .A2(n6048), .ZN(n6043) );
  NAND2_X1 U6172 ( .A1(n6047), .A2(n4839), .ZN(n6048) );
  NAND2_X1 U6173 ( .A1(n6091), .A2(n6090), .ZN(n7410) );
  XNOR2_X1 U6174 ( .A(n5635), .B(SI_30_), .ZN(n8244) );
  NAND2_X1 U6175 ( .A1(n5481), .A2(n5480), .ZN(n5483) );
  XNOR2_X1 U6176 ( .A(n5481), .B(n5480), .ZN(n7865) );
  AND2_X1 U6177 ( .A1(n5634), .A2(n5633), .ZN(n5647) );
  OAI21_X1 U6178 ( .B1(n9135), .B2(n9318), .A(n9134), .ZN(n9136) );
  INV_X1 U6179 ( .A(n8492), .ZN(n5594) );
  NAND2_X1 U6180 ( .A1(n5594), .A2(n7272), .ZN(n5802) );
  NAND2_X1 U6181 ( .A1(n8952), .A2(n9014), .ZN(n9016) );
  INV_X1 U6182 ( .A(n7302), .ZN(n7753) );
  XNOR2_X1 U6183 ( .A(n5457), .B(n5456), .ZN(n7847) );
  NAND2_X2 U6184 ( .A1(n5348), .A2(n8433), .ZN(n8437) );
  INV_X1 U6185 ( .A(n6088), .ZN(n6091) );
  NAND2_X1 U6186 ( .A1(n6806), .A2(n6805), .ZN(n6804) );
  INV_X1 U6187 ( .A(n6478), .ZN(n6455) );
  NAND2_X1 U6188 ( .A1(n6478), .A2(n9204), .ZN(n6557) );
  NAND2_X1 U6189 ( .A1(n7302), .A2(n5683), .ZN(n7314) );
  NAND2_X1 U6190 ( .A1(n5678), .A2(n5683), .ZN(n7302) );
  AOI21_X1 U6191 ( .B1(n5854), .B2(n5853), .A(n9517), .ZN(n5858) );
  INV_X1 U6192 ( .A(n9118), .ZN(n9394) );
  INV_X1 U6193 ( .A(n5007), .ZN(n4968) );
  INV_X1 U6194 ( .A(n5899), .ZN(n5900) );
  NAND2_X1 U6195 ( .A1(n5077), .A2(n8295), .ZN(n8298) );
  AOI21_X2 U6196 ( .B1(n7580), .B2(n5812), .A(n5599), .ZN(n7674) );
  INV_X1 U6197 ( .A(n8262), .ZN(n5011) );
  AND2_X1 U6198 ( .A1(n8287), .A2(n8288), .ZN(n8368) );
  INV_X1 U6199 ( .A(n5898), .ZN(n8245) );
  NAND2_X1 U6200 ( .A1(n9126), .A2(n8231), .ZN(n8233) );
  AOI21_X2 U6201 ( .B1(n9367), .B2(n8187), .A(n8186), .ZN(n9348) );
  INV_X1 U6202 ( .A(n7562), .ZN(n7564) );
  INV_X1 U6203 ( .A(n8277), .ZN(n8799) );
  AND2_X1 U6204 ( .A1(n5650), .A2(n7016), .ZN(n4822) );
  AND2_X1 U6205 ( .A1(n8071), .A2(n7396), .ZN(n4823) );
  AND2_X1 U6206 ( .A1(n5120), .A2(n5119), .ZN(n4824) );
  NAND2_X1 U6207 ( .A1(n6506), .A2(n6505), .ZN(n4825) );
  OR2_X2 U6208 ( .A1(n7046), .A2(n7291), .ZN(n4826) );
  OR2_X1 U6209 ( .A1(n5410), .A2(n5409), .ZN(n4827) );
  OR2_X1 U6210 ( .A1(n8720), .A2(n8551), .ZN(n4829) );
  AND2_X1 U6211 ( .A1(n8690), .A2(n8671), .ZN(n4830) );
  AND2_X1 U6212 ( .A1(n9517), .A2(n5855), .ZN(n4831) );
  NAND2_X1 U6213 ( .A1(n5087), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4833) );
  INV_X1 U6214 ( .A(n8028), .ZN(n7382) );
  INV_X1 U6215 ( .A(n9796), .ZN(n7556) );
  AND2_X1 U6216 ( .A1(n4877), .A2(n4876), .ZN(n4834) );
  NAND2_X1 U6217 ( .A1(n6549), .A2(n6548), .ZN(n9725) );
  INV_X1 U6218 ( .A(n9725), .ZN(n9318) );
  AND2_X1 U6219 ( .A1(n6447), .A2(n6446), .ZN(n9152) );
  INV_X1 U6220 ( .A(n9152), .ZN(n9043) );
  INV_X1 U6221 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5875) );
  AND2_X1 U6222 ( .A1(n4897), .A2(n4896), .ZN(n4836) );
  AND2_X1 U6223 ( .A1(n9719), .A2(n9731), .ZN(n4837) );
  NOR2_X1 U6224 ( .A1(n6219), .A2(n7721), .ZN(n4838) );
  AND2_X1 U6225 ( .A1(n7423), .A2(n6042), .ZN(n4839) );
  AND2_X1 U6226 ( .A1(n8488), .A2(n9818), .ZN(n4840) );
  AND2_X1 U6227 ( .A1(n6262), .A2(n6261), .ZN(n4841) );
  AND2_X1 U6228 ( .A1(n5024), .A2(n5023), .ZN(n4842) );
  INV_X1 U6229 ( .A(n5052), .ZN(n5012) );
  NAND2_X1 U6230 ( .A1(n7313), .A2(n7290), .ZN(n4843) );
  NAND2_X1 U6231 ( .A1(n5596), .A2(n7290), .ZN(n5597) );
  NAND2_X1 U6232 ( .A1(n5779), .A2(n5790), .ZN(n5775) );
  INV_X1 U6233 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4959) );
  AND2_X1 U6234 ( .A1(n7294), .A2(n7291), .ZN(n7292) );
  INV_X1 U6235 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4966) );
  NOR2_X1 U6236 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5845) );
  OAI21_X1 U6237 ( .B1(n8492), .B2(n7272), .A(n7254), .ZN(n7008) );
  INV_X1 U6238 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4977) );
  INV_X1 U6239 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5873) );
  INV_X1 U6240 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5199) );
  INV_X1 U6241 ( .A(n5373), .ZN(n4999) );
  OR2_X1 U6242 ( .A1(n7362), .A2(n5794), .ZN(n7262) );
  NAND2_X1 U6243 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  INV_X1 U6244 ( .A(n6351), .ZN(n6349) );
  INV_X1 U6245 ( .A(n6171), .ZN(n5906) );
  INV_X1 U6246 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6093) );
  INV_X1 U6247 ( .A(n7148), .ZN(n7159) );
  NAND2_X1 U6248 ( .A1(n9049), .A2(n9760), .ZN(n7997) );
  INV_X1 U6249 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5878) );
  INV_X1 U6250 ( .A(n5332), .ZN(n4920) );
  AND2_X1 U6251 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  INV_X1 U6252 ( .A(n5465), .ZN(n5464) );
  INV_X1 U6253 ( .A(n5426), .ZN(n5416) );
  XNOR2_X1 U6254 ( .A(n4268), .B(n9885), .ZN(n5038) );
  AND2_X1 U6255 ( .A1(n6870), .A2(n5587), .ZN(n7076) );
  INV_X1 U6256 ( .A(n4284), .ZN(n5518) );
  OAI22_X1 U6257 ( .A1(n8579), .A2(n8277), .B1(n8578), .B2(n8577), .ZN(n8580)
         );
  INV_X1 U6258 ( .A(n9833), .ZN(n5541) );
  NOR2_X1 U6259 ( .A1(n4838), .A2(n6222), .ZN(n6223) );
  NAND2_X1 U6260 ( .A1(n7084), .A2(n7085), .ZN(n7083) );
  INV_X1 U6261 ( .A(n6089), .ZN(n6090) );
  INV_X1 U6262 ( .A(n6997), .ZN(n5976) );
  INV_X1 U6263 ( .A(n9013), .ZN(n9014) );
  NAND2_X1 U6264 ( .A1(n6349), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6360) );
  OR2_X1 U6265 ( .A1(n6232), .A2(n6231), .ZN(n6248) );
  INV_X1 U6266 ( .A(n9401), .ZN(n8201) );
  NAND2_X1 U6267 ( .A1(n6478), .A2(n8172), .ZN(n8166) );
  NAND2_X1 U6268 ( .A1(n9043), .A2(n9720), .ZN(n8237) );
  OR2_X1 U6269 ( .A1(n8166), .A2(n6483), .ZN(n6485) );
  OR2_X1 U6270 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  NAND2_X1 U6271 ( .A1(n4889), .A2(n4888), .ZN(n4892) );
  NAND2_X1 U6272 ( .A1(n5464), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5513) );
  AND2_X1 U6273 ( .A1(n5514), .A2(n8571), .ZN(n8597) );
  OR2_X1 U6274 ( .A1(n5445), .A2(n8343), .ZN(n5465) );
  NAND2_X1 U6275 ( .A1(n8320), .A2(n5396), .ZN(n5410) );
  OR2_X1 U6276 ( .A1(n8445), .A2(n5496), .ZN(n8443) );
  OR2_X1 U6277 ( .A1(n5356), .A2(n5355), .ZN(n5373) );
  INV_X1 U6278 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7706) );
  INV_X1 U6279 ( .A(n9783), .ZN(n9787) );
  OR2_X1 U6280 ( .A1(n5513), .A2(n5512), .ZN(n8571) );
  AND2_X1 U6281 ( .A1(n5561), .A2(n5833), .ZN(n9929) );
  INV_X1 U6282 ( .A(n7575), .ZN(n7576) );
  AND2_X1 U6283 ( .A1(n7017), .A2(n7016), .ZN(n9570) );
  INV_X1 U6284 ( .A(n9868), .ZN(n5559) );
  OR2_X1 U6285 ( .A1(n6416), .A2(n6632), .ZN(n6440) );
  INV_X1 U6286 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6086) );
  OR2_X1 U6287 ( .A1(n4348), .A2(n7838), .ZN(n7872) );
  INV_X1 U6288 ( .A(n9033), .ZN(n9023) );
  INV_X1 U6289 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7530) );
  INV_X1 U6290 ( .A(n9108), .ZN(n9673) );
  INV_X1 U6291 ( .A(n9295), .ZN(n9258) );
  INV_X1 U6292 ( .A(n9455), .ZN(n9305) );
  INV_X1 U6293 ( .A(n9354), .ZN(n9319) );
  OR2_X1 U6294 ( .A1(n8166), .A2(n6753), .ZN(n9328) );
  AND2_X1 U6295 ( .A1(n6559), .A2(n6558), .ZN(n9723) );
  OR2_X1 U6296 ( .A1(n6840), .A2(n8175), .ZN(n9767) );
  NAND2_X1 U6297 ( .A1(n6455), .A2(n8054), .ZN(n6840) );
  AND2_X1 U6298 ( .A1(n4913), .A2(n4912), .ZN(n5281) );
  AND2_X1 U6299 ( .A1(n5465), .A2(n5446), .ZN(n8636) );
  AND2_X1 U6300 ( .A1(n5583), .A2(n5560), .ZN(n5575) );
  AND2_X1 U6301 ( .A1(n5588), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8454) );
  INV_X1 U6302 ( .A(n8445), .ZN(n8460) );
  AND4_X1 U6303 ( .A1(n5343), .A2(n5342), .A3(n5341), .A4(n5340), .ZN(n8764)
         );
  AND2_X1 U6304 ( .A1(n6879), .A2(n6878), .ZN(n9783) );
  INV_X1 U6305 ( .A(n9788), .ZN(n9784) );
  INV_X1 U6306 ( .A(n9570), .ZN(n9803) );
  INV_X1 U6307 ( .A(n8539), .ZN(n9812) );
  OR2_X1 U6308 ( .A1(n9832), .A2(n7003), .ZN(n8678) );
  AND2_X1 U6309 ( .A1(n9865), .A2(n5553), .ZN(n7024) );
  INV_X1 U6310 ( .A(n9947), .ZN(n9909) );
  AND2_X1 U6311 ( .A1(n7005), .A2(n7255), .ZN(n7025) );
  NAND2_X1 U6312 ( .A1(n6870), .A2(n5559), .ZN(n9832) );
  AND2_X1 U6313 ( .A1(n5231), .A2(n5247), .ZN(n7702) );
  INV_X1 U6314 ( .A(n9027), .ZN(n9038) );
  INV_X1 U6315 ( .A(n7244), .ZN(n8175) );
  AND4_X1 U6316 ( .A1(n6279), .A2(n6278), .A3(n6277), .A4(n6276), .ZN(n8941)
         );
  AND2_X1 U6317 ( .A1(n9673), .A2(n6753), .ZN(n9702) );
  INV_X1 U6318 ( .A(n9704), .ZN(n9641) );
  INV_X1 U6319 ( .A(n9204), .ZN(n9736) );
  NAND2_X1 U6320 ( .A1(n8149), .A2(n8060), .ZN(n9155) );
  AOI22_X1 U6321 ( .A1(n9223), .A2(n8195), .B1(n9244), .B2(n9230), .ZN(n9209)
         );
  AND2_X1 U6322 ( .A1(n9289), .A2(n9291), .ZN(n9307) );
  AND2_X1 U6323 ( .A1(n6560), .A2(n6753), .ZN(n9720) );
  INV_X1 U6324 ( .A(n9343), .ZN(n9558) );
  INV_X1 U6325 ( .A(n9487), .ZN(n9765) );
  AND2_X1 U6326 ( .A1(n9723), .A2(n9491), .ZN(n9562) );
  OR2_X1 U6327 ( .A1(n8158), .A2(n8175), .ZN(n9491) );
  INV_X1 U6328 ( .A(n9491), .ZN(n9772) );
  AND2_X1 U6329 ( .A1(n6832), .A2(n6831), .ZN(n6843) );
  AND2_X1 U6330 ( .A1(n6512), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6477) );
  INV_X1 U6331 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5882) );
  INV_X1 U6332 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6226) );
  XNOR2_X1 U6333 ( .A(n5111), .B(n5112), .ZN(n6032) );
  NAND2_X1 U6334 ( .A1(n5830), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9868) );
  INV_X1 U6335 ( .A(n8842), .ZN(n8655) );
  OR2_X1 U6336 ( .A1(n8452), .A2(n8765), .ZN(n8466) );
  OR2_X1 U6337 ( .A1(n8452), .A2(n8277), .ZN(n8465) );
  INV_X1 U6338 ( .A(n8552), .ZN(n8694) );
  INV_X1 U6339 ( .A(n7318), .ZN(n8485) );
  INV_X1 U6340 ( .A(n8529), .ZN(n9786) );
  INV_X2 U6341 ( .A(n9829), .ZN(n9831) );
  NAND2_X1 U6342 ( .A1(n9829), .A2(n9828), .ZN(n8808) );
  INV_X1 U6343 ( .A(n9967), .ZN(n9965) );
  INV_X1 U6344 ( .A(n9951), .ZN(n9949) );
  AND2_X2 U6345 ( .A1(n7025), .A2(n7256), .ZN(n9951) );
  NOR2_X1 U6346 ( .A1(n9833), .A2(n9832), .ZN(n9848) );
  CLKBUF_X1 U6347 ( .A(n9848), .Z(n9869) );
  NAND2_X1 U6348 ( .A1(n5523), .A2(n5526), .ZN(n7870) );
  INV_X1 U6349 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6738) );
  INV_X1 U6350 ( .A(n9415), .ZN(n9182) );
  INV_X1 U6351 ( .A(n9031), .ZN(n9000) );
  INV_X1 U6352 ( .A(n8198), .ZN(n9186) );
  INV_X1 U6353 ( .A(n8941), .ZN(n9309) );
  INV_X1 U6354 ( .A(n9702), .ZN(n9688) );
  OR2_X1 U6355 ( .A1(P1_U3083), .A2(n6539), .ZN(n9112) );
  NAND2_X1 U6356 ( .A1(n9740), .A2(n7143), .ZN(n9365) );
  NAND2_X1 U6357 ( .A1(n7165), .A2(n9142), .ZN(n9740) );
  INV_X1 U6358 ( .A(n9782), .ZN(n9779) );
  OR3_X1 U6359 ( .A1(n9484), .A2(n9483), .A3(n9482), .ZN(n9513) );
  INV_X1 U6360 ( .A(n9774), .ZN(n9773) );
  NAND2_X1 U6361 ( .A1(n9515), .A2(n6734), .ZN(n9748) );
  AND2_X1 U6362 ( .A1(n6513), .A2(n6477), .ZN(n9515) );
  NAND2_X1 U6363 ( .A1(n5887), .A2(n5886), .ZN(n7850) );
  INV_X1 U6364 ( .A(n8172), .ZN(n8054) );
  INV_X1 U6365 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6869) );
  INV_X1 U6366 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6733) );
  INV_X1 U6367 ( .A(n6601), .ZN(n9522) );
  NOR2_X1 U6368 ( .A1(n10003), .A2(n10002), .ZN(n10001) );
  NOR2_X1 U6369 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  NOR2_X2 U6370 ( .A1(n6870), .A2(n9868), .ZN(P2_U3966) );
  AND2_X1 U6371 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4845) );
  AND2_X1 U6372 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4847) );
  INV_X1 U6373 ( .A(SI_1_), .ZN(n4848) );
  NAND2_X1 U6374 ( .A1(n4849), .A2(SI_1_), .ZN(n4850) );
  INV_X1 U6375 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6589) );
  XNOR2_X1 U6376 ( .A(n4852), .B(SI_2_), .ZN(n5044) );
  INV_X1 U6377 ( .A(n4852), .ZN(n4853) );
  NAND2_X1 U6378 ( .A1(n4853), .A2(SI_2_), .ZN(n4854) );
  INV_X1 U6379 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6592) );
  INV_X1 U6380 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6577) );
  XNOR2_X1 U6381 ( .A(n4855), .B(SI_3_), .ZN(n5068) );
  INV_X1 U6382 ( .A(n4855), .ZN(n4856) );
  NAND2_X1 U6383 ( .A1(n4856), .A2(SI_3_), .ZN(n4857) );
  INV_X1 U6384 ( .A(n4858), .ZN(n4859) );
  INV_X1 U6385 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4860) );
  MUX2_X1 U6386 ( .A(n6579), .B(n4860), .S(n6581), .Z(n4861) );
  INV_X1 U6387 ( .A(n4861), .ZN(n4862) );
  MUX2_X1 U6388 ( .A(n6580), .B(n6598), .S(n6581), .Z(n4863) );
  XNOR2_X1 U6389 ( .A(n4863), .B(SI_6_), .ZN(n5112) );
  INV_X1 U6390 ( .A(n4863), .ZN(n4864) );
  MUX2_X1 U6391 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6581), .Z(n4866) );
  XNOR2_X1 U6392 ( .A(n4866), .B(SI_7_), .ZN(n5133) );
  INV_X1 U6393 ( .A(n5133), .ZN(n4865) );
  NAND2_X1 U6394 ( .A1(n4866), .A2(SI_7_), .ZN(n4867) );
  MUX2_X1 U6395 ( .A(n6599), .B(n6086), .S(n6581), .Z(n4869) );
  INV_X1 U6396 ( .A(SI_8_), .ZN(n4868) );
  NAND2_X1 U6397 ( .A1(n4869), .A2(n4868), .ZN(n4872) );
  INV_X1 U6398 ( .A(n4869), .ZN(n4870) );
  NAND2_X1 U6399 ( .A1(n4870), .A2(SI_8_), .ZN(n4871) );
  NAND2_X1 U6400 ( .A1(n4872), .A2(n4871), .ZN(n5150) );
  MUX2_X1 U6401 ( .A(n6730), .B(n6728), .S(n6581), .Z(n4874) );
  INV_X1 U6402 ( .A(SI_9_), .ZN(n4873) );
  NAND2_X1 U6403 ( .A1(n4874), .A2(n4873), .ZN(n4877) );
  INV_X1 U6404 ( .A(n4874), .ZN(n4875) );
  NAND2_X1 U6405 ( .A1(n4875), .A2(SI_9_), .ZN(n4876) );
  MUX2_X1 U6406 ( .A(n6738), .B(n6733), .S(n6581), .Z(n4879) );
  INV_X1 U6407 ( .A(SI_10_), .ZN(n4878) );
  NAND2_X1 U6408 ( .A1(n4879), .A2(n4878), .ZN(n4882) );
  INV_X1 U6409 ( .A(n4879), .ZN(n4880) );
  NAND2_X1 U6410 ( .A1(n4880), .A2(SI_10_), .ZN(n4881) );
  NAND2_X1 U6411 ( .A1(n5192), .A2(n4832), .ZN(n4883) );
  MUX2_X1 U6412 ( .A(n6743), .B(n6741), .S(n6581), .Z(n4884) );
  XNOR2_X1 U6413 ( .A(n4884), .B(SI_11_), .ZN(n5208) );
  INV_X1 U6414 ( .A(n5208), .ZN(n4887) );
  INV_X1 U6415 ( .A(n4884), .ZN(n4885) );
  NAND2_X1 U6416 ( .A1(n4885), .A2(SI_11_), .ZN(n4886) );
  MUX2_X1 U6417 ( .A(n6747), .B(n6749), .S(n6581), .Z(n4889) );
  INV_X1 U6418 ( .A(SI_12_), .ZN(n4888) );
  INV_X1 U6419 ( .A(n4889), .ZN(n4890) );
  NAND2_X1 U6420 ( .A1(n4890), .A2(SI_12_), .ZN(n4891) );
  NAND2_X1 U6421 ( .A1(n4892), .A2(n4891), .ZN(n5225) );
  MUX2_X1 U6422 ( .A(n6792), .B(n6791), .S(n6581), .Z(n4894) );
  INV_X1 U6423 ( .A(SI_13_), .ZN(n4893) );
  INV_X1 U6424 ( .A(n4894), .ZN(n4895) );
  NAND2_X1 U6425 ( .A1(n4895), .A2(SI_13_), .ZN(n4896) );
  MUX2_X1 U6426 ( .A(n6797), .B(n6795), .S(n6581), .Z(n4900) );
  XNOR2_X1 U6427 ( .A(n4900), .B(SI_14_), .ZN(n5261) );
  INV_X1 U6428 ( .A(n5261), .ZN(n4899) );
  INV_X1 U6429 ( .A(n4900), .ZN(n4901) );
  NAND2_X1 U6430 ( .A1(n4901), .A2(SI_14_), .ZN(n4902) );
  MUX2_X1 U6431 ( .A(n6829), .B(n6828), .S(n6581), .Z(n4904) );
  INV_X1 U6432 ( .A(SI_15_), .ZN(n4903) );
  NAND2_X1 U6433 ( .A1(n4904), .A2(n4903), .ZN(n4907) );
  INV_X1 U6434 ( .A(n4904), .ZN(n4905) );
  NAND2_X1 U6435 ( .A1(n4905), .A2(SI_15_), .ZN(n4906) );
  NAND2_X1 U6436 ( .A1(n4907), .A2(n4906), .ZN(n5302) );
  INV_X1 U6437 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n4908) );
  MUX2_X1 U6438 ( .A(n4908), .B(n6869), .S(n6581), .Z(n4910) );
  INV_X1 U6439 ( .A(SI_16_), .ZN(n4909) );
  INV_X1 U6440 ( .A(n4910), .ZN(n4911) );
  NAND2_X1 U6441 ( .A1(n4911), .A2(SI_16_), .ZN(n4912) );
  NAND2_X1 U6442 ( .A1(n4914), .A2(n4913), .ZN(n5316) );
  INV_X1 U6443 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4915) );
  MUX2_X1 U6444 ( .A(n6993), .B(n4915), .S(n6581), .Z(n4916) );
  XNOR2_X1 U6445 ( .A(n4916), .B(SI_17_), .ZN(n5315) );
  INV_X1 U6446 ( .A(n5315), .ZN(n4919) );
  INV_X1 U6447 ( .A(n4916), .ZN(n4917) );
  NAND2_X1 U6448 ( .A1(n4917), .A2(SI_17_), .ZN(n4918) );
  MUX2_X1 U6449 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6581), .Z(n4921) );
  XNOR2_X1 U6450 ( .A(n4921), .B(SI_18_), .ZN(n5332) );
  NAND2_X1 U6451 ( .A1(n5333), .A2(n4920), .ZN(n4923) );
  NAND2_X1 U6452 ( .A1(n4921), .A2(SI_18_), .ZN(n4922) );
  MUX2_X1 U6453 ( .A(n7138), .B(n7141), .S(n6581), .Z(n4925) );
  INV_X1 U6454 ( .A(SI_19_), .ZN(n4924) );
  NAND2_X1 U6455 ( .A1(n4925), .A2(n4924), .ZN(n4928) );
  INV_X1 U6456 ( .A(n4925), .ZN(n4926) );
  NAND2_X1 U6457 ( .A1(n4926), .A2(SI_19_), .ZN(n4927) );
  NAND2_X1 U6458 ( .A1(n4928), .A2(n4927), .ZN(n5349) );
  MUX2_X1 U6459 ( .A(n7252), .B(n7243), .S(n6581), .Z(n4930) );
  INV_X1 U6460 ( .A(SI_20_), .ZN(n4929) );
  NAND2_X1 U6461 ( .A1(n4930), .A2(n4929), .ZN(n4933) );
  INV_X1 U6462 ( .A(n4930), .ZN(n4931) );
  NAND2_X1 U6463 ( .A1(n4931), .A2(SI_20_), .ZN(n4932) );
  MUX2_X1 U6464 ( .A(n7360), .B(n7333), .S(n6581), .Z(n4934) );
  XNOR2_X1 U6465 ( .A(n4934), .B(SI_21_), .ZN(n5384) );
  INV_X1 U6466 ( .A(n4934), .ZN(n4935) );
  NAND2_X1 U6467 ( .A1(n4935), .A2(SI_21_), .ZN(n4936) );
  MUX2_X1 U6468 ( .A(n7464), .B(n7463), .S(n6581), .Z(n4939) );
  INV_X1 U6469 ( .A(SI_22_), .ZN(n4938) );
  NAND2_X1 U6470 ( .A1(n4939), .A2(n4938), .ZN(n4942) );
  INV_X1 U6471 ( .A(n4939), .ZN(n4940) );
  NAND2_X1 U6472 ( .A1(n4940), .A2(SI_22_), .ZN(n4941) );
  NAND2_X1 U6473 ( .A1(n4942), .A2(n4941), .ZN(n5397) );
  INV_X1 U6474 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7596) );
  INV_X1 U6475 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n4943) );
  MUX2_X1 U6476 ( .A(n7596), .B(n4943), .S(n6581), .Z(n4945) );
  INV_X1 U6477 ( .A(SI_23_), .ZN(n4944) );
  NAND2_X1 U6478 ( .A1(n4945), .A2(n4944), .ZN(n4948) );
  INV_X1 U6479 ( .A(n4945), .ZN(n4946) );
  NAND2_X1 U6480 ( .A1(n4946), .A2(SI_23_), .ZN(n4947) );
  MUX2_X1 U6481 ( .A(n7783), .B(n7781), .S(n6581), .Z(n5433) );
  XNOR2_X1 U6482 ( .A(n5433), .B(SI_24_), .ZN(n5432) );
  NAND2_X1 U6483 ( .A1(n5284), .A2(n4955), .ZN(n4978) );
  INV_X1 U6484 ( .A(n4978), .ZN(n4958) );
  NOR2_X1 U6485 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4957) );
  NOR2_X1 U6486 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4956) );
  NAND4_X1 U6487 ( .A1(n4958), .A2(n4957), .A3(n4956), .A4(n5535), .ZN(n4961)
         );
  NAND4_X1 U6488 ( .A1(n6633), .A2(n5532), .A3(n4959), .A4(n4988), .ZN(n4960)
         );
  NOR2_X1 U6489 ( .A1(n4961), .A2(n4960), .ZN(n4962) );
  NOR2_X1 U6490 ( .A1(n4968), .A2(n4967), .ZN(n4969) );
  NAND2_X1 U6491 ( .A1(n4970), .A2(n4969), .ZN(n5576) );
  NAND2_X1 U6492 ( .A1(n5523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4971) );
  NAND2_X1 U6493 ( .A1(n7780), .A2(n5489), .ZN(n4975) );
  OR2_X1 U6494 ( .A1(n5097), .A2(n7783), .ZN(n4974) );
  NOR2_X1 U6495 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4979) );
  INV_X1 U6496 ( .A(n4983), .ZN(n4980) );
  NAND2_X1 U6497 ( .A1(n4980), .A2(n4959), .ZN(n4981) );
  NAND2_X1 U6498 ( .A1(n4983), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6499 ( .A1(n5829), .A2(n7362), .ZN(n4990) );
  NAND2_X1 U6500 ( .A1(n4986), .A2(n4985), .ZN(n4987) );
  INV_X1 U6501 ( .A(n5562), .ZN(n5794) );
  XNOR2_X1 U6502 ( .A(n8842), .B(n5049), .ZN(n5428) );
  INV_X1 U6503 ( .A(n5428), .ZN(n8369) );
  NAND3_X1 U6504 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5121) );
  INV_X1 U6505 ( .A(n5121), .ZN(n4991) );
  NAND2_X1 U6506 ( .A1(n4991), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5142) );
  INV_X1 U6507 ( .A(n5142), .ZN(n4992) );
  NAND2_X1 U6508 ( .A1(n4992), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5160) );
  INV_X1 U6509 ( .A(n5160), .ZN(n4993) );
  NAND2_X1 U6510 ( .A1(n4993), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5180) );
  INV_X1 U6511 ( .A(n5235), .ZN(n4995) );
  NAND2_X1 U6512 ( .A1(n4995), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5251) );
  INV_X1 U6513 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5294) );
  INV_X1 U6514 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8363) );
  INV_X1 U6515 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5355) );
  INV_X1 U6516 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8324) );
  INV_X1 U6517 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8415) );
  INV_X1 U6518 ( .A(n5419), .ZN(n5001) );
  INV_X1 U6519 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5002) );
  NAND2_X1 U6520 ( .A1(n5419), .A2(n5002), .ZN(n5003) );
  NAND2_X1 U6521 ( .A1(n5445), .A2(n5003), .ZN(n8652) );
  INV_X1 U6522 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5004) );
  INV_X1 U6523 ( .A(n5006), .ZN(n8916) );
  NAND2_X1 U6524 ( .A1(n5007), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5008) );
  OR2_X1 U6525 ( .A1(n8652), .A2(n5467), .ZN(n5017) );
  INV_X1 U6526 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U6527 ( .A1(n5010), .A2(n8916), .ZN(n7906) );
  NAND2_X1 U6528 ( .A1(n5011), .A2(n7906), .ZN(n5050) );
  NAND2_X1 U6529 ( .A1(n5087), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5014) );
  AND2_X2 U6530 ( .A1(n8262), .A2(n7906), .ZN(n5052) );
  NAND2_X1 U6531 ( .A1(n5629), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5013) );
  OAI211_X1 U6532 ( .C1(n5518), .C2(n6699), .A(n5014), .B(n5013), .ZN(n5015)
         );
  INV_X1 U6533 ( .A(n5015), .ZN(n5016) );
  NOR2_X1 U6534 ( .A1(n8672), .A2(n5496), .ZN(n5429) );
  INV_X1 U6535 ( .A(n5429), .ZN(n8372) );
  XNOR2_X1 U6536 ( .A(n5019), .B(n5018), .ZN(n6583) );
  NAND2_X1 U6537 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5020) );
  INV_X1 U6538 ( .A(n5021), .ZN(n5022) );
  NAND2_X1 U6539 ( .A1(n5051), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5024) );
  NAND2_X1 U6540 ( .A1(n5052), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5023) );
  NAND2_X1 U6541 ( .A1(n5087), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U6542 ( .A1(n5072), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5025) );
  CLKBUF_X1 U6543 ( .A(n5594), .Z(n7606) );
  XNOR2_X1 U6544 ( .A(n5038), .B(n5036), .ZN(n7074) );
  INV_X1 U6545 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6546 ( .A1(n5028), .A2(n5027), .ZN(n5030) );
  AND2_X1 U6547 ( .A1(n5030), .A2(n5029), .ZN(n8921) );
  MUX2_X1 U6548 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8921), .S(n6877), .Z(n9874) );
  OR2_X1 U6549 ( .A1(n4269), .A2(n9874), .ZN(n5035) );
  NAND2_X1 U6550 ( .A1(n5052), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U6551 ( .A1(n5072), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U6552 ( .A1(n4283), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6553 ( .A1(n5087), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5031) );
  NAND4_X1 U6554 ( .A1(n5034), .A2(n5033), .A3(n5032), .A4(n5031), .ZN(n5593)
         );
  AND2_X1 U6555 ( .A1(n5593), .A2(n9874), .ZN(n7254) );
  NAND2_X1 U6556 ( .A1(n7254), .A2(n5650), .ZN(n8254) );
  AND2_X1 U6557 ( .A1(n5035), .A2(n8254), .ZN(n7075) );
  INV_X1 U6558 ( .A(n5036), .ZN(n5037) );
  NAND2_X1 U6559 ( .A1(n5038), .A2(n5037), .ZN(n5039) );
  NOR2_X1 U6560 ( .A1(n5021), .A2(n5528), .ZN(n5040) );
  MUX2_X1 U6561 ( .A(n5528), .B(n5040), .S(P2_IR_REG_2__SCAN_IN), .Z(n5041) );
  INV_X1 U6562 ( .A(n5041), .ZN(n5043) );
  INV_X1 U6563 ( .A(n5066), .ZN(n5042) );
  NAND2_X1 U6564 ( .A1(n5043), .A2(n5042), .ZN(n6991) );
  XNOR2_X1 U6565 ( .A(n5045), .B(n5044), .ZN(n6588) );
  OR2_X1 U6566 ( .A1(n5046), .A2(n6588), .ZN(n5048) );
  XNOR2_X1 U6567 ( .A(n4269), .B(n4267), .ZN(n5057) );
  NAND2_X1 U6568 ( .A1(n5072), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5056) );
  INV_X1 U6569 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7613) );
  OR2_X1 U6570 ( .A1(n5050), .A2(n7613), .ZN(n5055) );
  NAND2_X1 U6571 ( .A1(n4284), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5054) );
  NOR2_X1 U6572 ( .A1(n4835), .A2(n5496), .ZN(n5058) );
  NAND2_X1 U6573 ( .A1(n5057), .A2(n5058), .ZN(n5062) );
  INV_X1 U6574 ( .A(n5057), .ZN(n8294) );
  INV_X1 U6575 ( .A(n5058), .ZN(n5059) );
  NAND2_X1 U6576 ( .A1(n8294), .A2(n5059), .ZN(n5060) );
  NAND2_X1 U6577 ( .A1(n5062), .A2(n5060), .ZN(n8247) );
  NAND2_X1 U6578 ( .A1(n8296), .A2(n5062), .ZN(n5077) );
  NOR2_X1 U6579 ( .A1(n5066), .A2(n5528), .ZN(n5063) );
  MUX2_X1 U6580 ( .A(n5528), .B(n5063), .S(P2_IR_REG_3__SCAN_IN), .Z(n5064) );
  INV_X1 U6581 ( .A(n5064), .ZN(n5067) );
  INV_X1 U6582 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U6583 ( .A1(n5066), .A2(n5065), .ZN(n5156) );
  NAND2_X1 U6584 ( .A1(n5067), .A2(n5156), .ZN(n6965) );
  XNOR2_X1 U6585 ( .A(n5069), .B(n5068), .ZN(n6591) );
  OR2_X1 U6586 ( .A1(n5046), .A2(n6591), .ZN(n5071) );
  OR2_X1 U6587 ( .A1(n4285), .A2(n6577), .ZN(n5070) );
  OAI211_X1 U6588 ( .C1(n6877), .C2(n6965), .A(n5071), .B(n5070), .ZN(n8301)
         );
  XNOR2_X1 U6589 ( .A(n4269), .B(n7492), .ZN(n5078) );
  NAND2_X1 U6590 ( .A1(n4283), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5076) );
  INV_X1 U6591 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8303) );
  NAND2_X1 U6592 ( .A1(n5072), .A2(n8303), .ZN(n5075) );
  NAND2_X1 U6593 ( .A1(n5052), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U6594 ( .A1(n5087), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5073) );
  NOR2_X1 U6595 ( .A1(n7607), .A2(n5496), .ZN(n5079) );
  XNOR2_X1 U6596 ( .A(n5078), .B(n5079), .ZN(n8295) );
  INV_X1 U6597 ( .A(n5078), .ZN(n5080) );
  NAND2_X1 U6598 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  NAND2_X1 U6599 ( .A1(n5156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5082) );
  XNOR2_X1 U6600 ( .A(n5082), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6888) );
  INV_X1 U6601 ( .A(n6888), .ZN(n6950) );
  XNOR2_X1 U6602 ( .A(n5084), .B(n5083), .ZN(n6586) );
  OR2_X1 U6603 ( .A1(n5046), .A2(n6586), .ZN(n5086) );
  OR2_X1 U6604 ( .A1(n5097), .A2(n6578), .ZN(n5085) );
  OAI211_X1 U6605 ( .C1(n6877), .C2(n6950), .A(n5086), .B(n5085), .ZN(n8387)
         );
  XNOR2_X1 U6606 ( .A(n4269), .B(n8387), .ZN(n8378) );
  XNOR2_X1 U6607 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7520) );
  INV_X1 U6608 ( .A(n7520), .ZN(n8386) );
  NAND2_X1 U6609 ( .A1(n5072), .A2(n8386), .ZN(n5090) );
  NAND2_X1 U6610 ( .A1(n4284), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U6611 ( .A1(n5052), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5088) );
  NOR2_X1 U6612 ( .A1(n7224), .A2(n5496), .ZN(n5091) );
  AND2_X1 U6613 ( .A1(n8378), .A2(n5091), .ZN(n8380) );
  INV_X1 U6614 ( .A(n8378), .ZN(n5093) );
  INV_X1 U6615 ( .A(n5091), .ZN(n5092) );
  NAND2_X1 U6616 ( .A1(n5093), .A2(n5092), .ZN(n8379) );
  OR2_X1 U6617 ( .A1(n5156), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6618 ( .A1(n5094), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5115) );
  XNOR2_X1 U6619 ( .A(n5115), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6905) );
  INV_X1 U6620 ( .A(n6905), .ZN(n6898) );
  OR2_X1 U6621 ( .A1(n4285), .A2(n6579), .ZN(n5098) );
  INV_X1 U6622 ( .A(n9818), .ZN(n7295) );
  XNOR2_X1 U6623 ( .A(n4269), .B(n7295), .ZN(n5106) );
  NAND2_X1 U6624 ( .A1(n4284), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5105) );
  INV_X1 U6625 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U6626 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5099) );
  NAND2_X1 U6627 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  AND2_X1 U6628 ( .A1(n5121), .A2(n5101), .ZN(n9820) );
  NAND2_X1 U6629 ( .A1(n5072), .A2(n9820), .ZN(n5104) );
  NAND2_X1 U6630 ( .A1(n5087), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6631 ( .A1(n5052), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U6632 ( .A1(n8488), .A2(n5650), .ZN(n5107) );
  XNOR2_X1 U6633 ( .A(n5106), .B(n5107), .ZN(n7114) );
  INV_X1 U6634 ( .A(n7114), .ZN(n5110) );
  INV_X1 U6635 ( .A(n5106), .ZN(n5109) );
  INV_X1 U6636 ( .A(n5107), .ZN(n5108) );
  INV_X1 U6637 ( .A(n5046), .ZN(n5113) );
  OR2_X1 U6638 ( .A1(n4285), .A2(n6580), .ZN(n5120) );
  NAND2_X1 U6639 ( .A1(n5115), .A2(n5114), .ZN(n5116) );
  NAND2_X1 U6640 ( .A1(n5116), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5117) );
  INV_X1 U6641 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5154) );
  OR2_X1 U6642 ( .A1(n5117), .A2(n5154), .ZN(n5118) );
  NAND2_X1 U6643 ( .A1(n5117), .A2(n5154), .ZN(n5135) );
  INV_X1 U6644 ( .A(n6921), .ZN(n6913) );
  NAND2_X1 U6645 ( .A1(n5351), .A2(n6921), .ZN(n5119) );
  XNOR2_X1 U6646 ( .A(n4268), .B(n9900), .ZN(n5127) );
  NAND2_X1 U6647 ( .A1(n4283), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6648 ( .A1(n5087), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5124) );
  INV_X1 U6649 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7236) );
  NAND2_X1 U6650 ( .A1(n5121), .A2(n7236), .ZN(n5122) );
  AND2_X1 U6651 ( .A1(n5142), .A2(n5122), .ZN(n7237) );
  NAND2_X1 U6652 ( .A1(n5072), .A2(n7237), .ZN(n5123) );
  NAND2_X1 U6653 ( .A1(n5052), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5126) );
  INV_X1 U6654 ( .A(n8487), .ZN(n7319) );
  OR2_X1 U6655 ( .A1(n7319), .A2(n5496), .ZN(n5128) );
  NAND2_X1 U6656 ( .A1(n5127), .A2(n5128), .ZN(n5132) );
  INV_X1 U6657 ( .A(n5127), .ZN(n5130) );
  INV_X1 U6658 ( .A(n5128), .ZN(n5129) );
  NAND2_X1 U6659 ( .A1(n5130), .A2(n5129), .ZN(n5131) );
  AND2_X1 U6660 ( .A1(n5132), .A2(n5131), .ZN(n7233) );
  XNOR2_X1 U6661 ( .A(n5134), .B(n5133), .ZN(n6065) );
  NAND2_X1 U6662 ( .A1(n6065), .A2(n5113), .ZN(n5140) );
  INV_X1 U6663 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U6664 ( .A1(n5135), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5136) );
  XNOR2_X1 U6665 ( .A(n5136), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U6666 ( .A1(n5351), .A2(n6920), .ZN(n5137) );
  XNOR2_X1 U6667 ( .A(n4269), .B(n9904), .ZN(n5148) );
  NAND2_X1 U6668 ( .A1(n5577), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5147) );
  INV_X1 U6669 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6670 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  AND2_X1 U6671 ( .A1(n5160), .A2(n5143), .ZN(n7308) );
  NAND2_X1 U6672 ( .A1(n5072), .A2(n7308), .ZN(n5146) );
  NAND2_X1 U6673 ( .A1(n5628), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U6674 ( .A1(n5052), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5144) );
  NOR2_X1 U6675 ( .A1(n7553), .A2(n5496), .ZN(n5149) );
  XNOR2_X1 U6676 ( .A(n5148), .B(n5149), .ZN(n7245) );
  XNOR2_X1 U6677 ( .A(n5151), .B(n5150), .ZN(n6602) );
  NAND2_X1 U6678 ( .A1(n6602), .A2(n5489), .ZN(n5159) );
  INV_X1 U6679 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5153) );
  INV_X1 U6680 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5152) );
  NAND4_X1 U6681 ( .A1(n5114), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n5155)
         );
  OR2_X1 U6682 ( .A1(n5156), .A2(n5155), .ZN(n5172) );
  NAND2_X1 U6683 ( .A1(n5172), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5157) );
  XNOR2_X1 U6684 ( .A(n5157), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7030) );
  AOI22_X1 U6685 ( .A1(n5352), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5351), .B2(
        n7030), .ZN(n5158) );
  NAND2_X1 U6686 ( .A1(n5159), .A2(n5158), .ZN(n9806) );
  XNOR2_X1 U6687 ( .A(n5049), .B(n9914), .ZN(n5166) );
  NAND2_X1 U6688 ( .A1(n4284), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5165) );
  INV_X1 U6689 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6914) );
  NAND2_X1 U6690 ( .A1(n5160), .A2(n6914), .ZN(n5161) );
  AND2_X1 U6691 ( .A1(n5180), .A2(n5161), .ZN(n9804) );
  NAND2_X1 U6692 ( .A1(n5072), .A2(n9804), .ZN(n5164) );
  NAND2_X1 U6693 ( .A1(n5628), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U6694 ( .A1(n5052), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5162) );
  NOR2_X1 U6695 ( .A1(n7318), .A2(n5496), .ZN(n5167) );
  XNOR2_X1 U6696 ( .A(n5166), .B(n5167), .ZN(n7363) );
  INV_X1 U6697 ( .A(n5166), .ZN(n5168) );
  NAND2_X1 U6698 ( .A1(n5168), .A2(n5167), .ZN(n5169) );
  NAND2_X1 U6699 ( .A1(n5170), .A2(n5169), .ZN(n7687) );
  INV_X1 U6700 ( .A(n7687), .ZN(n5190) );
  XNOR2_X1 U6701 ( .A(n5171), .B(n4834), .ZN(n6727) );
  NAND2_X1 U6702 ( .A1(n6727), .A2(n5489), .ZN(n5178) );
  OAI21_X1 U6703 ( .B1(n5172), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5173) );
  MUX2_X1 U6704 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5173), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5176) );
  INV_X1 U6705 ( .A(n5174), .ZN(n5175) );
  AOI22_X1 U6706 ( .A1(n5352), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5351), .B2(
        n7128), .ZN(n5177) );
  NAND2_X1 U6707 ( .A1(n5178), .A2(n5177), .ZN(n7690) );
  XNOR2_X1 U6708 ( .A(n7690), .B(n4269), .ZN(n5187) );
  NAND2_X1 U6709 ( .A1(n5577), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6710 ( .A1(n5180), .A2(n5179), .ZN(n5181) );
  AND2_X1 U6711 ( .A1(n5200), .A2(n5181), .ZN(n7585) );
  NAND2_X1 U6712 ( .A1(n5072), .A2(n7585), .ZN(n5184) );
  NAND2_X1 U6713 ( .A1(n5628), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6714 ( .A1(n5052), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5182) );
  NOR2_X1 U6715 ( .A1(n7670), .A2(n5496), .ZN(n5186) );
  OR2_X1 U6716 ( .A1(n5187), .A2(n5186), .ZN(n5191) );
  NAND2_X1 U6717 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  NAND2_X1 U6718 ( .A1(n5191), .A2(n5188), .ZN(n7686) );
  INV_X1 U6719 ( .A(n7686), .ZN(n5189) );
  NAND2_X1 U6720 ( .A1(n6732), .A2(n5489), .ZN(n5198) );
  NOR2_X1 U6721 ( .A1(n5174), .A2(n5528), .ZN(n5194) );
  MUX2_X1 U6722 ( .A(n5528), .B(n5194), .S(P2_IR_REG_10__SCAN_IN), .Z(n5195)
         );
  INV_X1 U6723 ( .A(n5195), .ZN(n5196) );
  AND2_X1 U6724 ( .A1(n5193), .A2(n5196), .ZN(n7341) );
  AOI22_X1 U6725 ( .A1(n5352), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5351), .B2(
        n7341), .ZN(n5197) );
  XNOR2_X1 U6726 ( .A(n9928), .B(n4268), .ZN(n5207) );
  NAND2_X1 U6727 ( .A1(n4284), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6728 ( .A1(n5200), .A2(n5199), .ZN(n5201) );
  AND2_X1 U6729 ( .A1(n5214), .A2(n5201), .ZN(n7679) );
  NAND2_X1 U6730 ( .A1(n5072), .A2(n7679), .ZN(n5204) );
  NAND2_X1 U6731 ( .A1(n5628), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6732 ( .A1(n5052), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5202) );
  NOR2_X1 U6733 ( .A1(n7691), .A2(n5496), .ZN(n5206) );
  XNOR2_X1 U6734 ( .A(n5207), .B(n5206), .ZN(n7711) );
  XNOR2_X1 U6735 ( .A(n5209), .B(n5208), .ZN(n6740) );
  NAND2_X1 U6736 ( .A1(n6740), .A2(n5489), .ZN(n5212) );
  NAND2_X1 U6737 ( .A1(n5193), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5210) );
  XNOR2_X1 U6738 ( .A(n5210), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7473) );
  AOI22_X1 U6739 ( .A1(n5352), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5351), .B2(
        n7473), .ZN(n5211) );
  NAND2_X1 U6740 ( .A1(n5212), .A2(n5211), .ZN(n8427) );
  XNOR2_X1 U6741 ( .A(n8427), .B(n5444), .ZN(n5220) );
  NAND2_X1 U6742 ( .A1(n4284), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5219) );
  INV_X1 U6743 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6744 ( .A1(n5214), .A2(n5213), .ZN(n5215) );
  AND2_X1 U6745 ( .A1(n5235), .A2(n5215), .ZN(n8428) );
  NAND2_X1 U6746 ( .A1(n5072), .A2(n8428), .ZN(n5218) );
  NAND2_X1 U6747 ( .A1(n5629), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6748 ( .A1(n5628), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5216) );
  NOR2_X1 U6749 ( .A1(n8335), .A2(n5496), .ZN(n5221) );
  XNOR2_X1 U6750 ( .A(n5220), .B(n5221), .ZN(n8422) );
  INV_X1 U6751 ( .A(n5220), .ZN(n5222) );
  NAND2_X1 U6752 ( .A1(n5222), .A2(n5221), .ZN(n5223) );
  XNOR2_X1 U6753 ( .A(n5226), .B(n5225), .ZN(n6746) );
  NAND2_X1 U6754 ( .A1(n6746), .A2(n5489), .ZN(n5233) );
  NAND2_X1 U6755 ( .A1(n5227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5230) );
  INV_X1 U6756 ( .A(n5230), .ZN(n5228) );
  NAND2_X1 U6757 ( .A1(n5228), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6758 ( .A1(n5230), .A2(n5229), .ZN(n5247) );
  AOI22_X1 U6759 ( .A1(n5352), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5351), .B2(
        n7702), .ZN(n5232) );
  NAND2_X1 U6760 ( .A1(n5233), .A2(n5232), .ZN(n8338) );
  XNOR2_X1 U6761 ( .A(n8338), .B(n5444), .ZN(n5241) );
  NAND2_X1 U6762 ( .A1(n5577), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5240) );
  INV_X1 U6763 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6764 ( .A1(n5235), .A2(n5234), .ZN(n5236) );
  AND2_X1 U6765 ( .A1(n5251), .A2(n5236), .ZN(n7774) );
  NAND2_X1 U6766 ( .A1(n5072), .A2(n7774), .ZN(n5239) );
  NAND2_X1 U6767 ( .A1(n5628), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6768 ( .A1(n5629), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5237) );
  OR2_X1 U6769 ( .A1(n7830), .A2(n5496), .ZN(n5242) );
  NAND2_X1 U6770 ( .A1(n5241), .A2(n5242), .ZN(n8329) );
  NAND2_X1 U6771 ( .A1(n8331), .A2(n8329), .ZN(n5245) );
  INV_X1 U6772 ( .A(n5241), .ZN(n5244) );
  INV_X1 U6773 ( .A(n5242), .ZN(n5243) );
  NAND2_X1 U6774 ( .A1(n5244), .A2(n5243), .ZN(n8330) );
  NAND2_X1 U6775 ( .A1(n5245), .A2(n8330), .ZN(n8401) );
  NAND2_X1 U6776 ( .A1(n6790), .A2(n5489), .ZN(n5250) );
  NAND2_X1 U6777 ( .A1(n5247), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5248) );
  XNOR2_X1 U6778 ( .A(n5248), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7812) );
  AOI22_X1 U6779 ( .A1(n5352), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5351), .B2(
        n7812), .ZN(n5249) );
  XNOR2_X1 U6780 ( .A(n8894), .B(n5049), .ZN(n5257) );
  NAND2_X1 U6781 ( .A1(n4284), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6782 ( .A1(n5251), .A2(n7706), .ZN(n5252) );
  AND2_X1 U6783 ( .A1(n5269), .A2(n5252), .ZN(n8403) );
  NAND2_X1 U6784 ( .A1(n5072), .A2(n8403), .ZN(n5255) );
  NAND2_X1 U6785 ( .A1(n5629), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6786 ( .A1(n5628), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5253) );
  NOR2_X1 U6787 ( .A1(n8480), .A2(n5496), .ZN(n5258) );
  NAND2_X1 U6788 ( .A1(n5257), .A2(n5258), .ZN(n5275) );
  INV_X1 U6789 ( .A(n5257), .ZN(n8274) );
  INV_X1 U6790 ( .A(n5258), .ZN(n5259) );
  NAND2_X1 U6791 ( .A1(n8274), .A2(n5259), .ZN(n5260) );
  AND2_X1 U6792 ( .A1(n5275), .A2(n5260), .ZN(n8402) );
  XNOR2_X1 U6793 ( .A(n5262), .B(n5261), .ZN(n6794) );
  NAND2_X1 U6794 ( .A1(n6794), .A2(n5489), .ZN(n5267) );
  NOR2_X1 U6795 ( .A1(n5263), .A2(n5528), .ZN(n5264) );
  MUX2_X1 U6796 ( .A(n5528), .B(n5264), .S(P2_IR_REG_14__SCAN_IN), .Z(n5265)
         );
  NOR2_X1 U6797 ( .A1(n5265), .A2(n5304), .ZN(n7891) );
  AOI22_X1 U6798 ( .A1(n5352), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5351), .B2(
        n7891), .ZN(n5266) );
  XNOR2_X1 U6799 ( .A(n9576), .B(n5444), .ZN(n5279) );
  NAND2_X1 U6800 ( .A1(n4284), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5274) );
  INV_X1 U6801 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6802 ( .A1(n5269), .A2(n5268), .ZN(n5270) );
  AND2_X1 U6803 ( .A1(n5295), .A2(n5270), .ZN(n9575) );
  NAND2_X1 U6804 ( .A1(n5072), .A2(n9575), .ZN(n5273) );
  NAND2_X1 U6805 ( .A1(n5628), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6806 ( .A1(n5629), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5271) );
  NOR2_X1 U6807 ( .A1(n8479), .A2(n5496), .ZN(n5277) );
  XNOR2_X1 U6808 ( .A(n5279), .B(n5277), .ZN(n8285) );
  AND2_X1 U6809 ( .A1(n8285), .A2(n5275), .ZN(n5276) );
  INV_X1 U6810 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6811 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  XNOR2_X1 U6812 ( .A(n5282), .B(n5281), .ZN(n6823) );
  NAND2_X1 U6813 ( .A1(n6823), .A2(n5489), .ZN(n5288) );
  NAND2_X1 U6814 ( .A1(n5283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6815 ( .A1(n5285), .A2(n5284), .ZN(n5317) );
  OR2_X1 U6816 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  AOI22_X1 U6817 ( .A1(n5352), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5351), .B2(
        n8503), .ZN(n5287) );
  XNOR2_X1 U6818 ( .A(n8884), .B(n5049), .ZN(n8353) );
  NAND2_X1 U6819 ( .A1(n4284), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5293) );
  INV_X1 U6820 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8498) );
  NAND2_X1 U6821 ( .A1(n5297), .A2(n8498), .ZN(n5289) );
  AND2_X1 U6822 ( .A1(n5321), .A2(n5289), .ZN(n8781) );
  NAND2_X1 U6823 ( .A1(n5072), .A2(n8781), .ZN(n5292) );
  NAND2_X1 U6824 ( .A1(n5628), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6825 ( .A1(n5629), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5290) );
  NOR2_X1 U6826 ( .A1(n8763), .A2(n5496), .ZN(n5309) );
  NAND2_X1 U6827 ( .A1(n4284), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6828 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  AND2_X1 U6829 ( .A1(n5297), .A2(n5296), .ZN(n8793) );
  NAND2_X1 U6830 ( .A1(n5072), .A2(n8793), .ZN(n5300) );
  NAND2_X1 U6831 ( .A1(n5628), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6832 ( .A1(n5629), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5298) );
  NOR2_X1 U6833 ( .A1(n8546), .A2(n5496), .ZN(n8349) );
  XNOR2_X1 U6834 ( .A(n5303), .B(n5302), .ZN(n6827) );
  NAND2_X1 U6835 ( .A1(n6827), .A2(n5489), .ZN(n5307) );
  OR2_X1 U6836 ( .A1(n5304), .A2(n5528), .ZN(n5305) );
  XNOR2_X1 U6837 ( .A(n5305), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7911) );
  AOI22_X1 U6838 ( .A1(n5352), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5351), .B2(
        n7911), .ZN(n5306) );
  XNOR2_X1 U6839 ( .A(n8888), .B(n5049), .ZN(n8348) );
  OAI22_X1 U6840 ( .A1(n8353), .A2(n5309), .B1(n8349), .B2(n8348), .ZN(n5308)
         );
  INV_X1 U6841 ( .A(n8348), .ZN(n8351) );
  INV_X1 U6842 ( .A(n8349), .ZN(n5310) );
  INV_X1 U6843 ( .A(n5309), .ZN(n8352) );
  OAI21_X1 U6844 ( .B1(n8351), .B2(n5310), .A(n8352), .ZN(n5312) );
  NOR2_X1 U6845 ( .A1(n8352), .A2(n5310), .ZN(n5311) );
  AOI22_X1 U6846 ( .A1(n8353), .A2(n5312), .B1(n5311), .B2(n8348), .ZN(n5313)
         );
  NAND2_X1 U6847 ( .A1(n5314), .A2(n5313), .ZN(n8361) );
  XNOR2_X1 U6848 ( .A(n5316), .B(n5315), .ZN(n6951) );
  NAND2_X1 U6849 ( .A1(n6951), .A2(n5489), .ZN(n5320) );
  NAND2_X1 U6850 ( .A1(n5317), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5318) );
  XNOR2_X1 U6851 ( .A(n5318), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7924) );
  AOI22_X1 U6852 ( .A1(n5352), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5351), .B2(
        n7924), .ZN(n5319) );
  XNOR2_X1 U6853 ( .A(n8880), .B(n5049), .ZN(n5327) );
  NAND2_X1 U6854 ( .A1(n5577), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6855 ( .A1(n5321), .A2(n8363), .ZN(n5322) );
  AND2_X1 U6856 ( .A1(n5338), .A2(n5322), .ZN(n8769) );
  NAND2_X1 U6857 ( .A1(n5072), .A2(n8769), .ZN(n5325) );
  NAND2_X1 U6858 ( .A1(n5628), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6859 ( .A1(n5629), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5323) );
  NOR2_X1 U6860 ( .A1(n8749), .A2(n5496), .ZN(n5328) );
  NAND2_X1 U6861 ( .A1(n5327), .A2(n5328), .ZN(n5331) );
  INV_X1 U6862 ( .A(n5327), .ZN(n8436) );
  INV_X1 U6863 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U6864 ( .A1(n8436), .A2(n5329), .ZN(n5330) );
  AND2_X1 U6865 ( .A1(n5331), .A2(n5330), .ZN(n8362) );
  NAND2_X1 U6866 ( .A1(n8435), .A2(n5331), .ZN(n5348) );
  XNOR2_X1 U6867 ( .A(n5333), .B(n5332), .ZN(n7081) );
  NAND2_X1 U6868 ( .A1(n7081), .A2(n5489), .ZN(n5336) );
  NAND2_X1 U6869 ( .A1(n4357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5334) );
  XNOR2_X1 U6870 ( .A(n5334), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8530) );
  AOI22_X1 U6871 ( .A1(n5352), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5351), .B2(
        n8530), .ZN(n5335) );
  XNOR2_X1 U6872 ( .A(n8755), .B(n5444), .ZN(n5344) );
  INV_X1 U6873 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6874 ( .A1(n5338), .A2(n5337), .ZN(n5339) );
  AND2_X1 U6875 ( .A1(n5356), .A2(n5339), .ZN(n8752) );
  NAND2_X1 U6876 ( .A1(n8752), .A2(n5072), .ZN(n5343) );
  NAND2_X1 U6877 ( .A1(n5577), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6878 ( .A1(n5628), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6879 ( .A1(n5629), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5340) );
  NOR2_X1 U6880 ( .A1(n8764), .A2(n5496), .ZN(n5345) );
  NAND2_X1 U6881 ( .A1(n5344), .A2(n5345), .ZN(n5362) );
  INV_X1 U6882 ( .A(n5344), .ZN(n8307) );
  INV_X1 U6883 ( .A(n5345), .ZN(n5346) );
  NAND2_X1 U6884 ( .A1(n8307), .A2(n5346), .ZN(n5347) );
  AND2_X1 U6885 ( .A1(n5362), .A2(n5347), .ZN(n8433) );
  XNOR2_X1 U6886 ( .A(n5350), .B(n5349), .ZN(n7137) );
  NAND2_X1 U6887 ( .A1(n7137), .A2(n5489), .ZN(n5354) );
  AOI22_X1 U6888 ( .A1(n5352), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9823), .B2(
        n5351), .ZN(n5353) );
  XNOR2_X1 U6889 ( .A(n8869), .B(n5049), .ZN(n5364) );
  NAND2_X1 U6890 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U6891 ( .A1(n5373), .A2(n5357), .ZN(n8734) );
  NAND2_X1 U6892 ( .A1(n4284), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6893 ( .A1(n5628), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5358) );
  AND2_X1 U6894 ( .A1(n5359), .A2(n5358), .ZN(n5361) );
  NAND2_X1 U6895 ( .A1(n5629), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5360) );
  OAI211_X1 U6896 ( .C1(n8734), .C2(n5467), .A(n5361), .B(n5360), .ZN(n8549)
         );
  NAND2_X1 U6897 ( .A1(n8549), .A2(n5650), .ZN(n5365) );
  XNOR2_X1 U6898 ( .A(n5364), .B(n5365), .ZN(n8315) );
  AND2_X1 U6899 ( .A1(n8315), .A2(n5362), .ZN(n5363) );
  INV_X1 U6900 ( .A(n5364), .ZN(n5366) );
  NAND2_X1 U6901 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  XNOR2_X1 U6902 ( .A(n5369), .B(n5368), .ZN(n7242) );
  NAND2_X1 U6903 ( .A1(n7242), .A2(n5489), .ZN(n5371) );
  OR2_X1 U6904 ( .A1(n4285), .A2(n7252), .ZN(n5370) );
  XNOR2_X1 U6905 ( .A(n8863), .B(n5049), .ZN(n5378) );
  INV_X1 U6906 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6907 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  NAND2_X1 U6908 ( .A1(n5388), .A2(n5374), .ZN(n8717) );
  OR2_X1 U6909 ( .A1(n8717), .A2(n5467), .ZN(n5377) );
  AOI22_X1 U6910 ( .A1(n4284), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5087), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6911 ( .A1(n5629), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5375) );
  NOR2_X1 U6912 ( .A1(n8551), .A2(n5496), .ZN(n5379) );
  NAND2_X1 U6913 ( .A1(n5378), .A2(n5379), .ZN(n5383) );
  INV_X1 U6914 ( .A(n5378), .ZN(n8319) );
  INV_X1 U6915 ( .A(n5379), .ZN(n5380) );
  NAND2_X1 U6916 ( .A1(n8319), .A2(n5380), .ZN(n5381) );
  NAND2_X1 U6917 ( .A1(n5383), .A2(n5381), .ZN(n8396) );
  XNOR2_X1 U6918 ( .A(n5385), .B(n5384), .ZN(n7332) );
  NAND2_X1 U6919 ( .A1(n7332), .A2(n5489), .ZN(n5387) );
  OR2_X1 U6920 ( .A1(n5097), .A2(n7360), .ZN(n5386) );
  XNOR2_X1 U6921 ( .A(n8706), .B(n5444), .ZN(n5395) );
  NAND2_X1 U6922 ( .A1(n5388), .A2(n8324), .ZN(n5389) );
  NAND2_X1 U6923 ( .A1(n5400), .A2(n5389), .ZN(n8323) );
  OR2_X1 U6924 ( .A1(n8323), .A2(n5467), .ZN(n5392) );
  AOI22_X1 U6925 ( .A1(n4284), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5628), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6926 ( .A1(n5629), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6927 ( .A1(n8694), .A2(n5650), .ZN(n5393) );
  XNOR2_X1 U6928 ( .A(n5395), .B(n5393), .ZN(n8317) );
  INV_X1 U6929 ( .A(n5393), .ZN(n5394) );
  NAND2_X1 U6930 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  OR2_X1 U6931 ( .A1(n4285), .A2(n7464), .ZN(n5399) );
  XNOR2_X1 U6932 ( .A(n8853), .B(n5444), .ZN(n5408) );
  XNOR2_X1 U6933 ( .A(n5410), .B(n5408), .ZN(n8412) );
  NAND2_X1 U6934 ( .A1(n5400), .A2(n8415), .ZN(n5401) );
  NAND2_X1 U6935 ( .A1(n5417), .A2(n5401), .ZN(n8416) );
  INV_X1 U6936 ( .A(n8416), .ZN(n8688) );
  NAND2_X1 U6937 ( .A1(n8688), .A2(n5072), .ZN(n5407) );
  INV_X1 U6938 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6939 ( .A1(n5087), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6940 ( .A1(n5629), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5402) );
  OAI211_X1 U6941 ( .C1(n5518), .C2(n5404), .A(n5403), .B(n5402), .ZN(n5405)
         );
  INV_X1 U6942 ( .A(n5405), .ZN(n5406) );
  INV_X1 U6943 ( .A(n8671), .ZN(n8476) );
  NAND2_X1 U6944 ( .A1(n8476), .A2(n5650), .ZN(n8411) );
  NAND2_X1 U6945 ( .A1(n8412), .A2(n8411), .ZN(n5411) );
  INV_X1 U6946 ( .A(n5408), .ZN(n5409) );
  NAND2_X1 U6947 ( .A1(n7593), .A2(n5489), .ZN(n5415) );
  OR2_X1 U6948 ( .A1(n5097), .A2(n7596), .ZN(n5414) );
  XNOR2_X1 U6949 ( .A(n8848), .B(n5049), .ZN(n5426) );
  INV_X1 U6950 ( .A(n8672), .ZN(n8475) );
  INV_X1 U6951 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U6952 ( .A1(n5417), .A2(n8289), .ZN(n5418) );
  NAND2_X1 U6953 ( .A1(n5419), .A2(n5418), .ZN(n8679) );
  OR2_X1 U6954 ( .A1(n8679), .A2(n5467), .ZN(n5424) );
  INV_X1 U6955 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6678) );
  NAND2_X1 U6956 ( .A1(n5577), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6957 ( .A1(n5628), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5420) );
  OAI211_X1 U6958 ( .C1(n6678), .C2(n5012), .A(n5421), .B(n5420), .ZN(n5422)
         );
  INV_X1 U6959 ( .A(n5422), .ZN(n5423) );
  NAND2_X1 U6960 ( .A1(n5424), .A2(n5423), .ZN(n8695) );
  AND2_X1 U6961 ( .A1(n8695), .A2(n5650), .ZN(n8288) );
  NAND2_X1 U6962 ( .A1(n8287), .A2(n4352), .ZN(n5431) );
  OAI21_X1 U6963 ( .B1(n5429), .B2(n5428), .A(n8367), .ZN(n5430) );
  INV_X1 U6964 ( .A(n5432), .ZN(n5436) );
  INV_X1 U6965 ( .A(n5433), .ZN(n5434) );
  NAND2_X1 U6966 ( .A1(n5434), .A2(SI_24_), .ZN(n5435) );
  INV_X1 U6967 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7848) );
  INV_X1 U6968 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7852) );
  MUX2_X1 U6969 ( .A(n7848), .B(n7852), .S(n6581), .Z(n5439) );
  INV_X1 U6970 ( .A(SI_25_), .ZN(n5438) );
  NAND2_X1 U6971 ( .A1(n5439), .A2(n5438), .ZN(n5455) );
  INV_X1 U6972 ( .A(n5439), .ZN(n5440) );
  NAND2_X1 U6973 ( .A1(n5440), .A2(SI_25_), .ZN(n5441) );
  NAND2_X1 U6974 ( .A1(n5455), .A2(n5441), .ZN(n5456) );
  NAND2_X1 U6975 ( .A1(n7847), .A2(n5489), .ZN(n5443) );
  OR2_X1 U6976 ( .A1(n4285), .A2(n7848), .ZN(n5442) );
  XNOR2_X1 U6977 ( .A(n8838), .B(n5444), .ZN(n8444) );
  INV_X1 U6978 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U6979 ( .A1(n5445), .A2(n8343), .ZN(n5446) );
  NAND2_X1 U6980 ( .A1(n8636), .A2(n5072), .ZN(n5452) );
  INV_X1 U6981 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6982 ( .A1(n5087), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U6983 ( .A1(n5629), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5447) );
  OAI211_X1 U6984 ( .C1(n5518), .C2(n5449), .A(n5448), .B(n5447), .ZN(n5450)
         );
  INV_X1 U6985 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U6986 ( .A1(n8561), .A2(n5650), .ZN(n5453) );
  NOR2_X1 U6987 ( .A1(n8444), .A2(n5453), .ZN(n5454) );
  AOI21_X1 U6988 ( .B1(n8444), .B2(n5453), .A(n5454), .ZN(n8341) );
  INV_X1 U6989 ( .A(n5454), .ZN(n5478) );
  INV_X1 U6990 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7868) );
  INV_X1 U6991 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7866) );
  MUX2_X1 U6992 ( .A(n7868), .B(n7866), .S(n6581), .Z(n5459) );
  INV_X1 U6993 ( .A(SI_26_), .ZN(n5458) );
  NAND2_X1 U6994 ( .A1(n5459), .A2(n5458), .ZN(n5482) );
  INV_X1 U6995 ( .A(n5459), .ZN(n5460) );
  NAND2_X1 U6996 ( .A1(n5460), .A2(SI_26_), .ZN(n5461) );
  NAND2_X1 U6997 ( .A1(n7865), .A2(n5489), .ZN(n5463) );
  OR2_X1 U6998 ( .A1(n4285), .A2(n7868), .ZN(n5462) );
  XNOR2_X1 U6999 ( .A(n8834), .B(n5049), .ZN(n5474) );
  INV_X1 U7000 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U7001 ( .A1(n5465), .A2(n8451), .ZN(n5466) );
  NAND2_X1 U7002 ( .A1(n5513), .A2(n5466), .ZN(n8626) );
  INV_X1 U7003 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7004 ( .A1(n5087), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7005 ( .A1(n5629), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5468) );
  OAI211_X1 U7006 ( .C1(n5518), .C2(n5470), .A(n5469), .B(n5468), .ZN(n5471)
         );
  INV_X1 U7007 ( .A(n5471), .ZN(n5472) );
  NOR2_X1 U7008 ( .A1(n8563), .A2(n5496), .ZN(n5475) );
  NAND2_X1 U7009 ( .A1(n5474), .A2(n5475), .ZN(n5479) );
  INV_X1 U7010 ( .A(n5474), .ZN(n8265) );
  INV_X1 U7011 ( .A(n5475), .ZN(n5476) );
  NAND2_X1 U7012 ( .A1(n8265), .A2(n5476), .ZN(n5477) );
  NAND2_X1 U7013 ( .A1(n5479), .A2(n5477), .ZN(n8446) );
  INV_X1 U7014 ( .A(n5479), .ZN(n5502) );
  INV_X1 U7015 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7901) );
  INV_X1 U7016 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5484) );
  MUX2_X1 U7017 ( .A(n7901), .B(n5484), .S(n6581), .Z(n5486) );
  INV_X1 U7018 ( .A(SI_27_), .ZN(n5485) );
  NAND2_X1 U7019 ( .A1(n5486), .A2(n5485), .ZN(n5506) );
  INV_X1 U7020 ( .A(n5486), .ZN(n5487) );
  NAND2_X1 U7021 ( .A1(n5487), .A2(SI_27_), .ZN(n5488) );
  NAND2_X1 U7022 ( .A1(n7884), .A2(n5489), .ZN(n5491) );
  OR2_X1 U7023 ( .A1(n4285), .A2(n7901), .ZN(n5490) );
  XNOR2_X1 U7024 ( .A(n8828), .B(n5049), .ZN(n5497) );
  XNOR2_X1 U7025 ( .A(n5513), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8607) );
  INV_X1 U7026 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U7027 ( .A1(n5577), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7028 ( .A1(n5629), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5492) );
  OAI211_X1 U7029 ( .C1(n5494), .C2(n5050), .A(n5493), .B(n5492), .ZN(n5495)
         );
  NOR2_X1 U7030 ( .A1(n8588), .A2(n5496), .ZN(n5498) );
  NAND2_X1 U7031 ( .A1(n5497), .A2(n5498), .ZN(n5503) );
  INV_X1 U7032 ( .A(n5497), .ZN(n5500) );
  INV_X1 U7033 ( .A(n5498), .ZN(n5499) );
  NAND2_X1 U7034 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  INV_X1 U7035 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8242) );
  INV_X1 U7036 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5508) );
  MUX2_X1 U7037 ( .A(n8242), .B(n5508), .S(n6581), .Z(n5610) );
  XNOR2_X1 U7038 ( .A(n5610), .B(SI_28_), .ZN(n5607) );
  NAND2_X1 U7039 ( .A1(n7903), .A2(n5489), .ZN(n5510) );
  OR2_X1 U7040 ( .A1(n4285), .A2(n8242), .ZN(n5509) );
  INV_X1 U7041 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8269) );
  INV_X1 U7042 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5511) );
  OAI21_X1 U7043 ( .B1(n5513), .B2(n8269), .A(n5511), .ZN(n5514) );
  NAND2_X1 U7044 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5512) );
  NAND2_X1 U7045 ( .A1(n8597), .A2(n5072), .ZN(n5521) );
  INV_X1 U7046 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7047 ( .A1(n5628), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7048 ( .A1(n5629), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5515) );
  OAI211_X1 U7049 ( .C1(n5518), .C2(n5517), .A(n5516), .B(n5515), .ZN(n5519)
         );
  INV_X1 U7050 ( .A(n5519), .ZN(n5520) );
  NOR2_X1 U7051 ( .A1(n8579), .A2(n5496), .ZN(n5522) );
  XNOR2_X1 U7052 ( .A(n5522), .B(n5049), .ZN(n5567) );
  INV_X1 U7053 ( .A(n5567), .ZN(n5568) );
  NAND2_X1 U7054 ( .A1(n5524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5525) );
  MUX2_X1 U7055 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5525), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5526) );
  INV_X1 U7056 ( .A(n7870), .ZN(n5540) );
  NOR2_X1 U7057 ( .A1(n5527), .A2(n5528), .ZN(n5529) );
  MUX2_X1 U7058 ( .A(n5528), .B(n5529), .S(P2_IR_REG_25__SCAN_IN), .Z(n5530)
         );
  INV_X1 U7059 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U7060 ( .A1(n5531), .A2(n5524), .ZN(n7849) );
  INV_X1 U7061 ( .A(P2_B_REG_SCAN_IN), .ZN(n5537) );
  XOR2_X1 U7062 ( .A(n7785), .B(n5537), .Z(n5538) );
  NAND2_X1 U7063 ( .A1(n7849), .A2(n5538), .ZN(n5539) );
  NAND2_X1 U7064 ( .A1(n7849), .A2(n7870), .ZN(n9867) );
  NOR4_X1 U7065 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5550) );
  INV_X1 U7066 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9842) );
  INV_X1 U7067 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9840) );
  INV_X1 U7068 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9861) );
  INV_X1 U7069 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9864) );
  NAND4_X1 U7070 ( .A1(n9842), .A2(n9840), .A3(n9861), .A4(n9864), .ZN(n5547)
         );
  NOR4_X1 U7071 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5545) );
  NOR4_X1 U7072 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5544) );
  NOR4_X1 U7073 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5543) );
  NOR4_X1 U7074 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5542) );
  NAND4_X1 U7075 ( .A1(n5545), .A2(n5544), .A3(n5543), .A4(n5542), .ZN(n5546)
         );
  NOR4_X1 U7076 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n5547), .A4(n5546), .ZN(n5549) );
  NOR4_X1 U7077 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5548) );
  NAND3_X1 U7078 ( .A1(n5550), .A2(n5549), .A3(n5548), .ZN(n5551) );
  INV_X1 U7079 ( .A(n7259), .ZN(n5554) );
  NAND2_X1 U7080 ( .A1(n7785), .A2(n7870), .ZN(n9865) );
  INV_X1 U7081 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7082 ( .A1(n9833), .A2(n5552), .ZN(n5553) );
  NAND2_X1 U7083 ( .A1(n5554), .A2(n7024), .ZN(n5555) );
  NOR2_X1 U7084 ( .A1(n7255), .A2(n5555), .ZN(n5583) );
  OR2_X1 U7085 ( .A1(n5556), .A2(n6633), .ZN(n5557) );
  NAND2_X1 U7086 ( .A1(n5558), .A2(n5557), .ZN(n5830) );
  INV_X1 U7087 ( .A(n9832), .ZN(n5560) );
  AND2_X1 U7088 ( .A1(n5794), .A2(n5561), .ZN(n9819) );
  NAND2_X1 U7089 ( .A1(n5575), .A2(n9819), .ZN(n5563) );
  NAND2_X1 U7090 ( .A1(n9905), .A2(n9823), .ZN(n7003) );
  NOR3_X1 U7091 ( .A1(n8599), .A2(n8469), .A3(n5568), .ZN(n5564) );
  AOI21_X1 U7092 ( .B1(n8599), .B2(n5568), .A(n5564), .ZN(n5573) );
  INV_X1 U7093 ( .A(n5585), .ZN(n5833) );
  NAND2_X1 U7094 ( .A1(n5565), .A2(n5662), .ZN(n6750) );
  INV_X1 U7095 ( .A(n6750), .ZN(n6873) );
  NOR2_X1 U7096 ( .A1(n9929), .A2(n6873), .ZN(n5566) );
  OAI21_X1 U7097 ( .B1(n8599), .B2(n8458), .A(n8445), .ZN(n5572) );
  NOR3_X1 U7098 ( .A1(n8599), .A2(n5567), .A3(n8469), .ZN(n5570) );
  NOR2_X1 U7099 ( .A1(n8822), .A2(n5568), .ZN(n5569) );
  OAI211_X1 U7100 ( .C1(n5574), .C2(n5573), .A(n5572), .B(n5571), .ZN(n5592)
         );
  NAND2_X1 U7101 ( .A1(n5575), .A2(n5585), .ZN(n8452) );
  OR2_X2 U7102 ( .A1(n6750), .A2(n5576), .ZN(n8277) );
  INV_X1 U7103 ( .A(n8571), .ZN(n5581) );
  INV_X1 U7104 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U7105 ( .A1(n5577), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7106 ( .A1(n5629), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5578) );
  OAI211_X1 U7107 ( .C1(n8572), .C2(n5050), .A(n5579), .B(n5578), .ZN(n5580)
         );
  AOI21_X1 U7108 ( .B1(n5581), .B2(n5072), .A(n5580), .ZN(n8587) );
  OAI22_X1 U7109 ( .A1(n8588), .A2(n8465), .B1(n8466), .B2(n8587), .ZN(n5582)
         );
  INV_X1 U7110 ( .A(n5582), .ZN(n5590) );
  INV_X1 U7111 ( .A(n5583), .ZN(n5584) );
  NAND2_X1 U7112 ( .A1(n5584), .A2(n7003), .ZN(n7077) );
  OAI21_X1 U7113 ( .B1(n6750), .B2(n5585), .A(n5830), .ZN(n5586) );
  INV_X1 U7114 ( .A(n5586), .ZN(n5587) );
  NAND2_X1 U7115 ( .A1(n7077), .A2(n7076), .ZN(n5588) );
  AOI22_X1 U7116 ( .A1(n8454), .A2(n8597), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5589) );
  AND2_X1 U7117 ( .A1(n5590), .A2(n5589), .ZN(n5591) );
  NAND2_X1 U7118 ( .A1(n5592), .A2(n5591), .ZN(P2_U3222) );
  INV_X1 U7119 ( .A(n4835), .ZN(n8491) );
  NAND2_X1 U7120 ( .A1(n4835), .A2(n4267), .ZN(n5673) );
  INV_X1 U7121 ( .A(n5593), .ZN(n5659) );
  NAND2_X1 U7122 ( .A1(n9877), .A2(n5802), .ZN(n5661) );
  NAND2_X1 U7123 ( .A1(n7607), .A2(n8301), .ZN(n5668) );
  INV_X1 U7124 ( .A(n7607), .ZN(n8490) );
  NAND2_X1 U7125 ( .A1(n8490), .A2(n7492), .ZN(n5657) );
  NAND2_X1 U7126 ( .A1(n5668), .A2(n5657), .ZN(n7014) );
  INV_X1 U7127 ( .A(n7014), .ZN(n5808) );
  NAND2_X1 U7128 ( .A1(n7015), .A2(n5808), .ZN(n5595) );
  NAND2_X1 U7129 ( .A1(n5595), .A2(n5668), .ZN(n7046) );
  NAND2_X1 U7130 ( .A1(n7224), .A2(n8387), .ZN(n5669) );
  INV_X1 U7131 ( .A(n7224), .ZN(n8489) );
  NAND2_X1 U7132 ( .A1(n7215), .A2(n8489), .ZN(n7220) );
  NAND2_X1 U7133 ( .A1(n5669), .A2(n7220), .ZN(n7291) );
  NAND2_X1 U7134 ( .A1(n8488), .A2(n7295), .ZN(n7214) );
  INV_X1 U7135 ( .A(n7314), .ZN(n5596) );
  NAND2_X1 U7136 ( .A1(n7553), .A2(n9904), .ZN(n5684) );
  INV_X1 U7137 ( .A(n7553), .ZN(n8486) );
  NAND2_X1 U7138 ( .A1(n8486), .A2(n7552), .ZN(n5685) );
  INV_X1 U7139 ( .A(n8488), .ZN(n7296) );
  NAND2_X1 U7140 ( .A1(n7296), .A2(n9818), .ZN(n7746) );
  AND2_X1 U7141 ( .A1(n7746), .A2(n5683), .ZN(n7313) );
  NAND2_X1 U7142 ( .A1(n4843), .A2(n5597), .ZN(n5598) );
  NAND2_X1 U7143 ( .A1(n7318), .A2(n9806), .ZN(n5689) );
  NAND2_X1 U7144 ( .A1(n9914), .A2(n8485), .ZN(n5688) );
  NAND2_X1 U7145 ( .A1(n9794), .A2(n9796), .ZN(n9795) );
  NAND2_X1 U7146 ( .A1(n9795), .A2(n5689), .ZN(n7580) );
  OR2_X1 U7147 ( .A1(n7690), .A2(n7670), .ZN(n5698) );
  NAND2_X1 U7148 ( .A1(n7690), .A2(n7670), .ZN(n5692) );
  NAND2_X1 U7149 ( .A1(n5698), .A2(n5692), .ZN(n7579) );
  INV_X1 U7150 ( .A(n7579), .ZN(n5812) );
  INV_X1 U7151 ( .A(n5692), .ZN(n5599) );
  NAND2_X1 U7152 ( .A1(n9928), .A2(n7691), .ZN(n5696) );
  NAND2_X1 U7153 ( .A1(n5697), .A2(n5696), .ZN(n7668) );
  INV_X1 U7154 ( .A(n7668), .ZN(n7673) );
  NAND2_X1 U7155 ( .A1(n7674), .A2(n7673), .ZN(n7672) );
  NAND2_X1 U7156 ( .A1(n7672), .A2(n5697), .ZN(n7549) );
  NAND2_X1 U7157 ( .A1(n8427), .A2(n8335), .ZN(n5801) );
  NAND2_X1 U7158 ( .A1(n7549), .A2(n5801), .ZN(n7766) );
  OR2_X1 U7159 ( .A1(n8338), .A2(n7830), .ZN(n5800) );
  OR2_X1 U7160 ( .A1(n8427), .A2(n8335), .ZN(n7765) );
  AND2_X1 U7161 ( .A1(n5800), .A2(n7765), .ZN(n5705) );
  NAND2_X1 U7162 ( .A1(n7766), .A2(n5705), .ZN(n5600) );
  NAND2_X1 U7163 ( .A1(n8338), .A2(n7830), .ZN(n5799) );
  NAND2_X1 U7164 ( .A1(n5600), .A2(n5799), .ZN(n7828) );
  OR2_X1 U7165 ( .A1(n8894), .A2(n8480), .ZN(n5712) );
  NAND2_X1 U7166 ( .A1(n8894), .A2(n8480), .ZN(n5711) );
  XNOR2_X1 U7167 ( .A(n9576), .B(n8479), .ZN(n9578) );
  OR2_X1 U7168 ( .A1(n9576), .A2(n8479), .ZN(n5601) );
  NAND2_X2 U7169 ( .A1(n9573), .A2(n5601), .ZN(n8798) );
  OR2_X1 U7170 ( .A1(n8888), .A2(n8546), .ZN(n5721) );
  NAND2_X1 U7171 ( .A1(n8888), .A2(n8546), .ZN(n5722) );
  NAND2_X1 U7172 ( .A1(n5721), .A2(n5722), .ZN(n8797) );
  NAND2_X1 U7173 ( .A1(n8884), .A2(n8763), .ZN(n5724) );
  INV_X1 U7174 ( .A(n5724), .ZN(n5602) );
  OR2_X1 U7175 ( .A1(n8884), .A2(n8763), .ZN(n5725) );
  NAND2_X1 U7176 ( .A1(n8880), .A2(n8749), .ZN(n5732) );
  INV_X1 U7177 ( .A(n8764), .ZN(n8477) );
  NAND2_X1 U7178 ( .A1(n8875), .A2(n8764), .ZN(n5796) );
  OAI21_X2 U7179 ( .B1(n8747), .B2(n5798), .A(n5796), .ZN(n8738) );
  INV_X1 U7180 ( .A(n8549), .ZN(n8750) );
  OR2_X1 U7181 ( .A1(n8869), .A2(n8750), .ZN(n5740) );
  NAND2_X1 U7182 ( .A1(n8869), .A2(n8750), .ZN(n8722) );
  NAND2_X1 U7183 ( .A1(n8738), .A2(n8739), .ZN(n8721) );
  NAND2_X1 U7184 ( .A1(n8863), .A2(n8551), .ZN(n5743) );
  NAND2_X1 U7185 ( .A1(n5744), .A2(n5743), .ZN(n8726) );
  INV_X1 U7186 ( .A(n8722), .ZN(n5603) );
  NOR2_X1 U7187 ( .A1(n8726), .A2(n5603), .ZN(n5604) );
  NAND2_X1 U7188 ( .A1(n8721), .A2(n5604), .ZN(n8723) );
  XNOR2_X1 U7189 ( .A(n8859), .B(n8694), .ZN(n8707) );
  NAND2_X1 U7190 ( .A1(n8853), .A2(n8671), .ZN(n5752) );
  NAND2_X1 U7191 ( .A1(n5751), .A2(n5752), .ZN(n8554) );
  INV_X1 U7192 ( .A(n8668), .ZN(n5605) );
  XNOR2_X1 U7193 ( .A(n8848), .B(n8695), .ZN(n8555) );
  INV_X1 U7194 ( .A(n8695), .ZN(n8658) );
  NAND2_X1 U7195 ( .A1(n8848), .A2(n8658), .ZN(n5655) );
  NAND2_X1 U7196 ( .A1(n8842), .A2(n8672), .ZN(n5757) );
  NAND2_X1 U7197 ( .A1(n8661), .A2(n5756), .ZN(n8639) );
  NAND2_X1 U7198 ( .A1(n8838), .A2(n8659), .ZN(n5654) );
  NAND2_X1 U7199 ( .A1(n5760), .A2(n5654), .ZN(n8640) );
  INV_X1 U7200 ( .A(n8640), .ZN(n5819) );
  NAND2_X1 U7201 ( .A1(n8834), .A2(n8563), .ZN(n5769) );
  INV_X1 U7202 ( .A(n8610), .ZN(n5770) );
  OR2_X1 U7203 ( .A1(n8828), .A2(n8588), .ZN(n5768) );
  NAND2_X1 U7204 ( .A1(n8822), .A2(n8579), .ZN(n5765) );
  NAND2_X1 U7205 ( .A1(n5773), .A2(n5765), .ZN(n8593) );
  INV_X1 U7206 ( .A(n8593), .ZN(n5606) );
  NAND2_X1 U7207 ( .A1(n8585), .A2(n5606), .ZN(n8590) );
  NAND2_X1 U7208 ( .A1(n8590), .A2(n5773), .ZN(n8576) );
  INV_X1 U7209 ( .A(SI_28_), .ZN(n5609) );
  NAND2_X1 U7210 ( .A1(n5610), .A2(n5609), .ZN(n5611) );
  INV_X1 U7211 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7907) );
  INV_X1 U7212 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9525) );
  MUX2_X1 U7213 ( .A(n7907), .B(n9525), .S(n6581), .Z(n5618) );
  XNOR2_X1 U7214 ( .A(n5618), .B(SI_29_), .ZN(n5613) );
  NAND2_X1 U7215 ( .A1(n7947), .A2(n5489), .ZN(n5615) );
  OR2_X1 U7216 ( .A1(n5097), .A2(n7907), .ZN(n5614) );
  NAND2_X1 U7217 ( .A1(n8576), .A2(n5778), .ZN(n5616) );
  INV_X1 U7218 ( .A(SI_29_), .ZN(n5617) );
  AND2_X1 U7219 ( .A1(n5618), .A2(n5617), .ZN(n5621) );
  INV_X1 U7220 ( .A(n5618), .ZN(n5619) );
  NAND2_X1 U7221 ( .A1(n5619), .A2(SI_29_), .ZN(n5620) );
  NAND2_X1 U7222 ( .A1(n8244), .A2(n5489), .ZN(n5624) );
  INV_X1 U7223 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8260) );
  OR2_X1 U7224 ( .A1(n4285), .A2(n8260), .ZN(n5623) );
  NAND2_X1 U7225 ( .A1(n4284), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7226 ( .A1(n5628), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7227 ( .A1(n5629), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5625) );
  AND3_X1 U7228 ( .A1(n5627), .A2(n5626), .A3(n5625), .ZN(n8577) );
  NOR2_X1 U7229 ( .A1(n8811), .A2(n8577), .ZN(n5789) );
  NAND2_X1 U7230 ( .A1(n4283), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7231 ( .A1(n5628), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7232 ( .A1(n5629), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5630) );
  NAND3_X1 U7233 ( .A1(n5632), .A2(n5631), .A3(n5630), .ZN(n6744) );
  INV_X1 U7234 ( .A(n8811), .ZN(n5633) );
  INV_X1 U7235 ( .A(n5635), .ZN(n5636) );
  NAND2_X1 U7236 ( .A1(n5636), .A2(SI_30_), .ZN(n5640) );
  NAND2_X1 U7237 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  NAND2_X1 U7238 ( .A1(n5640), .A2(n5639), .ZN(n5643) );
  XNOR2_X1 U7239 ( .A(n5641), .B(SI_31_), .ZN(n5642) );
  INV_X1 U7240 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5644) );
  NOR2_X1 U7241 ( .A1(n4285), .A2(n5644), .ZN(n5645) );
  INV_X1 U7242 ( .A(n8810), .ZN(n5646) );
  INV_X1 U7243 ( .A(n6744), .ZN(n8536) );
  NAND2_X1 U7244 ( .A1(n8811), .A2(n8577), .ZN(n5782) );
  NOR2_X1 U7245 ( .A1(n8810), .A2(n6744), .ZN(n5791) );
  NAND2_X1 U7246 ( .A1(n5648), .A2(n4739), .ZN(n5649) );
  XNOR2_X1 U7247 ( .A(n5649), .B(n7139), .ZN(n5651) );
  OR2_X1 U7248 ( .A1(n7362), .A2(n5562), .ZN(n7016) );
  NAND2_X1 U7249 ( .A1(n5662), .A2(n9823), .ZN(n5652) );
  NAND2_X1 U7250 ( .A1(n4271), .A2(n5654), .ZN(n5759) );
  INV_X1 U7251 ( .A(n8848), .ZN(n8675) );
  AND2_X1 U7252 ( .A1(n7746), .A2(n5669), .ZN(n5656) );
  NAND2_X1 U7253 ( .A1(n7220), .A2(n5657), .ZN(n5658) );
  NAND2_X1 U7254 ( .A1(n5678), .A2(n7214), .ZN(n5810) );
  AOI21_X1 U7255 ( .B1(n5667), .B2(n5658), .A(n5810), .ZN(n5681) );
  INV_X1 U7256 ( .A(n5659), .ZN(n9872) );
  INV_X1 U7257 ( .A(n9874), .ZN(n9873) );
  NAND2_X1 U7258 ( .A1(n9872), .A2(n9873), .ZN(n7325) );
  INV_X1 U7259 ( .A(n7325), .ZN(n5804) );
  NOR2_X1 U7260 ( .A1(n5804), .A2(n5660), .ZN(n5664) );
  AOI21_X1 U7261 ( .B1(n5662), .B2(n7325), .A(n5661), .ZN(n5663) );
  MUX2_X1 U7262 ( .A(n5664), .B(n5663), .S(n4270), .Z(n5676) );
  OAI211_X1 U7263 ( .C1(n5676), .C2(n5665), .A(n4270), .B(n5673), .ZN(n5666)
         );
  NAND3_X1 U7264 ( .A1(n5666), .A2(n5808), .A3(n5667), .ZN(n5672) );
  NAND2_X1 U7265 ( .A1(n7746), .A2(n5683), .ZN(n5809) );
  OAI21_X1 U7266 ( .B1(n5670), .B2(n5809), .A(n4270), .ZN(n5671) );
  NAND2_X1 U7267 ( .A1(n5672), .A2(n5671), .ZN(n5679) );
  NAND2_X1 U7268 ( .A1(n5673), .A2(n5802), .ZN(n5675) );
  OAI211_X1 U7269 ( .C1(n5676), .C2(n5675), .A(n5790), .B(n5674), .ZN(n5677)
         );
  NAND3_X1 U7270 ( .A1(n5679), .A2(n5678), .A3(n5677), .ZN(n5680) );
  OAI21_X1 U7271 ( .B1(n5681), .B2(n4270), .A(n5680), .ZN(n5682) );
  OAI211_X1 U7272 ( .C1(n5683), .C2(n4270), .A(n5682), .B(n7290), .ZN(n5687)
         );
  MUX2_X1 U7273 ( .A(n5685), .B(n5684), .S(n4270), .Z(n5686) );
  NAND3_X1 U7274 ( .A1(n5687), .A2(n9796), .A3(n5686), .ZN(n5691) );
  MUX2_X1 U7275 ( .A(n5689), .B(n5688), .S(n4270), .Z(n5690) );
  NAND3_X1 U7276 ( .A1(n5691), .A2(n5692), .A3(n5690), .ZN(n5704) );
  NAND2_X1 U7277 ( .A1(n5696), .A2(n5692), .ZN(n5695) );
  INV_X1 U7278 ( .A(n5698), .ZN(n5694) );
  INV_X1 U7279 ( .A(n5697), .ZN(n5693) );
  AOI211_X1 U7280 ( .C1(n4270), .C2(n5695), .A(n5694), .B(n5693), .ZN(n5703)
         );
  NAND2_X1 U7281 ( .A1(n5801), .A2(n5696), .ZN(n5701) );
  INV_X1 U7282 ( .A(n5696), .ZN(n5699) );
  OAI211_X1 U7283 ( .C1(n5699), .C2(n5698), .A(n7765), .B(n5697), .ZN(n5700)
         );
  MUX2_X1 U7284 ( .A(n5701), .B(n5700), .S(n4270), .Z(n5702) );
  AOI21_X1 U7285 ( .B1(n5704), .B2(n5703), .A(n5702), .ZN(n5708) );
  INV_X1 U7286 ( .A(n5705), .ZN(n5706) );
  OAI21_X1 U7287 ( .B1(n5708), .B2(n5706), .A(n5799), .ZN(n5710) );
  NAND2_X1 U7288 ( .A1(n5799), .A2(n5801), .ZN(n5707) );
  OAI21_X1 U7289 ( .B1(n5708), .B2(n5707), .A(n5800), .ZN(n5709) );
  MUX2_X1 U7290 ( .A(n5710), .B(n5709), .S(n4270), .Z(n5716) );
  INV_X1 U7291 ( .A(n5711), .ZN(n5714) );
  INV_X1 U7292 ( .A(n5712), .ZN(n5713) );
  MUX2_X1 U7293 ( .A(n5714), .B(n5713), .S(n4270), .Z(n5715) );
  AOI211_X1 U7294 ( .C1(n5716), .C2(n7829), .A(n9578), .B(n5715), .ZN(n5720)
         );
  NOR2_X1 U7295 ( .A1(n9576), .A2(n4270), .ZN(n5718) );
  INV_X1 U7296 ( .A(n9576), .ZN(n9586) );
  NOR2_X1 U7297 ( .A1(n9586), .A2(n5790), .ZN(n5717) );
  MUX2_X1 U7298 ( .A(n5718), .B(n5717), .S(n8479), .Z(n5719) );
  NOR3_X1 U7299 ( .A1(n5720), .A2(n5719), .A3(n8797), .ZN(n5728) );
  NAND2_X1 U7300 ( .A1(n5725), .A2(n5724), .ZN(n8776) );
  INV_X1 U7301 ( .A(n8776), .ZN(n8784) );
  MUX2_X1 U7302 ( .A(n5722), .B(n5721), .S(n4270), .Z(n5723) );
  NAND2_X1 U7303 ( .A1(n8784), .A2(n5723), .ZN(n5727) );
  MUX2_X1 U7304 ( .A(n5725), .B(n5724), .S(n4270), .Z(n5726) );
  OAI211_X1 U7305 ( .C1(n5728), .C2(n5727), .A(n8760), .B(n5726), .ZN(n5734)
         );
  INV_X1 U7306 ( .A(n5729), .ZN(n5730) );
  NOR2_X1 U7307 ( .A1(n5798), .A2(n5730), .ZN(n5731) );
  MUX2_X1 U7308 ( .A(n5732), .B(n5731), .S(n4270), .Z(n5733) );
  NAND3_X1 U7309 ( .A1(n5734), .A2(n5796), .A3(n5733), .ZN(n5742) );
  INV_X1 U7310 ( .A(n5798), .ZN(n5735) );
  NAND3_X1 U7311 ( .A1(n5742), .A2(n5740), .A3(n5735), .ZN(n5737) );
  INV_X1 U7312 ( .A(n5744), .ZN(n5736) );
  AOI21_X1 U7313 ( .B1(n5737), .B2(n8722), .A(n5736), .ZN(n5739) );
  NAND2_X1 U7314 ( .A1(n4305), .A2(n5743), .ZN(n5738) );
  NAND2_X1 U7315 ( .A1(n8706), .A2(n8694), .ZN(n5745) );
  OAI211_X1 U7316 ( .C1(n5739), .C2(n5738), .A(n5745), .B(n5751), .ZN(n5750)
         );
  INV_X1 U7317 ( .A(n5740), .ZN(n5741) );
  AOI21_X1 U7318 ( .B1(n5742), .B2(n5796), .A(n5741), .ZN(n5747) );
  NAND2_X1 U7319 ( .A1(n5743), .A2(n8722), .ZN(n5746) );
  OAI211_X1 U7320 ( .C1(n5747), .C2(n5746), .A(n5745), .B(n5744), .ZN(n5748)
         );
  NAND3_X1 U7321 ( .A1(n5748), .A2(n5752), .A3(n4305), .ZN(n5749) );
  MUX2_X1 U7322 ( .A(n5750), .B(n5749), .S(n4270), .Z(n5754) );
  MUX2_X1 U7323 ( .A(n5752), .B(n5751), .S(n4270), .Z(n5753) );
  MUX2_X1 U7324 ( .A(n5757), .B(n5756), .S(n4270), .Z(n5758) );
  NOR2_X1 U7325 ( .A1(n8834), .A2(n8563), .ZN(n5763) );
  INV_X1 U7326 ( .A(n5760), .ZN(n5761) );
  NOR2_X1 U7327 ( .A1(n5763), .A2(n5761), .ZN(n5762) );
  OAI22_X2 U7328 ( .A1(n5764), .A2(n5763), .B1(n5762), .B2(n4270), .ZN(n5771)
         );
  INV_X1 U7329 ( .A(n8588), .ZN(n8474) );
  OAI21_X1 U7330 ( .B1(n8609), .B2(n8474), .A(n5765), .ZN(n5766) );
  AOI21_X1 U7331 ( .B1(n5771), .B2(n5770), .A(n5766), .ZN(n5767) );
  MUX2_X1 U7332 ( .A(n5768), .B(n5767), .S(n4270), .Z(n5774) );
  NAND3_X1 U7333 ( .A1(n5771), .A2(n5770), .A3(n5769), .ZN(n5772) );
  INV_X1 U7334 ( .A(n8579), .ZN(n8473) );
  INV_X1 U7335 ( .A(n5776), .ZN(n5785) );
  INV_X1 U7336 ( .A(n5778), .ZN(n5777) );
  NOR2_X1 U7337 ( .A1(n5777), .A2(n4270), .ZN(n5781) );
  NOR2_X1 U7338 ( .A1(n8575), .A2(n8579), .ZN(n5780) );
  MUX2_X1 U7339 ( .A(n5781), .B(n5780), .S(n8822), .Z(n5784) );
  INV_X1 U7340 ( .A(n5782), .ZN(n5783) );
  AOI211_X1 U7341 ( .C1(n5785), .C2(n5784), .A(n5783), .B(n5789), .ZN(n5787)
         );
  INV_X1 U7342 ( .A(n5823), .ZN(n5786) );
  NOR2_X1 U7343 ( .A1(n5791), .A2(n5789), .ZN(n5824) );
  INV_X1 U7344 ( .A(n5792), .ZN(n5793) );
  NAND2_X1 U7345 ( .A1(n5793), .A2(n4270), .ZN(n5795) );
  INV_X1 U7346 ( .A(n8575), .ZN(n5822) );
  INV_X1 U7347 ( .A(n8707), .ZN(n8701) );
  INV_X1 U7348 ( .A(n5796), .ZN(n5797) );
  NOR2_X1 U7349 ( .A1(n5798), .A2(n5797), .ZN(n8746) );
  NAND2_X1 U7350 ( .A1(n5800), .A2(n5799), .ZN(n7771) );
  NAND2_X1 U7351 ( .A1(n7765), .A2(n5801), .ZN(n7563) );
  INV_X1 U7352 ( .A(n9877), .ZN(n5803) );
  NOR4_X1 U7353 ( .A1(n5804), .A2(n7009), .A3(n5803), .A4(n5562), .ZN(n5807)
         );
  INV_X1 U7354 ( .A(n7291), .ZN(n5806) );
  NAND4_X1 U7355 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n7010), .ZN(n5811)
         );
  INV_X1 U7356 ( .A(n7290), .ZN(n7316) );
  NOR4_X1 U7357 ( .A1(n5811), .A2(n5810), .A3(n5809), .A4(n7316), .ZN(n5813)
         );
  NAND4_X1 U7358 ( .A1(n5813), .A2(n9796), .A3(n7673), .A4(n5812), .ZN(n5814)
         );
  OR4_X1 U7359 ( .A1(n4766), .A2(n7771), .A3(n7563), .A4(n5814), .ZN(n5815) );
  NOR4_X1 U7360 ( .A1(n8776), .A2(n9578), .A3(n8797), .A4(n5815), .ZN(n5816)
         );
  NAND4_X1 U7361 ( .A1(n8739), .A2(n8760), .A3(n8746), .A4(n5816), .ZN(n5817)
         );
  NOR4_X1 U7362 ( .A1(n8554), .A2(n8701), .A3(n8726), .A4(n5817), .ZN(n5818)
         );
  NAND4_X1 U7363 ( .A1(n5819), .A2(n8558), .A3(n5818), .A4(n8555), .ZN(n5820)
         );
  NOR4_X1 U7364 ( .A1(n8593), .A2(n8610), .A3(n5653), .A4(n5820), .ZN(n5821)
         );
  NAND4_X1 U7365 ( .A1(n5824), .A2(n5823), .A3(n5822), .A4(n5821), .ZN(n5825)
         );
  XNOR2_X1 U7366 ( .A(n5825), .B(n9823), .ZN(n5827) );
  AOI22_X1 U7367 ( .A1(n5827), .A2(n7362), .B1(n5826), .B2(n5562), .ZN(n5828)
         );
  OR2_X1 U7368 ( .A1(n5830), .A2(P2_U3152), .ZN(n7594) );
  INV_X1 U7369 ( .A(n7594), .ZN(n5831) );
  NOR4_X1 U7370 ( .A1(n9832), .A2(n8277), .A3(n5832), .A4(n5833), .ZN(n5835)
         );
  OAI21_X1 U7371 ( .B1(n7594), .B2(n5565), .A(P2_B_REG_SCAN_IN), .ZN(n5834) );
  OR2_X1 U7372 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  NOR2_X1 U7373 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5843) );
  NOR2_X1 U7374 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5842) );
  NOR2_X1 U7375 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5841) );
  NOR2_X1 U7376 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5840) );
  NOR2_X1 U7377 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5844) );
  NAND2_X1 U7378 ( .A1(n5884), .A2(n5846), .ZN(n5852) );
  NAND2_X1 U7379 ( .A1(n5848), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5849) );
  MUX2_X1 U7380 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5849), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5850) );
  INV_X1 U7381 ( .A(n5851), .ZN(n5854) );
  INV_X1 U7382 ( .A(n5852), .ZN(n5853) );
  INV_X2 U7383 ( .A(n5859), .ZN(n9620) );
  INV_X2 U7384 ( .A(n6067), .ZN(n6082) );
  NAND2_X1 U7385 ( .A1(n6951), .A2(n6082), .ZN(n5871) );
  OR2_X1 U7386 ( .A1(n6225), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U7387 ( .A1(n5865), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7388 ( .A1(n6244), .A2(n5873), .ZN(n5866) );
  NAND2_X1 U7389 ( .A1(n5866), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5868) );
  INV_X1 U7390 ( .A(n5868), .ZN(n5867) );
  NAND2_X1 U7391 ( .A1(n5867), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7392 ( .A1(n5868), .A2(n6642), .ZN(n6267) );
  AOI22_X1 U7393 ( .A1(n7939), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6282), .B2(
        n9104), .ZN(n5870) );
  INV_X1 U7394 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5872) );
  NAND4_X1 U7395 ( .A1(n6642), .A2(n6226), .A3(n5873), .A4(n5872), .ZN(n5874)
         );
  AOI21_X1 U7396 ( .B1(n5916), .B2(n5875), .A(n9517), .ZN(n5876) );
  NAND2_X1 U7397 ( .A1(n5881), .A2(n5882), .ZN(n5877) );
  NAND2_X1 U7398 ( .A1(n5851), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5885) );
  OR2_X1 U7399 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  INV_X1 U7400 ( .A(n5888), .ZN(n5889) );
  NAND2_X1 U7401 ( .A1(n5889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5891) );
  INV_X1 U7402 ( .A(n5895), .ZN(n9518) );
  NAND2_X1 U7403 ( .A1(n5893), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7404 ( .A1(n9518), .A2(n5897), .ZN(n5899) );
  NAND2_X1 U7405 ( .A1(n7942), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5913) );
  INV_X4 U7406 ( .A(n5989), .ZN(n6798) );
  NAND2_X1 U7407 ( .A1(n6798), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5912) );
  AND2_X2 U7408 ( .A1(n5898), .A2(n5900), .ZN(n6172) );
  NAND3_X1 U7409 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6023) );
  INV_X1 U7410 ( .A(n6023), .ZN(n5901) );
  NAND2_X1 U7411 ( .A1(n5901), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6058) );
  INV_X1 U7412 ( .A(n6058), .ZN(n5902) );
  NAND2_X1 U7413 ( .A1(n5902), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6075) );
  INV_X1 U7414 ( .A(n6075), .ZN(n5903) );
  NAND2_X1 U7415 ( .A1(n5903), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6094) );
  INV_X1 U7416 ( .A(n6189), .ZN(n5905) );
  NAND2_X1 U7417 ( .A1(n5905), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6191) );
  INV_X1 U7418 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6169) );
  INV_X1 U7419 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6231) );
  INV_X1 U7420 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7421 ( .A1(n6250), .A2(n5908), .ZN(n5909) );
  AND2_X1 U7422 ( .A1(n6273), .A2(n5909), .ZN(n9303) );
  NAND2_X1 U7423 ( .A1(n6172), .A2(n9303), .ZN(n5911) );
  NAND2_X2 U7424 ( .A1(n8245), .A2(n5899), .ZN(n6026) );
  NAND2_X1 U7425 ( .A1(n5941), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5910) );
  NAND4_X1 U7426 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(n9294)
         );
  XNOR2_X2 U7427 ( .A(n5915), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6478) );
  INV_X1 U7428 ( .A(n5916), .ZN(n5917) );
  NAND2_X1 U7429 ( .A1(n5917), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7430 ( .A1(n6455), .A2(n6483), .ZN(n6570) );
  AND2_X4 U7431 ( .A1(n5919), .A2(n6570), .ZN(n6452) );
  OAI22_X1 U7432 ( .A1(n9305), .A2(n6408), .B1(n9320), .B2(n6387), .ZN(n6263)
         );
  INV_X1 U7433 ( .A(n6263), .ZN(n6266) );
  INV_X2 U7434 ( .A(n6406), .ZN(n6388) );
  NAND2_X1 U7435 ( .A1(n9455), .A2(n6388), .ZN(n5921) );
  INV_X2 U7436 ( .A(n6012), .ZN(n6448) );
  NAND2_X1 U7437 ( .A1(n9294), .A2(n6448), .ZN(n5920) );
  NAND2_X1 U7438 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  NAND2_X4 U7439 ( .A1(n6557), .A2(n6499), .ZN(n7142) );
  XNOR2_X1 U7440 ( .A(n5922), .B(n7142), .ZN(n6264) );
  INV_X1 U7441 ( .A(n6264), .ZN(n6265) );
  INV_X2 U7442 ( .A(n6012), .ZN(n6343) );
  INV_X1 U7443 ( .A(SI_0_), .ZN(n5924) );
  INV_X1 U7444 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5923) );
  AND2_X1 U7445 ( .A1(n5926), .A2(n5925), .ZN(n9528) );
  MUX2_X1 U7446 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9528), .S(n6511), .Z(n9731) );
  INV_X1 U7447 ( .A(n6513), .ZN(n5936) );
  AOI22_X1 U7448 ( .A1(n6343), .A2(n9731), .B1(n5936), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5927) );
  INV_X1 U7449 ( .A(n5927), .ZN(n5934) );
  NAND2_X1 U7450 ( .A1(n6172), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5932) );
  INV_X1 U7451 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7452 ( .A1(n6798), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7453 ( .A1(n5941), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7454 ( .A1(n9719), .A2(n6343), .ZN(n5938) );
  AOI22_X1 U7455 ( .A1(n5919), .A2(n9731), .B1(n5936), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7456 ( .A1(n5938), .A2(n5937), .ZN(n6805) );
  INV_X1 U7457 ( .A(n6805), .ZN(n5939) );
  NAND2_X1 U7458 ( .A1(n5939), .A2(n7142), .ZN(n5940) );
  NAND2_X1 U7459 ( .A1(n6172), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5944) );
  INV_X1 U7460 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U7461 ( .A1(n6544), .A2(n6343), .ZN(n5951) );
  NAND2_X1 U7462 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5946) );
  MUX2_X1 U7463 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5946), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5949) );
  INV_X1 U7464 ( .A(n5947), .ZN(n5948) );
  NAND2_X1 U7465 ( .A1(n5949), .A2(n5948), .ZN(n6582) );
  INV_X1 U7466 ( .A(n6582), .ZN(n9608) );
  NAND2_X1 U7467 ( .A1(n6388), .A2(n9730), .ZN(n5950) );
  NAND2_X1 U7468 ( .A1(n5951), .A2(n5950), .ZN(n5952) );
  INV_X2 U7469 ( .A(n7142), .ZN(n6368) );
  XNOR2_X1 U7470 ( .A(n5952), .B(n6368), .ZN(n5956) );
  NAND2_X1 U7471 ( .A1(n6815), .A2(n5956), .ZN(n5955) );
  NAND2_X1 U7472 ( .A1(n6452), .A2(n6544), .ZN(n5954) );
  NAND2_X1 U7473 ( .A1(n9730), .A2(n6448), .ZN(n5953) );
  NAND2_X1 U7474 ( .A1(n5954), .A2(n5953), .ZN(n6814) );
  NAND2_X1 U7475 ( .A1(n5955), .A2(n6814), .ZN(n5959) );
  INV_X1 U7476 ( .A(n6815), .ZN(n5957) );
  INV_X1 U7477 ( .A(n5956), .ZN(n6816) );
  NAND2_X1 U7478 ( .A1(n5957), .A2(n6816), .ZN(n5958) );
  NAND2_X1 U7479 ( .A1(n5959), .A2(n5958), .ZN(n6996) );
  INV_X1 U7480 ( .A(n6996), .ZN(n5977) );
  NAND2_X1 U7481 ( .A1(n6172), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7482 ( .A1(n6798), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5964) );
  INV_X1 U7483 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5960) );
  OR2_X1 U7484 ( .A1(n6025), .A2(n5960), .ZN(n5963) );
  INV_X1 U7485 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5961) );
  OR2_X1 U7486 ( .A1(n6026), .A2(n5961), .ZN(n5962) );
  NAND2_X1 U7487 ( .A1(n6033), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5969) );
  NOR2_X1 U7488 ( .A1(n5947), .A2(n9517), .ZN(n5966) );
  NAND2_X1 U7489 ( .A1(n6282), .A2(n6527), .ZN(n5968) );
  OAI211_X1 U7490 ( .C1(n6067), .C2(n6588), .A(n5969), .B(n5968), .ZN(n6543)
         );
  OAI22_X1 U7491 ( .A1(n7101), .A2(n6408), .B1(n9755), .B2(n6406), .ZN(n5970)
         );
  XNOR2_X1 U7492 ( .A(n5970), .B(n6368), .ZN(n5972) );
  OAI22_X1 U7493 ( .A1(n7101), .A2(n6387), .B1(n9755), .B2(n6408), .ZN(n5973)
         );
  INV_X1 U7494 ( .A(n5973), .ZN(n5971) );
  NAND2_X1 U7495 ( .A1(n5972), .A2(n5971), .ZN(n5978) );
  INV_X1 U7496 ( .A(n5972), .ZN(n5974) );
  NAND2_X1 U7497 ( .A1(n5974), .A2(n5973), .ZN(n5975) );
  NAND2_X1 U7498 ( .A1(n5978), .A2(n5975), .ZN(n6997) );
  NAND2_X1 U7499 ( .A1(n5977), .A2(n5976), .ZN(n6994) );
  INV_X1 U7500 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7206) );
  NAND2_X1 U7501 ( .A1(n6172), .A2(n7206), .ZN(n5984) );
  NAND2_X1 U7502 ( .A1(n6798), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5983) );
  INV_X1 U7503 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5979) );
  OR2_X1 U7504 ( .A1(n6025), .A2(n5979), .ZN(n5982) );
  INV_X1 U7505 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5980) );
  OR2_X1 U7506 ( .A1(n6026), .A2(n5980), .ZN(n5981) );
  NAND2_X1 U7507 ( .A1(n6033), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7508 ( .A1(n5967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7509 ( .A(n5985), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U7510 ( .A1(n6282), .A2(n9529), .ZN(n5986) );
  INV_X1 U7511 ( .A(n7107), .ZN(n7209) );
  OAI22_X1 U7512 ( .A1(n7192), .A2(n6408), .B1(n7209), .B2(n6406), .ZN(n5988)
         );
  XNOR2_X1 U7513 ( .A(n5988), .B(n6368), .ZN(n6004) );
  OAI22_X1 U7514 ( .A1(n7192), .A2(n6387), .B1(n7209), .B2(n6408), .ZN(n6002)
         );
  XNOR2_X1 U7515 ( .A(n6004), .B(n6002), .ZN(n7085) );
  XNOR2_X1 U7516 ( .A(n7206), .B(P1_REG3_REG_4__SCAN_IN), .ZN(n7198) );
  NAND2_X1 U7517 ( .A1(n6172), .A2(n7198), .ZN(n5996) );
  INV_X1 U7518 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5990) );
  INV_X1 U7519 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5991) );
  OR2_X1 U7520 ( .A1(n6025), .A2(n5991), .ZN(n5994) );
  INV_X1 U7521 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5992) );
  OR2_X1 U7522 ( .A1(n6026), .A2(n5992), .ZN(n5993) );
  NAND2_X1 U7523 ( .A1(n6033), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7524 ( .A1(n5997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5998) );
  XNOR2_X1 U7525 ( .A(n5998), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U7526 ( .A1(n6282), .A2(n6526), .ZN(n5999) );
  OAI211_X1 U7527 ( .C1(n6067), .C2(n6586), .A(n6000), .B(n5999), .ZN(n7199)
         );
  INV_X1 U7528 ( .A(n7199), .ZN(n9760) );
  OAI22_X1 U7529 ( .A1(n7145), .A2(n6408), .B1(n9760), .B2(n6406), .ZN(n6001)
         );
  XNOR2_X1 U7530 ( .A(n6001), .B(n6368), .ZN(n6044) );
  OAI22_X1 U7531 ( .A1(n7145), .A2(n6387), .B1(n9760), .B2(n6408), .ZN(n6045)
         );
  XNOR2_X1 U7532 ( .A(n6044), .B(n6045), .ZN(n7182) );
  INV_X1 U7533 ( .A(n6002), .ZN(n6003) );
  NAND2_X1 U7534 ( .A1(n6004), .A2(n6003), .ZN(n7183) );
  AND2_X1 U7535 ( .A1(n7182), .A2(n7183), .ZN(n7181) );
  NAND2_X1 U7536 ( .A1(n7942), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7537 ( .A1(n6798), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6010) );
  INV_X1 U7538 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7539 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6005) );
  NAND2_X1 U7540 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  AND2_X1 U7541 ( .A1(n6023), .A2(n6007), .ZN(n7547) );
  NAND2_X1 U7542 ( .A1(n6172), .A2(n7547), .ZN(n6009) );
  NAND2_X1 U7543 ( .A1(n5941), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7544 ( .A1(n9048), .A2(n6448), .ZN(n6018) );
  NAND2_X1 U7545 ( .A1(n6033), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7546 ( .A1(n6013), .A2(n9517), .ZN(n6014) );
  XNOR2_X1 U7547 ( .A(n6014), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U7548 ( .A1(n6282), .A2(n9653), .ZN(n6015) );
  OAI211_X1 U7549 ( .C1(n6067), .C2(n6585), .A(n6016), .B(n6015), .ZN(n7376)
         );
  NAND2_X1 U7550 ( .A1(n5919), .A2(n7376), .ZN(n6017) );
  NAND2_X1 U7551 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  XNOR2_X1 U7552 ( .A(n6019), .B(n6368), .ZN(n7423) );
  INV_X1 U7553 ( .A(n7423), .ZN(n6022) );
  NAND2_X1 U7554 ( .A1(n6452), .A2(n9048), .ZN(n6021) );
  NAND2_X1 U7555 ( .A1(n7376), .A2(n6448), .ZN(n6020) );
  AND2_X1 U7556 ( .A1(n6021), .A2(n6020), .ZN(n6042) );
  INV_X1 U7557 ( .A(n6042), .ZN(n7543) );
  NAND2_X1 U7558 ( .A1(n6022), .A2(n7543), .ZN(n6041) );
  INV_X1 U7559 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U7560 ( .A1(n6023), .A2(n6765), .ZN(n6024) );
  AND2_X1 U7561 ( .A1(n6058), .A2(n6024), .ZN(n7443) );
  NAND2_X1 U7562 ( .A1(n6172), .A2(n7443), .ZN(n6031) );
  NAND2_X1 U7563 ( .A1(n6798), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6030) );
  INV_X1 U7564 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6520) );
  OR2_X1 U7565 ( .A1(n6025), .A2(n6520), .ZN(n6029) );
  INV_X1 U7566 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7567 ( .A1(n6033), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6040) );
  NOR2_X1 U7568 ( .A1(n6034), .A2(n9517), .ZN(n6035) );
  MUX2_X1 U7569 ( .A(n9517), .B(n6035), .S(P1_IR_REG_6__SCAN_IN), .Z(n6038) );
  INV_X1 U7570 ( .A(n6036), .ZN(n6037) );
  OR2_X1 U7571 ( .A1(n6038), .A2(n6037), .ZN(n6597) );
  INV_X1 U7572 ( .A(n6597), .ZN(n6771) );
  NAND2_X1 U7573 ( .A1(n6282), .A2(n6771), .ZN(n6039) );
  OAI22_X1 U7574 ( .A1(n7537), .A2(n6387), .B1(n9766), .B2(n6408), .ZN(n6054)
         );
  XNOR2_X1 U7575 ( .A(n6053), .B(n6054), .ZN(n7427) );
  AND2_X1 U7576 ( .A1(n6041), .A2(n7427), .ZN(n6047) );
  NAND2_X1 U7577 ( .A1(n7083), .A2(n6043), .ZN(n6052) );
  INV_X1 U7578 ( .A(n6044), .ZN(n6046) );
  NAND2_X1 U7579 ( .A1(n6046), .A2(n6045), .ZN(n7421) );
  AND2_X1 U7580 ( .A1(n7421), .A2(n6047), .ZN(n6050) );
  INV_X1 U7581 ( .A(n6048), .ZN(n6049) );
  INV_X1 U7582 ( .A(n6053), .ZN(n6055) );
  OR2_X1 U7583 ( .A1(n6055), .A2(n6054), .ZN(n6056) );
  INV_X1 U7584 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7585 ( .A1(n6058), .A2(n6057), .ZN(n6059) );
  AND2_X1 U7586 ( .A1(n6075), .A2(n6059), .ZN(n7403) );
  NAND2_X1 U7587 ( .A1(n6172), .A2(n7403), .ZN(n6064) );
  NAND2_X1 U7588 ( .A1(n6798), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6063) );
  INV_X1 U7589 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6060) );
  OR2_X1 U7590 ( .A1(n6026), .A2(n6060), .ZN(n6062) );
  INV_X1 U7591 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7400) );
  OR2_X1 U7592 ( .A1(n6025), .A2(n7400), .ZN(n6061) );
  NAND2_X1 U7593 ( .A1(n6036), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6066) );
  XNOR2_X1 U7594 ( .A(n6066), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6786) );
  OAI22_X1 U7595 ( .A1(n7380), .A2(n6408), .B1(n7405), .B2(n6406), .ZN(n6068)
         );
  XNOR2_X1 U7596 ( .A(n6068), .B(n6368), .ZN(n6071) );
  OAI22_X1 U7597 ( .A1(n7380), .A2(n6387), .B1(n7405), .B2(n6408), .ZN(n6072)
         );
  INV_X1 U7598 ( .A(n6072), .ZN(n6069) );
  AND2_X1 U7599 ( .A1(n6071), .A2(n6069), .ZN(n7352) );
  INV_X1 U7600 ( .A(n7352), .ZN(n6070) );
  INV_X1 U7601 ( .A(n6071), .ZN(n6073) );
  NAND2_X1 U7602 ( .A1(n6073), .A2(n6072), .ZN(n7353) );
  NAND2_X1 U7603 ( .A1(n6074), .A2(n7353), .ZN(n6088) );
  INV_X1 U7604 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7414) );
  NAND2_X1 U7605 ( .A1(n6075), .A2(n7414), .ZN(n6076) );
  AND2_X1 U7606 ( .A1(n6094), .A2(n6076), .ZN(n7413) );
  NAND2_X1 U7607 ( .A1(n6172), .A2(n7413), .ZN(n6081) );
  NAND2_X1 U7608 ( .A1(n6798), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6080) );
  INV_X1 U7609 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6077) );
  OR2_X1 U7610 ( .A1(n6026), .A2(n6077), .ZN(n6079) );
  INV_X1 U7611 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7384) );
  OR2_X1 U7612 ( .A1(n6025), .A2(n7384), .ZN(n6078) );
  NAND2_X1 U7613 ( .A1(n6082), .A2(n6602), .ZN(n6085) );
  NAND2_X1 U7614 ( .A1(n4350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6083) );
  XNOR2_X1 U7615 ( .A(n6083), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9665) );
  NAND2_X1 U7616 ( .A1(n6282), .A2(n9665), .ZN(n6084) );
  OAI211_X1 U7617 ( .C1(n4446), .C2(n6086), .A(n6085), .B(n6084), .ZN(n7598)
         );
  INV_X1 U7618 ( .A(n7598), .ZN(n7374) );
  OAI22_X1 U7619 ( .A1(n7373), .A2(n6387), .B1(n7374), .B2(n6408), .ZN(n6089)
         );
  NAND2_X1 U7620 ( .A1(n6088), .A2(n6089), .ZN(n7409) );
  OAI22_X1 U7621 ( .A1(n7373), .A2(n6408), .B1(n7374), .B2(n6406), .ZN(n6087)
         );
  XNOR2_X1 U7622 ( .A(n6087), .B(n6368), .ZN(n7411) );
  NAND2_X1 U7623 ( .A1(n7409), .A2(n7411), .ZN(n6092) );
  NAND2_X1 U7624 ( .A1(n6094), .A2(n6093), .ZN(n6095) );
  AND2_X1 U7625 ( .A1(n6112), .A2(n6095), .ZN(n7511) );
  NAND2_X1 U7626 ( .A1(n6172), .A2(n7511), .ZN(n6099) );
  NAND2_X1 U7627 ( .A1(n7942), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7628 ( .A1(n6798), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7629 ( .A1(n5941), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6096) );
  NAND4_X1 U7630 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n6096), .ZN(n9546)
         );
  NAND2_X1 U7631 ( .A1(n9546), .A2(n6448), .ZN(n6104) );
  NAND2_X1 U7632 ( .A1(n5860), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6100) );
  XNOR2_X1 U7633 ( .A(n6100), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6858) );
  INV_X1 U7634 ( .A(n6858), .ZN(n6729) );
  NAND2_X1 U7635 ( .A1(n6727), .A2(n6082), .ZN(n6102) );
  NAND2_X1 U7636 ( .A1(n7939), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n6101) );
  OAI211_X1 U7637 ( .C1(n6511), .C2(n6729), .A(n6102), .B(n6101), .ZN(n9486)
         );
  NAND2_X1 U7638 ( .A1(n6388), .A2(n9486), .ZN(n6103) );
  NAND2_X1 U7639 ( .A1(n6104), .A2(n6103), .ZN(n6105) );
  XNOR2_X1 U7640 ( .A(n6105), .B(n6368), .ZN(n6110) );
  NAND2_X1 U7641 ( .A1(n6452), .A2(n9546), .ZN(n6107) );
  NAND2_X1 U7642 ( .A1(n9486), .A2(n6448), .ZN(n6106) );
  NAND2_X1 U7643 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  XNOR2_X1 U7644 ( .A(n6110), .B(n6108), .ZN(n7494) );
  INV_X1 U7645 ( .A(n6108), .ZN(n6109) );
  AND2_X1 U7646 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  NAND2_X1 U7647 ( .A1(n6112), .A2(n7530), .ZN(n6113) );
  AND2_X1 U7648 ( .A1(n6138), .A2(n6113), .ZN(n9550) );
  NAND2_X1 U7649 ( .A1(n6172), .A2(n9550), .ZN(n6119) );
  NAND2_X1 U7650 ( .A1(n6798), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6118) );
  INV_X1 U7651 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6114) );
  OR2_X1 U7652 ( .A1(n6025), .A2(n6114), .ZN(n6117) );
  INV_X1 U7653 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6115) );
  OR2_X1 U7654 ( .A1(n6026), .A2(n6115), .ZN(n6116) );
  NAND2_X1 U7655 ( .A1(n6732), .A2(n6082), .ZN(n6125) );
  OR2_X1 U7656 ( .A1(n6120), .A2(n9517), .ZN(n6163) );
  INV_X1 U7657 ( .A(n6163), .ZN(n6121) );
  NAND2_X1 U7658 ( .A1(n6121), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6123) );
  INV_X1 U7659 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7660 ( .A1(n6163), .A2(n6122), .ZN(n6133) );
  AOI22_X1 U7661 ( .A1(n7939), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6282), .B2(
        n9695), .ZN(n6124) );
  NAND2_X1 U7662 ( .A1(n6125), .A2(n6124), .ZN(n9552) );
  NAND2_X1 U7663 ( .A1(n9552), .A2(n6388), .ZN(n6126) );
  OAI21_X1 U7664 ( .B1(n7734), .B2(n6408), .A(n6126), .ZN(n6127) );
  XNOR2_X1 U7665 ( .A(n6127), .B(n6368), .ZN(n7527) );
  INV_X1 U7666 ( .A(n7734), .ZN(n9045) );
  NAND2_X1 U7667 ( .A1(n9045), .A2(n6452), .ZN(n6129) );
  NAND2_X1 U7668 ( .A1(n9552), .A2(n6448), .ZN(n6128) );
  AND2_X1 U7669 ( .A1(n6129), .A2(n6128), .ZN(n6131) );
  NAND2_X1 U7670 ( .A1(n7527), .A2(n6131), .ZN(n6130) );
  INV_X1 U7671 ( .A(n7527), .ZN(n6132) );
  INV_X1 U7672 ( .A(n6131), .ZN(n7526) );
  NAND2_X1 U7673 ( .A1(n6132), .A2(n7526), .ZN(n6215) );
  NAND2_X1 U7674 ( .A1(n6740), .A2(n6082), .ZN(n6136) );
  NAND2_X1 U7675 ( .A1(n6133), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6134) );
  XNOR2_X1 U7676 ( .A(n6134), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6860) );
  AOI22_X1 U7677 ( .A1(n7939), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6282), .B2(
        n6860), .ZN(n6135) );
  NAND2_X1 U7678 ( .A1(n9479), .A2(n6388), .ZN(n6145) );
  NAND2_X1 U7679 ( .A1(n7942), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7680 ( .A1(n6798), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6142) );
  INV_X1 U7681 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7682 ( .A1(n6138), .A2(n6137), .ZN(n6139) );
  AND2_X1 U7683 ( .A1(n6189), .A2(n6139), .ZN(n7740) );
  NAND2_X1 U7684 ( .A1(n6172), .A2(n7740), .ZN(n6141) );
  NAND2_X1 U7685 ( .A1(n5941), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6140) );
  NAND4_X1 U7686 ( .A1(n6143), .A2(n6142), .A3(n6141), .A4(n6140), .ZN(n9545)
         );
  NAND2_X1 U7687 ( .A1(n9545), .A2(n6448), .ZN(n6144) );
  NAND2_X1 U7688 ( .A1(n6145), .A2(n6144), .ZN(n6146) );
  XNOR2_X1 U7689 ( .A(n6146), .B(n7142), .ZN(n6202) );
  AOI22_X1 U7690 ( .A1(n9479), .A2(n6343), .B1(n6452), .B2(n9545), .ZN(n6203)
         );
  XNOR2_X1 U7691 ( .A(n6202), .B(n6203), .ZN(n7721) );
  NAND2_X1 U7692 ( .A1(n6794), .A2(n6082), .ZN(n6152) );
  NOR2_X1 U7693 ( .A1(n6147), .A2(n9517), .ZN(n6148) );
  MUX2_X1 U7694 ( .A(n9517), .B(n6148), .S(P1_IR_REG_14__SCAN_IN), .Z(n6149)
         );
  INV_X1 U7695 ( .A(n6149), .ZN(n6150) );
  AND2_X1 U7696 ( .A1(n6150), .A2(n6225), .ZN(n7624) );
  AOI22_X1 U7697 ( .A1(n7939), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6282), .B2(
        n7624), .ZN(n6151) );
  NAND2_X1 U7698 ( .A1(n9359), .A2(n6388), .ZN(n6160) );
  NAND2_X1 U7699 ( .A1(n7942), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7700 ( .A1(n5941), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6157) );
  INV_X1 U7701 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7702 ( .A1(n6171), .A2(n6153), .ZN(n6154) );
  AND2_X1 U7703 ( .A1(n6232), .A2(n6154), .ZN(n9358) );
  NAND2_X1 U7704 ( .A1(n6172), .A2(n9358), .ZN(n6156) );
  NAND2_X1 U7705 ( .A1(n6798), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6155) );
  NAND4_X1 U7706 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n9373)
         );
  NAND2_X1 U7707 ( .A1(n9373), .A2(n6448), .ZN(n6159) );
  NAND2_X1 U7708 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  XNOR2_X1 U7709 ( .A(n6161), .B(n7142), .ZN(n6220) );
  NAND2_X1 U7710 ( .A1(n6790), .A2(n6082), .ZN(n6168) );
  OAI21_X1 U7711 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7712 ( .A1(n6163), .A2(n6162), .ZN(n6183) );
  INV_X1 U7713 ( .A(n6183), .ZN(n6165) );
  INV_X1 U7714 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7715 ( .A1(n6165), .A2(n6164), .ZN(n6185) );
  NAND2_X1 U7716 ( .A1(n6185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6166) );
  XNOR2_X1 U7717 ( .A(n6166), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7283) );
  AOI22_X1 U7718 ( .A1(n7939), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6282), .B2(
        n7283), .ZN(n6167) );
  NAND2_X1 U7719 ( .A1(n9470), .A2(n6388), .ZN(n6178) );
  NAND2_X1 U7720 ( .A1(n5941), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7721 ( .A1(n7942), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7722 ( .A1(n6191), .A2(n6169), .ZN(n6170) );
  AND2_X1 U7723 ( .A1(n6171), .A2(n6170), .ZN(n9381) );
  NAND2_X1 U7724 ( .A1(n6172), .A2(n9381), .ZN(n6174) );
  NAND2_X1 U7725 ( .A1(n6798), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6173) );
  NAND4_X1 U7726 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .ZN(n9353)
         );
  NAND2_X1 U7727 ( .A1(n9353), .A2(n6448), .ZN(n6177) );
  NAND2_X1 U7728 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  XNOR2_X1 U7729 ( .A(n6179), .B(n6368), .ZN(n6182) );
  AND2_X1 U7730 ( .A1(n6452), .A2(n9353), .ZN(n6180) );
  AOI21_X1 U7731 ( .B1(n9470), .B2(n6343), .A(n6180), .ZN(n6181) );
  NAND2_X1 U7732 ( .A1(n6746), .A2(n6082), .ZN(n6187) );
  NAND2_X1 U7733 ( .A1(n6183), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6184) );
  AOI22_X1 U7734 ( .A1(n7939), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6282), .B2(
        n7065), .ZN(n6186) );
  NAND2_X1 U7735 ( .A1(n9597), .A2(n6388), .ZN(n6199) );
  INV_X1 U7736 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7737 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  AND2_X1 U7738 ( .A1(n6191), .A2(n6190), .ZN(n7839) );
  NAND2_X1 U7739 ( .A1(n6172), .A2(n7839), .ZN(n6197) );
  NAND2_X1 U7740 ( .A1(n6798), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6196) );
  INV_X1 U7741 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6192) );
  OR2_X1 U7742 ( .A1(n6026), .A2(n6192), .ZN(n6195) );
  INV_X1 U7743 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6193) );
  OR2_X1 U7744 ( .A1(n6025), .A2(n6193), .ZN(n6194) );
  NAND2_X1 U7745 ( .A1(n9374), .A2(n6448), .ZN(n6198) );
  NAND2_X1 U7746 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  NOR2_X1 U7747 ( .A1(n7788), .A2(n6387), .ZN(n6201) );
  AOI21_X1 U7748 ( .B1(n9597), .B2(n6343), .A(n6201), .ZN(n6206) );
  INV_X1 U7749 ( .A(n6240), .ZN(n6212) );
  INV_X1 U7750 ( .A(n6202), .ZN(n6204) );
  OR2_X1 U7751 ( .A1(n6204), .A2(n6203), .ZN(n7835) );
  INV_X1 U7752 ( .A(n6205), .ZN(n6208) );
  INV_X1 U7753 ( .A(n6206), .ZN(n6207) );
  NAND2_X1 U7754 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  NAND2_X1 U7755 ( .A1(n7871), .A2(n6209), .ZN(n7838) );
  OR2_X1 U7756 ( .A1(n7838), .A2(n6210), .ZN(n6213) );
  NOR2_X1 U7757 ( .A1(n6213), .A2(n6220), .ZN(n6211) );
  AND2_X1 U7758 ( .A1(n7835), .A2(n6211), .ZN(n6239) );
  AOI22_X1 U7759 ( .A1(n9359), .A2(n6343), .B1(n6452), .B2(n9373), .ZN(n7856)
         );
  INV_X1 U7760 ( .A(n6213), .ZN(n6214) );
  AND2_X1 U7761 ( .A1(n6214), .A2(n7835), .ZN(n6218) );
  AND2_X1 U7762 ( .A1(n6215), .A2(n6218), .ZN(n6216) );
  NAND2_X1 U7763 ( .A1(n6217), .A2(n6216), .ZN(n6224) );
  INV_X1 U7764 ( .A(n6218), .ZN(n6219) );
  NAND2_X1 U7765 ( .A1(n6221), .A2(n6220), .ZN(n6222) );
  NAND2_X1 U7766 ( .A1(n6827), .A2(n6082), .ZN(n6230) );
  NAND2_X1 U7767 ( .A1(n6225), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6227) );
  XNOR2_X1 U7768 ( .A(n6227), .B(n6226), .ZN(n9071) );
  INV_X1 U7769 ( .A(n9071), .ZN(n6228) );
  AOI22_X1 U7770 ( .A1(n7939), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6282), .B2(
        n6228), .ZN(n6229) );
  NAND2_X1 U7771 ( .A1(n5941), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7772 ( .A1(n7942), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7773 ( .A1(n6232), .A2(n6231), .ZN(n6233) );
  AND2_X1 U7774 ( .A1(n6248), .A2(n6233), .ZN(n9339) );
  NAND2_X1 U7775 ( .A1(n6172), .A2(n9339), .ZN(n6235) );
  NAND2_X1 U7776 ( .A1(n6798), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6234) );
  NAND4_X1 U7777 ( .A1(n6237), .A2(n6236), .A3(n6235), .A4(n6234), .ZN(n9354)
         );
  OAI22_X1 U7778 ( .A1(n9342), .A2(n6406), .B1(n9319), .B2(n6408), .ZN(n6238)
         );
  XNOR2_X1 U7779 ( .A(n6238), .B(n7142), .ZN(n6242) );
  AOI22_X1 U7780 ( .A1(n9465), .A2(n6343), .B1(n6452), .B2(n9354), .ZN(n9029)
         );
  NAND2_X1 U7781 ( .A1(n7722), .A2(n7721), .ZN(n7836) );
  NAND2_X1 U7782 ( .A1(n7836), .A2(n6239), .ZN(n6241) );
  NAND2_X1 U7783 ( .A1(n6241), .A2(n6240), .ZN(n7853) );
  NAND2_X1 U7784 ( .A1(n6243), .A2(n6242), .ZN(n9028) );
  NAND2_X1 U7785 ( .A1(n6823), .A2(n6082), .ZN(n6246) );
  XNOR2_X1 U7786 ( .A(n6244), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9089) );
  AOI22_X1 U7787 ( .A1(n7939), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6282), .B2(
        n9089), .ZN(n6245) );
  NAND2_X1 U7788 ( .A1(n6798), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6256) );
  INV_X1 U7789 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7790 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  AND2_X1 U7791 ( .A1(n6250), .A2(n6249), .ZN(n9322) );
  NAND2_X1 U7792 ( .A1(n6172), .A2(n9322), .ZN(n6255) );
  INV_X1 U7793 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6251) );
  OR2_X1 U7794 ( .A1(n6025), .A2(n6251), .ZN(n6254) );
  INV_X1 U7795 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6252) );
  OR2_X1 U7796 ( .A1(n6026), .A2(n6252), .ZN(n6253) );
  AOI22_X1 U7797 ( .A1(n9462), .A2(n6343), .B1(n6452), .B2(n9308), .ZN(n6261)
         );
  NAND2_X1 U7798 ( .A1(n9462), .A2(n6388), .ZN(n6258) );
  NAND2_X1 U7799 ( .A1(n9308), .A2(n6343), .ZN(n6257) );
  NAND2_X1 U7800 ( .A1(n6258), .A2(n6257), .ZN(n6259) );
  XNOR2_X1 U7801 ( .A(n6259), .B(n7142), .ZN(n6260) );
  XOR2_X1 U7802 ( .A(n6261), .B(n6260), .Z(n8963) );
  INV_X1 U7803 ( .A(n6260), .ZN(n6262) );
  XNOR2_X1 U7804 ( .A(n6264), .B(n6263), .ZN(n8970) );
  NAND2_X1 U7805 ( .A1(n7081), .A2(n6082), .ZN(n6270) );
  NAND2_X1 U7806 ( .A1(n6267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6268) );
  XNOR2_X1 U7807 ( .A(n6268), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9703) );
  AOI22_X1 U7808 ( .A1(n7939), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9703), .B2(
        n6282), .ZN(n6269) );
  INV_X1 U7809 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7810 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  AND2_X1 U7811 ( .A1(n6287), .A2(n6274), .ZN(n9286) );
  NAND2_X1 U7812 ( .A1(n6172), .A2(n9286), .ZN(n6279) );
  NAND2_X1 U7813 ( .A1(n6798), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6278) );
  INV_X1 U7814 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n6275) );
  OR2_X1 U7815 ( .A1(n6025), .A2(n6275), .ZN(n6277) );
  INV_X1 U7816 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n6655) );
  OR2_X1 U7817 ( .A1(n6026), .A2(n6655), .ZN(n6276) );
  OAI22_X1 U7818 ( .A1(n9288), .A2(n6406), .B1(n8941), .B2(n6408), .ZN(n6280)
         );
  XOR2_X1 U7819 ( .A(n7142), .B(n6280), .Z(n9005) );
  INV_X1 U7820 ( .A(n9005), .ZN(n6281) );
  OAI22_X1 U7821 ( .A1(n9288), .A2(n6408), .B1(n8941), .B2(n6387), .ZN(n9004)
         );
  NAND2_X1 U7822 ( .A1(n7137), .A2(n6082), .ZN(n6284) );
  AOI22_X1 U7823 ( .A1(n7939), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9736), .B2(
        n6282), .ZN(n6283) );
  INV_X1 U7824 ( .A(n9446), .ZN(n9272) );
  NAND2_X1 U7825 ( .A1(n5941), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U7826 ( .A1(n7942), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6291) );
  INV_X1 U7827 ( .A(n6287), .ZN(n6285) );
  NAND2_X1 U7828 ( .A1(n6285), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6303) );
  INV_X1 U7829 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U7830 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  AND2_X1 U7831 ( .A1(n6303), .A2(n6288), .ZN(n9270) );
  NAND2_X1 U7832 ( .A1(n6172), .A2(n9270), .ZN(n6290) );
  NAND2_X1 U7833 ( .A1(n6798), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6289) );
  NAND4_X1 U7834 ( .A1(n6292), .A2(n6291), .A3(n6290), .A4(n6289), .ZN(n9295)
         );
  OAI22_X1 U7835 ( .A1(n9272), .A2(n6408), .B1(n9258), .B2(n6387), .ZN(n6297)
         );
  NAND2_X1 U7836 ( .A1(n9446), .A2(n6388), .ZN(n6294) );
  NAND2_X1 U7837 ( .A1(n9295), .A2(n6448), .ZN(n6293) );
  NAND2_X1 U7838 ( .A1(n6294), .A2(n6293), .ZN(n6295) );
  XNOR2_X1 U7839 ( .A(n6295), .B(n7142), .ZN(n6296) );
  XOR2_X1 U7840 ( .A(n6297), .B(n6296), .Z(n8938) );
  INV_X1 U7841 ( .A(n6296), .ZN(n6299) );
  INV_X1 U7842 ( .A(n6297), .ZN(n6298) );
  NAND2_X1 U7843 ( .A1(n7242), .A2(n6082), .ZN(n6301) );
  NAND2_X1 U7844 ( .A1(n7939), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7845 ( .A1(n9442), .A2(n6388), .ZN(n6310) );
  NAND2_X1 U7846 ( .A1(n7942), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U7847 ( .A1(n6798), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6307) );
  INV_X1 U7848 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7849 ( .A1(n6303), .A2(n6302), .ZN(n6304) );
  AND2_X1 U7850 ( .A1(n6318), .A2(n6304), .ZN(n9261) );
  NAND2_X1 U7851 ( .A1(n6172), .A2(n9261), .ZN(n6306) );
  NAND2_X1 U7852 ( .A1(n5941), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6305) );
  NAND4_X1 U7853 ( .A1(n6308), .A2(n6307), .A3(n6306), .A4(n6305), .ZN(n9276)
         );
  NAND2_X1 U7854 ( .A1(n9276), .A2(n6448), .ZN(n6309) );
  NAND2_X1 U7855 ( .A1(n6310), .A2(n6309), .ZN(n6311) );
  XNOR2_X1 U7856 ( .A(n6311), .B(n6368), .ZN(n6314) );
  AND2_X1 U7857 ( .A1(n6452), .A2(n9276), .ZN(n6312) );
  AOI21_X1 U7858 ( .B1(n9442), .B2(n6448), .A(n6312), .ZN(n6313) );
  NOR2_X1 U7859 ( .A1(n6314), .A2(n6313), .ZN(n8986) );
  INV_X1 U7860 ( .A(n8946), .ZN(n6331) );
  NAND2_X1 U7861 ( .A1(n7332), .A2(n6082), .ZN(n6316) );
  NAND2_X1 U7862 ( .A1(n7939), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7863 ( .A1(n9437), .A2(n5919), .ZN(n6327) );
  INV_X1 U7864 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U7865 ( .A1(n6318), .A2(n6317), .ZN(n6319) );
  AND2_X1 U7866 ( .A1(n6336), .A2(n6319), .ZN(n9248) );
  NAND2_X1 U7867 ( .A1(n9248), .A2(n6172), .ZN(n6325) );
  NAND2_X1 U7868 ( .A1(n6798), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6324) );
  INV_X1 U7869 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6320) );
  OR2_X1 U7870 ( .A1(n6025), .A2(n6320), .ZN(n6323) );
  INV_X1 U7871 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n6321) );
  OR2_X1 U7872 ( .A1(n6026), .A2(n6321), .ZN(n6322) );
  NAND2_X1 U7873 ( .A1(n9235), .A2(n6448), .ZN(n6326) );
  NAND2_X1 U7874 ( .A1(n6327), .A2(n6326), .ZN(n6328) );
  XNOR2_X1 U7875 ( .A(n6328), .B(n7142), .ZN(n6330) );
  INV_X1 U7876 ( .A(n9437), .ZN(n9251) );
  OAI22_X1 U7877 ( .A1(n9251), .A2(n6408), .B1(n9259), .B2(n6387), .ZN(n6329)
         );
  XNOR2_X1 U7878 ( .A(n6330), .B(n6329), .ZN(n8945) );
  OAI22_X1 U7879 ( .A1(n6331), .A2(n8945), .B1(n6330), .B2(n6329), .ZN(n6345)
         );
  NAND2_X1 U7880 ( .A1(n7462), .A2(n6082), .ZN(n6333) );
  NAND2_X1 U7881 ( .A1(n7939), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6332) );
  INV_X1 U7882 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6342) );
  INV_X1 U7883 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7884 ( .A1(n6336), .A2(n6335), .ZN(n6337) );
  NAND2_X1 U7885 ( .A1(n6351), .A2(n6337), .ZN(n9227) );
  INV_X1 U7886 ( .A(n6172), .ZN(n6491) );
  OR2_X1 U7887 ( .A1(n9227), .A2(n6491), .ZN(n6341) );
  NAND2_X1 U7888 ( .A1(n7942), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U7889 ( .A1(n6798), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6338) );
  AND2_X1 U7890 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  OAI211_X1 U7891 ( .C1(n6026), .C2(n6342), .A(n6341), .B(n6340), .ZN(n9217)
         );
  AOI22_X1 U7892 ( .A1(n9430), .A2(n6343), .B1(n6452), .B2(n9217), .ZN(n6346)
         );
  INV_X1 U7893 ( .A(n9217), .ZN(n9244) );
  OAI22_X1 U7894 ( .A1(n9230), .A2(n6406), .B1(n9244), .B2(n6408), .ZN(n6344)
         );
  XNOR2_X1 U7895 ( .A(n6344), .B(n7142), .ZN(n8997) );
  NAND2_X1 U7896 ( .A1(n7593), .A2(n6082), .ZN(n6348) );
  NAND2_X1 U7897 ( .A1(n7939), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6347) );
  INV_X1 U7898 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6355) );
  INV_X1 U7899 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7900 ( .A1(n6351), .A2(n6350), .ZN(n6352) );
  NAND2_X1 U7901 ( .A1(n6360), .A2(n6352), .ZN(n9212) );
  OR2_X1 U7902 ( .A1(n9212), .A2(n6491), .ZN(n6354) );
  AOI22_X1 U7903 ( .A1(n6798), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n7942), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n6353) );
  OAI211_X1 U7904 ( .C1(n6026), .C2(n6355), .A(n6354), .B(n6353), .ZN(n9234)
         );
  INV_X1 U7905 ( .A(n9234), .ZN(n8197) );
  OAI22_X1 U7906 ( .A1(n4452), .A2(n6406), .B1(n8197), .B2(n6408), .ZN(n6356)
         );
  XOR2_X1 U7907 ( .A(n7142), .B(n6356), .Z(n6378) );
  NAND2_X1 U7908 ( .A1(n6377), .A2(n6378), .ZN(n8929) );
  OAI22_X1 U7909 ( .A1(n4452), .A2(n6408), .B1(n8197), .B2(n6387), .ZN(n8931)
         );
  NAND2_X1 U7910 ( .A1(n8929), .A2(n8931), .ZN(n8979) );
  NAND2_X1 U7911 ( .A1(n7780), .A2(n6082), .ZN(n6358) );
  NAND2_X1 U7912 ( .A1(n7939), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6357) );
  INV_X1 U7913 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U7914 ( .A1(n6360), .A2(n6359), .ZN(n6361) );
  AND2_X1 U7915 ( .A1(n6398), .A2(n6361), .ZN(n9203) );
  NAND2_X1 U7916 ( .A1(n9203), .A2(n6172), .ZN(n6367) );
  INV_X1 U7917 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U7918 ( .A1(n7942), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U7919 ( .A1(n5941), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6362) );
  OAI211_X1 U7920 ( .C1(n6364), .C2(n5989), .A(n6363), .B(n6362), .ZN(n6365)
         );
  INV_X1 U7921 ( .A(n6365), .ZN(n6366) );
  OAI22_X1 U7922 ( .A1(n9192), .A2(n6406), .B1(n8957), .B2(n6408), .ZN(n6369)
         );
  XNOR2_X1 U7923 ( .A(n6369), .B(n6368), .ZN(n6372) );
  OR2_X1 U7924 ( .A1(n9192), .A2(n6408), .ZN(n6371) );
  NAND2_X1 U7925 ( .A1(n9218), .A2(n6452), .ZN(n6370) );
  NAND2_X1 U7926 ( .A1(n6372), .A2(n6373), .ZN(n6381) );
  INV_X1 U7927 ( .A(n6372), .ZN(n6375) );
  INV_X1 U7928 ( .A(n6373), .ZN(n6374) );
  NAND2_X1 U7929 ( .A1(n6375), .A2(n6374), .ZN(n6376) );
  AND2_X1 U7930 ( .A1(n6381), .A2(n6376), .ZN(n8977) );
  INV_X1 U7931 ( .A(n6378), .ZN(n6379) );
  NAND2_X1 U7932 ( .A1(n6380), .A2(n6379), .ZN(n8978) );
  NAND3_X1 U7933 ( .A1(n8979), .A2(n8977), .A3(n8978), .ZN(n8976) );
  NAND2_X1 U7934 ( .A1(n8976), .A2(n6381), .ZN(n8953) );
  NAND2_X1 U7935 ( .A1(n7847), .A2(n6082), .ZN(n6383) );
  NAND2_X1 U7936 ( .A1(n7939), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6382) );
  XNOR2_X1 U7937 ( .A(n6398), .B(P1_REG3_REG_25__SCAN_IN), .ZN(n9180) );
  INV_X1 U7938 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U7939 ( .A1(n6798), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U7940 ( .A1(n7942), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6384) );
  OAI211_X1 U7941 ( .C1(n6026), .C2(n6653), .A(n6385), .B(n6384), .ZN(n6386)
         );
  AOI21_X1 U7942 ( .B1(n9180), .B2(n6172), .A(n6386), .ZN(n9044) );
  OAI22_X1 U7943 ( .A1(n9182), .A2(n6408), .B1(n9044), .B2(n6387), .ZN(n6411)
         );
  NAND2_X1 U7944 ( .A1(n9415), .A2(n6388), .ZN(n6390) );
  OR2_X1 U7945 ( .A1(n9044), .A2(n6408), .ZN(n6389) );
  NAND2_X1 U7946 ( .A1(n6390), .A2(n6389), .ZN(n6391) );
  XNOR2_X1 U7947 ( .A(n6391), .B(n7142), .ZN(n6412) );
  XOR2_X1 U7948 ( .A(n6411), .B(n6412), .Z(n8954) );
  NAND2_X1 U7949 ( .A1(n7865), .A2(n6082), .ZN(n6393) );
  NAND2_X1 U7950 ( .A1(n7939), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6392) );
  INV_X1 U7951 ( .A(n6398), .ZN(n6395) );
  AND2_X1 U7952 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n6394) );
  NAND2_X1 U7953 ( .A1(n6395), .A2(n6394), .ZN(n6416) );
  INV_X1 U7954 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6397) );
  INV_X1 U7955 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6396) );
  OAI21_X1 U7956 ( .B1(n6398), .B2(n6397), .A(n6396), .ZN(n6399) );
  NAND2_X1 U7957 ( .A1(n6416), .A2(n6399), .ZN(n9020) );
  INV_X1 U7958 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U7959 ( .A1(n7942), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U7960 ( .A1(n5941), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6400) );
  OAI211_X1 U7961 ( .C1(n6402), .C2(n5989), .A(n6401), .B(n6400), .ZN(n6403)
         );
  INV_X1 U7962 ( .A(n6403), .ZN(n6404) );
  OAI22_X1 U7963 ( .A1(n9167), .A2(n6406), .B1(n8198), .B2(n6408), .ZN(n6407)
         );
  XNOR2_X1 U7964 ( .A(n6407), .B(n7142), .ZN(n6432) );
  OR2_X1 U7965 ( .A1(n9167), .A2(n6408), .ZN(n6410) );
  NAND2_X1 U7966 ( .A1(n9186), .A2(n6452), .ZN(n6409) );
  NAND2_X1 U7967 ( .A1(n6410), .A2(n6409), .ZN(n6431) );
  XNOR2_X1 U7968 ( .A(n6432), .B(n6431), .ZN(n9015) );
  NOR2_X1 U7969 ( .A1(n6412), .A2(n6411), .ZN(n9013) );
  NOR2_X1 U7970 ( .A1(n9015), .A2(n9013), .ZN(n6413) );
  NAND2_X1 U7971 ( .A1(n7884), .A2(n6082), .ZN(n6415) );
  NAND2_X1 U7972 ( .A1(n7939), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U7973 ( .A1(n9405), .A2(n6388), .ZN(n6425) );
  INV_X1 U7974 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U7975 ( .A1(n6416), .A2(n6632), .ZN(n6417) );
  NAND2_X1 U7976 ( .A1(n9149), .A2(n6172), .ZN(n6423) );
  INV_X1 U7977 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U7978 ( .A1(n6798), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U7979 ( .A1(n5941), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6418) );
  OAI211_X1 U7980 ( .C1(n6025), .C2(n6420), .A(n6419), .B(n6418), .ZN(n6421)
         );
  INV_X1 U7981 ( .A(n6421), .ZN(n6422) );
  NAND2_X1 U7982 ( .A1(n9173), .A2(n6448), .ZN(n6424) );
  NAND2_X1 U7983 ( .A1(n6425), .A2(n6424), .ZN(n6426) );
  XNOR2_X1 U7984 ( .A(n6426), .B(n7142), .ZN(n6430) );
  NAND2_X1 U7985 ( .A1(n9405), .A2(n6448), .ZN(n6428) );
  NAND2_X1 U7986 ( .A1(n9173), .A2(n6452), .ZN(n6427) );
  NAND2_X1 U7987 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  NOR2_X1 U7988 ( .A1(n6430), .A2(n6429), .ZN(n6480) );
  AOI21_X1 U7989 ( .B1(n6430), .B2(n6429), .A(n6480), .ZN(n8922) );
  INV_X1 U7990 ( .A(n8922), .ZN(n6434) );
  NAND2_X1 U7991 ( .A1(n6432), .A2(n6431), .ZN(n8923) );
  INV_X1 U7992 ( .A(n8923), .ZN(n6433) );
  NOR2_X1 U7993 ( .A1(n6434), .A2(n6433), .ZN(n6435) );
  NAND2_X1 U7994 ( .A1(n7903), .A2(n6082), .ZN(n6437) );
  NAND2_X1 U7995 ( .A1(n7939), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U7996 ( .A1(n9401), .A2(n6388), .ZN(n6450) );
  INV_X1 U7997 ( .A(n6440), .ZN(n6438) );
  NAND2_X1 U7998 ( .A1(n6438), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8202) );
  INV_X1 U7999 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8000 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  NAND2_X1 U8001 ( .A1(n8202), .A2(n6441), .ZN(n9141) );
  INV_X1 U8002 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8003 ( .A1(n7942), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U8004 ( .A1(n5941), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6442) );
  OAI211_X1 U8005 ( .C1(n6444), .C2(n5989), .A(n6443), .B(n6442), .ZN(n6445)
         );
  INV_X1 U8006 ( .A(n6445), .ZN(n6446) );
  NAND2_X1 U8007 ( .A1(n9043), .A2(n6448), .ZN(n6449) );
  NAND2_X1 U8008 ( .A1(n6450), .A2(n6449), .ZN(n6451) );
  XNOR2_X1 U8009 ( .A(n6451), .B(n7142), .ZN(n6454) );
  AOI22_X1 U8010 ( .A1(n9401), .A2(n6343), .B1(n6452), .B2(n9043), .ZN(n6453)
         );
  XNOR2_X1 U8011 ( .A(n6454), .B(n6453), .ZN(n6481) );
  INV_X1 U8012 ( .A(n6840), .ZN(n6458) );
  INV_X1 U8013 ( .A(n6483), .ZN(n6457) );
  NAND2_X1 U8014 ( .A1(n7850), .A2(P1_B_REG_SCAN_IN), .ZN(n6460) );
  INV_X1 U8015 ( .A(n7782), .ZN(n6459) );
  MUX2_X1 U8016 ( .A(n6460), .B(P1_B_REG_SCAN_IN), .S(n6459), .Z(n6461) );
  INV_X1 U8017 ( .A(n7850), .ZN(n6462) );
  OAI22_X1 U8018 ( .A1(n6734), .A2(P1_D_REG_1__SCAN_IN), .B1(n6473), .B2(n6462), .ZN(n6831) );
  NOR4_X1 U8019 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6466) );
  NOR4_X1 U8020 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6465) );
  NOR4_X1 U8021 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6464) );
  NOR4_X1 U8022 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6463) );
  AND4_X1 U8023 ( .A1(n6466), .A2(n6465), .A3(n6464), .A4(n6463), .ZN(n6472)
         );
  NOR2_X1 U8024 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .ZN(
        n6470) );
  NOR4_X1 U8025 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6469) );
  NOR4_X1 U8026 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6468) );
  NOR4_X1 U8027 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6467) );
  AND4_X1 U8028 ( .A1(n6470), .A2(n6469), .A3(n6468), .A4(n6467), .ZN(n6471)
         );
  NAND2_X1 U8029 ( .A1(n6472), .A2(n6471), .ZN(n6564) );
  INV_X1 U8030 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6737) );
  NOR2_X1 U8031 ( .A1(n6564), .A2(n6737), .ZN(n6474) );
  INV_X1 U8032 ( .A(n6473), .ZN(n7867) );
  NAND2_X1 U8033 ( .A1(n7867), .A2(n7782), .ZN(n6735) );
  OAI21_X1 U8034 ( .B1(n6734), .B2(n6474), .A(n6735), .ZN(n6833) );
  OR2_X1 U8035 ( .A1(n6831), .A2(n6833), .ZN(n6486) );
  OAI21_X1 U8036 ( .B1(n6475), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6476) );
  INV_X1 U8037 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6701) );
  INV_X1 U8038 ( .A(n9515), .ZN(n8177) );
  NOR2_X1 U8039 ( .A1(n6486), .A2(n8177), .ZN(n6498) );
  AND2_X1 U8040 ( .A1(n6498), .A2(n8166), .ZN(n6479) );
  AND2_X1 U8041 ( .A1(n6481), .A2(n9018), .ZN(n6507) );
  NAND3_X1 U8042 ( .A1(n6481), .A2(n9018), .A3(n6480), .ZN(n6506) );
  AND2_X1 U8043 ( .A1(n6486), .A2(n9515), .ZN(n6482) );
  NOR2_X1 U8044 ( .A1(n6840), .A2(n7244), .ZN(n9727) );
  NAND2_X1 U8045 ( .A1(n6482), .A2(n9727), .ZN(n6810) );
  NOR2_X1 U8046 ( .A1(n9765), .A2(n6834), .ZN(n6484) );
  AND3_X1 U8047 ( .A1(n6485), .A2(n6513), .A3(n6512), .ZN(n6488) );
  INV_X1 U8048 ( .A(n6486), .ZN(n6487) );
  OR2_X1 U8049 ( .A1(n9487), .A2(n6487), .ZN(n6808) );
  NAND2_X1 U8050 ( .A1(n6488), .A2(n6808), .ZN(n6489) );
  NAND2_X1 U8051 ( .A1(n6489), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6490) );
  OR2_X1 U8052 ( .A1(n8202), .A2(n6491), .ZN(n6497) );
  INV_X1 U8053 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U8054 ( .A1(n7942), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U8055 ( .A1(n5941), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6492) );
  OAI211_X1 U8056 ( .C1(n6494), .C2(n5989), .A(n6493), .B(n6492), .ZN(n6495)
         );
  INV_X1 U8057 ( .A(n6495), .ZN(n6496) );
  INV_X1 U8058 ( .A(n9131), .ZN(n9042) );
  INV_X1 U8059 ( .A(n6498), .ZN(n6500) );
  OR2_X1 U8060 ( .A1(n6499), .A2(n6557), .ZN(n8178) );
  NOR2_X1 U8061 ( .A1(n6500), .A2(n8178), .ZN(n6501) );
  NAND2_X1 U8062 ( .A1(n6501), .A2(n9624), .ZN(n9036) );
  AOI22_X1 U8063 ( .A1(n9042), .A2(n9021), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6503) );
  NAND2_X1 U8064 ( .A1(n9173), .A2(n9033), .ZN(n6502) );
  OAI211_X1 U8065 ( .C1(n9000), .C2(n9141), .A(n6503), .B(n6502), .ZN(n6504)
         );
  AOI21_X1 U8066 ( .B1(n9401), .B2(n9038), .A(n6504), .ZN(n6505) );
  AOI21_X1 U8067 ( .B1(n8924), .B2(n6507), .A(n4825), .ZN(n6508) );
  NAND2_X1 U8068 ( .A1(n6509), .A2(n6508), .ZN(P1_U3218) );
  NAND2_X1 U8069 ( .A1(n8166), .A2(n6513), .ZN(n6510) );
  NAND2_X1 U8070 ( .A1(n6510), .A2(n6512), .ZN(n6537) );
  NAND2_X1 U8071 ( .A1(n6537), .A2(n6511), .ZN(n6757) );
  NAND2_X1 U8072 ( .A1(n6757), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8073 ( .A(n6512), .ZN(n7572) );
  AND2_X1 U8074 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7495) );
  MUX2_X1 U8075 ( .A(n7400), .B(P1_REG2_REG_7__SCAN_IN), .S(n6786), .Z(n6779)
         );
  NAND2_X1 U8076 ( .A1(n6771), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U8077 ( .A1(n9529), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U8078 ( .A1(n6527), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6515) );
  INV_X1 U8079 ( .A(n6514), .ZN(n9628) );
  XNOR2_X1 U8080 ( .A(n6582), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9610) );
  NAND3_X1 U8081 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .A3(n9610), .ZN(n9609) );
  OAI21_X1 U8082 ( .B1(n6582), .B2(n9742), .A(n9609), .ZN(n9627) );
  NAND2_X1 U8083 ( .A1(n9628), .A2(n9627), .ZN(n9626) );
  NAND2_X1 U8084 ( .A1(n6515), .A2(n9626), .ZN(n9531) );
  INV_X1 U8085 ( .A(n9529), .ZN(n6590) );
  INV_X1 U8086 ( .A(n6517), .ZN(n6516) );
  AOI21_X1 U8087 ( .B1(n5979), .B2(n6590), .A(n6516), .ZN(n9532) );
  NAND2_X1 U8088 ( .A1(n9531), .A2(n9532), .ZN(n9530) );
  NAND2_X1 U8089 ( .A1(n6517), .A2(n9530), .ZN(n9639) );
  INV_X1 U8090 ( .A(n6526), .ZN(n9640) );
  AOI22_X1 U8091 ( .A1(n6526), .A2(n5991), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n9640), .ZN(n9638) );
  INV_X1 U8092 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6518) );
  MUX2_X1 U8093 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6518), .S(n9653), .Z(n6519)
         );
  INV_X1 U8094 ( .A(n6519), .ZN(n9655) );
  MUX2_X1 U8095 ( .A(n6520), .B(P1_REG2_REG_6__SCAN_IN), .S(n6597), .Z(n6773)
         );
  NAND2_X1 U8096 ( .A1(n6774), .A2(n6773), .ZN(n6772) );
  NAND2_X1 U8097 ( .A1(n6521), .A2(n6772), .ZN(n6780) );
  NOR2_X1 U8098 ( .A1(n9676), .A2(n7384), .ZN(n9672) );
  OAI22_X1 U8099 ( .A1(n9672), .A2(n9665), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n6522), .ZN(n9678) );
  NAND2_X1 U8100 ( .A1(n6858), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6523) );
  OAI21_X1 U8101 ( .B1(n6858), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6523), .ZN(
        n6524) );
  NOR2_X1 U8102 ( .A1(n9620), .A2(P1_U3084), .ZN(n7885) );
  NAND2_X1 U8103 ( .A1(n6537), .A2(n7885), .ZN(n9108) );
  AOI211_X1 U8104 ( .C1(n9678), .C2(n6524), .A(n6857), .B(n9688), .ZN(n6542)
         );
  NOR2_X1 U8105 ( .A1(n6771), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8106 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9653), .ZN(n6531) );
  INV_X1 U8107 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6525) );
  MUX2_X1 U8108 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6525), .S(n9653), .Z(n9659)
         );
  NOR2_X1 U8109 ( .A1(n6526), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6530) );
  MUX2_X1 U8110 ( .A(n5990), .B(P1_REG1_REG_4__SCAN_IN), .S(n6526), .Z(n9645)
         );
  INV_X1 U8111 ( .A(n6527), .ZN(n9630) );
  INV_X1 U8112 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9776) );
  XNOR2_X1 U8113 ( .A(n9630), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U8114 ( .A1(n9608), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6529) );
  INV_X1 U8115 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6528) );
  MUX2_X1 U8116 ( .A(n6528), .B(P1_REG1_REG_1__SCAN_IN), .S(n6582), .Z(n9613)
         );
  NAND3_X1 U8117 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n9613), .ZN(n9612) );
  NAND2_X1 U8118 ( .A1(n6529), .A2(n9612), .ZN(n9634) );
  NAND2_X1 U8119 ( .A1(n9633), .A2(n9634), .ZN(n9632) );
  OAI21_X1 U8120 ( .B1(n9630), .B2(n9776), .A(n9632), .ZN(n9535) );
  MUX2_X1 U8121 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7111), .S(n9529), .Z(n9534)
         );
  NAND2_X1 U8122 ( .A1(n9535), .A2(n9534), .ZN(n9533) );
  OAI21_X1 U8123 ( .B1(n7111), .B2(n6590), .A(n9533), .ZN(n9646) );
  NOR2_X1 U8124 ( .A1(n9645), .A2(n9646), .ZN(n9644) );
  NOR2_X1 U8125 ( .A1(n6530), .A2(n9644), .ZN(n9660) );
  NAND2_X1 U8126 ( .A1(n9659), .A2(n9660), .ZN(n9658) );
  NAND2_X1 U8127 ( .A1(n6531), .A2(n9658), .ZN(n6768) );
  INV_X1 U8128 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9780) );
  AOI22_X1 U8129 ( .A1(n6771), .A2(n9780), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6597), .ZN(n6767) );
  NOR2_X1 U8130 ( .A1(n6768), .A2(n6767), .ZN(n6766) );
  NOR2_X1 U8131 ( .A1(n6532), .A2(n6766), .ZN(n6783) );
  INV_X1 U8132 ( .A(n6786), .ZN(n6593) );
  INV_X1 U8133 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7461) );
  AOI22_X1 U8134 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6593), .B1(n6786), .B2(
        n7461), .ZN(n6782) );
  NOR2_X1 U8135 ( .A1(n6783), .A2(n6782), .ZN(n6781) );
  NOR2_X1 U8136 ( .A1(n6786), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6533) );
  NOR2_X1 U8137 ( .A1(n6781), .A2(n6533), .ZN(n9680) );
  AND2_X1 U8138 ( .A1(n9665), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9679) );
  OAI22_X1 U8139 ( .A1(n9680), .A2(n9679), .B1(n9665), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n9669) );
  INV_X1 U8140 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6534) );
  MUX2_X1 U8141 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6534), .S(n6858), .Z(n6535)
         );
  NAND2_X1 U8142 ( .A1(n6535), .A2(n9669), .ZN(n6850) );
  OAI21_X1 U8143 ( .B1(n9669), .B2(n6535), .A(n6850), .ZN(n6538) );
  NOR2_X1 U8144 ( .A1(n9624), .A2(P1_U3084), .ZN(n7904) );
  AND2_X1 U8145 ( .A1(n7904), .A2(n9620), .ZN(n6536) );
  AND2_X1 U8146 ( .A1(n6538), .A2(n9712), .ZN(n6541) );
  INV_X1 U8147 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10002) );
  OAI22_X1 U8148 ( .A1(n9641), .A2(n6729), .B1(n9112), .B2(n10002), .ZN(n6540)
         );
  OR4_X1 U8149 ( .A1(n7495), .A2(n6542), .A3(n6541), .A4(n6540), .ZN(P1_U3250)
         );
  NAND2_X1 U8150 ( .A1(n7101), .A2(n6543), .ZN(n7989) );
  NAND2_X1 U8151 ( .A1(n6818), .A2(n9755), .ZN(n7991) );
  NAND2_X1 U8152 ( .A1(n7989), .A2(n7991), .ZN(n8022) );
  INV_X1 U8153 ( .A(n8022), .ZN(n6554) );
  NAND2_X1 U8154 ( .A1(n6545), .A2(n6553), .ZN(n6551) );
  INV_X1 U8155 ( .A(n9731), .ZN(n6841) );
  INV_X1 U8156 ( .A(n6544), .ZN(n6838) );
  NAND2_X1 U8157 ( .A1(n6838), .A2(n9730), .ZN(n6546) );
  NAND2_X1 U8158 ( .A1(n7994), .A2(n6554), .ZN(n7102) );
  OAI21_X1 U8159 ( .B1(n6554), .B2(n7994), .A(n7102), .ZN(n6550) );
  NAND2_X1 U8160 ( .A1(n6478), .A2(n9736), .ZN(n6549) );
  NAND2_X1 U8161 ( .A1(n8172), .A2(n8175), .ZN(n6548) );
  NAND2_X1 U8162 ( .A1(n6550), .A2(n9725), .ZN(n6563) );
  AND2_X1 U8163 ( .A1(n8022), .A2(n6553), .ZN(n6552) );
  INV_X1 U8164 ( .A(n6551), .ZN(n9718) );
  NAND2_X1 U8165 ( .A1(n6552), .A2(n9717), .ZN(n7100) );
  NAND2_X1 U8166 ( .A1(n9717), .A2(n6553), .ZN(n6555) );
  NAND2_X1 U8167 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  NAND2_X1 U8168 ( .A1(n7100), .A2(n6556), .ZN(n9759) );
  OR2_X1 U8169 ( .A1(n9735), .A2(n6557), .ZN(n6559) );
  OR2_X1 U8170 ( .A1(n6570), .A2(n8054), .ZN(n6558) );
  INV_X1 U8171 ( .A(n9723), .ZN(n9549) );
  NAND2_X1 U8172 ( .A1(n9759), .A2(n9549), .ZN(n6562) );
  INV_X1 U8173 ( .A(n8166), .ZN(n6560) );
  AOI22_X1 U8174 ( .A1(n9050), .A2(n9721), .B1(n9720), .B2(n6544), .ZN(n6561)
         );
  NAND3_X1 U8175 ( .A1(n6563), .A2(n6562), .A3(n6561), .ZN(n9757) );
  INV_X1 U8176 ( .A(n6564), .ZN(n6566) );
  OAI21_X1 U8177 ( .B1(n6734), .B2(P1_D_REG_0__SCAN_IN), .A(n6735), .ZN(n6565)
         );
  OAI21_X1 U8178 ( .B1(n6566), .B2(n6734), .A(n6565), .ZN(n6567) );
  INV_X1 U8179 ( .A(n6831), .ZN(n9516) );
  NAND2_X1 U8180 ( .A1(n6844), .A2(n9516), .ZN(n7165) );
  NAND2_X1 U8181 ( .A1(n9515), .A2(n9736), .ZN(n6568) );
  MUX2_X1 U8182 ( .A(n9757), .B(P1_REG2_REG_2__SCAN_IN), .S(n9743), .Z(n6575)
         );
  INV_X1 U8183 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6569) );
  OAI22_X1 U8184 ( .A1(n9341), .A2(n9755), .B1(n9142), .B2(n6569), .ZN(n6574)
         );
  INV_X1 U8185 ( .A(n9759), .ZN(n6572) );
  NAND3_X1 U8186 ( .A1(n9740), .A2(n9736), .A3(n9735), .ZN(n9343) );
  NOR2_X1 U8187 ( .A1(n6570), .A2(n8172), .ZN(n6571) );
  INV_X1 U8188 ( .A(n9346), .ZN(n9384) );
  NAND2_X1 U8189 ( .A1(n9729), .A2(n9755), .ZN(n7106) );
  OAI21_X1 U8190 ( .B1(n9729), .B2(n9755), .A(n7106), .ZN(n9756) );
  OAI22_X1 U8191 ( .A1(n6572), .A2(n9343), .B1(n9384), .B2(n9756), .ZN(n6573)
         );
  OR3_X1 U8192 ( .A1(n6575), .A2(n6574), .A3(n6573), .ZN(P1_U3289) );
  INV_X2 U8193 ( .A(n7592), .ZN(n8920) );
  INV_X1 U8194 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6576) );
  INV_X2 U8195 ( .A(n8918), .ZN(n8259) );
  OAI222_X1 U8196 ( .A1(n6978), .A2(P2_U3152), .B1(n8920), .B2(n6583), .C1(
        n6576), .C2(n8259), .ZN(P2_U3357) );
  OAI222_X1 U8197 ( .A1(n6991), .A2(P2_U3152), .B1(n8920), .B2(n6588), .C1(
        n4479), .C2(n8259), .ZN(P2_U3356) );
  OAI222_X1 U8198 ( .A1(n6965), .A2(P2_U3152), .B1(n8920), .B2(n6591), .C1(
        n6577), .C2(n8259), .ZN(P2_U3355) );
  OAI222_X1 U8199 ( .A1(n6950), .A2(P2_U3152), .B1(n8920), .B2(n6586), .C1(
        n6578), .C2(n8259), .ZN(P2_U3354) );
  OAI222_X1 U8200 ( .A1(n6898), .A2(P2_U3152), .B1(n8920), .B2(n6585), .C1(
        n6579), .C2(n8259), .ZN(P2_U3353) );
  NAND2_X1 U8201 ( .A1(n6581), .A2(P1_U3084), .ZN(n9527) );
  OAI222_X1 U8202 ( .A1(n9524), .A2(n4445), .B1(n9527), .B2(n6583), .C1(
        P1_U3084), .C2(n6582), .ZN(P1_U3352) );
  INV_X1 U8203 ( .A(n9527), .ZN(n6601) );
  INV_X1 U8204 ( .A(n9524), .ZN(n9520) );
  AOI22_X1 U8205 ( .A1(n9653), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9520), .ZN(n6584) );
  OAI21_X1 U8206 ( .B1(n6585), .B2(n9522), .A(n6584), .ZN(P1_U3348) );
  OAI222_X1 U8207 ( .A1(n9524), .A2(n6587), .B1(n9522), .B2(n6586), .C1(
        P1_U3084), .C2(n9640), .ZN(P1_U3349) );
  OAI222_X1 U8208 ( .A1(n9524), .A2(n6589), .B1(n9522), .B2(n6588), .C1(
        P1_U3084), .C2(n9630), .ZN(P1_U3351) );
  OAI222_X1 U8209 ( .A1(n9524), .A2(n6592), .B1(n9522), .B2(n6591), .C1(
        P1_U3084), .C2(n6590), .ZN(P1_U3350) );
  INV_X1 U8210 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6594) );
  OAI222_X1 U8211 ( .A1(n9524), .A2(n6594), .B1(n9522), .B2(n6596), .C1(
        P1_U3084), .C2(n6593), .ZN(P1_U3346) );
  INV_X1 U8212 ( .A(n6920), .ZN(n6939) );
  OAI222_X1 U8213 ( .A1(n6939), .A2(P2_U3152), .B1(n8920), .B2(n6596), .C1(
        n6595), .C2(n8259), .ZN(P2_U3351) );
  INV_X1 U8214 ( .A(n7030), .ZN(n7039) );
  INV_X1 U8215 ( .A(n6602), .ZN(n6600) );
  OAI222_X1 U8216 ( .A1(n7039), .A2(P2_U3152), .B1(n8920), .B2(n6600), .C1(
        n6599), .C2(n8259), .ZN(P2_U3350) );
  AOI222_X1 U8217 ( .A1(n6602), .A2(n6601), .B1(P2_DATAO_REG_8__SCAN_IN), .B2(
        n9520), .C1(P1_STATE_REG_SCAN_IN), .C2(n9665), .ZN(n6726) );
  NOR2_X1 U8218 ( .A1(keyinput20), .A2(keyinput5), .ZN(n6603) );
  NAND3_X1 U8219 ( .A1(keyinput7), .A2(keyinput12), .A3(n6603), .ZN(n6615) );
  NAND4_X1 U8220 ( .A1(keyinput39), .A2(keyinput33), .A3(keyinput63), .A4(
        keyinput54), .ZN(n6614) );
  NOR4_X1 U8221 ( .A1(keyinput55), .A2(keyinput47), .A3(keyinput29), .A4(
        keyinput32), .ZN(n6605) );
  NOR2_X1 U8222 ( .A1(keyinput4), .A2(keyinput19), .ZN(n6604) );
  NAND4_X1 U8223 ( .A1(n6605), .A2(keyinput52), .A3(keyinput34), .A4(n6604), 
        .ZN(n6613) );
  NOR3_X1 U8224 ( .A1(keyinput43), .A2(keyinput6), .A3(keyinput35), .ZN(n6611)
         );
  INV_X1 U8225 ( .A(keyinput17), .ZN(n6606) );
  NOR4_X1 U8226 ( .A1(keyinput42), .A2(keyinput21), .A3(keyinput11), .A4(n6606), .ZN(n6610) );
  NAND2_X1 U8227 ( .A1(keyinput13), .A2(keyinput22), .ZN(n6608) );
  NAND4_X1 U8228 ( .A1(keyinput15), .A2(keyinput1), .A3(keyinput41), .A4(
        keyinput23), .ZN(n6607) );
  NOR4_X1 U8229 ( .A1(keyinput3), .A2(keyinput38), .A3(n6608), .A4(n6607), 
        .ZN(n6609) );
  NAND4_X1 U8230 ( .A1(keyinput14), .A2(n6611), .A3(n6610), .A4(n6609), .ZN(
        n6612) );
  NOR4_X1 U8231 ( .A1(n6615), .A2(n6614), .A3(n6613), .A4(n6612), .ZN(n6724)
         );
  NAND3_X1 U8232 ( .A1(keyinput26), .A2(keyinput40), .A3(keyinput59), .ZN(
        n6629) );
  NOR3_X1 U8233 ( .A1(keyinput18), .A2(keyinput50), .A3(keyinput9), .ZN(n6620)
         );
  NAND2_X1 U8234 ( .A1(keyinput16), .A2(keyinput25), .ZN(n6616) );
  NOR3_X1 U8235 ( .A1(keyinput51), .A2(keyinput28), .A3(n6616), .ZN(n6619) );
  NAND2_X1 U8236 ( .A1(keyinput48), .A2(keyinput56), .ZN(n6617) );
  NOR3_X1 U8237 ( .A1(keyinput45), .A2(keyinput2), .A3(n6617), .ZN(n6618) );
  NAND4_X1 U8238 ( .A1(keyinput61), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(
        n6628) );
  NOR2_X1 U8239 ( .A1(keyinput60), .A2(keyinput30), .ZN(n6626) );
  NAND2_X1 U8240 ( .A1(keyinput24), .A2(keyinput57), .ZN(n6624) );
  NOR3_X1 U8241 ( .A1(keyinput27), .A2(keyinput31), .A3(keyinput53), .ZN(n6622) );
  NOR3_X1 U8242 ( .A1(keyinput46), .A2(keyinput62), .A3(keyinput58), .ZN(n6621) );
  NAND4_X1 U8243 ( .A1(keyinput0), .A2(n6622), .A3(keyinput36), .A4(n6621), 
        .ZN(n6623) );
  NOR4_X1 U8244 ( .A1(keyinput10), .A2(keyinput8), .A3(n6624), .A4(n6623), 
        .ZN(n6625) );
  NAND4_X1 U8245 ( .A1(keyinput37), .A2(keyinput44), .A3(n6626), .A4(n6625), 
        .ZN(n6627) );
  NOR4_X1 U8246 ( .A1(keyinput49), .A2(n6629), .A3(n6628), .A4(n6627), .ZN(
        n6723) );
  AOI22_X1 U8247 ( .A1(n8498), .A2(keyinput49), .B1(n6420), .B2(keyinput26), 
        .ZN(n6630) );
  OAI221_X1 U8248 ( .B1(n8498), .B2(keyinput49), .C1(n6420), .C2(keyinput26), 
        .A(n6630), .ZN(n6640) );
  AOI22_X1 U8249 ( .A1(n6633), .A2(keyinput61), .B1(n6632), .B2(keyinput18), 
        .ZN(n6631) );
  OAI221_X1 U8250 ( .B1(n6633), .B2(keyinput61), .C1(n6632), .C2(keyinput18), 
        .A(n6631), .ZN(n6639) );
  XOR2_X1 U8251 ( .A(n5961), .B(keyinput50), .Z(n6637) );
  XNOR2_X1 U8252 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput9), .ZN(n6636) );
  XNOR2_X1 U8253 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput40), .ZN(n6635) );
  XNOR2_X1 U8254 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput59), .ZN(n6634) );
  NAND4_X1 U8255 ( .A1(n6637), .A2(n6636), .A3(n6635), .A4(n6634), .ZN(n6638)
         );
  NOR3_X1 U8256 ( .A1(n6640), .A2(n6639), .A3(n6638), .ZN(n6676) );
  AOI22_X1 U8257 ( .A1(n5928), .A2(keyinput51), .B1(n6642), .B2(keyinput25), 
        .ZN(n6641) );
  OAI221_X1 U8258 ( .B1(n5928), .B2(keyinput51), .C1(n6642), .C2(keyinput25), 
        .A(n6641), .ZN(n6650) );
  INV_X1 U8259 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6799) );
  INV_X1 U8260 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9744) );
  AOI22_X1 U8261 ( .A1(n6799), .A2(keyinput16), .B1(n9744), .B2(keyinput28), 
        .ZN(n6643) );
  OAI221_X1 U8262 ( .B1(n6799), .B2(keyinput16), .C1(n9744), .C2(keyinput28), 
        .A(n6643), .ZN(n6649) );
  AOI22_X1 U8263 ( .A1(n6193), .A2(keyinput45), .B1(n6137), .B2(keyinput2), 
        .ZN(n6644) );
  OAI221_X1 U8264 ( .B1(n6193), .B2(keyinput45), .C1(n6137), .C2(keyinput2), 
        .A(n6644), .ZN(n6648) );
  INV_X1 U8265 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6646) );
  AOI22_X1 U8266 ( .A1(n6646), .A2(keyinput56), .B1(n6829), .B2(keyinput48), 
        .ZN(n6645) );
  OAI221_X1 U8267 ( .B1(n6646), .B2(keyinput56), .C1(n6829), .C2(keyinput48), 
        .A(n6645), .ZN(n6647) );
  NOR4_X1 U8268 ( .A1(n6650), .A2(n6649), .A3(n6648), .A4(n6647), .ZN(n6675)
         );
  INV_X1 U8269 ( .A(P1_RD_REG_SCAN_IN), .ZN(n9607) );
  INV_X1 U8270 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6848) );
  AOI22_X1 U8271 ( .A1(n9607), .A2(keyinput60), .B1(keyinput30), .B2(n6848), 
        .ZN(n6651) );
  OAI221_X1 U8272 ( .B1(n9607), .B2(keyinput60), .C1(n6848), .C2(keyinput30), 
        .A(n6651), .ZN(n6662) );
  INV_X1 U8273 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9746) );
  AOI22_X1 U8274 ( .A1(n6653), .A2(keyinput37), .B1(n9746), .B2(keyinput44), 
        .ZN(n6652) );
  OAI221_X1 U8275 ( .B1(n6653), .B2(keyinput37), .C1(n9746), .C2(keyinput44), 
        .A(n6652), .ZN(n6661) );
  INV_X1 U8276 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6656) );
  AOI22_X1 U8277 ( .A1(n6656), .A2(keyinput27), .B1(keyinput31), .B2(n6655), 
        .ZN(n6654) );
  OAI221_X1 U8278 ( .B1(n6656), .B2(keyinput27), .C1(n6655), .C2(keyinput31), 
        .A(n6654), .ZN(n6660) );
  INV_X1 U8279 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6658) );
  INV_X1 U8280 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U8281 ( .A1(n6658), .A2(keyinput53), .B1(n9955), .B2(keyinput0), 
        .ZN(n6657) );
  OAI221_X1 U8282 ( .B1(n6658), .B2(keyinput53), .C1(n9955), .C2(keyinput0), 
        .A(n6657), .ZN(n6659) );
  NOR4_X1 U8283 ( .A1(n6662), .A2(n6661), .A3(n6660), .A4(n6659), .ZN(n6674)
         );
  INV_X1 U8284 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7614) );
  AOI22_X1 U8285 ( .A1(n9776), .A2(keyinput57), .B1(keyinput8), .B2(n7614), 
        .ZN(n6663) );
  OAI221_X1 U8286 ( .B1(n9776), .B2(keyinput57), .C1(n7614), .C2(keyinput8), 
        .A(n6663), .ZN(n6672) );
  AOI22_X1 U8287 ( .A1(n9842), .A2(keyinput24), .B1(n6791), .B2(keyinput10), 
        .ZN(n6664) );
  OAI221_X1 U8288 ( .B1(n9842), .B2(keyinput24), .C1(n6791), .C2(keyinput10), 
        .A(n6664), .ZN(n6671) );
  INV_X1 U8289 ( .A(SI_17_), .ZN(n6666) );
  AOI22_X1 U8290 ( .A1(n6666), .A2(keyinput36), .B1(n7781), .B2(keyinput58), 
        .ZN(n6665) );
  OAI221_X1 U8291 ( .B1(n6666), .B2(keyinput36), .C1(n7781), .C2(keyinput58), 
        .A(n6665), .ZN(n6670) );
  XNOR2_X1 U8292 ( .A(P2_IR_REG_30__SCAN_IN), .B(keyinput62), .ZN(n6668) );
  XNOR2_X1 U8293 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput46), .ZN(n6667) );
  NAND2_X1 U8294 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  NOR4_X1 U8295 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n6673)
         );
  NAND4_X1 U8296 ( .A1(n6676), .A2(n6675), .A3(n6674), .A4(n6673), .ZN(n6722)
         );
  AOI22_X1 U8297 ( .A1(n6520), .A2(keyinput19), .B1(keyinput34), .B2(n6678), 
        .ZN(n6677) );
  OAI221_X1 U8298 ( .B1(n6520), .B2(keyinput19), .C1(n6678), .C2(keyinput34), 
        .A(n6677), .ZN(n6686) );
  INV_X1 U8299 ( .A(SI_18_), .ZN(n6680) );
  AOI22_X1 U8300 ( .A1(n6730), .A2(keyinput4), .B1(n6680), .B2(keyinput52), 
        .ZN(n6679) );
  OAI221_X1 U8301 ( .B1(n6730), .B2(keyinput4), .C1(n6680), .C2(keyinput52), 
        .A(n6679), .ZN(n6685) );
  AOI22_X1 U8302 ( .A1(n6027), .A2(keyinput63), .B1(keyinput54), .B2(n9840), 
        .ZN(n6681) );
  OAI221_X1 U8303 ( .B1(n6027), .B2(keyinput63), .C1(n9840), .C2(keyinput54), 
        .A(n6681), .ZN(n6684) );
  INV_X1 U8304 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9102) );
  INV_X1 U8305 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7637) );
  AOI22_X1 U8306 ( .A1(n9102), .A2(keyinput39), .B1(keyinput33), .B2(n7637), 
        .ZN(n6682) );
  OAI221_X1 U8307 ( .B1(n9102), .B2(keyinput39), .C1(n7637), .C2(keyinput33), 
        .A(n6682), .ZN(n6683) );
  NOR4_X1 U8308 ( .A1(n6686), .A2(n6685), .A3(n6684), .A4(n6683), .ZN(n6720)
         );
  INV_X1 U8309 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7804) );
  AOI22_X1 U8310 ( .A1(n5494), .A2(keyinput29), .B1(keyinput32), .B2(n7804), 
        .ZN(n6687) );
  OAI221_X1 U8311 ( .B1(n5494), .B2(keyinput29), .C1(n7804), .C2(keyinput32), 
        .A(n6687), .ZN(n6696) );
  INV_X1 U8312 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n6689) );
  AOI22_X1 U8313 ( .A1(n6689), .A2(keyinput20), .B1(n6439), .B2(keyinput7), 
        .ZN(n6688) );
  OAI221_X1 U8314 ( .B1(n6689), .B2(keyinput20), .C1(n6439), .C2(keyinput7), 
        .A(n6688), .ZN(n6695) );
  XNOR2_X1 U8315 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput55), .ZN(n6693) );
  XNOR2_X1 U8316 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput47), .ZN(n6692) );
  XNOR2_X1 U8317 ( .A(P1_REG1_REG_31__SCAN_IN), .B(keyinput5), .ZN(n6691) );
  XNOR2_X1 U8318 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput12), .ZN(n6690) );
  NAND4_X1 U8319 ( .A1(n6693), .A2(n6692), .A3(n6691), .A4(n6690), .ZN(n6694)
         );
  NOR3_X1 U8320 ( .A1(n6696), .A2(n6695), .A3(n6694), .ZN(n6719) );
  AOI22_X1 U8321 ( .A1(n7414), .A2(keyinput41), .B1(keyinput23), .B2(n5644), 
        .ZN(n6697) );
  OAI221_X1 U8322 ( .B1(n7414), .B2(keyinput41), .C1(n5644), .C2(keyinput23), 
        .A(n6697), .ZN(n6707) );
  INV_X1 U8323 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9745) );
  AOI22_X1 U8324 ( .A1(n9745), .A2(keyinput15), .B1(keyinput1), .B2(n6699), 
        .ZN(n6698) );
  OAI221_X1 U8325 ( .B1(n9745), .B2(keyinput15), .C1(n6699), .C2(keyinput1), 
        .A(n6698), .ZN(n6706) );
  AOI22_X1 U8326 ( .A1(n6701), .A2(keyinput42), .B1(keyinput11), .B2(n5908), 
        .ZN(n6700) );
  OAI221_X1 U8327 ( .B1(n6701), .B2(keyinput42), .C1(n5908), .C2(keyinput11), 
        .A(n6700), .ZN(n6705) );
  INV_X1 U8328 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7893) );
  INV_X1 U8329 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6703) );
  AOI22_X1 U8330 ( .A1(n7893), .A2(keyinput17), .B1(keyinput21), .B2(n6703), 
        .ZN(n6702) );
  OAI221_X1 U8331 ( .B1(n7893), .B2(keyinput17), .C1(n6703), .C2(keyinput21), 
        .A(n6702), .ZN(n6704) );
  NOR4_X1 U8332 ( .A1(n6707), .A2(n6706), .A3(n6705), .A4(n6704), .ZN(n6718)
         );
  INV_X1 U8333 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U8334 ( .A1(n7252), .A2(keyinput38), .B1(keyinput22), .B2(n9959), 
        .ZN(n6708) );
  OAI221_X1 U8335 ( .B1(n7252), .B2(keyinput38), .C1(n9959), .C2(keyinput22), 
        .A(n6708), .ZN(n6716) );
  AOI22_X1 U8336 ( .A1(n5114), .A2(keyinput43), .B1(keyinput6), .B2(n9861), 
        .ZN(n6709) );
  OAI221_X1 U8337 ( .B1(n5114), .B2(keyinput43), .C1(n9861), .C2(keyinput6), 
        .A(n6709), .ZN(n6715) );
  XOR2_X1 U8338 ( .A(n8572), .B(keyinput3), .Z(n6713) );
  INV_X1 U8339 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7052) );
  XOR2_X1 U8340 ( .A(n7052), .B(keyinput14), .Z(n6712) );
  XNOR2_X1 U8341 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput13), .ZN(n6711) );
  XNOR2_X1 U8342 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput35), .ZN(n6710) );
  NAND4_X1 U8343 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6714)
         );
  NOR3_X1 U8344 ( .A1(n6716), .A2(n6715), .A3(n6714), .ZN(n6717) );
  NAND4_X1 U8345 ( .A1(n6720), .A2(n6719), .A3(n6718), .A4(n6717), .ZN(n6721)
         );
  AOI211_X1 U8346 ( .C1(n6724), .C2(n6723), .A(n6722), .B(n6721), .ZN(n6725)
         );
  XNOR2_X1 U8347 ( .A(n6726), .B(n6725), .ZN(P1_U3345) );
  INV_X1 U8348 ( .A(n6727), .ZN(n6731) );
  OAI222_X1 U8349 ( .A1(n9527), .A2(n6731), .B1(n6729), .B2(P1_U3084), .C1(
        n6728), .C2(n9524), .ZN(P1_U3344) );
  INV_X1 U8350 ( .A(n7128), .ZN(n7044) );
  OAI222_X1 U8351 ( .A1(P2_U3152), .A2(n7044), .B1(n8920), .B2(n6731), .C1(
        n6730), .C2(n8259), .ZN(P2_U3349) );
  INV_X1 U8352 ( .A(n6732), .ZN(n6739) );
  INV_X1 U8353 ( .A(n9695), .ZN(n6849) );
  OAI222_X1 U8354 ( .A1(n9527), .A2(n6739), .B1(n6849), .B2(P1_U3084), .C1(
        n6733), .C2(n9524), .ZN(P1_U3343) );
  INV_X1 U8355 ( .A(n9748), .ZN(n9747) );
  OAI21_X1 U8356 ( .B1(n9747), .B2(P1_D_REG_0__SCAN_IN), .A(n6735), .ZN(n6736)
         );
  OAI21_X1 U8357 ( .B1(n9515), .B2(n6737), .A(n6736), .ZN(P1_U3440) );
  INV_X1 U8358 ( .A(n7341), .ZN(n7136) );
  OAI222_X1 U8359 ( .A1(P2_U3152), .A2(n7136), .B1(n8920), .B2(n6739), .C1(
        n6738), .C2(n8259), .ZN(P2_U3348) );
  INV_X1 U8360 ( .A(n6740), .ZN(n6742) );
  INV_X1 U8361 ( .A(n6860), .ZN(n9054) );
  OAI222_X1 U8362 ( .A1(n9522), .A2(n6742), .B1(n9054), .B2(P1_U3084), .C1(
        n6741), .C2(n9524), .ZN(P1_U3342) );
  INV_X1 U8363 ( .A(n7473), .ZN(n7468) );
  OAI222_X1 U8364 ( .A1(n8259), .A2(n6743), .B1(n8920), .B2(n6742), .C1(
        P2_U3152), .C2(n7468), .ZN(P2_U3347) );
  NAND2_X1 U8365 ( .A1(n6744), .A2(P2_U3966), .ZN(n6745) );
  OAI21_X1 U8366 ( .B1(P2_U3966), .B2(n4391), .A(n6745), .ZN(P2_U3583) );
  INV_X1 U8367 ( .A(n6746), .ZN(n6748) );
  INV_X1 U8368 ( .A(n7702), .ZN(n7483) );
  OAI222_X1 U8369 ( .A1(n8259), .A2(n6747), .B1(n8920), .B2(n6748), .C1(n7483), 
        .C2(P2_U3152), .ZN(P2_U3346) );
  INV_X1 U8370 ( .A(n7065), .ZN(n6855) );
  OAI222_X1 U8371 ( .A1(n9524), .A2(n6749), .B1(n9527), .B2(n6748), .C1(
        P1_U3084), .C2(n6855), .ZN(P1_U3341) );
  OAI21_X1 U8372 ( .B1(n9832), .B2(n6750), .A(n6877), .ZN(n6752) );
  NAND2_X1 U8373 ( .A1(n9832), .A2(n7594), .ZN(n6751) );
  NAND2_X1 U8374 ( .A1(n6752), .A2(n6751), .ZN(n8527) );
  INV_X1 U8375 ( .A(n8527), .ZN(n9785) );
  NOR2_X1 U8376 ( .A1(n9785), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8377 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6761) );
  AND2_X1 U8378 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9619) );
  INV_X1 U8379 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9611) );
  OAI22_X1 U8380 ( .A1(n9620), .A2(n9619), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n9611), .ZN(n6755) );
  OAI21_X1 U8381 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n9620), .A(n6753), .ZN(
        n6754) );
  NAND2_X1 U8382 ( .A1(n6754), .A2(n4431), .ZN(n9623) );
  OAI211_X1 U8383 ( .C1(n9624), .C2(n6755), .A(n9623), .B(P1_STATE_REG_SCAN_IN), .ZN(n6756) );
  NOR2_X1 U8384 ( .A1(n6757), .A2(n6756), .ZN(n6759) );
  AND3_X1 U8385 ( .A1(n9712), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9611), .ZN(n6758) );
  AOI211_X1 U8386 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n6759), .B(
        n6758), .ZN(n6760) );
  OAI21_X1 U8387 ( .B1(n9112), .B2(n6761), .A(n6760), .ZN(P1_U3241) );
  NAND2_X1 U8388 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n8493), .ZN(n6762) );
  OAI21_X1 U8389 ( .B1(n8749), .B2(n8493), .A(n6762), .ZN(P2_U3569) );
  NAND2_X1 U8390 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n8493), .ZN(n6763) );
  OAI21_X1 U8391 ( .B1(n8551), .B2(n8493), .A(n6763), .ZN(P2_U3572) );
  NAND2_X1 U8392 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n8493), .ZN(n6764) );
  OAI21_X1 U8393 ( .B1(n8577), .B2(n8493), .A(n6764), .ZN(P2_U3582) );
  INV_X1 U8394 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6777) );
  NOR2_X1 U8395 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6765), .ZN(n7431) );
  INV_X1 U8396 ( .A(n9712), .ZN(n9648) );
  AOI21_X1 U8397 ( .B1(n6768), .B2(n6767), .A(n6766), .ZN(n6769) );
  NOR2_X1 U8398 ( .A1(n9648), .A2(n6769), .ZN(n6770) );
  AOI211_X1 U8399 ( .C1(n9704), .C2(n6771), .A(n7431), .B(n6770), .ZN(n6776)
         );
  OAI211_X1 U8400 ( .C1(n6774), .C2(n6773), .A(n9702), .B(n6772), .ZN(n6775)
         );
  OAI211_X1 U8401 ( .C1(n6777), .C2(n9112), .A(n6776), .B(n6775), .ZN(P1_U3247) );
  AOI21_X1 U8402 ( .B1(n6780), .B2(n6779), .A(n6778), .ZN(n6789) );
  AND2_X1 U8403 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7349) );
  AOI21_X1 U8404 ( .B1(n6783), .B2(n6782), .A(n6781), .ZN(n6784) );
  NOR2_X1 U8405 ( .A1(n9648), .A2(n6784), .ZN(n6785) );
  AOI211_X1 U8406 ( .C1(n9704), .C2(n6786), .A(n7349), .B(n6785), .ZN(n6788)
         );
  INV_X1 U8407 ( .A(n9112), .ZN(n9711) );
  NAND2_X1 U8408 ( .A1(n9711), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6787) );
  OAI211_X1 U8409 ( .C1(n6789), .C2(n9688), .A(n6788), .B(n6787), .ZN(P1_U3248) );
  INV_X1 U8410 ( .A(n6790), .ZN(n6793) );
  INV_X1 U8411 ( .A(n7283), .ZN(n7063) );
  OAI222_X1 U8412 ( .A1(n9522), .A2(n6793), .B1(n7063), .B2(P1_U3084), .C1(
        n6791), .C2(n9524), .ZN(P1_U3340) );
  INV_X1 U8413 ( .A(n7812), .ZN(n7805) );
  OAI222_X1 U8414 ( .A1(P2_U3152), .A2(n7805), .B1(n8920), .B2(n6793), .C1(
        n6792), .C2(n8259), .ZN(P2_U3345) );
  INV_X1 U8415 ( .A(n6794), .ZN(n6796) );
  INV_X1 U8416 ( .A(n7624), .ZN(n7617) );
  OAI222_X1 U8417 ( .A1(n9522), .A2(n6796), .B1(n7617), .B2(P1_U3084), .C1(
        n6795), .C2(n9524), .ZN(P1_U3339) );
  INV_X1 U8418 ( .A(n7891), .ZN(n7807) );
  OAI222_X1 U8419 ( .A1(n8259), .A2(n6797), .B1(n8920), .B2(n6796), .C1(
        P2_U3152), .C2(n7807), .ZN(P2_U3344) );
  INV_X1 U8420 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U8421 ( .A1(n6798), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6801) );
  OR2_X1 U8422 ( .A1(n6026), .A2(n6799), .ZN(n6800) );
  OAI211_X1 U8423 ( .C1(n6025), .C2(n6802), .A(n6801), .B(n6800), .ZN(n9113)
         );
  NAND2_X1 U8424 ( .A1(n9113), .A2(P1_U4006), .ZN(n6803) );
  OAI21_X1 U8425 ( .B1(P1_U4006), .B2(n5644), .A(n6803), .ZN(P1_U3586) );
  OAI21_X1 U8426 ( .B1(n6806), .B2(n6805), .A(n6804), .ZN(n9621) );
  INV_X1 U8427 ( .A(n9621), .ZN(n6813) );
  INV_X1 U8428 ( .A(n6834), .ZN(n6807) );
  AND2_X1 U8429 ( .A1(n6808), .A2(n6807), .ZN(n6809) );
  NAND2_X1 U8430 ( .A1(n6810), .A2(n6809), .ZN(n7000) );
  OAI22_X1 U8431 ( .A1(n9027), .A2(n6841), .B1(n6838), .B2(n9036), .ZN(n6811)
         );
  AOI21_X1 U8432 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7000), .A(n6811), .ZN(
        n6812) );
  OAI21_X1 U8433 ( .B1(n6813), .B2(n4371), .A(n6812), .ZN(P1_U3230) );
  XNOR2_X1 U8434 ( .A(n6815), .B(n6814), .ZN(n6817) );
  XNOR2_X1 U8435 ( .A(n6817), .B(n6816), .ZN(n6822) );
  NAND2_X1 U8436 ( .A1(n9487), .A2(n9730), .ZN(n9752) );
  AOI22_X1 U8437 ( .A1(n9021), .A2(n6818), .B1(n9033), .B2(n9719), .ZN(n6819)
         );
  OAI21_X1 U8438 ( .B1(n7000), .B2(n9752), .A(n6819), .ZN(n6820) );
  AOI21_X1 U8439 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n7000), .A(n6820), .ZN(
        n6821) );
  OAI21_X1 U8440 ( .B1(n6822), .B2(n4371), .A(n6821), .ZN(P1_U3220) );
  INV_X1 U8441 ( .A(n6823), .ZN(n6868) );
  AOI22_X1 U8442 ( .A1(n8503), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8918), .ZN(n6824) );
  OAI21_X1 U8443 ( .B1(n6868), .B2(n8920), .A(n6824), .ZN(P2_U3342) );
  NAND2_X1 U8444 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8493), .ZN(n6825) );
  OAI21_X1 U8445 ( .B1(n8587), .B2(n8493), .A(n6825), .ZN(P2_U3581) );
  NAND2_X1 U8446 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n8493), .ZN(n6826) );
  OAI21_X1 U8447 ( .B1(n8563), .B2(n8493), .A(n6826), .ZN(P2_U3578) );
  INV_X1 U8448 ( .A(n6827), .ZN(n6830) );
  OAI222_X1 U8449 ( .A1(n9524), .A2(n6828), .B1(n9527), .B2(n6830), .C1(
        P1_U3084), .C2(n9071), .ZN(P1_U3338) );
  INV_X1 U8450 ( .A(n7911), .ZN(n7921) );
  OAI222_X1 U8451 ( .A1(n7921), .A2(P2_U3152), .B1(n8920), .B2(n6830), .C1(
        n6829), .C2(n8259), .ZN(P2_U3343) );
  OR2_X1 U8452 ( .A1(n9767), .A2(n9204), .ZN(n6832) );
  NOR2_X1 U8453 ( .A1(n6834), .A2(n6833), .ZN(n6835) );
  INV_X1 U8454 ( .A(n9716), .ZN(n6836) );
  NAND2_X1 U8455 ( .A1(n9719), .A2(n6841), .ZN(n7988) );
  NAND2_X1 U8456 ( .A1(n6836), .A2(n7988), .ZN(n8023) );
  NAND3_X1 U8457 ( .A1(n8023), .A2(n8178), .A3(n6840), .ZN(n6837) );
  OAI21_X1 U8458 ( .B1(n6838), .B2(n9328), .A(n6837), .ZN(n7093) );
  INV_X1 U8459 ( .A(n7093), .ZN(n6839) );
  OAI21_X1 U8460 ( .B1(n6841), .B2(n6840), .A(n6839), .ZN(n6845) );
  NAND2_X1 U8461 ( .A1(n6845), .A2(n9782), .ZN(n6842) );
  OAI21_X1 U8462 ( .B1(n9782), .B2(n9611), .A(n6842), .ZN(P1_U3523) );
  INV_X1 U8463 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6847) );
  NAND2_X1 U8464 ( .A1(n6845), .A2(n9774), .ZN(n6846) );
  OAI21_X1 U8465 ( .B1(n9774), .B2(n6847), .A(n6846), .ZN(P1_U3454) );
  AOI22_X1 U8466 ( .A1(n6860), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n6848), .B2(
        n9054), .ZN(n9059) );
  INV_X1 U8467 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9568) );
  AOI22_X1 U8468 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n9695), .B1(n6849), .B2(
        n9568), .ZN(n9687) );
  OAI21_X1 U8469 ( .B1(n6858), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6850), .ZN(
        n9686) );
  NAND2_X1 U8470 ( .A1(n9687), .A2(n9686), .ZN(n9685) );
  OAI21_X1 U8471 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9695), .A(n9685), .ZN(
        n9058) );
  NAND2_X1 U8472 ( .A1(n9059), .A2(n9058), .ZN(n9057) );
  OAI21_X1 U8473 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6860), .A(n9057), .ZN(
        n6853) );
  INV_X1 U8474 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6851) );
  MUX2_X1 U8475 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6851), .S(n7065), .Z(n6852)
         );
  NAND2_X1 U8476 ( .A1(n6852), .A2(n6853), .ZN(n7058) );
  OAI21_X1 U8477 ( .B1(n6853), .B2(n6852), .A(n7058), .ZN(n6866) );
  NAND2_X1 U8478 ( .A1(n9711), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6854) );
  NAND2_X1 U8479 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7840) );
  OAI211_X1 U8480 ( .C1(n9641), .C2(n6855), .A(n6854), .B(n7840), .ZN(n6865)
         );
  NOR2_X1 U8481 ( .A1(n6860), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6856) );
  AOI21_X1 U8482 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6860), .A(n6856), .ZN(
        n9052) );
  NAND2_X1 U8483 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n9695), .ZN(n6859) );
  OAI21_X1 U8484 ( .B1(n9695), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6859), .ZN(
        n9690) );
  NAND2_X1 U8485 ( .A1(n9052), .A2(n4318), .ZN(n9051) );
  OAI21_X1 U8486 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6860), .A(n9051), .ZN(
        n6863) );
  NAND2_X1 U8487 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7065), .ZN(n6861) );
  OAI21_X1 U8488 ( .B1(n7065), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6861), .ZN(
        n6862) );
  NOR2_X1 U8489 ( .A1(n6862), .A2(n6863), .ZN(n7064) );
  AOI211_X1 U8490 ( .C1(n6863), .C2(n6862), .A(n7064), .B(n9688), .ZN(n6864)
         );
  AOI211_X1 U8491 ( .C1(n9712), .C2(n6866), .A(n6865), .B(n6864), .ZN(n6867)
         );
  INV_X1 U8492 ( .A(n6867), .ZN(P1_U3253) );
  INV_X1 U8493 ( .A(n9089), .ZN(n9078) );
  OAI222_X1 U8494 ( .A1(n9524), .A2(n6869), .B1(n9078), .B2(P1_U3084), .C1(
        n9522), .C2(n6868), .ZN(P1_U3337) );
  INV_X1 U8495 ( .A(n6870), .ZN(n6871) );
  NAND2_X1 U8496 ( .A1(n6871), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6872) );
  OAI211_X1 U8497 ( .C1(n9832), .C2(n6873), .A(n7594), .B(n6872), .ZN(n6879)
         );
  NAND2_X1 U8498 ( .A1(n6879), .A2(n6877), .ZN(n6874) );
  NAND2_X1 U8499 ( .A1(n6874), .A2(n8493), .ZN(n6893) );
  NOR2_X1 U8500 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5100), .ZN(n7116) );
  INV_X1 U8501 ( .A(n6965), .ZN(n6887) );
  INV_X1 U8502 ( .A(n6991), .ZN(n6886) );
  INV_X1 U8503 ( .A(n6978), .ZN(n6885) );
  NAND2_X1 U8504 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6968) );
  NOR2_X1 U8505 ( .A1(n6967), .A2(n6968), .ZN(n6966) );
  AOI21_X1 U8506 ( .B1(n6885), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6966), .ZN(
        n6982) );
  XOR2_X1 U8507 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6991), .Z(n6981) );
  NOR2_X1 U8508 ( .A1(n6982), .A2(n6981), .ZN(n6980) );
  AOI21_X1 U8509 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n6886), .A(n6980), .ZN(
        n6955) );
  XOR2_X1 U8510 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6965), .Z(n6954) );
  NOR2_X1 U8511 ( .A1(n6955), .A2(n6954), .ZN(n6953) );
  NAND2_X1 U8512 ( .A1(n6888), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6875) );
  OAI21_X1 U8513 ( .B1(n6888), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6875), .ZN(
        n6941) );
  NAND2_X1 U8514 ( .A1(n6905), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6876) );
  OAI21_X1 U8515 ( .B1(n6905), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6876), .ZN(
        n6880) );
  AND2_X1 U8516 ( .A1(n6877), .A2(n5832), .ZN(n6878) );
  AOI211_X1 U8517 ( .C1(n6881), .C2(n6880), .A(n6899), .B(n9787), .ZN(n6882)
         );
  AOI211_X1 U8518 ( .C1(n9785), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7116), .B(
        n6882), .ZN(n6897) );
  NAND2_X1 U8519 ( .A1(n6888), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6890) );
  INV_X1 U8520 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7268) );
  MUX2_X1 U8521 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7268), .S(n6978), .Z(n6884)
         );
  INV_X1 U8522 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6883) );
  INV_X1 U8523 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6971) );
  AOI21_X1 U8524 ( .B1(n6885), .B2(P2_REG2_REG_1__SCAN_IN), .A(n6972), .ZN(
        n6986) );
  MUX2_X1 U8525 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n7613), .S(n6991), .Z(n6985)
         );
  OR2_X1 U8526 ( .A1(n6986), .A2(n6985), .ZN(n6988) );
  NAND2_X1 U8527 ( .A1(n6886), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6960) );
  INV_X1 U8528 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7484) );
  MUX2_X1 U8529 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7484), .S(n6965), .Z(n6959)
         );
  AOI21_X1 U8530 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n6887), .A(n6958), .ZN(
        n6945) );
  INV_X1 U8531 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7519) );
  MUX2_X1 U8532 ( .A(n7519), .B(P2_REG2_REG_4__SCAN_IN), .S(n6888), .Z(n6946)
         );
  NAND2_X1 U8533 ( .A1(n6890), .A2(n6889), .ZN(n6895) );
  INV_X1 U8534 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6891) );
  MUX2_X1 U8535 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6891), .S(n6905), .Z(n6894)
         );
  NOR2_X1 U8536 ( .A1(n5576), .A2(n5832), .ZN(n6892) );
  NAND2_X1 U8537 ( .A1(n6894), .A2(n6895), .ZN(n6906) );
  OAI211_X1 U8538 ( .C1(n6895), .C2(n6894), .A(n9784), .B(n6906), .ZN(n6896)
         );
  OAI211_X1 U8539 ( .C1(n9786), .C2(n6898), .A(n6897), .B(n6896), .ZN(P2_U3250) );
  NOR2_X1 U8540 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7236), .ZN(n6904) );
  AOI21_X1 U8541 ( .B1(n6905), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6899), .ZN(
        n6902) );
  NAND2_X1 U8542 ( .A1(n6921), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6900) );
  OAI21_X1 U8543 ( .B1(n6921), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6900), .ZN(
        n6901) );
  NOR2_X1 U8544 ( .A1(n6902), .A2(n6901), .ZN(n6915) );
  AOI211_X1 U8545 ( .C1(n6902), .C2(n6901), .A(n6915), .B(n9787), .ZN(n6903)
         );
  AOI211_X1 U8546 ( .C1(n9785), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6904), .B(
        n6903), .ZN(n6912) );
  NAND2_X1 U8547 ( .A1(n6905), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U8548 ( .A1(n6907), .A2(n6906), .ZN(n6910) );
  INV_X1 U8549 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6908) );
  MUX2_X1 U8550 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6908), .S(n6921), .Z(n6909)
         );
  NAND2_X1 U8551 ( .A1(n6909), .A2(n6910), .ZN(n6922) );
  OAI211_X1 U8552 ( .C1(n6910), .C2(n6909), .A(n9784), .B(n6922), .ZN(n6911)
         );
  OAI211_X1 U8553 ( .C1(n9786), .C2(n6913), .A(n6912), .B(n6911), .ZN(P2_U3251) );
  NOR2_X1 U8554 ( .A1(n6914), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7368) );
  MUX2_X1 U8555 ( .A(n9959), .B(P2_REG1_REG_7__SCAN_IN), .S(n6920), .Z(n6931)
         );
  INV_X1 U8556 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6916) );
  MUX2_X1 U8557 ( .A(n6916), .B(P2_REG1_REG_8__SCAN_IN), .S(n7030), .Z(n6917)
         );
  AOI211_X1 U8558 ( .C1(n6918), .C2(n6917), .A(n7029), .B(n9787), .ZN(n6919)
         );
  AOI211_X1 U8559 ( .C1(n9785), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7368), .B(
        n6919), .ZN(n6929) );
  INV_X1 U8560 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6924) );
  MUX2_X1 U8561 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6924), .S(n6920), .Z(n6935)
         );
  NAND2_X1 U8562 ( .A1(n6921), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8563 ( .A1(n6923), .A2(n6922), .ZN(n6936) );
  INV_X1 U8564 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6925) );
  MUX2_X1 U8565 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6925), .S(n7030), .Z(n6926)
         );
  NAND2_X1 U8566 ( .A1(n6926), .A2(n6927), .ZN(n7038) );
  OAI211_X1 U8567 ( .C1(n6927), .C2(n6926), .A(n9784), .B(n7038), .ZN(n6928)
         );
  OAI211_X1 U8568 ( .C1(n9786), .C2(n7039), .A(n6929), .B(n6928), .ZN(P2_U3253) );
  AND2_X1 U8569 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7248) );
  AOI211_X1 U8570 ( .C1(n6932), .C2(n6931), .A(n6930), .B(n9787), .ZN(n6933)
         );
  AOI211_X1 U8571 ( .C1(n9785), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7248), .B(
        n6933), .ZN(n6938) );
  OAI211_X1 U8572 ( .C1(n6936), .C2(n6935), .A(n9784), .B(n6934), .ZN(n6937)
         );
  OAI211_X1 U8573 ( .C1(n9786), .C2(n6939), .A(n6938), .B(n6937), .ZN(P2_U3252) );
  AND2_X1 U8574 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6944) );
  AOI211_X1 U8575 ( .C1(n6942), .C2(n6941), .A(n6940), .B(n9787), .ZN(n6943)
         );
  AOI211_X1 U8576 ( .C1(n9785), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6944), .B(
        n6943), .ZN(n6949) );
  XOR2_X1 U8577 ( .A(n6946), .B(n6945), .Z(n6947) );
  NAND2_X1 U8578 ( .A1(n9784), .A2(n6947), .ZN(n6948) );
  OAI211_X1 U8579 ( .C1(n9786), .C2(n6950), .A(n6949), .B(n6948), .ZN(P2_U3249) );
  INV_X1 U8580 ( .A(n6951), .ZN(n6992) );
  AOI22_X1 U8581 ( .A1(n9104), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9520), .ZN(n6952) );
  OAI21_X1 U8582 ( .B1(n6992), .B2(n9522), .A(n6952), .ZN(P1_U3336) );
  AND2_X1 U8583 ( .A1(P2_U3152), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6957) );
  AOI211_X1 U8584 ( .C1(n6955), .C2(n6954), .A(n6953), .B(n9787), .ZN(n6956)
         );
  AOI211_X1 U8585 ( .C1(n9785), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6957), .B(
        n6956), .ZN(n6964) );
  INV_X1 U8586 ( .A(n6958), .ZN(n6962) );
  NAND3_X1 U8587 ( .A1(n6988), .A2(n6960), .A3(n6959), .ZN(n6961) );
  NAND3_X1 U8588 ( .A1(n9784), .A2(n6962), .A3(n6961), .ZN(n6963) );
  OAI211_X1 U8589 ( .C1(n9786), .C2(n6965), .A(n6964), .B(n6963), .ZN(P2_U3248) );
  AND2_X1 U8590 ( .A1(P2_U3152), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6970) );
  AOI211_X1 U8591 ( .C1(n6968), .C2(n6967), .A(n6966), .B(n9787), .ZN(n6969)
         );
  AOI211_X1 U8592 ( .C1(n9785), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6970), .B(
        n6969), .ZN(n6977) );
  NOR2_X1 U8593 ( .A1(n6971), .A2(n6883), .ZN(n6975) );
  MUX2_X1 U8594 ( .A(n7268), .B(P2_REG2_REG_1__SCAN_IN), .S(n6978), .Z(n6974)
         );
  INV_X1 U8595 ( .A(n6972), .ZN(n6973) );
  OAI211_X1 U8596 ( .C1(n6975), .C2(n6974), .A(n9784), .B(n6973), .ZN(n6976)
         );
  OAI211_X1 U8597 ( .C1(n9786), .C2(n6978), .A(n6977), .B(n6976), .ZN(P2_U3246) );
  INV_X1 U8598 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6979) );
  NOR2_X1 U8599 ( .A1(n8527), .A2(n6979), .ZN(n6984) );
  AOI211_X1 U8600 ( .C1(n6982), .C2(n6981), .A(n6980), .B(n9787), .ZN(n6983)
         );
  AOI211_X1 U8601 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(P2_U3152), .A(n6984), .B(
        n6983), .ZN(n6990) );
  NAND2_X1 U8602 ( .A1(n6986), .A2(n6985), .ZN(n6987) );
  NAND3_X1 U8603 ( .A1(n9784), .A2(n6988), .A3(n6987), .ZN(n6989) );
  OAI211_X1 U8604 ( .C1(n9786), .C2(n6991), .A(n6990), .B(n6989), .ZN(P2_U3247) );
  INV_X1 U8605 ( .A(n7924), .ZN(n8518) );
  OAI222_X1 U8606 ( .A1(n8259), .A2(n6993), .B1(n8920), .B2(n6992), .C1(
        P2_U3152), .C2(n8518), .ZN(P2_U3341) );
  INV_X1 U8607 ( .A(n6994), .ZN(n6995) );
  AOI21_X1 U8608 ( .B1(n6997), .B2(n6996), .A(n6995), .ZN(n7002) );
  AOI22_X1 U8609 ( .A1(n9021), .A2(n9050), .B1(n9033), .B2(n6544), .ZN(n6998)
         );
  OAI21_X1 U8610 ( .B1(n9755), .B2(n9027), .A(n6998), .ZN(n6999) );
  AOI21_X1 U8611 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7000), .A(n6999), .ZN(
        n7001) );
  OAI21_X1 U8612 ( .B1(n7002), .B2(n4371), .A(n7001), .ZN(P1_U3235) );
  NAND3_X1 U8613 ( .A1(n7076), .A2(P2_STATE_REG_SCAN_IN), .A3(n7003), .ZN(
        n7004) );
  NOR2_X1 U8614 ( .A1(n7259), .A2(n7004), .ZN(n7005) );
  INV_X1 U8615 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7023) );
  XNOR2_X1 U8616 ( .A(n5565), .B(n7262), .ZN(n7006) );
  NAND2_X1 U8617 ( .A1(n7006), .A2(n7139), .ZN(n9799) );
  NAND2_X1 U8618 ( .A1(n5562), .A2(n9823), .ZN(n7007) );
  OR2_X1 U8619 ( .A1(n5565), .A2(n7007), .ZN(n9931) );
  OAI22_X1 U8620 ( .A1(n7610), .A2(n7010), .B1(n4267), .B2(n8491), .ZN(n7011)
         );
  NAND2_X1 U8621 ( .A1(n7271), .A2(n4266), .ZN(n9890) );
  NAND2_X1 U8622 ( .A1(n9890), .A2(n8301), .ZN(n7012) );
  NAND2_X1 U8623 ( .A1(n7012), .A2(n9905), .ZN(n7013) );
  OR2_X1 U8624 ( .A1(n7050), .A2(n7013), .ZN(n7485) );
  OAI21_X1 U8625 ( .B1(n7492), .B2(n9941), .A(n7485), .ZN(n7021) );
  XNOR2_X1 U8626 ( .A(n7015), .B(n7014), .ZN(n7020) );
  OR2_X1 U8627 ( .A1(n7224), .A2(n8765), .ZN(n7018) );
  OAI21_X1 U8628 ( .B1(n4835), .B2(n8277), .A(n7018), .ZN(n8302) );
  INV_X1 U8629 ( .A(n8302), .ZN(n7019) );
  OAI21_X1 U8630 ( .B1(n7020), .B2(n9570), .A(n7019), .ZN(n7488) );
  AOI211_X1 U8631 ( .C1(n9947), .C2(n7489), .A(n7021), .B(n7488), .ZN(n7026)
         );
  OR2_X1 U8632 ( .A1(n7026), .A2(n9949), .ZN(n7022) );
  OAI21_X1 U8633 ( .B1(n9951), .B2(n7023), .A(n7022), .ZN(P2_U3460) );
  INV_X1 U8634 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7028) );
  OR2_X1 U8635 ( .A1(n7026), .A2(n9965), .ZN(n7027) );
  OAI21_X1 U8636 ( .B1(n9967), .B2(n7028), .A(n7027), .ZN(P2_U3523) );
  NAND2_X1 U8637 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7688) );
  INV_X1 U8638 ( .A(n7688), .ZN(n7035) );
  AOI21_X1 U8639 ( .B1(n7030), .B2(P2_REG1_REG_8__SCAN_IN), .A(n7029), .ZN(
        n7033) );
  INV_X1 U8640 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7031) );
  MUX2_X1 U8641 ( .A(n7031), .B(P2_REG1_REG_9__SCAN_IN), .S(n7128), .Z(n7032)
         );
  NOR2_X1 U8642 ( .A1(n7033), .A2(n7032), .ZN(n7122) );
  AOI211_X1 U8643 ( .C1(n7033), .C2(n7032), .A(n7122), .B(n9787), .ZN(n7034)
         );
  AOI211_X1 U8644 ( .C1(n9785), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7035), .B(
        n7034), .ZN(n7043) );
  INV_X1 U8645 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7036) );
  MUX2_X1 U8646 ( .A(n7036), .B(P2_REG2_REG_9__SCAN_IN), .S(n7128), .Z(n7037)
         );
  INV_X1 U8647 ( .A(n7037), .ZN(n7041) );
  NAND2_X1 U8648 ( .A1(n7041), .A2(n7040), .ZN(n7129) );
  OAI211_X1 U8649 ( .C1(n7041), .C2(n7040), .A(n9784), .B(n7129), .ZN(n7042)
         );
  OAI211_X1 U8650 ( .C1(n9786), .C2(n7044), .A(n7043), .B(n7042), .ZN(P2_U3254) );
  NAND2_X1 U8651 ( .A1(n7607), .A2(n7492), .ZN(n7045) );
  NAND2_X1 U8652 ( .A1(n7293), .A2(n7291), .ZN(n7216) );
  OAI21_X1 U8653 ( .B1(n7293), .B2(n7291), .A(n7216), .ZN(n7517) );
  AOI21_X1 U8654 ( .B1(n7046), .B2(n7291), .A(n9570), .ZN(n7049) );
  OR2_X1 U8655 ( .A1(n7607), .A2(n8277), .ZN(n7048) );
  NAND2_X1 U8656 ( .A1(n8488), .A2(n8801), .ZN(n7047) );
  NAND2_X1 U8657 ( .A1(n7048), .A2(n7047), .ZN(n8385) );
  AOI21_X1 U8658 ( .B1(n7049), .B2(n4826), .A(n8385), .ZN(n7525) );
  NAND2_X1 U8659 ( .A1(n7050), .A2(n7215), .ZN(n7218) );
  OAI211_X1 U8660 ( .C1(n7050), .C2(n7215), .A(n9905), .B(n7218), .ZN(n7518)
         );
  OAI211_X1 U8661 ( .C1(n7215), .C2(n9941), .A(n7525), .B(n7518), .ZN(n7051)
         );
  AOI21_X1 U8662 ( .B1(n9947), .B2(n7517), .A(n7051), .ZN(n7056) );
  OR2_X1 U8663 ( .A1(n9951), .A2(n7052), .ZN(n7053) );
  OAI21_X1 U8664 ( .B1(n7056), .B2(n9949), .A(n7053), .ZN(P2_U3463) );
  INV_X1 U8665 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7054) );
  OR2_X1 U8666 ( .A1(n9967), .A2(n7054), .ZN(n7055) );
  OAI21_X1 U8667 ( .B1(n7056), .B2(n9965), .A(n7055), .ZN(P2_U3524) );
  NAND2_X1 U8668 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7877) );
  INV_X1 U8669 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7057) );
  MUX2_X1 U8670 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7057), .S(n7283), .Z(n7060)
         );
  OAI21_X1 U8671 ( .B1(n7065), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7058), .ZN(
        n7059) );
  NAND2_X1 U8672 ( .A1(n7060), .A2(n7059), .ZN(n7276) );
  OAI21_X1 U8673 ( .B1(n7060), .B2(n7059), .A(n7276), .ZN(n7061) );
  NAND2_X1 U8674 ( .A1(n9712), .A2(n7061), .ZN(n7062) );
  OAI211_X1 U8675 ( .C1(n9641), .C2(n7063), .A(n7877), .B(n7062), .ZN(n7071)
         );
  INV_X1 U8676 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7066) );
  MUX2_X1 U8677 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n7066), .S(n7283), .Z(n7067)
         );
  INV_X1 U8678 ( .A(n7067), .ZN(n7068) );
  AOI211_X1 U8679 ( .C1(n7069), .C2(n7068), .A(n7282), .B(n9688), .ZN(n7070)
         );
  AOI211_X1 U8680 ( .C1(P1_ADDR_REG_13__SCAN_IN), .C2(n9711), .A(n7071), .B(
        n7070), .ZN(n7072) );
  INV_X1 U8681 ( .A(n7072), .ZN(P1_U3254) );
  INV_X1 U8682 ( .A(n8466), .ZN(n8251) );
  INV_X1 U8683 ( .A(n8465), .ZN(n7718) );
  AOI22_X1 U8684 ( .A1(n8251), .A2(n8491), .B1(n7718), .B2(n9872), .ZN(n7080)
         );
  OAI21_X1 U8685 ( .B1(n7075), .B2(n7074), .A(n7073), .ZN(n7078) );
  AND2_X1 U8686 ( .A1(n7076), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7257) );
  NAND2_X1 U8687 ( .A1(n7077), .A2(n7257), .ZN(n8256) );
  AOI22_X1 U8688 ( .A1(n8460), .A2(n7078), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8256), .ZN(n7079) );
  OAI211_X1 U8689 ( .C1(n9885), .C2(n8458), .A(n7080), .B(n7079), .ZN(P2_U3224) );
  INV_X1 U8690 ( .A(n7081), .ZN(n7097) );
  AOI22_X1 U8691 ( .A1(n8530), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8918), .ZN(n7082) );
  OAI21_X1 U8692 ( .B1(n7097), .B2(n8920), .A(n7082), .ZN(P2_U3340) );
  OAI21_X1 U8693 ( .B1(n7085), .B2(n7084), .A(n7083), .ZN(n7086) );
  NAND2_X1 U8694 ( .A1(n7086), .A2(n9018), .ZN(n7092) );
  NAND2_X1 U8695 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9538) );
  INV_X1 U8696 ( .A(n9538), .ZN(n7087) );
  AOI21_X1 U8697 ( .B1(n9033), .B2(n6818), .A(n7087), .ZN(n7089) );
  OR2_X1 U8698 ( .A1(n9036), .A2(n7145), .ZN(n7088) );
  OAI211_X1 U8699 ( .C1(n9027), .C2(n7209), .A(n7089), .B(n7088), .ZN(n7090)
         );
  INV_X1 U8700 ( .A(n7090), .ZN(n7091) );
  OAI211_X1 U8701 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9000), .A(n7092), .B(
        n7091), .ZN(P1_U3216) );
  INV_X2 U8702 ( .A(n9142), .ZN(n9728) );
  AOI21_X1 U8703 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9728), .A(n7093), .ZN(
        n7096) );
  NAND2_X1 U8704 ( .A1(n9743), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7095) );
  OAI21_X1 U8705 ( .B1(n9551), .B2(n9346), .A(n9731), .ZN(n7094) );
  OAI211_X1 U8706 ( .C1(n7096), .C2(n9743), .A(n7095), .B(n7094), .ZN(P1_U3291) );
  INV_X1 U8707 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7098) );
  INV_X1 U8708 ( .A(n9703), .ZN(n9101) );
  OAI222_X1 U8709 ( .A1(n9524), .A2(n7098), .B1(n9527), .B2(n7097), .C1(
        P1_U3084), .C2(n9101), .ZN(P1_U3335) );
  INV_X1 U8710 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U8711 ( .A1(n7101), .A2(n9755), .ZN(n7099) );
  NAND2_X1 U8712 ( .A1(n7100), .A2(n7099), .ZN(n7146) );
  NAND2_X1 U8713 ( .A1(n7192), .A2(n7107), .ZN(n7995) );
  NAND2_X1 U8714 ( .A1(n9050), .A2(n7209), .ZN(n7992) );
  NAND2_X1 U8715 ( .A1(n7995), .A2(n7992), .ZN(n7157) );
  NAND2_X1 U8716 ( .A1(n7146), .A2(n7157), .ZN(n7144) );
  OAI21_X1 U8717 ( .B1(n7146), .B2(n7157), .A(n7144), .ZN(n7211) );
  INV_X1 U8718 ( .A(n7211), .ZN(n7109) );
  NAND2_X1 U8719 ( .A1(n6455), .A2(n9736), .ZN(n8158) );
  INV_X1 U8720 ( .A(n9720), .ZN(n9330) );
  OAI22_X1 U8721 ( .A1(n7101), .A2(n9330), .B1(n7145), .B2(n9328), .ZN(n7105)
         );
  XNOR2_X1 U8722 ( .A(n7158), .B(n7157), .ZN(n7103) );
  NOR2_X1 U8723 ( .A1(n7103), .A2(n9318), .ZN(n7104) );
  AOI211_X1 U8724 ( .C1(n9549), .C2(n7211), .A(n7105), .B(n7104), .ZN(n7213)
         );
  OR2_X1 U8725 ( .A1(n7106), .A2(n7107), .ZN(n7163) );
  INV_X1 U8726 ( .A(n7163), .ZN(n7197) );
  AOI21_X1 U8727 ( .B1(n7107), .B2(n7106), .A(n7197), .ZN(n7205) );
  AOI22_X1 U8728 ( .A1(n7205), .A2(n9554), .B1(n9487), .B2(n7107), .ZN(n7108)
         );
  OAI211_X1 U8729 ( .C1(n7109), .C2(n9491), .A(n7213), .B(n7108), .ZN(n7112)
         );
  NAND2_X1 U8730 ( .A1(n7112), .A2(n9782), .ZN(n7110) );
  OAI21_X1 U8731 ( .B1(n9782), .B2(n7111), .A(n7110), .ZN(P1_U3526) );
  NAND2_X1 U8732 ( .A1(n7112), .A2(n9774), .ZN(n7113) );
  OAI21_X1 U8733 ( .B1(n9774), .B2(n5980), .A(n7113), .ZN(P1_U3463) );
  XOR2_X1 U8734 ( .A(n7115), .B(n7114), .Z(n7120) );
  AOI22_X1 U8735 ( .A1(n8251), .A2(n8487), .B1(n9818), .B2(n8469), .ZN(n7118)
         );
  AOI21_X1 U8736 ( .B1(n8454), .B2(n9820), .A(n7116), .ZN(n7117) );
  OAI211_X1 U8737 ( .C1(n7224), .C2(n8465), .A(n7118), .B(n7117), .ZN(n7119)
         );
  AOI21_X1 U8738 ( .B1(n8460), .B2(n7120), .A(n7119), .ZN(n7121) );
  INV_X1 U8739 ( .A(n7121), .ZN(P2_U3229) );
  NAND2_X1 U8740 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7713) );
  INV_X1 U8741 ( .A(n7713), .ZN(n7127) );
  INV_X1 U8742 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7123) );
  MUX2_X1 U8743 ( .A(n7123), .B(P2_REG1_REG_10__SCAN_IN), .S(n7341), .Z(n7124)
         );
  AOI211_X1 U8744 ( .C1(n7125), .C2(n7124), .A(n7340), .B(n9787), .ZN(n7126)
         );
  AOI211_X1 U8745 ( .C1(n9785), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7127), .B(
        n7126), .ZN(n7135) );
  NAND2_X1 U8746 ( .A1(n7128), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7130) );
  NAND2_X1 U8747 ( .A1(n7130), .A2(n7129), .ZN(n7133) );
  INV_X1 U8748 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7131) );
  MUX2_X1 U8749 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7131), .S(n7341), .Z(n7132)
         );
  NAND2_X1 U8750 ( .A1(n7132), .A2(n7133), .ZN(n7334) );
  OAI211_X1 U8751 ( .C1(n7133), .C2(n7132), .A(n9784), .B(n7334), .ZN(n7134)
         );
  OAI211_X1 U8752 ( .C1(n9786), .C2(n7136), .A(n7135), .B(n7134), .ZN(P2_U3255) );
  INV_X1 U8753 ( .A(n7137), .ZN(n7140) );
  OAI222_X1 U8754 ( .A1(n7139), .A2(P2_U3152), .B1(n8920), .B2(n7140), .C1(
        n7138), .C2(n8259), .ZN(P2_U3339) );
  OAI222_X1 U8755 ( .A1(n9524), .A2(n7141), .B1(n9527), .B2(n7140), .C1(n9204), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  AND2_X1 U8756 ( .A1(n8178), .A2(n7142), .ZN(n7143) );
  NAND2_X1 U8757 ( .A1(n7192), .A2(n7209), .ZN(n7149) );
  NAND2_X1 U8758 ( .A1(n7144), .A2(n7149), .ZN(n7191) );
  NAND2_X1 U8759 ( .A1(n7145), .A2(n7199), .ZN(n7999) );
  NAND2_X1 U8760 ( .A1(n7997), .A2(n7999), .ZN(n7148) );
  NAND2_X1 U8761 ( .A1(n7191), .A2(n7148), .ZN(n7190) );
  NAND2_X1 U8762 ( .A1(n7145), .A2(n9760), .ZN(n7150) );
  AND2_X1 U8763 ( .A1(n7190), .A2(n7150), .ZN(n7156) );
  XNOR2_X1 U8764 ( .A(n9048), .B(n7376), .ZN(n7161) );
  AND2_X1 U8765 ( .A1(n7157), .A2(n7148), .ZN(n7147) );
  NAND2_X1 U8766 ( .A1(n7147), .A2(n7146), .ZN(n7155) );
  NOR2_X1 U8767 ( .A1(n7159), .A2(n7149), .ZN(n7153) );
  INV_X1 U8768 ( .A(n7161), .ZN(n7151) );
  NAND2_X1 U8769 ( .A1(n7151), .A2(n7150), .ZN(n7152) );
  NOR2_X1 U8770 ( .A1(n7153), .A2(n7152), .ZN(n7154) );
  NAND2_X1 U8771 ( .A1(n7155), .A2(n7154), .ZN(n7378) );
  OAI21_X1 U8772 ( .B1(n7156), .B2(n7151), .A(n7378), .ZN(n7173) );
  INV_X1 U8773 ( .A(n7157), .ZN(n8024) );
  XNOR2_X1 U8774 ( .A(n7161), .B(n7371), .ZN(n7162) );
  AOI222_X1 U8775 ( .A1(n9725), .A2(n7162), .B1(n4681), .B2(n9721), .C1(n9049), 
        .C2(n9720), .ZN(n7172) );
  MUX2_X1 U8776 ( .A(n6518), .B(n7172), .S(n9740), .Z(n7169) );
  INV_X1 U8777 ( .A(n7164), .ZN(n7196) );
  INV_X1 U8778 ( .A(n7376), .ZN(n7540) );
  AOI211_X1 U8779 ( .C1(n7376), .C2(n7196), .A(n9767), .B(n7440), .ZN(n7170)
         );
  NOR2_X1 U8780 ( .A1(n7165), .A2(n9736), .ZN(n9557) );
  INV_X1 U8781 ( .A(n7547), .ZN(n7166) );
  OAI22_X1 U8782 ( .A1(n9341), .A2(n7540), .B1(n9142), .B2(n7166), .ZN(n7167)
         );
  AOI21_X1 U8783 ( .B1(n7170), .B2(n9557), .A(n7167), .ZN(n7168) );
  OAI211_X1 U8784 ( .C1(n9365), .C2(n7173), .A(n7169), .B(n7168), .ZN(P1_U3286) );
  AOI21_X1 U8785 ( .B1(n9487), .B2(n7376), .A(n7170), .ZN(n7171) );
  OAI211_X1 U8786 ( .C1(n9562), .C2(n7173), .A(n7172), .B(n7171), .ZN(n7175)
         );
  NAND2_X1 U8787 ( .A1(n7175), .A2(n9782), .ZN(n7174) );
  OAI21_X1 U8788 ( .B1(n9782), .B2(n6525), .A(n7174), .ZN(P1_U3528) );
  INV_X1 U8789 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7177) );
  NAND2_X1 U8790 ( .A1(n7175), .A2(n9774), .ZN(n7176) );
  OAI21_X1 U8791 ( .B1(n9774), .B2(n7177), .A(n7176), .ZN(P1_U3469) );
  NAND2_X1 U8792 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9651) );
  INV_X1 U8793 ( .A(n9651), .ZN(n7178) );
  AOI21_X1 U8794 ( .B1(n9033), .B2(n9050), .A(n7178), .ZN(n7180) );
  INV_X1 U8795 ( .A(n9048), .ZN(n7433) );
  OR2_X1 U8796 ( .A1(n9036), .A2(n7433), .ZN(n7179) );
  OAI211_X1 U8797 ( .C1(n9027), .C2(n9760), .A(n7180), .B(n7179), .ZN(n7187)
         );
  NAND2_X1 U8798 ( .A1(n7083), .A2(n7181), .ZN(n7422) );
  INV_X1 U8799 ( .A(n7422), .ZN(n7185) );
  AOI21_X1 U8800 ( .B1(n7083), .B2(n7183), .A(n7182), .ZN(n7184) );
  NOR3_X1 U8801 ( .A1(n7185), .A2(n7184), .A3(n4371), .ZN(n7186) );
  AOI211_X1 U8802 ( .C1(n7198), .C2(n9031), .A(n7187), .B(n7186), .ZN(n7188)
         );
  INV_X1 U8803 ( .A(n7188), .ZN(P1_U3228) );
  XNOR2_X1 U8804 ( .A(n7189), .B(n7148), .ZN(n7195) );
  OAI21_X1 U8805 ( .B1(n7191), .B2(n7148), .A(n7190), .ZN(n9764) );
  OAI22_X1 U8806 ( .A1(n7433), .A2(n9328), .B1(n7192), .B2(n9330), .ZN(n7193)
         );
  AOI21_X1 U8807 ( .B1(n9764), .B2(n9549), .A(n7193), .ZN(n7194) );
  OAI21_X1 U8808 ( .B1(n9318), .B2(n7195), .A(n7194), .ZN(n9762) );
  INV_X1 U8809 ( .A(n9762), .ZN(n7204) );
  OAI21_X1 U8810 ( .B1(n9760), .B2(n7197), .A(n7196), .ZN(n9761) );
  AOI22_X1 U8811 ( .A1(n9743), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7198), .B2(
        n9728), .ZN(n7201) );
  NAND2_X1 U8812 ( .A1(n9551), .A2(n7199), .ZN(n7200) );
  OAI211_X1 U8813 ( .C1(n9761), .C2(n9384), .A(n7201), .B(n7200), .ZN(n7202)
         );
  AOI21_X1 U8814 ( .B1(n9764), .B2(n9558), .A(n7202), .ZN(n7203) );
  OAI21_X1 U8815 ( .B1(n7204), .B2(n9743), .A(n7203), .ZN(P1_U3287) );
  NAND2_X1 U8816 ( .A1(n7205), .A2(n9346), .ZN(n7208) );
  AOI22_X1 U8817 ( .A1(n9743), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9728), .B2(
        n7206), .ZN(n7207) );
  OAI211_X1 U8818 ( .C1(n7209), .C2(n9341), .A(n7208), .B(n7207), .ZN(n7210)
         );
  AOI21_X1 U8819 ( .B1(n9558), .B2(n7211), .A(n7210), .ZN(n7212) );
  OAI21_X1 U8820 ( .B1(n7213), .B2(n9743), .A(n7212), .ZN(P1_U3288) );
  INV_X1 U8821 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U8822 ( .A1(n7746), .A2(n7214), .ZN(n7222) );
  NAND2_X1 U8823 ( .A1(n7224), .A2(n7215), .ZN(n7297) );
  NAND2_X1 U8824 ( .A1(n7216), .A2(n7297), .ZN(n7217) );
  XOR2_X1 U8825 ( .A(n7222), .B(n7217), .Z(n9816) );
  AOI21_X1 U8826 ( .B1(n7218), .B2(n9818), .A(n9943), .ZN(n7219) );
  OR2_X1 U8827 ( .A1(n7218), .A2(n9818), .ZN(n7755) );
  AND2_X1 U8828 ( .A1(n7219), .A2(n7755), .ZN(n9817) );
  NAND2_X1 U8829 ( .A1(n4826), .A2(n7220), .ZN(n7221) );
  XOR2_X1 U8830 ( .A(n7222), .B(n7221), .Z(n7223) );
  OAI222_X1 U8831 ( .A1(n8765), .A2(n7319), .B1(n8277), .B2(n7224), .C1(n9570), 
        .C2(n7223), .ZN(n9825) );
  AOI211_X1 U8832 ( .C1(n9929), .C2(n9818), .A(n9817), .B(n9825), .ZN(n7225)
         );
  OAI21_X1 U8833 ( .B1(n9909), .B2(n9816), .A(n7225), .ZN(n7228) );
  NAND2_X1 U8834 ( .A1(n7228), .A2(n9951), .ZN(n7226) );
  OAI21_X1 U8835 ( .B1(n9951), .B2(n7227), .A(n7226), .ZN(P2_U3466) );
  INV_X1 U8836 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7230) );
  NAND2_X1 U8837 ( .A1(n7228), .A2(n9967), .ZN(n7229) );
  OAI21_X1 U8838 ( .B1(n9967), .B2(n7230), .A(n7229), .ZN(P2_U3525) );
  OAI21_X1 U8839 ( .B1(n7233), .B2(n7232), .A(n7231), .ZN(n7240) );
  OR2_X1 U8840 ( .A1(n7553), .A2(n8765), .ZN(n7235) );
  NAND2_X1 U8841 ( .A1(n8488), .A2(n8799), .ZN(n7234) );
  AND2_X1 U8842 ( .A1(n7235), .A2(n7234), .ZN(n7749) );
  OAI22_X1 U8843 ( .A1(n8452), .A2(n7749), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7236), .ZN(n7239) );
  INV_X1 U8844 ( .A(n7237), .ZN(n7758) );
  OAI22_X1 U8845 ( .A1(n8458), .A2(n9900), .B1(n8464), .B2(n7758), .ZN(n7238)
         );
  AOI211_X1 U8846 ( .C1(n7240), .C2(n8460), .A(n7239), .B(n7238), .ZN(n7241)
         );
  INV_X1 U8847 ( .A(n7241), .ZN(P2_U3241) );
  INV_X1 U8848 ( .A(n7242), .ZN(n7253) );
  OAI222_X1 U8849 ( .A1(n9527), .A2(n7253), .B1(P1_U3084), .B2(n7244), .C1(
        n7243), .C2(n9524), .ZN(P1_U3333) );
  XNOR2_X1 U8850 ( .A(n7246), .B(n7245), .ZN(n7251) );
  AOI22_X1 U8851 ( .A1(n8251), .A2(n8485), .B1(n9904), .B2(n8469), .ZN(n7250)
         );
  NOR2_X1 U8852 ( .A1(n8465), .A2(n7319), .ZN(n7247) );
  AOI211_X1 U8853 ( .C1(n8454), .C2(n7308), .A(n7248), .B(n7247), .ZN(n7249)
         );
  OAI211_X1 U8854 ( .C1(n7251), .C2(n8445), .A(n7250), .B(n7249), .ZN(P2_U3215) );
  OAI222_X1 U8855 ( .A1(P2_U3152), .A2(n5562), .B1(n8920), .B2(n7253), .C1(
        n7252), .C2(n8259), .ZN(P2_U3338) );
  XNOR2_X1 U8856 ( .A(n7009), .B(n7254), .ZN(n9881) );
  INV_X1 U8857 ( .A(n7255), .ZN(n7261) );
  NAND2_X1 U8858 ( .A1(n7257), .A2(n7256), .ZN(n7258) );
  NOR2_X1 U8859 ( .A1(n7259), .A2(n7258), .ZN(n7260) );
  NAND2_X1 U8860 ( .A1(n7261), .A2(n7260), .ZN(n7270) );
  INV_X1 U8861 ( .A(n7262), .ZN(n7263) );
  NAND2_X1 U8862 ( .A1(n7263), .A2(n9823), .ZN(n7577) );
  NAND2_X1 U8863 ( .A1(n9799), .A2(n7577), .ZN(n9828) );
  XNOR2_X1 U8864 ( .A(n7009), .B(n9877), .ZN(n7264) );
  NAND2_X1 U8865 ( .A1(n7264), .A2(n9803), .ZN(n7266) );
  AOI22_X1 U8866 ( .A1(n8491), .A2(n8801), .B1(n8799), .B2(n9872), .ZN(n7265)
         );
  NAND2_X1 U8867 ( .A1(n7266), .A2(n7265), .ZN(n9886) );
  INV_X1 U8868 ( .A(n8678), .ZN(n9821) );
  AOI22_X1 U8869 ( .A1(n9829), .A2(n9886), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9821), .ZN(n7267) );
  OAI21_X1 U8870 ( .B1(n7268), .B2(n9829), .A(n7267), .ZN(n7269) );
  AOI21_X1 U8871 ( .B1(n9805), .B2(n7272), .A(n7269), .ZN(n7274) );
  OR2_X1 U8872 ( .A1(n7270), .A2(n9823), .ZN(n8539) );
  INV_X1 U8873 ( .A(n7271), .ZN(n9883) );
  NAND2_X1 U8874 ( .A1(n7272), .A2(n9874), .ZN(n9882) );
  NAND3_X1 U8875 ( .A1(n8806), .A2(n9883), .A3(n9882), .ZN(n7273) );
  OAI211_X1 U8876 ( .C1(n9881), .C2(n8808), .A(n7274), .B(n7273), .ZN(P2_U3295) );
  INV_X1 U8877 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7289) );
  INV_X1 U8878 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7275) );
  MUX2_X1 U8879 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7275), .S(n7624), .Z(n7279)
         );
  OR2_X1 U8880 ( .A1(n7283), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7277) );
  NAND2_X1 U8881 ( .A1(n7277), .A2(n7276), .ZN(n7278) );
  NAND2_X1 U8882 ( .A1(n7279), .A2(n7278), .ZN(n7623) );
  OAI21_X1 U8883 ( .B1(n7279), .B2(n7278), .A(n7623), .ZN(n7280) );
  NAND2_X1 U8884 ( .A1(n9712), .A2(n7280), .ZN(n7281) );
  NAND2_X1 U8885 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U8886 ( .A1(n7281), .A2(n7858), .ZN(n7287) );
  INV_X1 U8887 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7284) );
  NOR2_X1 U8888 ( .A1(n7284), .A2(n7285), .ZN(n7619) );
  AOI211_X1 U8889 ( .C1(n7285), .C2(n7284), .A(n7619), .B(n9688), .ZN(n7286)
         );
  AOI211_X1 U8890 ( .C1(n9704), .C2(n7624), .A(n7287), .B(n7286), .ZN(n7288)
         );
  OAI21_X1 U8891 ( .B1(n9112), .B2(n7289), .A(n7288), .ZN(P1_U3255) );
  INV_X1 U8892 ( .A(n7316), .ZN(n7307) );
  INV_X1 U8893 ( .A(n4840), .ZN(n7294) );
  NAND2_X1 U8894 ( .A1(n7293), .A2(n7292), .ZN(n7301) );
  NAND2_X1 U8895 ( .A1(n7296), .A2(n7295), .ZN(n7298) );
  AND2_X1 U8896 ( .A1(n7298), .A2(n7297), .ZN(n7299) );
  OR2_X1 U8897 ( .A1(n4840), .A2(n7299), .ZN(n7300) );
  NAND2_X1 U8898 ( .A1(n7301), .A2(n7300), .ZN(n7752) );
  INV_X1 U8899 ( .A(n7752), .ZN(n7303) );
  NAND2_X1 U8900 ( .A1(n8487), .A2(n7754), .ZN(n7304) );
  INV_X1 U8901 ( .A(n7555), .ZN(n7305) );
  AOI21_X1 U8902 ( .B1(n7307), .B2(n7306), .A(n7305), .ZN(n9910) );
  INV_X1 U8903 ( .A(n8806), .ZN(n8683) );
  OR2_X1 U8904 ( .A1(n7755), .A2(n7754), .ZN(n7756) );
  AOI21_X1 U8905 ( .B1(n9904), .B2(n7756), .A(n9810), .ZN(n9906) );
  INV_X1 U8906 ( .A(n9906), .ZN(n7310) );
  INV_X1 U8907 ( .A(n7308), .ZN(n7309) );
  OAI22_X1 U8908 ( .A1(n8683), .A2(n7310), .B1(n7309), .B2(n8678), .ZN(n7311)
         );
  AOI21_X1 U8909 ( .B1(n9805), .B2(n9904), .A(n7311), .ZN(n7324) );
  NAND2_X1 U8910 ( .A1(n4826), .A2(n7312), .ZN(n7747) );
  NAND2_X1 U8911 ( .A1(n7747), .A2(n7313), .ZN(n7315) );
  AND2_X1 U8912 ( .A1(n7315), .A2(n7314), .ZN(n7317) );
  AOI21_X1 U8913 ( .B1(n7317), .B2(n7316), .A(n9570), .ZN(n7322) );
  OAI22_X1 U8914 ( .A1(n7319), .A2(n8277), .B1(n7318), .B2(n8765), .ZN(n7320)
         );
  AOI21_X1 U8915 ( .B1(n7322), .B2(n7321), .A(n7320), .ZN(n9908) );
  MUX2_X1 U8916 ( .A(n9908), .B(n6924), .S(n9831), .Z(n7323) );
  OAI211_X1 U8917 ( .C1(n9910), .C2(n8808), .A(n7324), .B(n7323), .ZN(P2_U3289) );
  NAND2_X1 U8918 ( .A1(n9877), .A2(n7325), .ZN(n7326) );
  INV_X1 U8919 ( .A(n7326), .ZN(n7331) );
  AOI22_X1 U8920 ( .A1(n7326), .A2(n9803), .B1(n8801), .B2(n8492), .ZN(n9871)
         );
  INV_X1 U8921 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7327) );
  OAI22_X1 U8922 ( .A1(n9831), .A2(n9871), .B1(n7327), .B2(n8678), .ZN(n7328)
         );
  AOI21_X1 U8923 ( .B1(n9831), .B2(P2_REG2_REG_0__SCAN_IN), .A(n7328), .ZN(
        n7330) );
  OAI21_X1 U8924 ( .B1(n8806), .B2(n9805), .A(n9874), .ZN(n7329) );
  OAI211_X1 U8925 ( .C1(n7331), .C2(n8808), .A(n7330), .B(n7329), .ZN(P2_U3296) );
  INV_X1 U8926 ( .A(n7332), .ZN(n7361) );
  OAI222_X1 U8927 ( .A1(n9527), .A2(n7361), .B1(P1_U3084), .B2(n8054), .C1(
        n7333), .C2(n9524), .ZN(P1_U3332) );
  NAND2_X1 U8928 ( .A1(n7341), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7335) );
  NAND2_X1 U8929 ( .A1(n7335), .A2(n7334), .ZN(n7339) );
  INV_X1 U8930 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7336) );
  MUX2_X1 U8931 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7336), .S(n7473), .Z(n7337)
         );
  INV_X1 U8932 ( .A(n7337), .ZN(n7338) );
  NOR2_X1 U8933 ( .A1(n7339), .A2(n7338), .ZN(n7467) );
  AOI21_X1 U8934 ( .B1(n7339), .B2(n7338), .A(n7467), .ZN(n7348) );
  AND2_X1 U8935 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8424) );
  INV_X1 U8936 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7342) );
  MUX2_X1 U8937 ( .A(n7342), .B(P2_REG1_REG_11__SCAN_IN), .S(n7473), .Z(n7343)
         );
  AOI211_X1 U8938 ( .C1(n7344), .C2(n7343), .A(n7472), .B(n9787), .ZN(n7345)
         );
  AOI211_X1 U8939 ( .C1(n9785), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n8424), .B(
        n7345), .ZN(n7347) );
  NAND2_X1 U8940 ( .A1(n8529), .A2(n7473), .ZN(n7346) );
  OAI211_X1 U8941 ( .C1(n7348), .C2(n9788), .A(n7347), .B(n7346), .ZN(P2_U3256) );
  AOI21_X1 U8942 ( .B1(n9021), .B2(n9046), .A(n7349), .ZN(n7351) );
  NAND2_X1 U8943 ( .A1(n9033), .A2(n4681), .ZN(n7350) );
  OAI211_X1 U8944 ( .C1(n7405), .C2(n9027), .A(n7351), .B(n7350), .ZN(n7358)
         );
  NAND2_X1 U8945 ( .A1(n6070), .A2(n7353), .ZN(n7354) );
  XNOR2_X1 U8946 ( .A(n7355), .B(n7354), .ZN(n7356) );
  NOR2_X1 U8947 ( .A1(n7356), .A2(n4371), .ZN(n7357) );
  AOI211_X1 U8948 ( .C1(n7403), .C2(n9031), .A(n7358), .B(n7357), .ZN(n7359)
         );
  INV_X1 U8949 ( .A(n7359), .ZN(P1_U3211) );
  OAI222_X1 U8950 ( .A1(P2_U3152), .A2(n7362), .B1(n8920), .B2(n7361), .C1(
        n7360), .C2(n8259), .ZN(P2_U3337) );
  XNOR2_X1 U8951 ( .A(n7364), .B(n7363), .ZN(n7370) );
  INV_X1 U8952 ( .A(n8452), .ZN(n8426) );
  OR2_X1 U8953 ( .A1(n7670), .A2(n8765), .ZN(n7365) );
  OAI21_X1 U8954 ( .B1(n7553), .B2(n8277), .A(n7365), .ZN(n9801) );
  INV_X1 U8955 ( .A(n9804), .ZN(n7366) );
  OAI22_X1 U8956 ( .A1(n8458), .A2(n9914), .B1(n8464), .B2(n7366), .ZN(n7367)
         );
  AOI211_X1 U8957 ( .C1(n8426), .C2(n9801), .A(n7368), .B(n7367), .ZN(n7369)
         );
  OAI21_X1 U8958 ( .B1(n7370), .B2(n8445), .A(n7369), .ZN(P2_U3223) );
  NOR2_X1 U8959 ( .A1(n9048), .A2(n7540), .ZN(n8000) );
  NAND2_X1 U8960 ( .A1(n9048), .A2(n7540), .ZN(n7395) );
  NAND2_X1 U8961 ( .A1(n7537), .A2(n7444), .ZN(n8067) );
  NAND2_X1 U8962 ( .A1(n4681), .A2(n9766), .ZN(n7396) );
  NAND2_X1 U8963 ( .A1(n8067), .A2(n7396), .ZN(n8069) );
  INV_X1 U8964 ( .A(n8069), .ZN(n7446) );
  NAND2_X1 U8965 ( .A1(n7372), .A2(n4823), .ZN(n8081) );
  NAND2_X1 U8966 ( .A1(n7380), .A2(n7454), .ZN(n8068) );
  NAND2_X1 U8967 ( .A1(n8081), .A2(n8068), .ZN(n7504) );
  NAND2_X1 U8968 ( .A1(n7373), .A2(n7598), .ZN(n8073) );
  NAND2_X1 U8969 ( .A1(n9046), .A2(n7374), .ZN(n7962) );
  AND2_X1 U8970 ( .A1(n8073), .A2(n7962), .ZN(n8028) );
  XNOR2_X1 U8971 ( .A(n7504), .B(n8028), .ZN(n7375) );
  AOI222_X1 U8972 ( .A1(n9725), .A2(n7375), .B1(n9546), .B2(n9721), .C1(n9047), 
        .C2(n9720), .ZN(n7600) );
  NAND2_X1 U8973 ( .A1(n9048), .A2(n7376), .ZN(n7377) );
  NAND2_X1 U8974 ( .A1(n7439), .A2(n8069), .ZN(n7438) );
  NAND2_X1 U8975 ( .A1(n7537), .A2(n9766), .ZN(n7379) );
  NAND2_X1 U8976 ( .A1(n7438), .A2(n7379), .ZN(n7393) );
  NAND2_X1 U8977 ( .A1(n8068), .A2(n8071), .ZN(n8026) );
  NAND2_X1 U8978 ( .A1(n7393), .A2(n8026), .ZN(n7392) );
  NAND2_X1 U8979 ( .A1(n7380), .A2(n7405), .ZN(n7381) );
  OAI21_X1 U8980 ( .B1(n4361), .B2(n7382), .A(n7502), .ZN(n7601) );
  INV_X1 U8981 ( .A(n7413), .ZN(n7383) );
  OAI22_X1 U8982 ( .A1(n9740), .A2(n7384), .B1(n7383), .B2(n9142), .ZN(n7385)
         );
  AOI21_X1 U8983 ( .B1(n9551), .B2(n7598), .A(n7385), .ZN(n7389) );
  NAND2_X1 U8984 ( .A1(n7401), .A2(n7598), .ZN(n7386) );
  NAND2_X1 U8985 ( .A1(n7386), .A2(n9554), .ZN(n7387) );
  NOR2_X1 U8986 ( .A1(n7509), .A2(n7387), .ZN(n7597) );
  NAND2_X1 U8987 ( .A1(n7597), .A2(n9557), .ZN(n7388) );
  OAI211_X1 U8988 ( .C1(n7601), .C2(n9365), .A(n7389), .B(n7388), .ZN(n7390)
         );
  INV_X1 U8989 ( .A(n7390), .ZN(n7391) );
  OAI21_X1 U8990 ( .B1(n9743), .B2(n7600), .A(n7391), .ZN(P1_U3283) );
  OAI21_X1 U8991 ( .B1(n7393), .B2(n8026), .A(n7392), .ZN(n7394) );
  INV_X1 U8992 ( .A(n7394), .ZN(n7457) );
  AND2_X1 U8993 ( .A1(n7396), .A2(n7395), .ZN(n8002) );
  NAND2_X1 U8994 ( .A1(n7397), .A2(n8002), .ZN(n7398) );
  NAND2_X1 U8995 ( .A1(n7398), .A2(n8067), .ZN(n8043) );
  XOR2_X1 U8996 ( .A(n8026), .B(n8043), .Z(n7399) );
  AOI222_X1 U8997 ( .A1(n9725), .A2(n7399), .B1(n9046), .B2(n9721), .C1(n4681), 
        .C2(n9720), .ZN(n7456) );
  MUX2_X1 U8998 ( .A(n7400), .B(n7456), .S(n9740), .Z(n7408) );
  INV_X1 U8999 ( .A(n7401), .ZN(n7402) );
  AOI211_X1 U9000 ( .C1(n7454), .C2(n7442), .A(n9767), .B(n7402), .ZN(n7453)
         );
  INV_X1 U9001 ( .A(n7403), .ZN(n7404) );
  OAI22_X1 U9002 ( .A1(n9341), .A2(n7405), .B1(n7404), .B2(n9142), .ZN(n7406)
         );
  AOI21_X1 U9003 ( .B1(n7453), .B2(n9557), .A(n7406), .ZN(n7407) );
  OAI211_X1 U9004 ( .C1(n7457), .C2(n9365), .A(n7408), .B(n7407), .ZN(P1_U3284) );
  NAND2_X1 U9005 ( .A1(n7410), .A2(n7409), .ZN(n7412) );
  XNOR2_X1 U9006 ( .A(n7412), .B(n7411), .ZN(n7420) );
  INV_X1 U9007 ( .A(n9546), .ZN(n7417) );
  NAND2_X1 U9008 ( .A1(n9031), .A2(n7413), .ZN(n7416) );
  NOR2_X1 U9009 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7414), .ZN(n9671) );
  AOI21_X1 U9010 ( .B1(n9033), .B2(n9047), .A(n9671), .ZN(n7415) );
  OAI211_X1 U9011 ( .C1(n7417), .C2(n9036), .A(n7416), .B(n7415), .ZN(n7418)
         );
  AOI21_X1 U9012 ( .B1(n9038), .B2(n7598), .A(n7418), .ZN(n7419) );
  OAI21_X1 U9013 ( .B1(n7420), .B2(n4371), .A(n7419), .ZN(P1_U3219) );
  INV_X1 U9014 ( .A(n7443), .ZN(n7437) );
  AND2_X1 U9015 ( .A1(n7422), .A2(n7421), .ZN(n7424) );
  NAND2_X1 U9016 ( .A1(n7424), .A2(n7423), .ZN(n7425) );
  OAI21_X1 U9017 ( .B1(n7424), .B2(n7423), .A(n7425), .ZN(n7542) );
  NOR2_X1 U9018 ( .A1(n7542), .A2(n7543), .ZN(n7541) );
  INV_X1 U9019 ( .A(n7425), .ZN(n7426) );
  NOR3_X1 U9020 ( .A1(n7541), .A2(n7427), .A3(n7426), .ZN(n7430) );
  INV_X1 U9021 ( .A(n7428), .ZN(n7429) );
  OAI21_X1 U9022 ( .B1(n7430), .B2(n7429), .A(n9018), .ZN(n7436) );
  AOI21_X1 U9023 ( .B1(n9021), .B2(n9047), .A(n7431), .ZN(n7432) );
  OAI21_X1 U9024 ( .B1(n7433), .B2(n9023), .A(n7432), .ZN(n7434) );
  AOI21_X1 U9025 ( .B1(n9038), .B2(n7444), .A(n7434), .ZN(n7435) );
  OAI211_X1 U9026 ( .C1(n9000), .C2(n7437), .A(n7436), .B(n7435), .ZN(P1_U3237) );
  OAI21_X1 U9027 ( .B1(n7439), .B2(n8069), .A(n7438), .ZN(n9771) );
  OR2_X1 U9028 ( .A1(n7440), .A2(n9766), .ZN(n7441) );
  NAND2_X1 U9029 ( .A1(n7442), .A2(n7441), .ZN(n9768) );
  AOI22_X1 U9030 ( .A1(n9551), .A2(n7444), .B1(n7443), .B2(n9728), .ZN(n7445)
         );
  OAI21_X1 U9031 ( .B1(n9768), .B2(n9384), .A(n7445), .ZN(n7451) );
  XNOR2_X1 U9032 ( .A(n8070), .B(n7446), .ZN(n7449) );
  NAND2_X1 U9033 ( .A1(n9771), .A2(n9549), .ZN(n7448) );
  AOI22_X1 U9034 ( .A1(n9047), .A2(n9721), .B1(n9720), .B2(n9048), .ZN(n7447)
         );
  OAI211_X1 U9035 ( .C1(n9318), .C2(n7449), .A(n7448), .B(n7447), .ZN(n9769)
         );
  MUX2_X1 U9036 ( .A(n9769), .B(P1_REG2_REG_6__SCAN_IN), .S(n9743), .Z(n7450)
         );
  AOI211_X1 U9037 ( .C1(n9558), .C2(n9771), .A(n7451), .B(n7450), .ZN(n7452)
         );
  INV_X1 U9038 ( .A(n7452), .ZN(P1_U3285) );
  AOI21_X1 U9039 ( .B1(n9487), .B2(n7454), .A(n7453), .ZN(n7455) );
  OAI211_X1 U9040 ( .C1(n9562), .C2(n7457), .A(n7456), .B(n7455), .ZN(n7459)
         );
  NAND2_X1 U9041 ( .A1(n7459), .A2(n9774), .ZN(n7458) );
  OAI21_X1 U9042 ( .B1(n9774), .B2(n6060), .A(n7458), .ZN(P1_U3475) );
  NAND2_X1 U9043 ( .A1(n7459), .A2(n9782), .ZN(n7460) );
  OAI21_X1 U9044 ( .B1(n9782), .B2(n7461), .A(n7460), .ZN(P1_U3530) );
  INV_X1 U9045 ( .A(n7462), .ZN(n7465) );
  OAI222_X1 U9046 ( .A1(n9524), .A2(n7463), .B1(n9527), .B2(n7465), .C1(n6455), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  INV_X1 U9047 ( .A(n5565), .ZN(n7466) );
  OAI222_X1 U9048 ( .A1(n7466), .A2(P2_U3152), .B1(n8920), .B2(n7465), .C1(
        n7464), .C2(n8259), .ZN(P2_U3336) );
  INV_X1 U9049 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7469) );
  MUX2_X1 U9050 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7469), .S(n7702), .Z(n7470)
         );
  NAND2_X1 U9051 ( .A1(n7470), .A2(n7471), .ZN(n7696) );
  OAI211_X1 U9052 ( .C1(n7471), .C2(n7470), .A(n9784), .B(n7696), .ZN(n7482)
         );
  AOI21_X1 U9053 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7473), .A(n7472), .ZN(
        n7476) );
  INV_X1 U9054 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7474) );
  MUX2_X1 U9055 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7474), .S(n7702), .Z(n7475)
         );
  NAND2_X1 U9056 ( .A1(n7476), .A2(n7475), .ZN(n7701) );
  OAI21_X1 U9057 ( .B1(n7476), .B2(n7475), .A(n7701), .ZN(n7480) );
  NAND2_X1 U9058 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8333) );
  INV_X1 U9059 ( .A(n8333), .ZN(n7479) );
  INV_X1 U9060 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7477) );
  NOR2_X1 U9061 ( .A1(n8527), .A2(n7477), .ZN(n7478) );
  AOI211_X1 U9062 ( .C1(n9783), .C2(n7480), .A(n7479), .B(n7478), .ZN(n7481)
         );
  OAI211_X1 U9063 ( .C1(n9786), .C2(n7483), .A(n7482), .B(n7481), .ZN(P2_U3257) );
  NOR2_X1 U9064 ( .A1(n9829), .A2(n7484), .ZN(n7487) );
  OAI22_X1 U9065 ( .A1(n8539), .A2(n7485), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8678), .ZN(n7486) );
  AOI211_X1 U9066 ( .C1(n9829), .C2(n7488), .A(n7487), .B(n7486), .ZN(n7491)
         );
  NAND2_X1 U9067 ( .A1(n9581), .A2(n7489), .ZN(n7490) );
  OAI211_X1 U9068 ( .C1(n7492), .C2(n8795), .A(n7491), .B(n7490), .ZN(P2_U3293) );
  XOR2_X1 U9069 ( .A(n7494), .B(n7493), .Z(n7500) );
  NAND2_X1 U9070 ( .A1(n9031), .A2(n7511), .ZN(n7497) );
  AOI21_X1 U9071 ( .B1(n9033), .B2(n9046), .A(n7495), .ZN(n7496) );
  OAI211_X1 U9072 ( .C1(n7734), .C2(n9036), .A(n7497), .B(n7496), .ZN(n7498)
         );
  AOI21_X1 U9073 ( .B1(n9038), .B2(n9486), .A(n7498), .ZN(n7499) );
  OAI21_X1 U9074 ( .B1(n7500), .B2(n4371), .A(n7499), .ZN(P1_U3229) );
  NAND2_X1 U9075 ( .A1(n9046), .A2(n7598), .ZN(n7501) );
  INV_X1 U9076 ( .A(n9486), .ZN(n7514) );
  NOR2_X1 U9077 ( .A1(n9546), .A2(n7514), .ZN(n8075) );
  NAND2_X1 U9078 ( .A1(n9546), .A2(n7514), .ZN(n9541) );
  INV_X1 U9079 ( .A(n9541), .ZN(n7503) );
  NOR2_X1 U9080 ( .A1(n8075), .A2(n7503), .ZN(n8029) );
  XNOR2_X1 U9081 ( .A(n7729), .B(n8029), .ZN(n9485) );
  NAND2_X1 U9082 ( .A1(n7504), .A2(n7962), .ZN(n7505) );
  XOR2_X1 U9083 ( .A(n8029), .B(n7732), .Z(n7507) );
  AOI22_X1 U9084 ( .A1(n9720), .A2(n9046), .B1(n9045), .B2(n9721), .ZN(n7506)
         );
  OAI21_X1 U9085 ( .B1(n7507), .B2(n9318), .A(n7506), .ZN(n7508) );
  AOI21_X1 U9086 ( .B1(n9485), .B2(n9549), .A(n7508), .ZN(n9490) );
  INV_X1 U9087 ( .A(n7509), .ZN(n7510) );
  AOI21_X1 U9088 ( .B1(n9486), .B2(n7510), .A(n9555), .ZN(n9488) );
  NAND2_X1 U9089 ( .A1(n9488), .A2(n9346), .ZN(n7513) );
  AOI22_X1 U9090 ( .A1(n9743), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7511), .B2(
        n9728), .ZN(n7512) );
  OAI211_X1 U9091 ( .C1(n7514), .C2(n9341), .A(n7513), .B(n7512), .ZN(n7515)
         );
  AOI21_X1 U9092 ( .B1(n9485), .B2(n9558), .A(n7515), .ZN(n7516) );
  OAI21_X1 U9093 ( .B1(n9490), .B2(n9743), .A(n7516), .ZN(P1_U3282) );
  AOI22_X1 U9094 ( .A1(n9581), .A2(n7517), .B1(n9805), .B2(n8387), .ZN(n7524)
         );
  INV_X1 U9095 ( .A(n7518), .ZN(n7522) );
  OAI22_X1 U9096 ( .A1(n8678), .A2(n7520), .B1(n7519), .B2(n9829), .ZN(n7521)
         );
  AOI21_X1 U9097 ( .B1(n9812), .B2(n7522), .A(n7521), .ZN(n7523) );
  OAI211_X1 U9098 ( .C1(n9831), .C2(n7525), .A(n7524), .B(n7523), .ZN(P2_U3292) );
  XNOR2_X1 U9099 ( .A(n7527), .B(n7526), .ZN(n7528) );
  XNOR2_X1 U9100 ( .A(n7529), .B(n7528), .ZN(n7535) );
  INV_X1 U9101 ( .A(n9545), .ZN(n7790) );
  NAND2_X1 U9102 ( .A1(n9031), .A2(n9550), .ZN(n7532) );
  NOR2_X1 U9103 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7530), .ZN(n9693) );
  AOI21_X1 U9104 ( .B1(n9033), .B2(n9546), .A(n9693), .ZN(n7531) );
  OAI211_X1 U9105 ( .C1(n7790), .C2(n9036), .A(n7532), .B(n7531), .ZN(n7533)
         );
  AOI21_X1 U9106 ( .B1(n9038), .B2(n9552), .A(n7533), .ZN(n7534) );
  OAI21_X1 U9107 ( .B1(n7535), .B2(n4371), .A(n7534), .ZN(P1_U3215) );
  NAND2_X1 U9108 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9663) );
  INV_X1 U9109 ( .A(n9663), .ZN(n7536) );
  AOI21_X1 U9110 ( .B1(n9033), .B2(n9049), .A(n7536), .ZN(n7539) );
  OR2_X1 U9111 ( .A1(n9036), .A2(n7537), .ZN(n7538) );
  OAI211_X1 U9112 ( .C1(n9027), .C2(n7540), .A(n7539), .B(n7538), .ZN(n7546)
         );
  AOI21_X1 U9113 ( .B1(n7543), .B2(n7542), .A(n7541), .ZN(n7544) );
  NOR2_X1 U9114 ( .A1(n7544), .A2(n4371), .ZN(n7545) );
  AOI211_X1 U9115 ( .C1(n7547), .C2(n9031), .A(n7546), .B(n7545), .ZN(n7548)
         );
  INV_X1 U9116 ( .A(n7548), .ZN(P1_U3225) );
  XNOR2_X1 U9117 ( .A(n7549), .B(n7563), .ZN(n7551) );
  OR2_X1 U9118 ( .A1(n7830), .A2(n8765), .ZN(n7550) );
  OAI21_X1 U9119 ( .B1(n7691), .B2(n8277), .A(n7550), .ZN(n8425) );
  AOI21_X1 U9120 ( .B1(n7551), .B2(n9803), .A(n8425), .ZN(n9937) );
  NAND2_X1 U9121 ( .A1(n7553), .A2(n7552), .ZN(n7554) );
  NAND2_X1 U9122 ( .A1(n9806), .A2(n8485), .ZN(n7557) );
  INV_X1 U9123 ( .A(n7691), .ZN(n8483) );
  NAND2_X1 U9124 ( .A1(n9928), .A2(n8483), .ZN(n7558) );
  INV_X1 U9125 ( .A(n7558), .ZN(n7559) );
  INV_X1 U9126 ( .A(n7670), .ZN(n8484) );
  OR2_X1 U9127 ( .A1(n7690), .A2(n8484), .ZN(n7664) );
  AND2_X1 U9128 ( .A1(n7668), .A2(n7664), .ZN(n7665) );
  OR2_X1 U9129 ( .A1(n7559), .A2(n7665), .ZN(n7560) );
  OAI21_X1 U9130 ( .B1(n7575), .B2(n4328), .A(n7560), .ZN(n7562) );
  NOR2_X1 U9131 ( .A1(n7564), .A2(n7563), .ZN(n7565) );
  NAND2_X1 U9132 ( .A1(n9810), .A2(n9914), .ZN(n9809) );
  INV_X1 U9133 ( .A(n8427), .ZN(n9938) );
  OAI21_X1 U9134 ( .B1(n7677), .B2(n9938), .A(n9905), .ZN(n7566) );
  OR2_X1 U9135 ( .A1(n7566), .A2(n7773), .ZN(n9936) );
  INV_X1 U9136 ( .A(n8428), .ZN(n7567) );
  OAI22_X1 U9137 ( .A1(n9829), .A2(n7336), .B1(n7567), .B2(n8678), .ZN(n7568)
         );
  AOI21_X1 U9138 ( .B1(n9805), .B2(n8427), .A(n7568), .ZN(n7569) );
  OAI21_X1 U9139 ( .B1(n9936), .B2(n8539), .A(n7569), .ZN(n7570) );
  AOI21_X1 U9140 ( .B1(n4359), .B2(n9581), .A(n7570), .ZN(n7571) );
  OAI21_X1 U9141 ( .B1(n9831), .B2(n9937), .A(n7571), .ZN(P2_U3285) );
  INV_X1 U9142 ( .A(n7593), .ZN(n7574) );
  NAND2_X1 U9143 ( .A1(n7572), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8181) );
  NAND2_X1 U9144 ( .A1(n9520), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7573) );
  OAI211_X1 U9145 ( .C1(n7574), .C2(n9522), .A(n8181), .B(n7573), .ZN(P1_U3330) );
  NAND2_X1 U9146 ( .A1(n7576), .A2(n7579), .ZN(n7666) );
  OAI21_X1 U9147 ( .B1(n7576), .B2(n7579), .A(n7666), .ZN(n9924) );
  INV_X1 U9148 ( .A(n9924), .ZN(n7591) );
  INV_X1 U9149 ( .A(n7577), .ZN(n7578) );
  NAND2_X1 U9150 ( .A1(n9829), .A2(n7578), .ZN(n9808) );
  XNOR2_X1 U9151 ( .A(n7580), .B(n7579), .ZN(n7584) );
  INV_X1 U9152 ( .A(n9799), .ZN(n7581) );
  NAND2_X1 U9153 ( .A1(n9924), .A2(n7581), .ZN(n7583) );
  AOI22_X1 U9154 ( .A1(n8799), .A2(n8485), .B1(n8483), .B2(n8801), .ZN(n7582)
         );
  OAI211_X1 U9155 ( .C1(n9570), .C2(n7584), .A(n7583), .B(n7582), .ZN(n9922)
         );
  NAND2_X1 U9156 ( .A1(n9922), .A2(n9829), .ZN(n7590) );
  INV_X1 U9157 ( .A(n7585), .ZN(n7689) );
  OAI22_X1 U9158 ( .A1(n9829), .A2(n7036), .B1(n7689), .B2(n8678), .ZN(n7588)
         );
  NAND2_X1 U9159 ( .A1(n9809), .A2(n7690), .ZN(n7586) );
  NAND2_X1 U9160 ( .A1(n7678), .A2(n7586), .ZN(n9921) );
  NOR2_X1 U9161 ( .A1(n8683), .A2(n9921), .ZN(n7587) );
  AOI211_X1 U9162 ( .C1(n9805), .C2(n7690), .A(n7588), .B(n7587), .ZN(n7589)
         );
  OAI211_X1 U9163 ( .C1(n7591), .C2(n9808), .A(n7590), .B(n7589), .ZN(P2_U3287) );
  NAND2_X1 U9164 ( .A1(n7593), .A2(n7592), .ZN(n7595) );
  OAI211_X1 U9165 ( .C1(n7596), .C2(n8259), .A(n7595), .B(n7594), .ZN(P2_U3335) );
  INV_X1 U9166 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9666) );
  AOI21_X1 U9167 ( .B1(n9487), .B2(n7598), .A(n7597), .ZN(n7599) );
  OAI211_X1 U9168 ( .C1(n7601), .C2(n9562), .A(n7600), .B(n7599), .ZN(n7603)
         );
  NAND2_X1 U9169 ( .A1(n7603), .A2(n9782), .ZN(n7602) );
  OAI21_X1 U9170 ( .B1(n9782), .B2(n9666), .A(n7602), .ZN(P1_U3531) );
  NAND2_X1 U9171 ( .A1(n7603), .A2(n9774), .ZN(n7604) );
  OAI21_X1 U9172 ( .B1(n9774), .B2(n6077), .A(n7604), .ZN(P1_U3478) );
  XNOR2_X1 U9173 ( .A(n7605), .B(n5805), .ZN(n7609) );
  OAI22_X1 U9174 ( .A1(n7607), .A2(n8765), .B1(n7606), .B2(n8277), .ZN(n7608)
         );
  AOI21_X1 U9175 ( .B1(n7609), .B2(n9803), .A(n7608), .ZN(n9893) );
  XNOR2_X1 U9176 ( .A(n7010), .B(n7610), .ZN(n9895) );
  AOI22_X1 U9177 ( .A1(n9895), .A2(n9581), .B1(n9805), .B2(n4267), .ZN(n7612)
         );
  NAND2_X1 U9178 ( .A1(n9883), .A2(n4267), .ZN(n9891) );
  NAND3_X1 U9179 ( .A1(n8806), .A2(n9890), .A3(n9891), .ZN(n7611) );
  OAI211_X1 U9180 ( .C1(n9831), .C2(n9893), .A(n7612), .B(n7611), .ZN(n7616)
         );
  OAI22_X1 U9181 ( .A1(n8678), .A2(n7614), .B1(n7613), .B2(n9829), .ZN(n7615)
         );
  OR2_X1 U9182 ( .A1(n7616), .A2(n7615), .ZN(P2_U3294) );
  NOR2_X1 U9183 ( .A1(n7618), .A2(n7617), .ZN(n7620) );
  NOR2_X1 U9184 ( .A1(n7620), .A2(n7619), .ZN(n9064) );
  XNOR2_X1 U9185 ( .A(n9064), .B(n9071), .ZN(n7622) );
  INV_X1 U9186 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7621) );
  NOR2_X1 U9187 ( .A1(n7621), .A2(n7622), .ZN(n9065) );
  AOI211_X1 U9188 ( .C1(n7622), .C2(n7621), .A(n9065), .B(n9688), .ZN(n7631)
         );
  NAND2_X1 U9189 ( .A1(n9711), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7629) );
  OAI21_X1 U9190 ( .B1(n7624), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7623), .ZN(
        n9070) );
  XNOR2_X1 U9191 ( .A(n9071), .B(n9070), .ZN(n7626) );
  INV_X1 U9192 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7625) );
  NOR2_X1 U9193 ( .A1(n7625), .A2(n7626), .ZN(n9072) );
  AOI21_X1 U9194 ( .B1(n7626), .B2(n7625), .A(n9072), .ZN(n7627) );
  AND2_X1 U9195 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9032) );
  AOI21_X1 U9196 ( .B1(n9712), .B2(n7627), .A(n9032), .ZN(n7628) );
  OAI211_X1 U9197 ( .C1(n9641), .C2(n9071), .A(n7629), .B(n7628), .ZN(n7630)
         );
  OR2_X1 U9198 ( .A1(n7631), .A2(n7630), .ZN(P1_U3256) );
  INV_X1 U9199 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10006) );
  NOR2_X1 U9200 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7632) );
  AOI21_X1 U9201 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7632), .ZN(n9975) );
  NOR2_X1 U9202 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7633) );
  AOI21_X1 U9203 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7633), .ZN(n9978) );
  NOR2_X1 U9204 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7634) );
  AOI21_X1 U9205 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7634), .ZN(n9981) );
  NOR2_X1 U9206 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7635) );
  AOI21_X1 U9207 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7635), .ZN(n9984) );
  NOR2_X1 U9208 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7636) );
  AOI21_X1 U9209 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7636), .ZN(n9987) );
  NOR2_X1 U9210 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7643) );
  XNOR2_X1 U9211 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10015) );
  NAND2_X1 U9212 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7641) );
  XNOR2_X1 U9213 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n7637), .ZN(n10013) );
  NAND2_X1 U9214 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7639) );
  XOR2_X1 U9215 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10011) );
  AOI21_X1 U9216 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9968) );
  INV_X1 U9217 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9972) );
  NAND3_X1 U9218 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9970) );
  OAI21_X1 U9219 ( .B1(n9968), .B2(n9972), .A(n9970), .ZN(n10010) );
  NAND2_X1 U9220 ( .A1(n10011), .A2(n10010), .ZN(n7638) );
  NAND2_X1 U9221 ( .A1(n7639), .A2(n7638), .ZN(n10012) );
  NAND2_X1 U9222 ( .A1(n10013), .A2(n10012), .ZN(n7640) );
  NAND2_X1 U9223 ( .A1(n7641), .A2(n7640), .ZN(n10014) );
  NOR2_X1 U9224 ( .A1(n10015), .A2(n10014), .ZN(n7642) );
  NOR2_X1 U9225 ( .A1(n7643), .A2(n7642), .ZN(n7644) );
  NOR2_X1 U9226 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7644), .ZN(n9998) );
  AND2_X1 U9227 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7644), .ZN(n9997) );
  NOR2_X1 U9228 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9997), .ZN(n7645) );
  NOR2_X1 U9229 ( .A1(n9998), .A2(n7645), .ZN(n7646) );
  NAND2_X1 U9230 ( .A1(n7646), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7648) );
  XOR2_X1 U9231 ( .A(n7646), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10000) );
  NAND2_X1 U9232 ( .A1(n10000), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7647) );
  NAND2_X1 U9233 ( .A1(n7648), .A2(n7647), .ZN(n7649) );
  NAND2_X1 U9234 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7649), .ZN(n7651) );
  XOR2_X1 U9235 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7649), .Z(n10009) );
  NAND2_X1 U9236 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10009), .ZN(n7650) );
  NAND2_X1 U9237 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  NAND2_X1 U9238 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7652), .ZN(n7654) );
  XOR2_X1 U9239 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7652), .Z(n10008) );
  NAND2_X1 U9240 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10008), .ZN(n7653) );
  NAND2_X1 U9241 ( .A1(n7654), .A2(n7653), .ZN(n7655) );
  AND2_X1 U9242 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7655), .ZN(n7656) );
  XNOR2_X1 U9243 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7655), .ZN(n10003) );
  NAND2_X1 U9244 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7657) );
  OAI21_X1 U9245 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7657), .ZN(n9995) );
  NAND2_X1 U9246 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7658) );
  OAI21_X1 U9247 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7658), .ZN(n9992) );
  AOI21_X1 U9248 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9991), .ZN(n9990) );
  NOR2_X1 U9249 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7659) );
  AOI21_X1 U9250 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7659), .ZN(n9989) );
  NAND2_X1 U9251 ( .A1(n9990), .A2(n9989), .ZN(n9988) );
  OAI21_X1 U9252 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9988), .ZN(n9986) );
  NAND2_X1 U9253 ( .A1(n9987), .A2(n9986), .ZN(n9985) );
  OAI21_X1 U9254 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9985), .ZN(n9983) );
  NAND2_X1 U9255 ( .A1(n9984), .A2(n9983), .ZN(n9982) );
  OAI21_X1 U9256 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9982), .ZN(n9980) );
  NAND2_X1 U9257 ( .A1(n9981), .A2(n9980), .ZN(n9979) );
  OAI21_X1 U9258 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9979), .ZN(n9977) );
  NAND2_X1 U9259 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  OAI21_X1 U9260 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9976), .ZN(n9974) );
  NAND2_X1 U9261 ( .A1(n9975), .A2(n9974), .ZN(n9973) );
  OAI21_X1 U9262 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9973), .ZN(n10005) );
  NOR2_X1 U9263 ( .A1(n10006), .A2(n10005), .ZN(n7660) );
  NAND2_X1 U9264 ( .A1(n10006), .A2(n10005), .ZN(n10004) );
  OAI21_X1 U9265 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7660), .A(n10004), .ZN(
        n7663) );
  XNOR2_X1 U9266 ( .A(n7661), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7662) );
  XNOR2_X1 U9267 ( .A(n7663), .B(n7662), .ZN(ADD_1071_U4) );
  AND2_X1 U9268 ( .A1(n7666), .A2(n7664), .ZN(n7669) );
  NAND2_X1 U9269 ( .A1(n7666), .A2(n7665), .ZN(n7667) );
  OAI21_X1 U9270 ( .B1(n7669), .B2(n7668), .A(n7667), .ZN(n9932) );
  OAI22_X1 U9271 ( .A1(n8335), .A2(n8765), .B1(n7670), .B2(n8277), .ZN(n7671)
         );
  INV_X1 U9272 ( .A(n7671), .ZN(n7676) );
  OAI211_X1 U9273 ( .C1(n7674), .C2(n7673), .A(n7672), .B(n9803), .ZN(n7675)
         );
  OAI211_X1 U9274 ( .C1(n9932), .C2(n9799), .A(n7676), .B(n7675), .ZN(n9934)
         );
  NAND2_X1 U9275 ( .A1(n9934), .A2(n9829), .ZN(n7683) );
  AOI211_X1 U9276 ( .C1(n9928), .C2(n7678), .A(n9943), .B(n7677), .ZN(n9927)
         );
  INV_X1 U9277 ( .A(n9928), .ZN(n7715) );
  NOR2_X1 U9278 ( .A1(n8795), .A2(n7715), .ZN(n7681) );
  INV_X1 U9279 ( .A(n7679), .ZN(n7714) );
  OAI22_X1 U9280 ( .A1(n9829), .A2(n7131), .B1(n7714), .B2(n8678), .ZN(n7680)
         );
  AOI211_X1 U9281 ( .C1(n9927), .C2(n9812), .A(n7681), .B(n7680), .ZN(n7682)
         );
  OAI211_X1 U9282 ( .C1(n9932), .C2(n9808), .A(n7683), .B(n7682), .ZN(P2_U3286) );
  INV_X1 U9283 ( .A(n7684), .ZN(n7685) );
  AOI21_X1 U9284 ( .B1(n7687), .B2(n7686), .A(n7685), .ZN(n7695) );
  OAI21_X1 U9285 ( .B1(n8464), .B2(n7689), .A(n7688), .ZN(n7693) );
  INV_X1 U9286 ( .A(n7690), .ZN(n9920) );
  OAI22_X1 U9287 ( .A1(n8458), .A2(n9920), .B1(n8466), .B2(n7691), .ZN(n7692)
         );
  AOI211_X1 U9288 ( .C1(n7718), .C2(n8485), .A(n7693), .B(n7692), .ZN(n7694)
         );
  OAI21_X1 U9289 ( .B1(n7695), .B2(n8445), .A(n7694), .ZN(P2_U3233) );
  NAND2_X1 U9290 ( .A1(n7702), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U9291 ( .A1(n7697), .A2(n7696), .ZN(n7699) );
  AOI22_X1 U9292 ( .A1(n7812), .A2(n7804), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7805), .ZN(n7698) );
  NOR2_X1 U9293 ( .A1(n7699), .A2(n7698), .ZN(n7803) );
  AOI21_X1 U9294 ( .B1(n7699), .B2(n7698), .A(n7803), .ZN(n7710) );
  INV_X1 U9295 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7700) );
  AOI22_X1 U9296 ( .A1(n7812), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n7700), .B2(
        n7805), .ZN(n7704) );
  OAI21_X1 U9297 ( .B1(n7702), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7701), .ZN(
        n7703) );
  NAND2_X1 U9298 ( .A1(n7704), .A2(n7703), .ZN(n7811) );
  OAI21_X1 U9299 ( .B1(n7704), .B2(n7703), .A(n7811), .ZN(n7705) );
  NAND2_X1 U9300 ( .A1(n7705), .A2(n9783), .ZN(n7709) );
  NOR2_X1 U9301 ( .A1(n7706), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8406) );
  NOR2_X1 U9302 ( .A1(n9786), .A2(n7805), .ZN(n7707) );
  AOI211_X1 U9303 ( .C1(n9785), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n8406), .B(
        n7707), .ZN(n7708) );
  OAI211_X1 U9304 ( .C1(n7710), .C2(n9788), .A(n7709), .B(n7708), .ZN(P2_U3258) );
  XNOR2_X1 U9305 ( .A(n7712), .B(n7711), .ZN(n7720) );
  OAI21_X1 U9306 ( .B1(n8464), .B2(n7714), .A(n7713), .ZN(n7717) );
  OAI22_X1 U9307 ( .A1(n8458), .A2(n7715), .B1(n8466), .B2(n8335), .ZN(n7716)
         );
  AOI211_X1 U9308 ( .C1(n7718), .C2(n8484), .A(n7717), .B(n7716), .ZN(n7719)
         );
  OAI21_X1 U9309 ( .B1(n7720), .B2(n8445), .A(n7719), .ZN(P2_U3219) );
  XNOR2_X1 U9310 ( .A(n7722), .B(n7721), .ZN(n7727) );
  NAND2_X1 U9311 ( .A1(n9031), .A2(n7740), .ZN(n7724) );
  NOR2_X1 U9312 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6137), .ZN(n9056) );
  AOI21_X1 U9313 ( .B1(n9021), .B2(n9374), .A(n9056), .ZN(n7723) );
  OAI211_X1 U9314 ( .C1(n7734), .C2(n9023), .A(n7724), .B(n7723), .ZN(n7725)
         );
  AOI21_X1 U9315 ( .B1(n9038), .B2(n9479), .A(n7725), .ZN(n7726) );
  OAI21_X1 U9316 ( .B1(n7727), .B2(n4371), .A(n7726), .ZN(P1_U3234) );
  AND2_X1 U9317 ( .A1(n9546), .A2(n9486), .ZN(n7728) );
  NAND2_X1 U9318 ( .A1(n7734), .A2(n9552), .ZN(n8078) );
  NAND2_X1 U9319 ( .A1(n9565), .A2(n9045), .ZN(n7957) );
  NAND2_X1 U9320 ( .A1(n8078), .A2(n7957), .ZN(n9543) );
  NAND2_X1 U9321 ( .A1(n9540), .A2(n9543), .ZN(n7731) );
  NAND2_X1 U9322 ( .A1(n7734), .A2(n9565), .ZN(n7730) );
  XNOR2_X1 U9323 ( .A(n9479), .B(n7790), .ZN(n8033) );
  XNOR2_X1 U9324 ( .A(n7787), .B(n8033), .ZN(n9478) );
  NAND2_X1 U9325 ( .A1(n9478), .A2(n9549), .ZN(n7738) );
  AND2_X1 U9326 ( .A1(n7957), .A2(n9541), .ZN(n8074) );
  INV_X1 U9327 ( .A(n8033), .ZN(n8087) );
  XNOR2_X1 U9328 ( .A(n8208), .B(n8087), .ZN(n7736) );
  OAI22_X1 U9329 ( .A1(n7734), .A2(n9330), .B1(n7788), .B2(n9328), .ZN(n7735)
         );
  AOI21_X1 U9330 ( .B1(n7736), .B2(n9725), .A(n7735), .ZN(n7737) );
  NAND2_X1 U9331 ( .A1(n7738), .A2(n7737), .ZN(n9484) );
  INV_X1 U9332 ( .A(n9484), .ZN(n7745) );
  NAND2_X1 U9333 ( .A1(n9555), .A2(n9565), .ZN(n9553) );
  NAND2_X1 U9334 ( .A1(n9553), .A2(n9479), .ZN(n7739) );
  NAND2_X1 U9335 ( .A1(n7797), .A2(n7739), .ZN(n9481) );
  AOI22_X1 U9336 ( .A1(n9743), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7740), .B2(
        n9728), .ZN(n7742) );
  NAND2_X1 U9337 ( .A1(n9551), .A2(n9479), .ZN(n7741) );
  OAI211_X1 U9338 ( .C1(n9481), .C2(n9384), .A(n7742), .B(n7741), .ZN(n7743)
         );
  AOI21_X1 U9339 ( .B1(n9478), .B2(n9558), .A(n7743), .ZN(n7744) );
  OAI21_X1 U9340 ( .B1(n7745), .B2(n9743), .A(n7744), .ZN(P1_U3280) );
  NAND2_X1 U9341 ( .A1(n7747), .A2(n7746), .ZN(n7748) );
  XOR2_X1 U9342 ( .A(n7753), .B(n7748), .Z(n7750) );
  OAI21_X1 U9343 ( .B1(n7750), .B2(n9570), .A(n7749), .ZN(n9901) );
  INV_X1 U9344 ( .A(n9901), .ZN(n7764) );
  NAND2_X1 U9345 ( .A1(n7752), .A2(n7753), .ZN(n9897) );
  AND3_X1 U9346 ( .A1(n7751), .A2(n9581), .A3(n9897), .ZN(n7762) );
  NOR2_X1 U9347 ( .A1(n8795), .A2(n9900), .ZN(n7761) );
  NOR2_X1 U9348 ( .A1(n9829), .A2(n6908), .ZN(n7760) );
  AOI21_X1 U9349 ( .B1(n7755), .B2(n7754), .A(n9943), .ZN(n7757) );
  NAND2_X1 U9350 ( .A1(n7757), .A2(n7756), .ZN(n9898) );
  OAI22_X1 U9351 ( .A1(n8539), .A2(n9898), .B1(n7758), .B2(n8678), .ZN(n7759)
         );
  NOR4_X1 U9352 ( .A1(n7762), .A2(n7761), .A3(n7760), .A4(n7759), .ZN(n7763)
         );
  OAI21_X1 U9353 ( .B1(n9831), .B2(n7764), .A(n7763), .ZN(P2_U3290) );
  NAND2_X1 U9354 ( .A1(n7766), .A2(n7765), .ZN(n7767) );
  XOR2_X1 U9355 ( .A(n7771), .B(n7767), .Z(n7768) );
  OAI222_X1 U9356 ( .A1(n8765), .A2(n8480), .B1(n8277), .B2(n8335), .C1(n9570), 
        .C2(n7768), .ZN(n9945) );
  INV_X1 U9357 ( .A(n9945), .ZN(n7779) );
  INV_X1 U9358 ( .A(n8335), .ZN(n8482) );
  OAI21_X1 U9359 ( .B1(n7772), .B2(n7771), .A(n7822), .ZN(n9948) );
  INV_X1 U9360 ( .A(n8338), .ZN(n9942) );
  OAI21_X1 U9361 ( .B1(n7773), .B2(n9942), .A(n7825), .ZN(n9944) );
  INV_X1 U9362 ( .A(n7774), .ZN(n8334) );
  OAI22_X1 U9363 ( .A1(n9829), .A2(n7469), .B1(n8334), .B2(n8678), .ZN(n7775)
         );
  AOI21_X1 U9364 ( .B1(n9805), .B2(n8338), .A(n7775), .ZN(n7776) );
  OAI21_X1 U9365 ( .B1(n9944), .B2(n8683), .A(n7776), .ZN(n7777) );
  AOI21_X1 U9366 ( .B1(n9948), .B2(n9581), .A(n7777), .ZN(n7778) );
  OAI21_X1 U9367 ( .B1(n9831), .B2(n7779), .A(n7778), .ZN(P2_U3284) );
  INV_X1 U9368 ( .A(n7780), .ZN(n7784) );
  OAI222_X1 U9369 ( .A1(n9527), .A2(n7784), .B1(P1_U3084), .B2(n7782), .C1(
        n7781), .C2(n9524), .ZN(P1_U3329) );
  OAI222_X1 U9370 ( .A1(n7785), .A2(P2_U3152), .B1(n8920), .B2(n7784), .C1(
        n7783), .C2(n8259), .ZN(P2_U3334) );
  NAND2_X1 U9371 ( .A1(n9479), .A2(n9545), .ZN(n7786) );
  OR2_X1 U9372 ( .A1(n9597), .A2(n7788), .ZN(n8092) );
  NAND2_X1 U9373 ( .A1(n9597), .A2(n7788), .ZN(n8091) );
  NAND2_X1 U9374 ( .A1(n8092), .A2(n8091), .ZN(n8183) );
  INV_X1 U9375 ( .A(n8183), .ZN(n7789) );
  XNOR2_X1 U9376 ( .A(n8184), .B(n7789), .ZN(n9601) );
  NAND2_X1 U9377 ( .A1(n9479), .A2(n7790), .ZN(n8090) );
  INV_X1 U9378 ( .A(n8090), .ZN(n7791) );
  OR2_X1 U9379 ( .A1(n7790), .A2(n9479), .ZN(n7965) );
  OAI21_X1 U9380 ( .B1(n8208), .B2(n7791), .A(n7965), .ZN(n7792) );
  XNOR2_X1 U9381 ( .A(n7792), .B(n8183), .ZN(n7793) );
  NAND2_X1 U9382 ( .A1(n7793), .A2(n9725), .ZN(n7795) );
  AOI22_X1 U9383 ( .A1(n9721), .A2(n9353), .B1(n9545), .B2(n9720), .ZN(n7794)
         );
  NAND2_X1 U9384 ( .A1(n7795), .A2(n7794), .ZN(n7796) );
  AOI21_X1 U9385 ( .B1(n9601), .B2(n9549), .A(n7796), .ZN(n9603) );
  AOI21_X1 U9386 ( .B1(n7797), .B2(n9597), .A(n9767), .ZN(n7798) );
  NAND2_X1 U9387 ( .A1(n7798), .A2(n9378), .ZN(n9598) );
  INV_X1 U9388 ( .A(n9557), .ZN(n9362) );
  AOI22_X1 U9389 ( .A1(n9743), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7839), .B2(
        n9728), .ZN(n7800) );
  NAND2_X1 U9390 ( .A1(n9551), .A2(n9597), .ZN(n7799) );
  OAI211_X1 U9391 ( .C1(n9598), .C2(n9362), .A(n7800), .B(n7799), .ZN(n7801)
         );
  AOI21_X1 U9392 ( .B1(n9601), .B2(n9558), .A(n7801), .ZN(n7802) );
  OAI21_X1 U9393 ( .B1(n9603), .B2(n9743), .A(n7802), .ZN(P1_U3279) );
  INV_X1 U9394 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7808) );
  NOR2_X1 U9395 ( .A1(n7891), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7888) );
  INV_X1 U9396 ( .A(n7888), .ZN(n7806) );
  OAI21_X1 U9397 ( .B1(n7808), .B2(n7807), .A(n7806), .ZN(n7809) );
  NOR2_X1 U9398 ( .A1(n7810), .A2(n7809), .ZN(n7887) );
  AOI21_X1 U9399 ( .B1(n7810), .B2(n7809), .A(n7887), .ZN(n7821) );
  INV_X1 U9400 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7813) );
  MUX2_X1 U9401 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7813), .S(n7891), .Z(n7814)
         );
  OAI21_X1 U9402 ( .B1(n7815), .B2(n7814), .A(n7890), .ZN(n7816) );
  NAND2_X1 U9403 ( .A1(n7816), .A2(n9783), .ZN(n7820) );
  INV_X1 U9404 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7817) );
  NAND2_X1 U9405 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8279) );
  OAI21_X1 U9406 ( .B1(n8527), .B2(n7817), .A(n8279), .ZN(n7818) );
  AOI21_X1 U9407 ( .B1(n8529), .B2(n7891), .A(n7818), .ZN(n7819) );
  OAI211_X1 U9408 ( .C1(n7821), .C2(n9788), .A(n7820), .B(n7819), .ZN(P2_U3259) );
  INV_X1 U9409 ( .A(n7830), .ZN(n8481) );
  AOI21_X1 U9410 ( .B1(n7829), .B2(n7823), .A(n4353), .ZN(n7824) );
  INV_X1 U9411 ( .A(n7824), .ZN(n8897) );
  AOI211_X1 U9412 ( .C1(n8894), .C2(n7825), .A(n9943), .B(n4347), .ZN(n8893)
         );
  INV_X1 U9413 ( .A(n8894), .ZN(n8410) );
  AOI22_X1 U9414 ( .A1(n9831), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8403), .B2(
        n9821), .ZN(n7826) );
  OAI21_X1 U9415 ( .B1(n8410), .B2(n8795), .A(n7826), .ZN(n7833) );
  OAI21_X1 U9416 ( .B1(n7829), .B2(n7828), .A(n7827), .ZN(n7831) );
  OAI22_X1 U9417 ( .A1(n7830), .A2(n8277), .B1(n8479), .B2(n8765), .ZN(n8407)
         );
  AOI21_X1 U9418 ( .B1(n7831), .B2(n9803), .A(n8407), .ZN(n8896) );
  NOR2_X1 U9419 ( .A1(n8896), .A2(n9831), .ZN(n7832) );
  AOI211_X1 U9420 ( .C1(n8893), .C2(n9812), .A(n7833), .B(n7832), .ZN(n7834)
         );
  OAI21_X1 U9421 ( .B1(n8897), .B2(n8808), .A(n7834), .ZN(P2_U3283) );
  INV_X1 U9422 ( .A(n7872), .ZN(n7837) );
  AOI21_X1 U9423 ( .B1(n7838), .B2(n4348), .A(n7837), .ZN(n7846) );
  INV_X1 U9424 ( .A(n9353), .ZN(n7967) );
  NAND2_X1 U9425 ( .A1(n9031), .A2(n7839), .ZN(n7843) );
  INV_X1 U9426 ( .A(n7840), .ZN(n7841) );
  AOI21_X1 U9427 ( .B1(n9033), .B2(n9545), .A(n7841), .ZN(n7842) );
  OAI211_X1 U9428 ( .C1(n7967), .C2(n9036), .A(n7843), .B(n7842), .ZN(n7844)
         );
  AOI21_X1 U9429 ( .B1(n9038), .B2(n9597), .A(n7844), .ZN(n7845) );
  OAI21_X1 U9430 ( .B1(n7846), .B2(n4371), .A(n7845), .ZN(P1_U3222) );
  INV_X1 U9431 ( .A(n7847), .ZN(n7851) );
  OAI222_X1 U9432 ( .A1(P2_U3152), .A2(n7849), .B1(n8920), .B2(n7851), .C1(
        n7848), .C2(n8259), .ZN(P2_U3333) );
  OAI222_X1 U9433 ( .A1(n9524), .A2(n7852), .B1(n9527), .B2(n7851), .C1(n7850), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9434 ( .A(n7853), .ZN(n7855) );
  NAND2_X1 U9435 ( .A1(n7855), .A2(n7854), .ZN(n7857) );
  XNOR2_X1 U9436 ( .A(n7857), .B(n7856), .ZN(n7864) );
  NAND2_X1 U9437 ( .A1(n9031), .A2(n9358), .ZN(n7861) );
  INV_X1 U9438 ( .A(n7858), .ZN(n7859) );
  AOI21_X1 U9439 ( .B1(n9033), .B2(n9353), .A(n7859), .ZN(n7860) );
  OAI211_X1 U9440 ( .C1(n9319), .C2(n9036), .A(n7861), .B(n7860), .ZN(n7862)
         );
  AOI21_X1 U9441 ( .B1(n9359), .B2(n9038), .A(n7862), .ZN(n7863) );
  OAI21_X1 U9442 ( .B1(n7864), .B2(n4371), .A(n7863), .ZN(P1_U3213) );
  INV_X1 U9443 ( .A(n7865), .ZN(n7869) );
  OAI222_X1 U9444 ( .A1(n9527), .A2(n7869), .B1(P1_U3084), .B2(n7867), .C1(
        n7866), .C2(n9524), .ZN(P1_U3327) );
  OAI222_X1 U9445 ( .A1(n7870), .A2(P2_U3152), .B1(n8920), .B2(n7869), .C1(
        n7868), .C2(n8259), .ZN(P2_U3332) );
  NAND2_X1 U9446 ( .A1(n7872), .A2(n7871), .ZN(n7876) );
  NAND2_X1 U9447 ( .A1(n7874), .A2(n7873), .ZN(n7875) );
  XNOR2_X1 U9448 ( .A(n7876), .B(n7875), .ZN(n7883) );
  NAND2_X1 U9449 ( .A1(n9031), .A2(n9381), .ZN(n7880) );
  INV_X1 U9450 ( .A(n7877), .ZN(n7878) );
  AOI21_X1 U9451 ( .B1(n9033), .B2(n9374), .A(n7878), .ZN(n7879) );
  OAI211_X1 U9452 ( .C1(n9331), .C2(n9036), .A(n7880), .B(n7879), .ZN(n7881)
         );
  AOI21_X1 U9453 ( .B1(n9038), .B2(n9470), .A(n7881), .ZN(n7882) );
  OAI21_X1 U9454 ( .B1(n7883), .B2(n4371), .A(n7882), .ZN(P1_U3232) );
  INV_X1 U9455 ( .A(n7884), .ZN(n7902) );
  AOI21_X1 U9456 ( .B1(n9520), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7885), .ZN(
        n7886) );
  OAI21_X1 U9457 ( .B1(n7902), .B2(n9522), .A(n7886), .ZN(P1_U3326) );
  XNOR2_X1 U9458 ( .A(n7911), .B(n7910), .ZN(n7889) );
  NOR2_X1 U9459 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7889), .ZN(n7912) );
  AOI21_X1 U9460 ( .B1(n7889), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7912), .ZN(
        n7900) );
  INV_X1 U9461 ( .A(n7892), .ZN(n7895) );
  NOR2_X1 U9462 ( .A1(n7893), .A2(n7892), .ZN(n7922) );
  INV_X1 U9463 ( .A(n7922), .ZN(n7894) );
  OAI211_X1 U9464 ( .C1(n7895), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9783), .B(
        n7894), .ZN(n7899) );
  NOR2_X1 U9465 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5294), .ZN(n7897) );
  NOR2_X1 U9466 ( .A1(n9786), .A2(n7921), .ZN(n7896) );
  AOI211_X1 U9467 ( .C1(n9785), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n7897), .B(
        n7896), .ZN(n7898) );
  OAI211_X1 U9468 ( .C1(n7900), .C2(n9788), .A(n7899), .B(n7898), .ZN(P2_U3260) );
  OAI222_X1 U9469 ( .A1(P2_U3152), .A2(n5832), .B1(n8920), .B2(n7902), .C1(
        n7901), .C2(n8259), .ZN(P2_U3331) );
  INV_X1 U9470 ( .A(n7903), .ZN(n8243) );
  AOI21_X1 U9471 ( .B1(n9520), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n7904), .ZN(
        n7905) );
  OAI21_X1 U9472 ( .B1(n8243), .B2(n9522), .A(n7905), .ZN(P1_U3325) );
  INV_X1 U9473 ( .A(n7947), .ZN(n9526) );
  OAI222_X1 U9474 ( .A1(P2_U3152), .A2(n7906), .B1(n8920), .B2(n9526), .C1(
        n7907), .C2(n8259), .ZN(P2_U3329) );
  NAND2_X1 U9475 ( .A1(n7924), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7915) );
  XOR2_X1 U9476 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n7924), .Z(n8509) );
  NAND2_X1 U9477 ( .A1(n8503), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7914) );
  INV_X1 U9478 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7908) );
  MUX2_X1 U9479 ( .A(n7908), .B(P2_REG2_REG_16__SCAN_IN), .S(n8503), .Z(n7909)
         );
  INV_X1 U9480 ( .A(n7909), .ZN(n8501) );
  NOR2_X1 U9481 ( .A1(n7911), .A2(n7910), .ZN(n7913) );
  NAND2_X1 U9482 ( .A1(n8501), .A2(n8502), .ZN(n8500) );
  NAND2_X1 U9483 ( .A1(n7914), .A2(n8500), .ZN(n8510) );
  NAND2_X1 U9484 ( .A1(n8509), .A2(n8510), .ZN(n8508) );
  NAND2_X1 U9485 ( .A1(n7915), .A2(n8508), .ZN(n7916) );
  NOR2_X1 U9486 ( .A1(n7916), .A2(n8530), .ZN(n7917) );
  NOR2_X1 U9487 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8520), .ZN(n8519) );
  NOR2_X1 U9488 ( .A1(n8519), .A2(n7917), .ZN(n7918) );
  XOR2_X1 U9489 ( .A(n7918), .B(P2_REG2_REG_19__SCAN_IN), .Z(n7928) );
  INV_X1 U9490 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7919) );
  XNOR2_X1 U9491 ( .A(n8530), .B(n7919), .ZN(n8522) );
  XNOR2_X1 U9492 ( .A(n7924), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8512) );
  XOR2_X1 U9493 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8503), .Z(n8495) );
  NOR2_X1 U9494 ( .A1(n7921), .A2(n7920), .ZN(n7923) );
  NOR2_X1 U9495 ( .A1(n7923), .A2(n7922), .ZN(n8496) );
  NAND2_X1 U9496 ( .A1(n8495), .A2(n8496), .ZN(n8494) );
  NOR2_X1 U9497 ( .A1(n8530), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7925) );
  XNOR2_X1 U9498 ( .A(n7926), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n7930) );
  INV_X1 U9499 ( .A(n7930), .ZN(n7927) );
  AOI22_X1 U9500 ( .A1(n7928), .A2(n9784), .B1(n7927), .B2(n9783), .ZN(n7932)
         );
  NOR2_X1 U9501 ( .A1(n7928), .A2(n9788), .ZN(n7929) );
  AOI211_X1 U9502 ( .C1(n9783), .C2(n7930), .A(n8529), .B(n7929), .ZN(n7931)
         );
  MUX2_X1 U9503 ( .A(n7932), .B(n7931), .S(n9823), .Z(n7934) );
  NAND2_X1 U9504 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n7933) );
  OAI211_X1 U9505 ( .C1(n7661), .C2(n8527), .A(n7934), .B(n7933), .ZN(P2_U3264) );
  NAND2_X1 U9506 ( .A1(n7935), .A2(n6082), .ZN(n7937) );
  NAND2_X1 U9507 ( .A1(n7939), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7936) );
  INV_X1 U9508 ( .A(n9113), .ZN(n7938) );
  AND2_X1 U9509 ( .A1(n8015), .A2(n7938), .ZN(n8058) );
  NAND2_X1 U9510 ( .A1(n8244), .A2(n6082), .ZN(n7941) );
  NAND2_X1 U9511 ( .A1(n7939), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7940) );
  INV_X1 U9512 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U9513 ( .A1(n7942), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U9514 ( .A1(n5941), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7943) );
  OAI211_X1 U9515 ( .C1(n5989), .C2(n7945), .A(n7944), .B(n7943), .ZN(n9041)
         );
  INV_X1 U9516 ( .A(n9041), .ZN(n7946) );
  NOR2_X1 U9517 ( .A1(n9118), .A2(n7946), .ZN(n8040) );
  NOR2_X1 U9518 ( .A1(n8058), .A2(n8040), .ZN(n8038) );
  AND2_X1 U9519 ( .A1(n9118), .A2(n7946), .ZN(n8037) );
  INV_X1 U9520 ( .A(n8037), .ZN(n8014) );
  NAND2_X1 U9521 ( .A1(n7947), .A2(n6082), .ZN(n7949) );
  NAND2_X1 U9522 ( .A1(n7939), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U9523 ( .A1(n9396), .A2(n9131), .ZN(n8160) );
  OR2_X1 U9524 ( .A1(n9410), .A2(n8198), .ZN(n8062) );
  NAND2_X1 U9525 ( .A1(n8062), .A2(n9168), .ZN(n8229) );
  AND2_X1 U9526 ( .A1(n4576), .A2(n8149), .ZN(n8050) );
  NAND2_X1 U9527 ( .A1(n9401), .A2(n9152), .ZN(n8231) );
  NAND2_X1 U9528 ( .A1(n9405), .A2(n9130), .ZN(n8060) );
  AND2_X1 U9529 ( .A1(n8231), .A2(n8060), .ZN(n8150) );
  INV_X1 U9530 ( .A(n8150), .ZN(n7952) );
  NAND2_X1 U9531 ( .A1(n9410), .A2(n8198), .ZN(n8228) );
  INV_X1 U9532 ( .A(n8228), .ZN(n7950) );
  AND2_X1 U9533 ( .A1(n8149), .A2(n7950), .ZN(n7951) );
  OR2_X1 U9534 ( .A1(n7952), .A2(n7951), .ZN(n8048) );
  NAND2_X1 U9535 ( .A1(n8159), .A2(n8152), .ZN(n8052) );
  INV_X1 U9536 ( .A(n8052), .ZN(n8012) );
  NAND2_X1 U9537 ( .A1(n9425), .A2(n8197), .ZN(n8133) );
  INV_X1 U9538 ( .A(n8019), .ZN(n8219) );
  AND2_X1 U9539 ( .A1(n8133), .A2(n8219), .ZN(n7955) );
  NAND2_X1 U9540 ( .A1(n9430), .A2(n9244), .ZN(n8018) );
  NAND2_X1 U9541 ( .A1(n9437), .A2(n9259), .ZN(n8222) );
  NAND2_X1 U9542 ( .A1(n8018), .A2(n8222), .ZN(n8066) );
  INV_X1 U9543 ( .A(n9276), .ZN(n9245) );
  AND2_X1 U9544 ( .A1(n9442), .A2(n9245), .ZN(n8221) );
  AND2_X1 U9545 ( .A1(n8123), .A2(n8221), .ZN(n7953) );
  OR2_X1 U9546 ( .A1(n8066), .A2(n7953), .ZN(n8129) );
  INV_X1 U9547 ( .A(n8129), .ZN(n7954) );
  NAND2_X1 U9548 ( .A1(n7955), .A2(n7954), .ZN(n8045) );
  NAND2_X1 U9549 ( .A1(n9450), .A2(n8941), .ZN(n8217) );
  NAND2_X1 U9550 ( .A1(n9455), .A2(n9320), .ZN(n9291) );
  AND2_X1 U9551 ( .A1(n8217), .A2(n9291), .ZN(n8218) );
  NAND2_X1 U9552 ( .A1(n9462), .A2(n9329), .ZN(n8213) );
  NAND2_X1 U9553 ( .A1(n9359), .A2(n9331), .ZN(n7969) );
  NAND2_X1 U9554 ( .A1(n9470), .A2(n7967), .ZN(n8209) );
  NAND2_X1 U9555 ( .A1(n7969), .A2(n8209), .ZN(n8102) );
  INV_X1 U9556 ( .A(n8078), .ZN(n7956) );
  OR2_X1 U9557 ( .A1(n7956), .A2(n8075), .ZN(n7958) );
  AND2_X1 U9558 ( .A1(n7958), .A2(n7957), .ZN(n8082) );
  INV_X1 U9559 ( .A(n8082), .ZN(n7964) );
  AND2_X1 U9560 ( .A1(n8073), .A2(n8068), .ZN(n8080) );
  NAND4_X1 U9561 ( .A1(n7964), .A2(n8091), .A3(n8080), .A4(n8090), .ZN(n7959)
         );
  NOR2_X1 U9562 ( .A1(n8102), .A2(n7959), .ZN(n7960) );
  NAND2_X1 U9563 ( .A1(n9465), .A2(n9319), .ZN(n8212) );
  AND3_X1 U9564 ( .A1(n8213), .A2(n7960), .A3(n8212), .ZN(n7961) );
  NAND2_X1 U9565 ( .A1(n8218), .A2(n7961), .ZN(n8044) );
  AND2_X1 U9566 ( .A1(n9342), .A2(n9354), .ZN(n8211) );
  AND2_X1 U9567 ( .A1(n8074), .A2(n7962), .ZN(n8083) );
  INV_X1 U9568 ( .A(n8083), .ZN(n7963) );
  AND3_X1 U9569 ( .A1(n7964), .A2(n8090), .A3(n7963), .ZN(n7966) );
  NAND2_X1 U9570 ( .A1(n8092), .A2(n7965), .ZN(n8088) );
  OAI21_X1 U9571 ( .B1(n7966), .B2(n8088), .A(n8091), .ZN(n7972) );
  OR2_X1 U9572 ( .A1(n9470), .A2(n7967), .ZN(n8089) );
  INV_X1 U9573 ( .A(n8089), .ZN(n7968) );
  NAND2_X1 U9574 ( .A1(n7969), .A2(n7968), .ZN(n7970) );
  OR2_X1 U9575 ( .A1(n9359), .A2(n9331), .ZN(n8210) );
  NAND2_X1 U9576 ( .A1(n7970), .A2(n8210), .ZN(n8101) );
  INV_X1 U9577 ( .A(n8101), .ZN(n7971) );
  OAI21_X1 U9578 ( .B1(n8102), .B2(n7972), .A(n7971), .ZN(n7973) );
  NAND2_X1 U9579 ( .A1(n7973), .A2(n8212), .ZN(n7974) );
  NAND3_X1 U9580 ( .A1(n8215), .A2(n4580), .A3(n7974), .ZN(n7975) );
  NAND3_X1 U9581 ( .A1(n8218), .A2(n8213), .A3(n7975), .ZN(n7976) );
  OAI21_X1 U9582 ( .B1(n8044), .B2(n8071), .A(n7976), .ZN(n7977) );
  INV_X1 U9583 ( .A(n7977), .ZN(n7978) );
  OR2_X1 U9584 ( .A1(n8045), .A2(n7978), .ZN(n7985) );
  OR2_X1 U9585 ( .A1(n9450), .A2(n8941), .ZN(n8115) );
  OR2_X1 U9586 ( .A1(n9455), .A2(n9320), .ZN(n9289) );
  NAND2_X1 U9587 ( .A1(n8115), .A2(n9289), .ZN(n8216) );
  INV_X1 U9588 ( .A(n8216), .ZN(n8111) );
  INV_X1 U9589 ( .A(n8217), .ZN(n7979) );
  NOR2_X1 U9590 ( .A1(n8019), .A2(n7979), .ZN(n8126) );
  INV_X1 U9591 ( .A(n8126), .ZN(n7980) );
  NOR2_X1 U9592 ( .A1(n9446), .A2(n9258), .ZN(n8020) );
  INV_X1 U9593 ( .A(n8020), .ZN(n8114) );
  AND2_X1 U9594 ( .A1(n8220), .A2(n8114), .ZN(n8122) );
  OAI211_X1 U9595 ( .C1(n8111), .C2(n7980), .A(n8123), .B(n8122), .ZN(n7981)
         );
  INV_X1 U9596 ( .A(n7981), .ZN(n7982) );
  OAI21_X1 U9597 ( .B1(n8129), .B2(n7982), .A(n8127), .ZN(n7983) );
  NAND2_X1 U9598 ( .A1(n7983), .A2(n8133), .ZN(n7984) );
  NAND4_X1 U9599 ( .A1(n7985), .A2(n7984), .A3(n8224), .A4(n8137), .ZN(n8047)
         );
  INV_X1 U9600 ( .A(n8067), .ZN(n8007) );
  INV_X1 U9601 ( .A(n9730), .ZN(n7986) );
  NAND2_X1 U9602 ( .A1(n6544), .A2(n7986), .ZN(n7987) );
  NAND3_X1 U9603 ( .A1(n7988), .A2(n8172), .A3(n7987), .ZN(n7990) );
  NAND2_X1 U9604 ( .A1(n7990), .A2(n7989), .ZN(n7993) );
  OAI211_X1 U9605 ( .C1(n7994), .C2(n7993), .A(n7992), .B(n7991), .ZN(n7996)
         );
  NAND2_X1 U9606 ( .A1(n7996), .A2(n7995), .ZN(n7998) );
  NAND2_X1 U9607 ( .A1(n7998), .A2(n7997), .ZN(n8005) );
  INV_X1 U9608 ( .A(n7999), .ZN(n8001) );
  NOR2_X1 U9609 ( .A1(n8001), .A2(n8000), .ZN(n8004) );
  INV_X1 U9610 ( .A(n8002), .ZN(n8003) );
  AOI21_X1 U9611 ( .B1(n8005), .B2(n8004), .A(n8003), .ZN(n8006) );
  OR3_X1 U9612 ( .A1(n8044), .A2(n8007), .A3(n8006), .ZN(n8008) );
  NOR2_X1 U9613 ( .A1(n8045), .A2(n8008), .ZN(n8009) );
  NAND2_X1 U9614 ( .A1(n9415), .A2(n9044), .ZN(n8063) );
  NAND2_X1 U9615 ( .A1(n9421), .A2(n8957), .ZN(n8136) );
  NAND2_X1 U9616 ( .A1(n8063), .A2(n8136), .ZN(n8227) );
  OAI21_X1 U9617 ( .B1(n8047), .B2(n8009), .A(n4577), .ZN(n8010) );
  OR2_X1 U9618 ( .A1(n8048), .A2(n8010), .ZN(n8011) );
  OAI211_X1 U9619 ( .C1(n8050), .C2(n8048), .A(n8012), .B(n8011), .ZN(n8013)
         );
  NAND3_X1 U9620 ( .A1(n8014), .A2(n8160), .A3(n8013), .ZN(n8016) );
  AOI21_X1 U9621 ( .B1(n8038), .B2(n8016), .A(n8170), .ZN(n8017) );
  XNOR2_X1 U9622 ( .A(n8017), .B(n9204), .ZN(n8176) );
  NAND2_X1 U9623 ( .A1(n8152), .A2(n8231), .ZN(n9124) );
  INV_X1 U9624 ( .A(n9124), .ZN(n9128) );
  NAND2_X1 U9625 ( .A1(n9168), .A2(n8063), .ZN(n9184) );
  NAND2_X1 U9626 ( .A1(n8137), .A2(n8136), .ZN(n9194) );
  NAND2_X1 U9627 ( .A1(n8224), .A2(n8133), .ZN(n9216) );
  NAND2_X1 U9628 ( .A1(n8127), .A2(n8018), .ZN(n9232) );
  NAND2_X1 U9629 ( .A1(n8123), .A2(n8222), .ZN(n9242) );
  INV_X1 U9630 ( .A(n8221), .ZN(n8116) );
  NAND2_X1 U9631 ( .A1(n8116), .A2(n8220), .ZN(n9255) );
  NOR2_X1 U9632 ( .A1(n8020), .A2(n8019), .ZN(n9275) );
  NAND2_X1 U9633 ( .A1(n8115), .A2(n8217), .ZN(n9281) );
  INV_X1 U9634 ( .A(n9281), .ZN(n9292) );
  NAND2_X1 U9635 ( .A1(n8215), .A2(n8213), .ZN(n9315) );
  INV_X1 U9636 ( .A(n8212), .ZN(n8021) );
  NAND2_X1 U9637 ( .A1(n8089), .A2(n8209), .ZN(n9368) );
  NOR3_X1 U9638 ( .A1(n8023), .A2(n7148), .A3(n8022), .ZN(n8025) );
  NOR4_X1 U9639 ( .A1(n8027), .A2(n7151), .A3(n8026), .A4(n8069), .ZN(n8031)
         );
  INV_X1 U9640 ( .A(n9543), .ZN(n8030) );
  NAND4_X1 U9641 ( .A1(n8031), .A2(n8030), .A3(n8029), .A4(n8028), .ZN(n8032)
         );
  OR4_X1 U9642 ( .A1(n9368), .A2(n8033), .A3(n8032), .A4(n8183), .ZN(n8034) );
  XNOR2_X1 U9643 ( .A(n9359), .B(n9331), .ZN(n9349) );
  XNOR2_X1 U9644 ( .A(n9167), .B(n9186), .ZN(n9161) );
  INV_X1 U9645 ( .A(n9161), .ZN(n9171) );
  NAND4_X1 U9646 ( .A1(n9128), .A2(n4570), .A3(n8035), .A4(n9171), .ZN(n8036)
         );
  AOI21_X1 U9647 ( .B1(n8039), .B2(n8038), .A(n8172), .ZN(n8168) );
  INV_X1 U9648 ( .A(n8168), .ZN(n8057) );
  INV_X1 U9649 ( .A(n8040), .ZN(n8041) );
  NAND2_X1 U9650 ( .A1(n8041), .A2(n9113), .ZN(n8042) );
  NAND2_X1 U9651 ( .A1(n8042), .A2(n8015), .ZN(n8163) );
  NOR3_X1 U9652 ( .A1(n8045), .A2(n8044), .A3(n8043), .ZN(n8046) );
  OAI21_X1 U9653 ( .B1(n8047), .B2(n8046), .A(n4577), .ZN(n8049) );
  AOI21_X1 U9654 ( .B1(n8050), .B2(n8049), .A(n8048), .ZN(n8053) );
  NAND2_X1 U9655 ( .A1(n9041), .A2(n9113), .ZN(n8051) );
  OAI211_X1 U9656 ( .C1(n8053), .C2(n8052), .A(n4304), .B(n8160), .ZN(n8055)
         );
  AOI211_X1 U9657 ( .C1(n8163), .C2(n8055), .A(n8054), .B(n8170), .ZN(n8056)
         );
  AND2_X1 U9658 ( .A1(n8060), .A2(n8228), .ZN(n8061) );
  INV_X1 U9659 ( .A(n8158), .ZN(n8100) );
  MUX2_X1 U9660 ( .A(n8062), .B(n8061), .S(n8100), .Z(n8147) );
  NAND2_X1 U9661 ( .A1(n8228), .A2(n8063), .ZN(n8064) );
  MUX2_X1 U9662 ( .A(n8064), .B(n8229), .S(n8100), .Z(n8065) );
  INV_X1 U9663 ( .A(n8065), .ZN(n8145) );
  INV_X1 U9664 ( .A(n8066), .ZN(n8120) );
  OAI211_X1 U9665 ( .C1(n8070), .C2(n8069), .A(n8068), .B(n8067), .ZN(n8072)
         );
  NAND3_X1 U9666 ( .A1(n8072), .A2(n8083), .A3(n8071), .ZN(n8079) );
  INV_X1 U9667 ( .A(n8073), .ZN(n8076) );
  OAI21_X1 U9668 ( .B1(n8076), .B2(n8075), .A(n8074), .ZN(n8077) );
  NAND4_X1 U9669 ( .A1(n8079), .A2(n8091), .A3(n8078), .A4(n8077), .ZN(n8086)
         );
  NAND2_X1 U9670 ( .A1(n8081), .A2(n8080), .ZN(n8084) );
  AOI21_X1 U9671 ( .B1(n8084), .B2(n8083), .A(n8082), .ZN(n8085) );
  MUX2_X1 U9672 ( .A(n8086), .B(n8085), .S(n8100), .Z(n8098) );
  NAND2_X1 U9673 ( .A1(n8092), .A2(n8087), .ZN(n8097) );
  NAND2_X1 U9674 ( .A1(n8210), .A2(n8158), .ZN(n8099) );
  NAND2_X1 U9675 ( .A1(n8088), .A2(n8091), .ZN(n8206) );
  NAND2_X1 U9676 ( .A1(n8206), .A2(n8089), .ZN(n8095) );
  NAND2_X1 U9677 ( .A1(n8091), .A2(n8090), .ZN(n8207) );
  AND2_X1 U9678 ( .A1(n8207), .A2(n8092), .ZN(n8093) );
  OR3_X1 U9679 ( .A1(n8102), .A2(n8093), .A3(n8158), .ZN(n8094) );
  OAI21_X1 U9680 ( .B1(n8099), .B2(n8095), .A(n8094), .ZN(n8096) );
  OAI21_X1 U9681 ( .B1(n8098), .B2(n8097), .A(n8096), .ZN(n8106) );
  INV_X1 U9682 ( .A(n9332), .ZN(n8105) );
  INV_X1 U9683 ( .A(n8099), .ZN(n8103) );
  AOI22_X1 U9684 ( .A1(n8103), .A2(n8102), .B1(n8101), .B2(n8100), .ZN(n8104)
         );
  NAND3_X1 U9685 ( .A1(n8106), .A2(n8105), .A3(n8104), .ZN(n8108) );
  MUX2_X1 U9686 ( .A(n8212), .B(n4580), .S(n8158), .Z(n8107) );
  NAND3_X1 U9687 ( .A1(n8108), .A2(n4814), .A3(n8107), .ZN(n8110) );
  MUX2_X1 U9688 ( .A(n8215), .B(n8213), .S(n8158), .Z(n8109) );
  NAND3_X1 U9689 ( .A1(n8110), .A2(n9307), .A3(n8109), .ZN(n8113) );
  MUX2_X1 U9690 ( .A(n8218), .B(n8111), .S(n8158), .Z(n8112) );
  NAND2_X1 U9691 ( .A1(n8113), .A2(n8112), .ZN(n8125) );
  NAND3_X1 U9692 ( .A1(n8125), .A2(n8115), .A3(n8114), .ZN(n8117) );
  NAND3_X1 U9693 ( .A1(n8117), .A2(n8116), .A3(n8219), .ZN(n8118) );
  NAND3_X1 U9694 ( .A1(n8118), .A2(n8123), .A3(n8220), .ZN(n8119) );
  INV_X1 U9695 ( .A(n8127), .ZN(n8223) );
  AOI21_X1 U9696 ( .B1(n8120), .B2(n8119), .A(n8223), .ZN(n8121) );
  NAND2_X1 U9697 ( .A1(n8137), .A2(n8121), .ZN(n8132) );
  NAND2_X1 U9698 ( .A1(n8123), .A2(n8122), .ZN(n8124) );
  AOI21_X1 U9699 ( .B1(n8126), .B2(n8125), .A(n8124), .ZN(n8128) );
  OAI21_X1 U9700 ( .B1(n8129), .B2(n8128), .A(n8127), .ZN(n8130) );
  NAND2_X1 U9701 ( .A1(n8130), .A2(n8133), .ZN(n8131) );
  MUX2_X1 U9702 ( .A(n8132), .B(n8131), .S(n8158), .Z(n8143) );
  NAND2_X1 U9703 ( .A1(n8136), .A2(n8224), .ZN(n8142) );
  INV_X1 U9704 ( .A(n8133), .ZN(n8134) );
  AND2_X1 U9705 ( .A1(n8137), .A2(n8134), .ZN(n8135) );
  NOR2_X1 U9706 ( .A1(n8227), .A2(n8135), .ZN(n8140) );
  INV_X1 U9707 ( .A(n8136), .ZN(n9183) );
  OAI211_X1 U9708 ( .C1(n9183), .C2(n8224), .A(n9168), .B(n8137), .ZN(n8138)
         );
  INV_X1 U9709 ( .A(n8138), .ZN(n8139) );
  MUX2_X1 U9710 ( .A(n8140), .B(n8139), .S(n8158), .Z(n8141) );
  OAI21_X1 U9711 ( .B1(n8143), .B2(n8142), .A(n8141), .ZN(n8144) );
  NAND2_X1 U9712 ( .A1(n8145), .A2(n8144), .ZN(n8146) );
  NAND2_X1 U9713 ( .A1(n8147), .A2(n8146), .ZN(n8151) );
  NAND3_X1 U9714 ( .A1(n8151), .A2(n8149), .A3(n8152), .ZN(n8148) );
  NAND2_X1 U9715 ( .A1(n8148), .A2(n8231), .ZN(n8155) );
  INV_X1 U9716 ( .A(n8149), .ZN(n8230) );
  OAI21_X1 U9717 ( .B1(n8151), .B2(n8230), .A(n8150), .ZN(n8153) );
  NAND2_X1 U9718 ( .A1(n8153), .A2(n8152), .ZN(n8154) );
  MUX2_X1 U9719 ( .A(n8155), .B(n8154), .S(n8158), .Z(n8157) );
  INV_X1 U9720 ( .A(n8232), .ZN(n8156) );
  NAND2_X1 U9721 ( .A1(n8157), .A2(n8156), .ZN(n8162) );
  MUX2_X1 U9722 ( .A(n8160), .B(n8159), .S(n8158), .Z(n8161) );
  NAND4_X1 U9723 ( .A1(n8163), .A2(n8162), .A3(n8161), .A4(n4304), .ZN(n8164)
         );
  NAND2_X1 U9724 ( .A1(n8165), .A2(n8164), .ZN(n8173) );
  NOR3_X1 U9725 ( .A1(n8173), .A2(n8170), .A3(n8166), .ZN(n8167) );
  NOR2_X1 U9726 ( .A1(n8168), .A2(n8167), .ZN(n8169) );
  INV_X1 U9727 ( .A(n8170), .ZN(n8171) );
  NAND4_X1 U9728 ( .A1(n8173), .A2(n8172), .A3(n8171), .A4(n6455), .ZN(n8174)
         );
  NOR4_X1 U9729 ( .A1(n8178), .A2(n8177), .A3(n9624), .A4(n9620), .ZN(n8180)
         );
  OAI21_X1 U9730 ( .B1(n6478), .B2(n8181), .A(P1_B_REG_SCAN_IN), .ZN(n8179) );
  OAI22_X1 U9731 ( .A1(n8182), .A2(n8181), .B1(n8180), .B2(n8179), .ZN(
        P1_U3240) );
  NAND2_X1 U9732 ( .A1(n9597), .A2(n9374), .ZN(n8185) );
  OR2_X1 U9733 ( .A1(n9470), .A2(n9353), .ZN(n8187) );
  AND2_X1 U9734 ( .A1(n9470), .A2(n9353), .ZN(n8186) );
  NAND2_X1 U9735 ( .A1(n9359), .A2(n9373), .ZN(n8189) );
  NOR2_X1 U9736 ( .A1(n9359), .A2(n9373), .ZN(n8188) );
  NOR2_X1 U9737 ( .A1(n9455), .A2(n9294), .ZN(n8191) );
  AOI22_X1 U9738 ( .A1(n9282), .A2(n9281), .B1(n9309), .B2(n9450), .ZN(n9267)
         );
  NAND2_X1 U9739 ( .A1(n9446), .A2(n9295), .ZN(n8192) );
  AOI22_X1 U9740 ( .A1(n9267), .A2(n8192), .B1(n9258), .B2(n9272), .ZN(n9254)
         );
  NAND2_X1 U9741 ( .A1(n9254), .A2(n8193), .ZN(n8194) );
  INV_X1 U9742 ( .A(n9442), .ZN(n9264) );
  NAND2_X1 U9743 ( .A1(n8194), .A2(n4828), .ZN(n9240) );
  AOI22_X1 U9744 ( .A1(n9240), .A2(n9242), .B1(n9437), .B2(n9235), .ZN(n9223)
         );
  NAND2_X1 U9745 ( .A1(n9430), .A2(n9217), .ZN(n8195) );
  OAI21_X1 U9746 ( .B1(n9425), .B2(n9234), .A(n9209), .ZN(n8196) );
  NAND2_X1 U9747 ( .A1(n9125), .A2(n9124), .ZN(n9123) );
  NAND2_X1 U9748 ( .A1(n9401), .A2(n9043), .ZN(n8199) );
  NAND2_X1 U9749 ( .A1(n9123), .A2(n8199), .ZN(n8200) );
  XNOR2_X1 U9750 ( .A(n8200), .B(n8232), .ZN(n9399) );
  INV_X1 U9751 ( .A(n9359), .ZN(n9592) );
  NAND2_X1 U9752 ( .A1(n9301), .A2(n9288), .ZN(n9283) );
  AND2_X2 U9753 ( .A1(n9179), .A2(n9167), .ZN(n9163) );
  AND2_X2 U9754 ( .A1(n9163), .A2(n9151), .ZN(n9147) );
  AOI211_X1 U9755 ( .C1(n9396), .C2(n9137), .A(n9767), .B(n9117), .ZN(n9395)
         );
  INV_X1 U9756 ( .A(n8202), .ZN(n8203) );
  AOI22_X1 U9757 ( .A1(n8203), .A2(n9728), .B1(n9743), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n8204) );
  OAI21_X1 U9758 ( .B1(n4440), .B2(n9341), .A(n8204), .ZN(n8205) );
  AOI21_X1 U9759 ( .B1(n9395), .B2(n9557), .A(n8205), .ZN(n8241) );
  INV_X1 U9760 ( .A(n8213), .ZN(n8214) );
  NAND2_X1 U9761 ( .A1(n9274), .A2(n9275), .ZN(n9273) );
  NAND2_X1 U9762 ( .A1(n9273), .A2(n8219), .ZN(n9256) );
  INV_X1 U9763 ( .A(n8222), .ZN(n9231) );
  NOR2_X1 U9764 ( .A1(n9215), .A2(n9216), .ZN(n9196) );
  INV_X1 U9765 ( .A(n9194), .ZN(n8225) );
  INV_X1 U9766 ( .A(n8224), .ZN(n9195) );
  NAND2_X1 U9767 ( .A1(n8225), .A2(n8224), .ZN(n8226) );
  NAND2_X1 U9768 ( .A1(n9127), .A2(n9128), .ZN(n9126) );
  XNOR2_X1 U9769 ( .A(n8233), .B(n8156), .ZN(n8239) );
  INV_X1 U9770 ( .A(P1_B_REG_SCAN_IN), .ZN(n8234) );
  NOR2_X1 U9771 ( .A1(n9620), .A2(n8234), .ZN(n8235) );
  NOR2_X1 U9772 ( .A1(n9328), .A2(n8235), .ZN(n9114) );
  NAND2_X1 U9773 ( .A1(n9114), .A2(n9041), .ZN(n8236) );
  OR2_X1 U9774 ( .A1(n9398), .A2(n9743), .ZN(n8240) );
  OAI211_X1 U9775 ( .C1(n9399), .C2(n9365), .A(n8241), .B(n8240), .ZN(P1_U3355) );
  OAI222_X1 U9776 ( .A1(P2_U3152), .A2(n5576), .B1(n8920), .B2(n8243), .C1(
        n8242), .C2(n8259), .ZN(P2_U3330) );
  INV_X1 U9777 ( .A(n8244), .ZN(n8261) );
  OAI222_X1 U9778 ( .A1(n9524), .A2(n4389), .B1(n9522), .B2(n8261), .C1(
        P1_U3084), .C2(n8245), .ZN(P1_U3323) );
  INV_X1 U9779 ( .A(n8296), .ZN(n8246) );
  AOI211_X1 U9780 ( .C1(n8248), .C2(n8247), .A(n8246), .B(n8445), .ZN(n8249)
         );
  AOI21_X1 U9781 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n8256), .A(n8249), .ZN(
        n8253) );
  AOI22_X1 U9782 ( .A1(n8251), .A2(n8490), .B1(n4267), .B2(n8469), .ZN(n8252)
         );
  OAI211_X1 U9783 ( .C1(n7606), .C2(n8465), .A(n8253), .B(n8252), .ZN(P2_U3239) );
  OAI22_X1 U9784 ( .A1(n8443), .A2(n5659), .B1(n9873), .B2(n8445), .ZN(n8255)
         );
  NAND2_X1 U9785 ( .A1(n8255), .A2(n8254), .ZN(n8258) );
  AOI22_X1 U9786 ( .A1(n8469), .A2(n9874), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8256), .ZN(n8257) );
  OAI211_X1 U9787 ( .C1(n7606), .C2(n8466), .A(n8258), .B(n8257), .ZN(P2_U3234) );
  OAI222_X1 U9788 ( .A1(n8262), .A2(P2_U3152), .B1(n8920), .B2(n8261), .C1(
        n8260), .C2(n8259), .ZN(P2_U3328) );
  INV_X1 U9789 ( .A(n8263), .ZN(n8264) );
  AOI21_X1 U9790 ( .B1(n8448), .B2(n8264), .A(n8445), .ZN(n8268) );
  NOR3_X1 U9791 ( .A1(n8265), .A2(n8563), .A3(n8443), .ZN(n8267) );
  OAI21_X1 U9792 ( .B1(n8268), .B2(n8267), .A(n8266), .ZN(n8273) );
  OAI22_X1 U9793 ( .A1(n8579), .A2(n8765), .B1(n8563), .B2(n8277), .ZN(n8612)
         );
  INV_X1 U9794 ( .A(n8612), .ZN(n8270) );
  OAI22_X1 U9795 ( .A1(n8270), .A2(n8452), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8269), .ZN(n8271) );
  AOI21_X1 U9796 ( .B1(n8607), .B2(n8454), .A(n8271), .ZN(n8272) );
  OAI211_X1 U9797 ( .C1(n8609), .C2(n8458), .A(n8273), .B(n8272), .ZN(P2_U3216) );
  INV_X1 U9798 ( .A(n8400), .ZN(n8276) );
  NOR3_X1 U9799 ( .A1(n8443), .A2(n8480), .A3(n8274), .ZN(n8275) );
  AOI21_X1 U9800 ( .B1(n8276), .B2(n8460), .A(n8275), .ZN(n8286) );
  INV_X1 U9801 ( .A(n9575), .ZN(n8280) );
  OAI22_X1 U9802 ( .A1(n8480), .A2(n8277), .B1(n8546), .B2(n8765), .ZN(n9572)
         );
  NAND2_X1 U9803 ( .A1(n8426), .A2(n9572), .ZN(n8278) );
  OAI211_X1 U9804 ( .C1(n8464), .C2(n8280), .A(n8279), .B(n8278), .ZN(n8283)
         );
  NOR2_X1 U9805 ( .A1(n8281), .A2(n8445), .ZN(n8282) );
  AOI211_X1 U9806 ( .C1(n9576), .C2(n8469), .A(n8283), .B(n8282), .ZN(n8284)
         );
  OAI21_X1 U9807 ( .B1(n8286), .B2(n8285), .A(n8284), .ZN(P2_U3217) );
  INV_X1 U9808 ( .A(n8443), .ZN(n8459) );
  AOI22_X1 U9809 ( .A1(n8287), .A2(n8460), .B1(n8459), .B2(n8695), .ZN(n8293)
         );
  OAI22_X1 U9810 ( .A1(n8464), .A2(n8679), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8289), .ZN(n8291) );
  OAI22_X1 U9811 ( .A1(n8671), .A2(n8465), .B1(n8466), .B2(n8672), .ZN(n8290)
         );
  AOI211_X1 U9812 ( .C1(n8848), .C2(n8469), .A(n8291), .B(n8290), .ZN(n8292)
         );
  OAI21_X1 U9813 ( .B1(n8293), .B2(n8368), .A(n8292), .ZN(P2_U3218) );
  NOR3_X1 U9814 ( .A1(n8443), .A2(n4835), .A3(n8294), .ZN(n8300) );
  INV_X1 U9815 ( .A(n8295), .ZN(n8297) );
  AOI21_X1 U9816 ( .B1(n8297), .B2(n8296), .A(n8445), .ZN(n8299) );
  OAI21_X1 U9817 ( .B1(n8300), .B2(n8299), .A(n8298), .ZN(n8306) );
  AOI22_X1 U9818 ( .A1(n8426), .A2(n8302), .B1(n8469), .B2(n8301), .ZN(n8305)
         );
  MUX2_X1 U9819 ( .A(P2_STATE_REG_SCAN_IN), .B(n8464), .S(n8303), .Z(n8304) );
  NAND3_X1 U9820 ( .A1(n8306), .A2(n8305), .A3(n8304), .ZN(P2_U3220) );
  INV_X1 U9821 ( .A(n8437), .ZN(n8309) );
  NOR3_X1 U9822 ( .A1(n8307), .A2(n8764), .A3(n8443), .ZN(n8308) );
  AOI21_X1 U9823 ( .B1(n8309), .B2(n8460), .A(n8308), .ZN(n8316) );
  OAI22_X1 U9824 ( .A1(n8551), .A2(n8765), .B1(n8764), .B2(n8277), .ZN(n8740)
         );
  AOI22_X1 U9825 ( .A1(n8426), .A2(n8740), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8310) );
  OAI21_X1 U9826 ( .B1(n8734), .B2(n8464), .A(n8310), .ZN(n8313) );
  NOR2_X1 U9827 ( .A1(n8311), .A2(n8445), .ZN(n8312) );
  AOI211_X1 U9828 ( .C1(n8869), .C2(n8469), .A(n8313), .B(n8312), .ZN(n8314)
         );
  OAI21_X1 U9829 ( .B1(n8316), .B2(n8315), .A(n8314), .ZN(P2_U3221) );
  INV_X1 U9830 ( .A(n8317), .ZN(n8318) );
  AOI21_X1 U9831 ( .B1(n8393), .B2(n8318), .A(n8445), .ZN(n8322) );
  NOR3_X1 U9832 ( .A1(n8319), .A2(n8551), .A3(n8443), .ZN(n8321) );
  OAI21_X1 U9833 ( .B1(n8322), .B2(n8321), .A(n8320), .ZN(n8328) );
  INV_X1 U9834 ( .A(n8323), .ZN(n8704) );
  OAI22_X1 U9835 ( .A1(n8671), .A2(n8765), .B1(n8551), .B2(n8277), .ZN(n8708)
         );
  INV_X1 U9836 ( .A(n8708), .ZN(n8325) );
  OAI22_X1 U9837 ( .A1(n8452), .A2(n8325), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8324), .ZN(n8326) );
  AOI21_X1 U9838 ( .B1(n8704), .B2(n8454), .A(n8326), .ZN(n8327) );
  OAI211_X1 U9839 ( .C1(n8706), .C2(n8458), .A(n8328), .B(n8327), .ZN(P2_U3225) );
  NAND2_X1 U9840 ( .A1(n8330), .A2(n8329), .ZN(n8332) );
  XOR2_X1 U9841 ( .A(n8332), .B(n8331), .Z(n8340) );
  OAI21_X1 U9842 ( .B1(n8464), .B2(n8334), .A(n8333), .ZN(n8337) );
  OAI22_X1 U9843 ( .A1(n8335), .A2(n8465), .B1(n8466), .B2(n8480), .ZN(n8336)
         );
  AOI211_X1 U9844 ( .C1(n8338), .C2(n8469), .A(n8337), .B(n8336), .ZN(n8339)
         );
  OAI21_X1 U9845 ( .B1(n8340), .B2(n8445), .A(n8339), .ZN(P2_U3226) );
  INV_X1 U9846 ( .A(n8838), .ZN(n8638) );
  OAI211_X1 U9847 ( .C1(n8342), .C2(n8341), .A(n8447), .B(n8460), .ZN(n8347)
         );
  OAI22_X1 U9848 ( .A1(n8563), .A2(n8765), .B1(n8672), .B2(n8277), .ZN(n8642)
         );
  INV_X1 U9849 ( .A(n8642), .ZN(n8344) );
  OAI22_X1 U9850 ( .A1(n8344), .A2(n8452), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8343), .ZN(n8345) );
  AOI21_X1 U9851 ( .B1(n8636), .B2(n8454), .A(n8345), .ZN(n8346) );
  OAI211_X1 U9852 ( .C1(n8638), .C2(n8458), .A(n8347), .B(n8346), .ZN(P2_U3227) );
  XNOR2_X1 U9853 ( .A(n8350), .B(n8348), .ZN(n8461) );
  NAND2_X1 U9854 ( .A1(n8461), .A2(n8349), .ZN(n8462) );
  OAI21_X1 U9855 ( .B1(n8351), .B2(n8350), .A(n8462), .ZN(n8355) );
  XNOR2_X1 U9856 ( .A(n8353), .B(n8352), .ZN(n8354) );
  XNOR2_X1 U9857 ( .A(n8355), .B(n8354), .ZN(n8360) );
  INV_X1 U9858 ( .A(n8781), .ZN(n8357) );
  OAI22_X1 U9859 ( .A1(n8749), .A2(n8765), .B1(n8546), .B2(n8277), .ZN(n8786)
         );
  AOI22_X1 U9860 ( .A1(n8426), .A2(n8786), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n8356) );
  OAI21_X1 U9861 ( .B1(n8357), .B2(n8464), .A(n8356), .ZN(n8358) );
  AOI21_X1 U9862 ( .B1(n8884), .B2(n8469), .A(n8358), .ZN(n8359) );
  OAI21_X1 U9863 ( .B1(n8360), .B2(n8445), .A(n8359), .ZN(P2_U3228) );
  INV_X1 U9864 ( .A(n8880), .ZN(n8772) );
  OAI211_X1 U9865 ( .C1(n8362), .C2(n8361), .A(n8435), .B(n8460), .ZN(n8366)
         );
  NOR2_X1 U9866 ( .A1(n8363), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8515) );
  OAI22_X1 U9867 ( .A1(n8763), .A2(n8465), .B1(n8466), .B2(n8764), .ZN(n8364)
         );
  AOI211_X1 U9868 ( .C1(n8454), .C2(n8769), .A(n8515), .B(n8364), .ZN(n8365)
         );
  OAI211_X1 U9869 ( .C1(n8772), .C2(n8458), .A(n8366), .B(n8365), .ZN(P2_U3230) );
  NOR2_X1 U9870 ( .A1(n8368), .A2(n8367), .ZN(n8370) );
  XNOR2_X1 U9871 ( .A(n8370), .B(n8369), .ZN(n8373) );
  OAI22_X1 U9872 ( .A1(n8373), .A2(n8445), .B1(n8672), .B2(n8443), .ZN(n8371)
         );
  OAI21_X1 U9873 ( .B1(n8373), .B2(n8372), .A(n8371), .ZN(n8377) );
  NOR2_X1 U9874 ( .A1(n8464), .A2(n8652), .ZN(n8375) );
  OAI22_X1 U9875 ( .A1(n8658), .A2(n8465), .B1(n8466), .B2(n8659), .ZN(n8374)
         );
  AOI211_X1 U9876 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3152), .A(n8375), 
        .B(n8374), .ZN(n8376) );
  OAI211_X1 U9877 ( .C1(n8655), .C2(n8458), .A(n8377), .B(n8376), .ZN(P2_U3231) );
  NAND4_X1 U9878 ( .A1(n8459), .A2(n8489), .A3(n8378), .A4(n8381), .ZN(n8391)
         );
  INV_X1 U9879 ( .A(n8379), .ZN(n8382) );
  NOR2_X1 U9880 ( .A1(n8382), .A2(n8380), .ZN(n8383) );
  MUX2_X1 U9881 ( .A(n8383), .B(n8382), .S(n8381), .Z(n8384) );
  NAND2_X1 U9882 ( .A1(n8384), .A2(n8460), .ZN(n8390) );
  AOI22_X1 U9883 ( .A1(n8426), .A2(n8385), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n8389) );
  AOI22_X1 U9884 ( .A1(n8469), .A2(n8387), .B1(n8454), .B2(n8386), .ZN(n8388)
         );
  NAND4_X1 U9885 ( .A1(n8391), .A2(n8390), .A3(n8389), .A4(n8388), .ZN(
        P2_U3232) );
  OAI22_X1 U9886 ( .A1(n8552), .A2(n8765), .B1(n8750), .B2(n8277), .ZN(n8727)
         );
  AOI22_X1 U9887 ( .A1(n8426), .A2(n8727), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8392) );
  OAI21_X1 U9888 ( .B1(n8717), .B2(n8464), .A(n8392), .ZN(n8398) );
  INV_X1 U9889 ( .A(n8393), .ZN(n8394) );
  AOI211_X1 U9890 ( .C1(n8396), .C2(n8395), .A(n8445), .B(n8394), .ZN(n8397)
         );
  AOI211_X1 U9891 ( .C1(n8863), .C2(n8469), .A(n8398), .B(n8397), .ZN(n8399)
         );
  INV_X1 U9892 ( .A(n8399), .ZN(P2_U3235) );
  OAI211_X1 U9893 ( .C1(n8402), .C2(n8401), .A(n8400), .B(n8460), .ZN(n8409)
         );
  INV_X1 U9894 ( .A(n8403), .ZN(n8404) );
  NOR2_X1 U9895 ( .A1(n8464), .A2(n8404), .ZN(n8405) );
  AOI211_X1 U9896 ( .C1(n8426), .C2(n8407), .A(n8406), .B(n8405), .ZN(n8408)
         );
  OAI211_X1 U9897 ( .C1(n8410), .C2(n8458), .A(n8409), .B(n8408), .ZN(P2_U3236) );
  NAND2_X1 U9898 ( .A1(n8459), .A2(n8476), .ZN(n8414) );
  NAND2_X1 U9899 ( .A1(n8460), .A2(n8411), .ZN(n8413) );
  MUX2_X1 U9900 ( .A(n8414), .B(n8413), .S(n8412), .Z(n8420) );
  OAI22_X1 U9901 ( .A1(n8464), .A2(n8416), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8415), .ZN(n8418) );
  OAI22_X1 U9902 ( .A1(n8552), .A2(n8465), .B1(n8466), .B2(n8658), .ZN(n8417)
         );
  AOI211_X1 U9903 ( .C1(n8853), .C2(n8469), .A(n8418), .B(n8417), .ZN(n8419)
         );
  NAND2_X1 U9904 ( .A1(n8420), .A2(n8419), .ZN(P2_U3237) );
  XOR2_X1 U9905 ( .A(n8422), .B(n8421), .Z(n8423) );
  NAND2_X1 U9906 ( .A1(n8423), .A2(n8460), .ZN(n8432) );
  AOI21_X1 U9907 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8431) );
  NAND2_X1 U9908 ( .A1(n8469), .A2(n8427), .ZN(n8430) );
  NAND2_X1 U9909 ( .A1(n8454), .A2(n8428), .ZN(n8429) );
  NAND4_X1 U9910 ( .A1(n8432), .A2(n8431), .A3(n8430), .A4(n8429), .ZN(
        P2_U3238) );
  INV_X1 U9911 ( .A(n8433), .ZN(n8434) );
  AOI21_X1 U9912 ( .B1(n8435), .B2(n8434), .A(n8445), .ZN(n8439) );
  NOR3_X1 U9913 ( .A1(n8436), .A2(n8749), .A3(n8443), .ZN(n8438) );
  OAI21_X1 U9914 ( .B1(n8439), .B2(n8438), .A(n8437), .ZN(n8442) );
  AND2_X1 U9915 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8524) );
  OAI22_X1 U9916 ( .A1(n8749), .A2(n8465), .B1(n8466), .B2(n8750), .ZN(n8440)
         );
  AOI211_X1 U9917 ( .C1(n8454), .C2(n8752), .A(n8524), .B(n8440), .ZN(n8441)
         );
  OAI211_X1 U9918 ( .C1(n8755), .C2(n8458), .A(n8442), .B(n8441), .ZN(P2_U3240) );
  NOR3_X1 U9919 ( .A1(n8444), .A2(n8659), .A3(n8443), .ZN(n8450) );
  AOI21_X1 U9920 ( .B1(n8447), .B2(n8446), .A(n8445), .ZN(n8449) );
  OAI21_X1 U9921 ( .B1(n8450), .B2(n8449), .A(n8448), .ZN(n8457) );
  INV_X1 U9922 ( .A(n8626), .ZN(n8455) );
  AOI22_X1 U9923 ( .A1(n8474), .A2(n8801), .B1(n8799), .B2(n8561), .ZN(n8623)
         );
  OAI22_X1 U9924 ( .A1(n8623), .A2(n8452), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8451), .ZN(n8453) );
  AOI21_X1 U9925 ( .B1(n8455), .B2(n8454), .A(n8453), .ZN(n8456) );
  OAI211_X1 U9926 ( .C1(n4485), .C2(n8458), .A(n8457), .B(n8456), .ZN(P2_U3242) );
  INV_X1 U9927 ( .A(n8546), .ZN(n8478) );
  AOI22_X1 U9928 ( .A1(n8461), .A2(n8460), .B1(n8459), .B2(n8478), .ZN(n8472)
         );
  INV_X1 U9929 ( .A(n8462), .ZN(n8471) );
  INV_X1 U9930 ( .A(n8793), .ZN(n8463) );
  OAI22_X1 U9931 ( .A1(n8464), .A2(n8463), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5294), .ZN(n8468) );
  OAI22_X1 U9932 ( .A1(n8763), .A2(n8466), .B1(n8465), .B2(n8479), .ZN(n8467)
         );
  AOI211_X1 U9933 ( .C1(n8888), .C2(n8469), .A(n8468), .B(n8467), .ZN(n8470)
         );
  OAI21_X1 U9934 ( .B1(n8472), .B2(n8471), .A(n8470), .ZN(P2_U3243) );
  MUX2_X1 U9935 ( .A(n8473), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8493), .Z(
        P2_U3580) );
  MUX2_X1 U9936 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8474), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9937 ( .A(n8561), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8493), .Z(
        P2_U3577) );
  MUX2_X1 U9938 ( .A(n8475), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8493), .Z(
        P2_U3576) );
  MUX2_X1 U9939 ( .A(n8695), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8493), .Z(
        P2_U3575) );
  MUX2_X1 U9940 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8476), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9941 ( .A(n8694), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8493), .Z(
        P2_U3573) );
  MUX2_X1 U9942 ( .A(n8549), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8493), .Z(
        P2_U3571) );
  MUX2_X1 U9943 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8477), .S(P2_U3966), .Z(
        P2_U3570) );
  INV_X1 U9944 ( .A(n8763), .ZN(n8802) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8802), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8478), .S(P2_U3966), .Z(
        P2_U3567) );
  INV_X1 U9947 ( .A(n8479), .ZN(n8800) );
  MUX2_X1 U9948 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8800), .S(P2_U3966), .Z(
        P2_U3566) );
  INV_X1 U9949 ( .A(n8480), .ZN(n8544) );
  MUX2_X1 U9950 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8544), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9951 ( .A(n8481), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8493), .Z(
        P2_U3564) );
  MUX2_X1 U9952 ( .A(n8482), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8493), .Z(
        P2_U3563) );
  MUX2_X1 U9953 ( .A(n8483), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8493), .Z(
        P2_U3562) );
  MUX2_X1 U9954 ( .A(n8484), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8493), .Z(
        P2_U3561) );
  MUX2_X1 U9955 ( .A(n8485), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8493), .Z(
        P2_U3560) );
  MUX2_X1 U9956 ( .A(n8486), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8493), .Z(
        P2_U3559) );
  MUX2_X1 U9957 ( .A(n8487), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8493), .Z(
        P2_U3558) );
  MUX2_X1 U9958 ( .A(n8488), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8493), .Z(
        P2_U3557) );
  MUX2_X1 U9959 ( .A(n8489), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8493), .Z(
        P2_U3556) );
  MUX2_X1 U9960 ( .A(n8490), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8493), .Z(
        P2_U3555) );
  MUX2_X1 U9961 ( .A(n8491), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8493), .Z(
        P2_U3554) );
  MUX2_X1 U9962 ( .A(n8492), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8493), .Z(
        P2_U3553) );
  MUX2_X1 U9963 ( .A(n9872), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8493), .Z(
        P2_U3552) );
  OAI21_X1 U9964 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(n8497) );
  NAND2_X1 U9965 ( .A1(n8497), .A2(n9783), .ZN(n8507) );
  NOR2_X1 U9966 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8498), .ZN(n8499) );
  AOI21_X1 U9967 ( .B1(n9785), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8499), .ZN(
        n8506) );
  OAI211_X1 U9968 ( .C1(n8502), .C2(n8501), .A(n9784), .B(n8500), .ZN(n8505)
         );
  NAND2_X1 U9969 ( .A1(n8529), .A2(n8503), .ZN(n8504) );
  NAND4_X1 U9970 ( .A1(n8507), .A2(n8506), .A3(n8505), .A4(n8504), .ZN(
        P2_U3261) );
  OAI211_X1 U9971 ( .C1(n8510), .C2(n8509), .A(n9784), .B(n8508), .ZN(n8517)
         );
  AOI211_X1 U9972 ( .C1(n8513), .C2(n8512), .A(n8511), .B(n9787), .ZN(n8514)
         );
  AOI211_X1 U9973 ( .C1(n9785), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8515), .B(
        n8514), .ZN(n8516) );
  OAI211_X1 U9974 ( .C1(n9786), .C2(n8518), .A(n8517), .B(n8516), .ZN(P2_U3262) );
  AOI21_X1 U9975 ( .B1(n8520), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8519), .ZN(
        n8532) );
  XNOR2_X1 U9976 ( .A(n8522), .B(n8521), .ZN(n8523) );
  NAND2_X1 U9977 ( .A1(n9783), .A2(n8523), .ZN(n8526) );
  INV_X1 U9978 ( .A(n8524), .ZN(n8525) );
  OAI211_X1 U9979 ( .C1(n10006), .C2(n8527), .A(n8526), .B(n8525), .ZN(n8528)
         );
  AOI21_X1 U9980 ( .B1(n8530), .B2(n8529), .A(n8528), .ZN(n8531) );
  OAI21_X1 U9981 ( .B1(n8532), .B2(n9788), .A(n8531), .ZN(P2_U3263) );
  INV_X1 U9982 ( .A(n8818), .ZN(n8570) );
  INV_X1 U9983 ( .A(n8888), .ZN(n8796) );
  INV_X1 U9984 ( .A(n8884), .ZN(n8783) );
  NAND2_X1 U9985 ( .A1(n8792), .A2(n8783), .ZN(n8778) );
  INV_X1 U9986 ( .A(n8863), .ZN(n8720) );
  NAND2_X1 U9987 ( .A1(n5633), .A2(n8568), .ZN(n8540) );
  XNOR2_X1 U9988 ( .A(n8810), .B(n8540), .ZN(n8533) );
  NAND2_X1 U9989 ( .A1(n8533), .A2(n9905), .ZN(n8809) );
  INV_X1 U9990 ( .A(n5832), .ZN(n8534) );
  NAND2_X1 U9991 ( .A1(n8534), .A2(P2_B_REG_SCAN_IN), .ZN(n8535) );
  NAND2_X1 U9992 ( .A1(n8801), .A2(n8535), .ZN(n8578) );
  OR2_X1 U9993 ( .A1(n8536), .A2(n8578), .ZN(n8813) );
  NOR2_X1 U9994 ( .A1(n9831), .A2(n8813), .ZN(n8542) );
  NOR2_X1 U9995 ( .A1(n8810), .A2(n8795), .ZN(n8537) );
  AOI211_X1 U9996 ( .C1(n9831), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8542), .B(
        n8537), .ZN(n8538) );
  OAI21_X1 U9997 ( .B1(n8539), .B2(n8809), .A(n8538), .ZN(P2_U3265) );
  OAI21_X1 U9998 ( .B1(n5633), .B2(n8568), .A(n8540), .ZN(n8814) );
  NOR2_X1 U9999 ( .A1(n5633), .A2(n8795), .ZN(n8541) );
  AOI211_X1 U10000 ( .C1(n9831), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8542), .B(
        n8541), .ZN(n8543) );
  OAI21_X1 U10001 ( .B1(n8814), .B2(n8683), .A(n8543), .ZN(P2_U3266) );
  INV_X1 U10002 ( .A(n8853), .ZN(n8690) );
  NAND2_X1 U10003 ( .A1(n9579), .A2(n9578), .ZN(n9577) );
  NAND2_X1 U10004 ( .A1(n9586), .A2(n8479), .ZN(n8545) );
  NAND2_X1 U10005 ( .A1(n8755), .A2(n8764), .ZN(n8548) );
  NOR2_X1 U10006 ( .A1(n8755), .A2(n8764), .ZN(n8547) );
  NAND2_X1 U10007 ( .A1(n8869), .A2(n8549), .ZN(n8550) );
  INV_X1 U10008 ( .A(n8869), .ZN(n8737) );
  NAND2_X1 U10009 ( .A1(n8706), .A2(n8552), .ZN(n8553) );
  INV_X1 U10010 ( .A(n8555), .ZN(n8556) );
  NAND2_X1 U10011 ( .A1(n8848), .A2(n8695), .ZN(n8557) );
  NAND2_X1 U10012 ( .A1(n8655), .A2(n8672), .ZN(n8559) );
  NAND2_X1 U10013 ( .A1(n8560), .A2(n8559), .ZN(n8632) );
  NAND2_X1 U10014 ( .A1(n8632), .A2(n8640), .ZN(n8631) );
  NAND2_X1 U10015 ( .A1(n4485), .A2(n8563), .ZN(n8564) );
  NAND2_X1 U10016 ( .A1(n8609), .A2(n8588), .ZN(n8565) );
  NAND2_X1 U10017 ( .A1(n8603), .A2(n8565), .ZN(n8594) );
  NAND2_X1 U10018 ( .A1(n8594), .A2(n8593), .ZN(n8592) );
  NAND2_X1 U10019 ( .A1(n8599), .A2(n8579), .ZN(n8566) );
  NAND2_X1 U10020 ( .A1(n8592), .A2(n8566), .ZN(n8567) );
  XNOR2_X1 U10021 ( .A(n8567), .B(n8575), .ZN(n8815) );
  INV_X1 U10022 ( .A(n8815), .ZN(n8584) );
  INV_X1 U10023 ( .A(n8595), .ZN(n8569) );
  AOI211_X1 U10024 ( .C1(n8818), .C2(n8569), .A(n9943), .B(n8568), .ZN(n8817)
         );
  NOR2_X1 U10025 ( .A1(n8570), .A2(n8795), .ZN(n8574) );
  OAI22_X1 U10026 ( .A1(n9829), .A2(n8572), .B1(n8571), .B2(n8678), .ZN(n8573)
         );
  AOI211_X1 U10027 ( .C1(n8817), .C2(n9812), .A(n8574), .B(n8573), .ZN(n8583)
         );
  INV_X1 U10028 ( .A(n8580), .ZN(n8581) );
  NAND2_X1 U10029 ( .A1(n8816), .A2(n9829), .ZN(n8582) );
  OAI211_X1 U10030 ( .C1(n8584), .C2(n8808), .A(n8583), .B(n8582), .ZN(
        P2_U3267) );
  INV_X1 U10031 ( .A(n8585), .ZN(n8586) );
  AOI21_X1 U10032 ( .B1(n8586), .B2(n8593), .A(n9570), .ZN(n8591) );
  OAI22_X1 U10033 ( .A1(n8588), .A2(n8277), .B1(n8587), .B2(n8765), .ZN(n8589)
         );
  AOI21_X1 U10034 ( .B1(n8591), .B2(n8590), .A(n8589), .ZN(n8825) );
  OAI21_X1 U10035 ( .B1(n8594), .B2(n8593), .A(n8592), .ZN(n8821) );
  NAND2_X1 U10036 ( .A1(n8821), .A2(n9581), .ZN(n8602) );
  INV_X1 U10037 ( .A(n8606), .ZN(n8596) );
  AOI21_X1 U10038 ( .B1(n8822), .B2(n8596), .A(n8595), .ZN(n8823) );
  AOI22_X1 U10039 ( .A1(n9831), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8597), .B2(
        n9821), .ZN(n8598) );
  OAI21_X1 U10040 ( .B1(n8599), .B2(n8795), .A(n8598), .ZN(n8600) );
  AOI21_X1 U10041 ( .B1(n8823), .B2(n8806), .A(n8600), .ZN(n8601) );
  OAI211_X1 U10042 ( .C1(n9831), .C2(n8825), .A(n8602), .B(n8601), .ZN(
        P2_U3268) );
  OAI21_X1 U10043 ( .B1(n8604), .B2(n8610), .A(n8603), .ZN(n8605) );
  INV_X1 U10044 ( .A(n8605), .ZN(n8831) );
  AOI211_X1 U10045 ( .C1(n8828), .C2(n4487), .A(n9943), .B(n8606), .ZN(n8827)
         );
  AOI22_X1 U10046 ( .A1(n9831), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8607), .B2(
        n9821), .ZN(n8608) );
  OAI21_X1 U10047 ( .B1(n8609), .B2(n8795), .A(n8608), .ZN(n8615) );
  AOI21_X1 U10048 ( .B1(n4325), .B2(n8610), .A(n9570), .ZN(n8613) );
  AOI21_X1 U10049 ( .B1(n8613), .B2(n8611), .A(n8612), .ZN(n8830) );
  NOR2_X1 U10050 ( .A1(n8830), .A2(n9831), .ZN(n8614) );
  AOI211_X1 U10051 ( .C1(n8827), .C2(n9812), .A(n8615), .B(n8614), .ZN(n8616)
         );
  OAI21_X1 U10052 ( .B1(n8831), .B2(n8808), .A(n8616), .ZN(P2_U3269) );
  OAI21_X1 U10053 ( .B1(n8618), .B2(n5653), .A(n8617), .ZN(n8619) );
  INV_X1 U10054 ( .A(n8619), .ZN(n8836) );
  AOI22_X1 U10055 ( .A1(n8834), .A2(n9805), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n9831), .ZN(n8630) );
  INV_X1 U10056 ( .A(n8620), .ZN(n8621) );
  AOI21_X1 U10057 ( .B1(n5653), .B2(n8622), .A(n8621), .ZN(n8624) );
  OAI21_X1 U10058 ( .B1(n8624), .B2(n9570), .A(n8623), .ZN(n8832) );
  AOI211_X1 U10059 ( .C1(n8834), .C2(n8634), .A(n9943), .B(n8625), .ZN(n8833)
         );
  INV_X1 U10060 ( .A(n8833), .ZN(n8627) );
  OAI22_X1 U10061 ( .A1(n8627), .A2(n9823), .B1(n8678), .B2(n8626), .ZN(n8628)
         );
  OAI21_X1 U10062 ( .B1(n8832), .B2(n8628), .A(n9829), .ZN(n8629) );
  OAI211_X1 U10063 ( .C1(n8836), .C2(n8808), .A(n8630), .B(n8629), .ZN(
        P2_U3270) );
  OAI21_X1 U10064 ( .B1(n8632), .B2(n8640), .A(n8631), .ZN(n8633) );
  INV_X1 U10065 ( .A(n8633), .ZN(n8841) );
  INV_X1 U10066 ( .A(n8634), .ZN(n8635) );
  AOI211_X1 U10067 ( .C1(n8838), .C2(n8649), .A(n9943), .B(n8635), .ZN(n8837)
         );
  NOR2_X1 U10068 ( .A1(n9831), .A2(n9823), .ZN(n8768) );
  AOI22_X1 U10069 ( .A1(n9831), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8636), .B2(
        n9821), .ZN(n8637) );
  OAI21_X1 U10070 ( .B1(n8638), .B2(n8795), .A(n8637), .ZN(n8646) );
  INV_X1 U10071 ( .A(n8639), .ZN(n8641) );
  AOI21_X1 U10072 ( .B1(n8641), .B2(n8640), .A(n9570), .ZN(n8644) );
  AOI21_X1 U10073 ( .B1(n8644), .B2(n8643), .A(n8642), .ZN(n8840) );
  NOR2_X1 U10074 ( .A1(n8840), .A2(n9831), .ZN(n8645) );
  AOI211_X1 U10075 ( .C1(n8837), .C2(n8768), .A(n8646), .B(n8645), .ZN(n8647)
         );
  OAI21_X1 U10076 ( .B1(n8841), .B2(n8808), .A(n8647), .ZN(P2_U3271) );
  XNOR2_X1 U10077 ( .A(n8648), .B(n8656), .ZN(n8846) );
  INV_X1 U10078 ( .A(n8677), .ZN(n8651) );
  INV_X1 U10079 ( .A(n8649), .ZN(n8650) );
  AOI21_X1 U10080 ( .B1(n8842), .B2(n8651), .A(n8650), .ZN(n8843) );
  INV_X1 U10081 ( .A(n8652), .ZN(n8653) );
  AOI22_X1 U10082 ( .A1(n9831), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8653), .B2(
        n9821), .ZN(n8654) );
  OAI21_X1 U10083 ( .B1(n8655), .B2(n8795), .A(n8654), .ZN(n8664) );
  AOI21_X1 U10084 ( .B1(n8657), .B2(n8656), .A(n9570), .ZN(n8662) );
  OAI22_X1 U10085 ( .A1(n8659), .A2(n8765), .B1(n8658), .B2(n8277), .ZN(n8660)
         );
  AOI21_X1 U10086 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8845) );
  NOR2_X1 U10087 ( .A1(n8845), .A2(n9831), .ZN(n8663) );
  AOI211_X1 U10088 ( .C1(n8843), .C2(n8806), .A(n8664), .B(n8663), .ZN(n8665)
         );
  OAI21_X1 U10089 ( .B1(n8846), .B2(n8808), .A(n8665), .ZN(P2_U3272) );
  OAI21_X1 U10090 ( .B1(n8667), .B2(n8556), .A(n8666), .ZN(n8852) );
  NAND2_X1 U10091 ( .A1(n8668), .A2(n8556), .ZN(n8669) );
  NAND2_X1 U10092 ( .A1(n8670), .A2(n8669), .ZN(n8674) );
  OAI22_X1 U10093 ( .A1(n8672), .A2(n8765), .B1(n8671), .B2(n8277), .ZN(n8673)
         );
  AOI21_X1 U10094 ( .B1(n8674), .B2(n9803), .A(n8673), .ZN(n8851) );
  INV_X1 U10095 ( .A(n8851), .ZN(n8685) );
  NOR2_X1 U10096 ( .A1(n8687), .A2(n8675), .ZN(n8676) );
  OR2_X1 U10097 ( .A1(n8677), .A2(n8676), .ZN(n8847) );
  INV_X1 U10098 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8680) );
  OAI22_X1 U10099 ( .A1(n9829), .A2(n8680), .B1(n8679), .B2(n8678), .ZN(n8681)
         );
  AOI21_X1 U10100 ( .B1(n8848), .B2(n9805), .A(n8681), .ZN(n8682) );
  OAI21_X1 U10101 ( .B1(n8847), .B2(n8683), .A(n8682), .ZN(n8684) );
  AOI21_X1 U10102 ( .B1(n8685), .B2(n9829), .A(n8684), .ZN(n8686) );
  OAI21_X1 U10103 ( .B1(n8852), .B2(n8808), .A(n8686), .ZN(P2_U3273) );
  XNOR2_X1 U10104 ( .A(n4336), .B(n8693), .ZN(n8857) );
  AOI21_X1 U10105 ( .B1(n8853), .B2(n8703), .A(n8687), .ZN(n8854) );
  AOI22_X1 U10106 ( .A1(n9831), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8688), .B2(
        n9821), .ZN(n8689) );
  OAI21_X1 U10107 ( .B1(n8690), .B2(n8795), .A(n8689), .ZN(n8699) );
  OAI211_X1 U10108 ( .C1(n8691), .C2(n8693), .A(n8692), .B(n9803), .ZN(n8697)
         );
  AOI22_X1 U10109 ( .A1(n8695), .A2(n8801), .B1(n8799), .B2(n8694), .ZN(n8696)
         );
  AND2_X1 U10110 ( .A1(n8697), .A2(n8696), .ZN(n8856) );
  NOR2_X1 U10111 ( .A1(n8856), .A2(n9831), .ZN(n8698) );
  AOI211_X1 U10112 ( .C1(n8854), .C2(n8806), .A(n8699), .B(n8698), .ZN(n8700)
         );
  OAI21_X1 U10113 ( .B1(n8857), .B2(n8808), .A(n8700), .ZN(P2_U3274) );
  XNOR2_X1 U10114 ( .A(n8702), .B(n8701), .ZN(n8862) );
  AOI211_X1 U10115 ( .C1(n8859), .C2(n8715), .A(n9943), .B(n4495), .ZN(n8858)
         );
  AOI22_X1 U10116 ( .A1(n9831), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8704), .B2(
        n9821), .ZN(n8705) );
  OAI21_X1 U10117 ( .B1(n8706), .B2(n8795), .A(n8705), .ZN(n8711) );
  XNOR2_X1 U10118 ( .A(n4335), .B(n8707), .ZN(n8709) );
  AOI21_X1 U10119 ( .B1(n8709), .B2(n9803), .A(n8708), .ZN(n8861) );
  NOR2_X1 U10120 ( .A1(n8861), .A2(n9831), .ZN(n8710) );
  AOI211_X1 U10121 ( .C1(n8858), .C2(n9812), .A(n8711), .B(n8710), .ZN(n8712)
         );
  OAI21_X1 U10122 ( .B1(n8862), .B2(n8808), .A(n8712), .ZN(P2_U3275) );
  OAI21_X1 U10123 ( .B1(n8714), .B2(n8726), .A(n8713), .ZN(n8867) );
  INV_X1 U10124 ( .A(n8733), .ZN(n8716) );
  AOI21_X1 U10125 ( .B1(n8863), .B2(n8716), .A(n4491), .ZN(n8864) );
  INV_X1 U10126 ( .A(n8717), .ZN(n8718) );
  AOI22_X1 U10127 ( .A1(n9831), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8718), .B2(
        n9821), .ZN(n8719) );
  OAI21_X1 U10128 ( .B1(n8720), .B2(n8795), .A(n8719), .ZN(n8730) );
  NAND2_X1 U10129 ( .A1(n8721), .A2(n8722), .ZN(n8725) );
  INV_X1 U10130 ( .A(n8723), .ZN(n8724) );
  AOI211_X1 U10131 ( .C1(n8726), .C2(n8725), .A(n9570), .B(n8724), .ZN(n8728)
         );
  NOR2_X1 U10132 ( .A1(n8728), .A2(n8727), .ZN(n8866) );
  NOR2_X1 U10133 ( .A1(n8866), .A2(n9831), .ZN(n8729) );
  AOI211_X1 U10134 ( .C1(n8864), .C2(n8806), .A(n8730), .B(n8729), .ZN(n8731)
         );
  OAI21_X1 U10135 ( .B1(n8867), .B2(n8808), .A(n8731), .ZN(P2_U3276) );
  XNOR2_X1 U10136 ( .A(n8732), .B(n8739), .ZN(n8872) );
  AOI211_X1 U10137 ( .C1(n8869), .C2(n8751), .A(n9943), .B(n8733), .ZN(n8868)
         );
  INV_X1 U10138 ( .A(n8734), .ZN(n8735) );
  AOI22_X1 U10139 ( .A1(n9831), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8735), .B2(
        n9821), .ZN(n8736) );
  OAI21_X1 U10140 ( .B1(n8737), .B2(n8795), .A(n8736), .ZN(n8743) );
  OAI21_X1 U10141 ( .B1(n8739), .B2(n8738), .A(n8721), .ZN(n8741) );
  AOI21_X1 U10142 ( .B1(n8741), .B2(n9803), .A(n8740), .ZN(n8871) );
  NOR2_X1 U10143 ( .A1(n8871), .A2(n9831), .ZN(n8742) );
  AOI211_X1 U10144 ( .C1(n8868), .C2(n8768), .A(n8743), .B(n8742), .ZN(n8744)
         );
  OAI21_X1 U10145 ( .B1(n8872), .B2(n8808), .A(n8744), .ZN(P2_U3277) );
  XOR2_X1 U10146 ( .A(n8746), .B(n8745), .Z(n8877) );
  XNOR2_X1 U10147 ( .A(n8747), .B(n8746), .ZN(n8748) );
  OAI222_X1 U10148 ( .A1(n8765), .A2(n8750), .B1(n8277), .B2(n8749), .C1(n9570), .C2(n8748), .ZN(n8873) );
  AOI211_X1 U10149 ( .C1(n8875), .C2(n8766), .A(n9943), .B(n4496), .ZN(n8874)
         );
  NAND2_X1 U10150 ( .A1(n8874), .A2(n9812), .ZN(n8754) );
  AOI22_X1 U10151 ( .A1(n9831), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8752), .B2(
        n9821), .ZN(n8753) );
  OAI211_X1 U10152 ( .C1(n8755), .C2(n8795), .A(n8754), .B(n8753), .ZN(n8756)
         );
  AOI21_X1 U10153 ( .B1(n8873), .B2(n9829), .A(n8756), .ZN(n8757) );
  OAI21_X1 U10154 ( .B1(n8877), .B2(n8808), .A(n8757), .ZN(P2_U3278) );
  AOI21_X1 U10155 ( .B1(n8760), .B2(n8759), .A(n8758), .ZN(n8882) );
  XNOR2_X1 U10156 ( .A(n8761), .B(n8760), .ZN(n8762) );
  OAI222_X1 U10157 ( .A1(n8765), .A2(n8764), .B1(n8277), .B2(n8763), .C1(n9570), .C2(n8762), .ZN(n8878) );
  INV_X1 U10158 ( .A(n8766), .ZN(n8767) );
  AOI211_X1 U10159 ( .C1(n8880), .C2(n8778), .A(n9943), .B(n8767), .ZN(n8879)
         );
  NAND2_X1 U10160 ( .A1(n8879), .A2(n8768), .ZN(n8771) );
  AOI22_X1 U10161 ( .A1(n9831), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8769), .B2(
        n9821), .ZN(n8770) );
  OAI211_X1 U10162 ( .C1(n8772), .C2(n8795), .A(n8771), .B(n8770), .ZN(n8773)
         );
  AOI21_X1 U10163 ( .B1(n8878), .B2(n9829), .A(n8773), .ZN(n8774) );
  OAI21_X1 U10164 ( .B1(n8882), .B2(n8808), .A(n8774), .ZN(P2_U3279) );
  OAI21_X1 U10165 ( .B1(n8777), .B2(n8776), .A(n8775), .ZN(n8887) );
  INV_X1 U10166 ( .A(n8792), .ZN(n8780) );
  INV_X1 U10167 ( .A(n8778), .ZN(n8779) );
  AOI211_X1 U10168 ( .C1(n8884), .C2(n8780), .A(n9943), .B(n8779), .ZN(n8883)
         );
  AOI22_X1 U10169 ( .A1(n9831), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8781), .B2(
        n9821), .ZN(n8782) );
  OAI21_X1 U10170 ( .B1(n8783), .B2(n8795), .A(n8782), .ZN(n8789) );
  XNOR2_X1 U10171 ( .A(n8785), .B(n8784), .ZN(n8787) );
  AOI21_X1 U10172 ( .B1(n8787), .B2(n9803), .A(n8786), .ZN(n8886) );
  NOR2_X1 U10173 ( .A1(n8886), .A2(n9831), .ZN(n8788) );
  AOI211_X1 U10174 ( .C1(n8883), .C2(n9812), .A(n8789), .B(n8788), .ZN(n8790)
         );
  OAI21_X1 U10175 ( .B1(n8887), .B2(n8808), .A(n8790), .ZN(P2_U3280) );
  XOR2_X1 U10176 ( .A(n8791), .B(n8797), .Z(n8892) );
  AOI21_X1 U10177 ( .B1(n8888), .B2(n4297), .A(n8792), .ZN(n8889) );
  AOI22_X1 U10178 ( .A1(n9831), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8793), .B2(
        n9821), .ZN(n8794) );
  OAI21_X1 U10179 ( .B1(n8796), .B2(n8795), .A(n8794), .ZN(n8805) );
  XNOR2_X1 U10180 ( .A(n8798), .B(n8797), .ZN(n8803) );
  AOI222_X1 U10181 ( .A1(n9803), .A2(n8803), .B1(n8802), .B2(n8801), .C1(n8800), .C2(n8799), .ZN(n8891) );
  NOR2_X1 U10182 ( .A1(n8891), .A2(n9831), .ZN(n8804) );
  AOI211_X1 U10183 ( .C1(n8889), .C2(n8806), .A(n8805), .B(n8804), .ZN(n8807)
         );
  OAI21_X1 U10184 ( .B1(n8892), .B2(n8808), .A(n8807), .ZN(P2_U3281) );
  OAI211_X1 U10185 ( .C1(n8810), .C2(n9941), .A(n8809), .B(n8813), .ZN(n8898)
         );
  MUX2_X1 U10186 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8898), .S(n9967), .Z(
        P2_U3551) );
  NAND2_X1 U10187 ( .A1(n8811), .A2(n9929), .ZN(n8812) );
  OAI211_X1 U10188 ( .C1(n8814), .C2(n9943), .A(n8813), .B(n8812), .ZN(n8899)
         );
  MUX2_X1 U10189 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8899), .S(n9967), .Z(
        P2_U3550) );
  NAND2_X1 U10190 ( .A1(n8815), .A2(n9947), .ZN(n8820) );
  NAND2_X1 U10191 ( .A1(n8820), .A2(n8819), .ZN(n8900) );
  MUX2_X1 U10192 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8900), .S(n9967), .Z(
        P2_U3549) );
  NAND2_X1 U10193 ( .A1(n8821), .A2(n9947), .ZN(n8826) );
  AOI22_X1 U10194 ( .A1(n8823), .A2(n9905), .B1(n9929), .B2(n8822), .ZN(n8824)
         );
  NAND3_X1 U10195 ( .A1(n8826), .A2(n8825), .A3(n8824), .ZN(n8901) );
  MUX2_X1 U10196 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8901), .S(n9967), .Z(
        P2_U3548) );
  AOI21_X1 U10197 ( .B1(n9929), .B2(n8828), .A(n8827), .ZN(n8829) );
  OAI211_X1 U10198 ( .C1(n8831), .C2(n9909), .A(n8830), .B(n8829), .ZN(n8902)
         );
  MUX2_X1 U10199 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8902), .S(n9967), .Z(
        P2_U3547) );
  AOI211_X1 U10200 ( .C1(n9929), .C2(n8834), .A(n8833), .B(n8832), .ZN(n8835)
         );
  OAI21_X1 U10201 ( .B1(n8836), .B2(n9909), .A(n8835), .ZN(n8903) );
  MUX2_X1 U10202 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8903), .S(n9967), .Z(
        P2_U3546) );
  AOI21_X1 U10203 ( .B1(n9929), .B2(n8838), .A(n8837), .ZN(n8839) );
  OAI211_X1 U10204 ( .C1(n8841), .C2(n9909), .A(n8840), .B(n8839), .ZN(n8904)
         );
  MUX2_X1 U10205 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8904), .S(n9967), .Z(
        P2_U3545) );
  AOI22_X1 U10206 ( .A1(n8843), .A2(n9905), .B1(n9929), .B2(n8842), .ZN(n8844)
         );
  OAI211_X1 U10207 ( .C1(n8846), .C2(n9909), .A(n8845), .B(n8844), .ZN(n8905)
         );
  MUX2_X1 U10208 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8905), .S(n9967), .Z(
        P2_U3544) );
  INV_X1 U10209 ( .A(n8847), .ZN(n8849) );
  AOI22_X1 U10210 ( .A1(n8849), .A2(n9905), .B1(n9929), .B2(n8848), .ZN(n8850)
         );
  OAI211_X1 U10211 ( .C1(n8852), .C2(n9909), .A(n8851), .B(n8850), .ZN(n8906)
         );
  MUX2_X1 U10212 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8906), .S(n9967), .Z(
        P2_U3543) );
  AOI22_X1 U10213 ( .A1(n8854), .A2(n9905), .B1(n9929), .B2(n8853), .ZN(n8855)
         );
  OAI211_X1 U10214 ( .C1(n8857), .C2(n9909), .A(n8856), .B(n8855), .ZN(n8907)
         );
  MUX2_X1 U10215 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8907), .S(n9967), .Z(
        P2_U3542) );
  AOI21_X1 U10216 ( .B1(n9929), .B2(n8859), .A(n8858), .ZN(n8860) );
  OAI211_X1 U10217 ( .C1(n8862), .C2(n9909), .A(n8861), .B(n8860), .ZN(n8908)
         );
  MUX2_X1 U10218 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8908), .S(n9967), .Z(
        P2_U3541) );
  AOI22_X1 U10219 ( .A1(n8864), .A2(n9905), .B1(n9929), .B2(n8863), .ZN(n8865)
         );
  OAI211_X1 U10220 ( .C1(n8867), .C2(n9909), .A(n8866), .B(n8865), .ZN(n8909)
         );
  MUX2_X1 U10221 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8909), .S(n9967), .Z(
        P2_U3540) );
  AOI21_X1 U10222 ( .B1(n9929), .B2(n8869), .A(n8868), .ZN(n8870) );
  OAI211_X1 U10223 ( .C1(n8872), .C2(n9909), .A(n8871), .B(n8870), .ZN(n8910)
         );
  MUX2_X1 U10224 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8910), .S(n9967), .Z(
        P2_U3539) );
  AOI211_X1 U10225 ( .C1(n9929), .C2(n8875), .A(n8874), .B(n8873), .ZN(n8876)
         );
  OAI21_X1 U10226 ( .B1(n8877), .B2(n9909), .A(n8876), .ZN(n8911) );
  MUX2_X1 U10227 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8911), .S(n9967), .Z(
        P2_U3538) );
  AOI211_X1 U10228 ( .C1(n9929), .C2(n8880), .A(n8879), .B(n8878), .ZN(n8881)
         );
  OAI21_X1 U10229 ( .B1(n8882), .B2(n9909), .A(n8881), .ZN(n8912) );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8912), .S(n9967), .Z(
        P2_U3537) );
  AOI21_X1 U10231 ( .B1(n9929), .B2(n8884), .A(n8883), .ZN(n8885) );
  OAI211_X1 U10232 ( .C1(n8887), .C2(n9909), .A(n8886), .B(n8885), .ZN(n8913)
         );
  MUX2_X1 U10233 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8913), .S(n9967), .Z(
        P2_U3536) );
  AOI22_X1 U10234 ( .A1(n8889), .A2(n9905), .B1(n9929), .B2(n8888), .ZN(n8890)
         );
  OAI211_X1 U10235 ( .C1(n8892), .C2(n9909), .A(n8891), .B(n8890), .ZN(n8914)
         );
  MUX2_X1 U10236 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8914), .S(n9967), .Z(
        P2_U3535) );
  AOI21_X1 U10237 ( .B1(n9929), .B2(n8894), .A(n8893), .ZN(n8895) );
  OAI211_X1 U10238 ( .C1(n8897), .C2(n9909), .A(n8896), .B(n8895), .ZN(n8915)
         );
  MUX2_X1 U10239 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8915), .S(n9967), .Z(
        P2_U3533) );
  MUX2_X1 U10240 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8898), .S(n9951), .Z(
        P2_U3519) );
  MUX2_X1 U10241 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8899), .S(n9951), .Z(
        P2_U3518) );
  MUX2_X1 U10242 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8900), .S(n9951), .Z(
        P2_U3517) );
  MUX2_X1 U10243 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8901), .S(n9951), .Z(
        P2_U3516) );
  MUX2_X1 U10244 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8902), .S(n9951), .Z(
        P2_U3515) );
  MUX2_X1 U10245 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8903), .S(n9951), .Z(
        P2_U3514) );
  MUX2_X1 U10246 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8904), .S(n9951), .Z(
        P2_U3513) );
  MUX2_X1 U10247 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8905), .S(n9951), .Z(
        P2_U3512) );
  MUX2_X1 U10248 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8906), .S(n9951), .Z(
        P2_U3511) );
  MUX2_X1 U10249 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8907), .S(n9951), .Z(
        P2_U3510) );
  MUX2_X1 U10250 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8908), .S(n9951), .Z(
        P2_U3509) );
  MUX2_X1 U10251 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8909), .S(n9951), .Z(
        P2_U3508) );
  MUX2_X1 U10252 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8910), .S(n9951), .Z(
        P2_U3507) );
  MUX2_X1 U10253 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8911), .S(n9951), .Z(
        P2_U3505) );
  MUX2_X1 U10254 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8912), .S(n9951), .Z(
        P2_U3502) );
  MUX2_X1 U10255 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8913), .S(n9951), .Z(
        P2_U3499) );
  MUX2_X1 U10256 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8914), .S(n9951), .Z(
        P2_U3496) );
  MUX2_X1 U10257 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8915), .S(n9951), .Z(
        P2_U3490) );
  INV_X1 U10258 ( .A(n7935), .ZN(n9523) );
  NOR4_X1 U10259 ( .A1(n8916), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n5528), .ZN(n8917) );
  AOI21_X1 U10260 ( .B1(n8918), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8917), .ZN(
        n8919) );
  OAI21_X1 U10261 ( .B1(n9523), .B2(n8920), .A(n8919), .ZN(P2_U3327) );
  MUX2_X1 U10262 ( .A(n8921), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  AOI22_X1 U10263 ( .A1(n9186), .A2(n9033), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8925) );
  OAI21_X1 U10264 ( .B1(n9152), .B2(n9036), .A(n8925), .ZN(n8927) );
  NOR2_X1 U10265 ( .A1(n9151), .A2(n9027), .ZN(n8926) );
  AOI211_X1 U10266 ( .C1(n9149), .C2(n9031), .A(n8927), .B(n8926), .ZN(n8928)
         );
  NAND2_X1 U10267 ( .A1(n8929), .A2(n8978), .ZN(n8930) );
  XOR2_X1 U10268 ( .A(n8931), .B(n8930), .Z(n8936) );
  AOI22_X1 U10269 ( .A1(n9033), .A2(n9217), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8933) );
  NAND2_X1 U10270 ( .A1(n9218), .A2(n9021), .ZN(n8932) );
  OAI211_X1 U10271 ( .C1(n9000), .C2(n9212), .A(n8933), .B(n8932), .ZN(n8934)
         );
  AOI21_X1 U10272 ( .B1(n9425), .B2(n9038), .A(n8934), .ZN(n8935) );
  OAI21_X1 U10273 ( .B1(n8936), .B2(n4371), .A(n8935), .ZN(P1_U3214) );
  XOR2_X1 U10274 ( .A(n8938), .B(n8937), .Z(n8944) );
  AOI22_X1 U10275 ( .A1(n9021), .A2(n9276), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3084), .ZN(n8940) );
  NAND2_X1 U10276 ( .A1(n9031), .A2(n9270), .ZN(n8939) );
  OAI211_X1 U10277 ( .C1(n8941), .C2(n9023), .A(n8940), .B(n8939), .ZN(n8942)
         );
  AOI21_X1 U10278 ( .B1(n9446), .B2(n9038), .A(n8942), .ZN(n8943) );
  OAI21_X1 U10279 ( .B1(n8944), .B2(n4371), .A(n8943), .ZN(P1_U3217) );
  XNOR2_X1 U10280 ( .A(n8946), .B(n8945), .ZN(n8951) );
  NAND2_X1 U10281 ( .A1(n9031), .A2(n9248), .ZN(n8948) );
  AOI22_X1 U10282 ( .A1(n9033), .A2(n9276), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8947) );
  OAI211_X1 U10283 ( .C1(n9244), .C2(n9036), .A(n8948), .B(n8947), .ZN(n8949)
         );
  AOI21_X1 U10284 ( .B1(n9437), .B2(n9038), .A(n8949), .ZN(n8950) );
  OAI21_X1 U10285 ( .B1(n8951), .B2(n4371), .A(n8950), .ZN(P1_U3221) );
  OAI21_X1 U10286 ( .B1(n8954), .B2(n8953), .A(n8952), .ZN(n8955) );
  NAND2_X1 U10287 ( .A1(n8955), .A2(n9018), .ZN(n8960) );
  AOI22_X1 U10288 ( .A1(n9186), .A2(n9021), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8956) );
  OAI21_X1 U10289 ( .B1(n8957), .B2(n9023), .A(n8956), .ZN(n8958) );
  AOI21_X1 U10290 ( .B1(n9180), .B2(n9031), .A(n8958), .ZN(n8959) );
  OAI211_X1 U10291 ( .C1(n9182), .C2(n9027), .A(n8960), .B(n8959), .ZN(
        P1_U3223) );
  AOI21_X1 U10292 ( .B1(n8963), .B2(n8962), .A(n8961), .ZN(n8968) );
  AOI22_X1 U10293 ( .A1(n9021), .A2(n9294), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8965) );
  NAND2_X1 U10294 ( .A1(n9031), .A2(n9322), .ZN(n8964) );
  OAI211_X1 U10295 ( .C1(n9319), .C2(n9023), .A(n8965), .B(n8964), .ZN(n8966)
         );
  AOI21_X1 U10296 ( .B1(n9462), .B2(n9038), .A(n8966), .ZN(n8967) );
  OAI21_X1 U10297 ( .B1(n8968), .B2(n4371), .A(n8967), .ZN(P1_U3224) );
  AOI21_X1 U10298 ( .B1(n4351), .B2(n8970), .A(n8969), .ZN(n8975) );
  AOI22_X1 U10299 ( .A1(n9021), .A2(n9309), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n8972) );
  NAND2_X1 U10300 ( .A1(n9031), .A2(n9303), .ZN(n8971) );
  OAI211_X1 U10301 ( .C1(n9329), .C2(n9023), .A(n8972), .B(n8971), .ZN(n8973)
         );
  AOI21_X1 U10302 ( .B1(n9455), .B2(n9038), .A(n8973), .ZN(n8974) );
  OAI21_X1 U10303 ( .B1(n8975), .B2(n4371), .A(n8974), .ZN(P1_U3226) );
  INV_X1 U10304 ( .A(n8976), .ZN(n8981) );
  AOI21_X1 U10305 ( .B1(n8979), .B2(n8978), .A(n8977), .ZN(n8980) );
  OAI21_X1 U10306 ( .B1(n8981), .B2(n8980), .A(n9018), .ZN(n8985) );
  AOI22_X1 U10307 ( .A1(n9033), .A2(n9234), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8982) );
  OAI21_X1 U10308 ( .B1(n9044), .B2(n9036), .A(n8982), .ZN(n8983) );
  AOI21_X1 U10309 ( .B1(n9203), .B2(n9031), .A(n8983), .ZN(n8984) );
  OAI211_X1 U10310 ( .C1(n9192), .C2(n9027), .A(n8985), .B(n8984), .ZN(
        P1_U3227) );
  NOR2_X1 U10311 ( .A1(n8986), .A2(n4360), .ZN(n8987) );
  XNOR2_X1 U10312 ( .A(n8988), .B(n8987), .ZN(n8993) );
  AOI22_X1 U10313 ( .A1(n9021), .A2(n9235), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8990) );
  NAND2_X1 U10314 ( .A1(n9031), .A2(n9261), .ZN(n8989) );
  OAI211_X1 U10315 ( .C1(n9258), .C2(n9023), .A(n8990), .B(n8989), .ZN(n8991)
         );
  AOI21_X1 U10316 ( .B1(n9442), .B2(n9038), .A(n8991), .ZN(n8992) );
  OAI21_X1 U10317 ( .B1(n8993), .B2(n4371), .A(n8992), .ZN(P1_U3231) );
  NAND2_X1 U10318 ( .A1(n8995), .A2(n8994), .ZN(n8996) );
  XOR2_X1 U10319 ( .A(n8997), .B(n8996), .Z(n9003) );
  AOI22_X1 U10320 ( .A1(n9033), .A2(n9235), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8999) );
  NAND2_X1 U10321 ( .A1(n9021), .A2(n9234), .ZN(n8998) );
  OAI211_X1 U10322 ( .C1(n9000), .C2(n9227), .A(n8999), .B(n8998), .ZN(n9001)
         );
  AOI21_X1 U10323 ( .B1(n9430), .B2(n9038), .A(n9001), .ZN(n9002) );
  OAI21_X1 U10324 ( .B1(n9003), .B2(n4371), .A(n9002), .ZN(P1_U3233) );
  XNOR2_X1 U10325 ( .A(n9005), .B(n9004), .ZN(n9006) );
  XNOR2_X1 U10326 ( .A(n9007), .B(n9006), .ZN(n9012) );
  NAND2_X1 U10327 ( .A1(n9033), .A2(n9294), .ZN(n9008) );
  NAND2_X1 U10328 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9705) );
  OAI211_X1 U10329 ( .C1(n9258), .C2(n9036), .A(n9008), .B(n9705), .ZN(n9010)
         );
  NOR2_X1 U10330 ( .A1(n9288), .A2(n9027), .ZN(n9009) );
  AOI211_X1 U10331 ( .C1(n9286), .C2(n9031), .A(n9010), .B(n9009), .ZN(n9011)
         );
  OAI21_X1 U10332 ( .B1(n9012), .B2(n4371), .A(n9011), .ZN(P1_U3236) );
  NAND3_X1 U10333 ( .A1(n9019), .A2(n9018), .A3(n9017), .ZN(n9026) );
  INV_X1 U10334 ( .A(n9020), .ZN(n9165) );
  AOI22_X1 U10335 ( .A1(n9173), .A2(n9021), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9022) );
  OAI21_X1 U10336 ( .B1(n9044), .B2(n9023), .A(n9022), .ZN(n9024) );
  AOI21_X1 U10337 ( .B1(n9165), .B2(n9031), .A(n9024), .ZN(n9025) );
  OAI211_X1 U10338 ( .C1(n9167), .C2(n9027), .A(n9026), .B(n9025), .ZN(
        P1_U3238) );
  NAND2_X1 U10339 ( .A1(n4692), .A2(n9028), .ZN(n9030) );
  XNOR2_X1 U10340 ( .A(n9030), .B(n9029), .ZN(n9040) );
  NAND2_X1 U10341 ( .A1(n9031), .A2(n9339), .ZN(n9035) );
  AOI21_X1 U10342 ( .B1(n9033), .B2(n9373), .A(n9032), .ZN(n9034) );
  OAI211_X1 U10343 ( .C1(n9329), .C2(n9036), .A(n9035), .B(n9034), .ZN(n9037)
         );
  AOI21_X1 U10344 ( .B1(n9465), .B2(n9038), .A(n9037), .ZN(n9039) );
  OAI21_X1 U10345 ( .B1(n9040), .B2(n4371), .A(n9039), .ZN(P1_U3239) );
  MUX2_X1 U10346 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9041), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10347 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9042), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10348 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9043), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9173), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10350 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9186), .S(P1_U4006), .Z(
        P1_U3581) );
  INV_X1 U10351 ( .A(n9044), .ZN(n9199) );
  MUX2_X1 U10352 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9199), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10353 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9218), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10354 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9234), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10355 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9217), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10356 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9235), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10357 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9276), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10358 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9295), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10359 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9309), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10360 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9294), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10361 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9308), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10362 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9354), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9373), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10364 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9353), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10365 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9374), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10366 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9545), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9045), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9546), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10369 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9046), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10370 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9047), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10371 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n4681), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10372 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9048), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9049), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10374 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9050), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10375 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6818), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10376 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6544), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9719), .S(P1_U4006), .Z(
        P1_U3555) );
  OAI21_X1 U10378 ( .B1(n9052), .B2(n4318), .A(n9051), .ZN(n9053) );
  NAND2_X1 U10379 ( .A1(n9053), .A2(n9702), .ZN(n9063) );
  NOR2_X1 U10380 ( .A1(n9641), .A2(n9054), .ZN(n9055) );
  AOI211_X1 U10381 ( .C1(n9711), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9056), .B(
        n9055), .ZN(n9062) );
  OAI21_X1 U10382 ( .B1(n9059), .B2(n9058), .A(n9057), .ZN(n9060) );
  NAND2_X1 U10383 ( .A1(n9060), .A2(n9712), .ZN(n9061) );
  NAND3_X1 U10384 ( .A1(n9063), .A2(n9062), .A3(n9061), .ZN(P1_U3252) );
  NOR2_X1 U10385 ( .A1(n9064), .A2(n9071), .ZN(n9066) );
  NAND2_X1 U10386 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9089), .ZN(n9067) );
  OAI21_X1 U10387 ( .B1(n9089), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9067), .ZN(
        n9068) );
  AOI211_X1 U10388 ( .C1(n9069), .C2(n9068), .A(n9088), .B(n9688), .ZN(n9081)
         );
  NOR2_X1 U10389 ( .A1(n9071), .A2(n9070), .ZN(n9073) );
  NOR2_X1 U10390 ( .A1(n9073), .A2(n9072), .ZN(n9075) );
  XNOR2_X1 U10391 ( .A(n9089), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9074) );
  NOR2_X1 U10392 ( .A1(n9075), .A2(n9074), .ZN(n9082) );
  AOI211_X1 U10393 ( .C1(n9075), .C2(n9074), .A(n9082), .B(n9648), .ZN(n9080)
         );
  NAND2_X1 U10394 ( .A1(n9711), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U10395 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n9076) );
  OAI211_X1 U10396 ( .C1(n9641), .C2(n9078), .A(n9077), .B(n9076), .ZN(n9079)
         );
  OR3_X1 U10397 ( .A1(n9081), .A2(n9080), .A3(n9079), .ZN(P1_U3257) );
  INV_X1 U10398 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9096) );
  XNOR2_X1 U10399 ( .A(n9104), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9084) );
  AOI21_X1 U10400 ( .B1(n9089), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9082), .ZN(
        n9083) );
  NOR2_X1 U10401 ( .A1(n9083), .A2(n9084), .ZN(n9103) );
  AOI21_X1 U10402 ( .B1(n9084), .B2(n9083), .A(n9103), .ZN(n9085) );
  NAND2_X1 U10403 ( .A1(n9712), .A2(n9085), .ZN(n9087) );
  NAND2_X1 U10404 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9086) );
  NAND2_X1 U10405 ( .A1(n9087), .A2(n9086), .ZN(n9094) );
  NAND2_X1 U10406 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9104), .ZN(n9090) );
  OAI21_X1 U10407 ( .B1(n9104), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9090), .ZN(
        n9091) );
  AOI211_X1 U10408 ( .C1(n9092), .C2(n9091), .A(n9097), .B(n9688), .ZN(n9093)
         );
  AOI211_X1 U10409 ( .C1(n9704), .C2(n9104), .A(n9094), .B(n9093), .ZN(n9095)
         );
  OAI21_X1 U10410 ( .B1(n9112), .B2(n9096), .A(n9095), .ZN(P1_U3258) );
  AOI21_X1 U10411 ( .B1(n9104), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9097), .ZN(
        n9699) );
  OR2_X1 U10412 ( .A1(n9703), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9099) );
  NAND2_X1 U10413 ( .A1(n9703), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U10414 ( .A1(n9099), .A2(n9098), .ZN(n9700) );
  NOR2_X1 U10415 ( .A1(n9699), .A2(n9700), .ZN(n9698) );
  AOI21_X1 U10416 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9703), .A(n9698), .ZN(
        n9100) );
  XNOR2_X1 U10417 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9100), .ZN(n9109) );
  AOI22_X1 U10418 ( .A1(n9703), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9102), .B2(
        n9101), .ZN(n9710) );
  AOI21_X1 U10419 ( .B1(n9104), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9103), .ZN(
        n9709) );
  NAND2_X1 U10420 ( .A1(n9710), .A2(n9709), .ZN(n9708) );
  OAI21_X1 U10421 ( .B1(n9703), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9708), .ZN(
        n9106) );
  INV_X1 U10422 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9105) );
  XOR2_X1 U10423 ( .A(n9106), .B(n9105), .Z(n9107) );
  AOI22_X1 U10424 ( .A1(n9109), .A2(n9702), .B1(n9712), .B2(n9107), .ZN(n9111)
         );
  INV_X1 U10425 ( .A(n9107), .ZN(n9110) );
  NAND2_X1 U10426 ( .A1(n9387), .A2(n9346), .ZN(n9116) );
  NAND2_X1 U10427 ( .A1(n9114), .A2(n9113), .ZN(n9392) );
  NOR2_X1 U10428 ( .A1(n9743), .A2(n9392), .ZN(n9120) );
  AOI21_X1 U10429 ( .B1(n9743), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9120), .ZN(
        n9115) );
  OAI211_X1 U10430 ( .C1(n9389), .C2(n9341), .A(n9116), .B(n9115), .ZN(
        P1_U3261) );
  INV_X1 U10431 ( .A(n9117), .ZN(n9119) );
  NAND2_X1 U10432 ( .A1(n9119), .A2(n9118), .ZN(n9391) );
  NAND3_X1 U10433 ( .A1(n9391), .A2(n9346), .A3(n9390), .ZN(n9122) );
  AOI21_X1 U10434 ( .B1(n9743), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9120), .ZN(
        n9121) );
  OAI211_X1 U10435 ( .C1(n9394), .C2(n9341), .A(n9122), .B(n9121), .ZN(
        P1_U3262) );
  OAI21_X1 U10436 ( .B1(n9125), .B2(n9124), .A(n9123), .ZN(n9404) );
  AOI22_X1 U10437 ( .A1(n9401), .A2(n9551), .B1(n9743), .B2(
        P1_REG2_REG_28__SCAN_IN), .ZN(n9145) );
  OAI21_X1 U10438 ( .B1(n9128), .B2(n9127), .A(n9126), .ZN(n9129) );
  INV_X1 U10439 ( .A(n9129), .ZN(n9135) );
  NOR2_X1 U10440 ( .A1(n9130), .A2(n9330), .ZN(n9133) );
  NOR2_X1 U10441 ( .A1(n9131), .A2(n9328), .ZN(n9132) );
  INV_X1 U10442 ( .A(n9136), .ZN(n9403) );
  INV_X1 U10443 ( .A(n9147), .ZN(n9139) );
  INV_X1 U10444 ( .A(n9137), .ZN(n9138) );
  AOI211_X1 U10445 ( .C1(n9401), .C2(n9139), .A(n9767), .B(n9138), .ZN(n9400)
         );
  NAND2_X1 U10446 ( .A1(n9400), .A2(n9204), .ZN(n9140) );
  OAI211_X1 U10447 ( .C1(n9142), .C2(n9141), .A(n9403), .B(n9140), .ZN(n9143)
         );
  NAND2_X1 U10448 ( .A1(n9143), .A2(n9740), .ZN(n9144) );
  OAI211_X1 U10449 ( .C1(n9404), .C2(n9365), .A(n9145), .B(n9144), .ZN(
        P1_U3263) );
  XOR2_X1 U10450 ( .A(n9155), .B(n9146), .Z(n9409) );
  INV_X1 U10451 ( .A(n9163), .ZN(n9148) );
  AOI21_X1 U10452 ( .B1(n9405), .B2(n9148), .A(n9147), .ZN(n9406) );
  AOI22_X1 U10453 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(n9743), .B1(n9149), .B2(
        n9728), .ZN(n9150) );
  OAI21_X1 U10454 ( .B1(n9151), .B2(n9341), .A(n9150), .ZN(n9159) );
  NOR2_X1 U10455 ( .A1(n9152), .A2(n9328), .ZN(n9157) );
  AOI211_X1 U10456 ( .C1(n9155), .C2(n9154), .A(n9318), .B(n9153), .ZN(n9156)
         );
  NOR2_X1 U10457 ( .A1(n9408), .A2(n9743), .ZN(n9158) );
  AOI211_X1 U10458 ( .C1(n9346), .C2(n9406), .A(n9159), .B(n9158), .ZN(n9160)
         );
  OAI21_X1 U10459 ( .B1(n9409), .B2(n9365), .A(n9160), .ZN(P1_U3264) );
  XNOR2_X1 U10460 ( .A(n9162), .B(n9161), .ZN(n9414) );
  INV_X1 U10461 ( .A(n9179), .ZN(n9164) );
  AOI21_X1 U10462 ( .B1(n9410), .B2(n9164), .A(n9163), .ZN(n9411) );
  AOI22_X1 U10463 ( .A1(n9743), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9165), .B2(
        n9728), .ZN(n9166) );
  OAI21_X1 U10464 ( .B1(n9167), .B2(n9341), .A(n9166), .ZN(n9176) );
  INV_X1 U10465 ( .A(n9168), .ZN(n9169) );
  NOR2_X1 U10466 ( .A1(n9170), .A2(n9169), .ZN(n9172) );
  XNOR2_X1 U10467 ( .A(n9172), .B(n9171), .ZN(n9174) );
  AOI222_X1 U10468 ( .A1(n9725), .A2(n9174), .B1(n9173), .B2(n9721), .C1(n9199), .C2(n9720), .ZN(n9413) );
  NOR2_X1 U10469 ( .A1(n9413), .A2(n9743), .ZN(n9175) );
  AOI211_X1 U10470 ( .C1(n9346), .C2(n9411), .A(n9176), .B(n9175), .ZN(n9177)
         );
  OAI21_X1 U10471 ( .B1(n9365), .B2(n9414), .A(n9177), .ZN(P1_U3265) );
  XOR2_X1 U10472 ( .A(n9178), .B(n9184), .Z(n9419) );
  AOI21_X1 U10473 ( .B1(n9415), .B2(n9201), .A(n9179), .ZN(n9416) );
  AOI22_X1 U10474 ( .A1(n9743), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9180), .B2(
        n9728), .ZN(n9181) );
  OAI21_X1 U10475 ( .B1(n9182), .B2(n9341), .A(n9181), .ZN(n9189) );
  NOR2_X1 U10476 ( .A1(n9193), .A2(n9183), .ZN(n9185) );
  XNOR2_X1 U10477 ( .A(n9185), .B(n9184), .ZN(n9187) );
  AOI222_X1 U10478 ( .A1(n9725), .A2(n9187), .B1(n9186), .B2(n9721), .C1(n9218), .C2(n9720), .ZN(n9418) );
  NOR2_X1 U10479 ( .A1(n9418), .A2(n9743), .ZN(n9188) );
  AOI211_X1 U10480 ( .C1(n9416), .C2(n9346), .A(n9189), .B(n9188), .ZN(n9190)
         );
  OAI21_X1 U10481 ( .B1(n9419), .B2(n9365), .A(n9190), .ZN(P1_U3266) );
  XNOR2_X1 U10482 ( .A(n9191), .B(n9194), .ZN(n9424) );
  NOR2_X1 U10483 ( .A1(n9192), .A2(n9341), .ZN(n9207) );
  INV_X1 U10484 ( .A(n9193), .ZN(n9198) );
  OAI21_X1 U10485 ( .B1(n9196), .B2(n9195), .A(n9194), .ZN(n9197) );
  NAND2_X1 U10486 ( .A1(n9198), .A2(n9197), .ZN(n9200) );
  AOI222_X1 U10487 ( .A1(n9725), .A2(n9200), .B1(n9199), .B2(n9721), .C1(n9234), .C2(n9720), .ZN(n9423) );
  INV_X1 U10488 ( .A(n9201), .ZN(n9202) );
  AOI211_X1 U10489 ( .C1(n9421), .C2(n9210), .A(n9767), .B(n9202), .ZN(n9420)
         );
  AOI22_X1 U10490 ( .A1(n9420), .A2(n9204), .B1(n9728), .B2(n9203), .ZN(n9205)
         );
  AOI21_X1 U10491 ( .B1(n9423), .B2(n9205), .A(n9743), .ZN(n9206) );
  AOI211_X1 U10492 ( .C1(n9743), .C2(P1_REG2_REG_24__SCAN_IN), .A(n9207), .B(
        n9206), .ZN(n9208) );
  OAI21_X1 U10493 ( .B1(n9365), .B2(n9424), .A(n9208), .ZN(P1_U3267) );
  XNOR2_X1 U10494 ( .A(n9209), .B(n9216), .ZN(n9429) );
  INV_X1 U10495 ( .A(n9210), .ZN(n9211) );
  AOI21_X1 U10496 ( .B1(n9425), .B2(n9224), .A(n9211), .ZN(n9426) );
  INV_X1 U10497 ( .A(n9212), .ZN(n9213) );
  AOI22_X1 U10498 ( .A1(n9743), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9213), .B2(
        n9728), .ZN(n9214) );
  OAI21_X1 U10499 ( .B1(n4452), .B2(n9341), .A(n9214), .ZN(n9221) );
  XOR2_X1 U10500 ( .A(n9216), .B(n9215), .Z(n9219) );
  AOI222_X1 U10501 ( .A1(n9725), .A2(n9219), .B1(n9218), .B2(n9721), .C1(n9217), .C2(n9720), .ZN(n9428) );
  NOR2_X1 U10502 ( .A1(n9428), .A2(n9743), .ZN(n9220) );
  AOI211_X1 U10503 ( .C1(n9426), .C2(n9346), .A(n9221), .B(n9220), .ZN(n9222)
         );
  OAI21_X1 U10504 ( .B1(n9429), .B2(n9365), .A(n9222), .ZN(P1_U3268) );
  XOR2_X1 U10505 ( .A(n9232), .B(n9223), .Z(n9434) );
  INV_X1 U10506 ( .A(n9246), .ZN(n9226) );
  INV_X1 U10507 ( .A(n9224), .ZN(n9225) );
  AOI21_X1 U10508 ( .B1(n9430), .B2(n9226), .A(n9225), .ZN(n9431) );
  INV_X1 U10509 ( .A(n9227), .ZN(n9228) );
  AOI22_X1 U10510 ( .A1(n9743), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9228), .B2(
        n9728), .ZN(n9229) );
  OAI21_X1 U10511 ( .B1(n9230), .B2(n9341), .A(n9229), .ZN(n9238) );
  NOR2_X1 U10512 ( .A1(n4312), .A2(n9231), .ZN(n9233) );
  XNOR2_X1 U10513 ( .A(n9233), .B(n9232), .ZN(n9236) );
  AOI222_X1 U10514 ( .A1(n9725), .A2(n9236), .B1(n9235), .B2(n9720), .C1(n9234), .C2(n9721), .ZN(n9433) );
  NOR2_X1 U10515 ( .A1(n9433), .A2(n9743), .ZN(n9237) );
  AOI211_X1 U10516 ( .C1(n9431), .C2(n9346), .A(n9238), .B(n9237), .ZN(n9239)
         );
  OAI21_X1 U10517 ( .B1(n9434), .B2(n9365), .A(n9239), .ZN(P1_U3269) );
  XNOR2_X1 U10518 ( .A(n9240), .B(n9242), .ZN(n9439) );
  AOI21_X1 U10519 ( .B1(n9242), .B2(n9241), .A(n4312), .ZN(n9243) );
  OAI222_X1 U10520 ( .A1(n9330), .A2(n9245), .B1(n9328), .B2(n9244), .C1(n9318), .C2(n9243), .ZN(n9435) );
  INV_X1 U10521 ( .A(n9260), .ZN(n9247) );
  AOI211_X1 U10522 ( .C1(n9437), .C2(n9247), .A(n9767), .B(n9246), .ZN(n9436)
         );
  NAND2_X1 U10523 ( .A1(n9436), .A2(n9557), .ZN(n9250) );
  AOI22_X1 U10524 ( .A1(n9743), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9248), .B2(
        n9728), .ZN(n9249) );
  OAI211_X1 U10525 ( .C1(n9251), .C2(n9341), .A(n9250), .B(n9249), .ZN(n9252)
         );
  AOI21_X1 U10526 ( .B1(n9435), .B2(n9740), .A(n9252), .ZN(n9253) );
  OAI21_X1 U10527 ( .B1(n9439), .B2(n9365), .A(n9253), .ZN(P1_U3270) );
  XNOR2_X1 U10528 ( .A(n9254), .B(n9255), .ZN(n9444) );
  XNOR2_X1 U10529 ( .A(n9256), .B(n9255), .ZN(n9257) );
  OAI222_X1 U10530 ( .A1(n9328), .A2(n9259), .B1(n9330), .B2(n9258), .C1(n9257), .C2(n9318), .ZN(n9440) );
  AOI211_X1 U10531 ( .C1(n9442), .C2(n9268), .A(n9767), .B(n9260), .ZN(n9441)
         );
  NAND2_X1 U10532 ( .A1(n9441), .A2(n9557), .ZN(n9263) );
  AOI22_X1 U10533 ( .A1(n9743), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9261), .B2(
        n9728), .ZN(n9262) );
  OAI211_X1 U10534 ( .C1(n9264), .C2(n9341), .A(n9263), .B(n9262), .ZN(n9265)
         );
  AOI21_X1 U10535 ( .B1(n9440), .B2(n9740), .A(n9265), .ZN(n9266) );
  OAI21_X1 U10536 ( .B1(n9444), .B2(n9365), .A(n9266), .ZN(P1_U3271) );
  XNOR2_X1 U10537 ( .A(n9267), .B(n9275), .ZN(n9449) );
  INV_X1 U10538 ( .A(n9268), .ZN(n9269) );
  AOI211_X1 U10539 ( .C1(n9446), .C2(n9283), .A(n9767), .B(n9269), .ZN(n9445)
         );
  AOI22_X1 U10540 ( .A1(n9743), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9270), .B2(
        n9728), .ZN(n9271) );
  OAI21_X1 U10541 ( .B1(n9272), .B2(n9341), .A(n9271), .ZN(n9279) );
  OAI21_X1 U10542 ( .B1(n9275), .B2(n9274), .A(n9273), .ZN(n9277) );
  AOI222_X1 U10543 ( .A1(n9725), .A2(n9277), .B1(n9276), .B2(n9721), .C1(n9309), .C2(n9720), .ZN(n9448) );
  NOR2_X1 U10544 ( .A1(n9448), .A2(n9743), .ZN(n9278) );
  AOI211_X1 U10545 ( .C1(n9445), .C2(n9557), .A(n9279), .B(n9278), .ZN(n9280)
         );
  OAI21_X1 U10546 ( .B1(n9365), .B2(n9449), .A(n9280), .ZN(P1_U3272) );
  XNOR2_X1 U10547 ( .A(n9282), .B(n9281), .ZN(n9454) );
  INV_X1 U10548 ( .A(n9301), .ZN(n9285) );
  INV_X1 U10549 ( .A(n9283), .ZN(n9284) );
  AOI21_X1 U10550 ( .B1(n9450), .B2(n9285), .A(n9284), .ZN(n9451) );
  AOI22_X1 U10551 ( .A1(n9743), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9286), .B2(
        n9728), .ZN(n9287) );
  OAI21_X1 U10552 ( .B1(n9288), .B2(n9341), .A(n9287), .ZN(n9298) );
  INV_X1 U10553 ( .A(n9289), .ZN(n9290) );
  AOI21_X1 U10554 ( .B1(n9306), .B2(n9291), .A(n9290), .ZN(n9293) );
  XNOR2_X1 U10555 ( .A(n9293), .B(n9292), .ZN(n9296) );
  AOI222_X1 U10556 ( .A1(n9725), .A2(n9296), .B1(n9295), .B2(n9721), .C1(n9294), .C2(n9720), .ZN(n9453) );
  NOR2_X1 U10557 ( .A1(n9453), .A2(n9743), .ZN(n9297) );
  AOI211_X1 U10558 ( .C1(n9451), .C2(n9346), .A(n9298), .B(n9297), .ZN(n9299)
         );
  OAI21_X1 U10559 ( .B1(n9365), .B2(n9454), .A(n9299), .ZN(P1_U3273) );
  XNOR2_X1 U10560 ( .A(n9300), .B(n9307), .ZN(n9459) );
  INV_X1 U10561 ( .A(n9321), .ZN(n9302) );
  AOI21_X1 U10562 ( .B1(n9455), .B2(n9302), .A(n9301), .ZN(n9456) );
  AOI22_X1 U10563 ( .A1(n9743), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9303), .B2(
        n9728), .ZN(n9304) );
  OAI21_X1 U10564 ( .B1(n9305), .B2(n9341), .A(n9304), .ZN(n9312) );
  XOR2_X1 U10565 ( .A(n9307), .B(n9306), .Z(n9310) );
  AOI222_X1 U10566 ( .A1(n9725), .A2(n9310), .B1(n9309), .B2(n9721), .C1(n9308), .C2(n9720), .ZN(n9458) );
  NOR2_X1 U10567 ( .A1(n9458), .A2(n9743), .ZN(n9311) );
  AOI211_X1 U10568 ( .C1(n9456), .C2(n9346), .A(n9312), .B(n9311), .ZN(n9313)
         );
  OAI21_X1 U10569 ( .B1(n9365), .B2(n9459), .A(n9313), .ZN(P1_U3274) );
  XNOR2_X1 U10570 ( .A(n9314), .B(n9315), .ZN(n9464) );
  XNOR2_X1 U10571 ( .A(n9316), .B(n9315), .ZN(n9317) );
  OAI222_X1 U10572 ( .A1(n9328), .A2(n9320), .B1(n9330), .B2(n9319), .C1(n9318), .C2(n9317), .ZN(n9460) );
  AOI211_X1 U10573 ( .C1(n9462), .C2(n9337), .A(n9767), .B(n9321), .ZN(n9461)
         );
  NAND2_X1 U10574 ( .A1(n9461), .A2(n9557), .ZN(n9324) );
  AOI22_X1 U10575 ( .A1(n9743), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9322), .B2(
        n9728), .ZN(n9323) );
  OAI211_X1 U10576 ( .C1(n4449), .C2(n9341), .A(n9324), .B(n9323), .ZN(n9325)
         );
  AOI21_X1 U10577 ( .B1(n9460), .B2(n9740), .A(n9325), .ZN(n9326) );
  OAI21_X1 U10578 ( .B1(n9464), .B2(n9365), .A(n9326), .ZN(P1_U3275) );
  XNOR2_X1 U10579 ( .A(n9327), .B(n9332), .ZN(n9336) );
  OAI22_X1 U10580 ( .A1(n9331), .A2(n9330), .B1(n9329), .B2(n9328), .ZN(n9335)
         );
  XNOR2_X1 U10581 ( .A(n9333), .B(n9332), .ZN(n9469) );
  NOR2_X1 U10582 ( .A1(n9469), .A2(n9723), .ZN(n9334) );
  AOI211_X1 U10583 ( .C1(n9725), .C2(n9336), .A(n9335), .B(n9334), .ZN(n9468)
         );
  INV_X1 U10584 ( .A(n9337), .ZN(n9338) );
  AOI21_X1 U10585 ( .B1(n9465), .B2(n9357), .A(n9338), .ZN(n9466) );
  AOI22_X1 U10586 ( .A1(n9743), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9339), .B2(
        n9728), .ZN(n9340) );
  OAI21_X1 U10587 ( .B1(n9342), .B2(n9341), .A(n9340), .ZN(n9345) );
  NOR2_X1 U10588 ( .A1(n9469), .A2(n9343), .ZN(n9344) );
  AOI211_X1 U10589 ( .C1(n9466), .C2(n9346), .A(n9345), .B(n9344), .ZN(n9347)
         );
  OAI21_X1 U10590 ( .B1(n9468), .B2(n9743), .A(n9347), .ZN(P1_U3276) );
  XNOR2_X1 U10591 ( .A(n9348), .B(n9349), .ZN(n9596) );
  INV_X1 U10592 ( .A(n9596), .ZN(n9366) );
  INV_X1 U10593 ( .A(n9349), .ZN(n9350) );
  XNOR2_X1 U10594 ( .A(n9351), .B(n9350), .ZN(n9352) );
  NAND2_X1 U10595 ( .A1(n9352), .A2(n9725), .ZN(n9356) );
  AOI22_X1 U10596 ( .A1(n9721), .A2(n9354), .B1(n9353), .B2(n9720), .ZN(n9355)
         );
  NAND2_X1 U10597 ( .A1(n9356), .A2(n9355), .ZN(n9594) );
  OAI211_X1 U10598 ( .C1(n9379), .C2(n9592), .A(n9357), .B(n9554), .ZN(n9591)
         );
  AOI22_X1 U10599 ( .A1(n9743), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9358), .B2(
        n9728), .ZN(n9361) );
  NAND2_X1 U10600 ( .A1(n9359), .A2(n9551), .ZN(n9360) );
  OAI211_X1 U10601 ( .C1(n9591), .C2(n9362), .A(n9361), .B(n9360), .ZN(n9363)
         );
  AOI21_X1 U10602 ( .B1(n9594), .B2(n9740), .A(n9363), .ZN(n9364) );
  OAI21_X1 U10603 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(P1_U3277) );
  XNOR2_X1 U10604 ( .A(n9367), .B(n4587), .ZN(n9474) );
  NAND2_X1 U10605 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  NAND2_X1 U10606 ( .A1(n9371), .A2(n9370), .ZN(n9372) );
  NAND2_X1 U10607 ( .A1(n9372), .A2(n9725), .ZN(n9376) );
  AOI22_X1 U10608 ( .A1(n9374), .A2(n9720), .B1(n9721), .B2(n9373), .ZN(n9375)
         );
  NAND2_X1 U10609 ( .A1(n9376), .A2(n9375), .ZN(n9377) );
  AOI21_X1 U10610 ( .B1(n9474), .B2(n9549), .A(n9377), .ZN(n9476) );
  AND2_X1 U10611 ( .A1(n9378), .A2(n9470), .ZN(n9380) );
  OR2_X1 U10612 ( .A1(n9380), .A2(n9379), .ZN(n9472) );
  AOI22_X1 U10613 ( .A1(n9743), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9381), .B2(
        n9728), .ZN(n9383) );
  NAND2_X1 U10614 ( .A1(n9551), .A2(n9470), .ZN(n9382) );
  OAI211_X1 U10615 ( .C1(n9472), .C2(n9384), .A(n9383), .B(n9382), .ZN(n9385)
         );
  AOI21_X1 U10616 ( .B1(n9474), .B2(n9558), .A(n9385), .ZN(n9386) );
  OAI21_X1 U10617 ( .B1(n9476), .B2(n9743), .A(n9386), .ZN(P1_U3278) );
  NAND2_X1 U10618 ( .A1(n9387), .A2(n9554), .ZN(n9388) );
  OAI211_X1 U10619 ( .C1(n9389), .C2(n9765), .A(n9388), .B(n9392), .ZN(n9493)
         );
  MUX2_X1 U10620 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9493), .S(n9782), .Z(
        P1_U3554) );
  NAND3_X1 U10621 ( .A1(n9391), .A2(n9554), .A3(n9390), .ZN(n9393) );
  OAI211_X1 U10622 ( .C1(n9394), .C2(n9765), .A(n9393), .B(n9392), .ZN(n9494)
         );
  MUX2_X1 U10623 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9494), .S(n9782), .Z(
        P1_U3553) );
  AOI21_X1 U10624 ( .B1(n9487), .B2(n9396), .A(n9395), .ZN(n9397) );
  OAI211_X1 U10625 ( .C1(n9399), .C2(n9562), .A(n9398), .B(n9397), .ZN(n9495)
         );
  MUX2_X1 U10626 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9495), .S(n9782), .Z(
        P1_U3552) );
  AOI21_X1 U10627 ( .B1(n9487), .B2(n9401), .A(n9400), .ZN(n9402) );
  OAI211_X1 U10628 ( .C1(n9404), .C2(n9562), .A(n9403), .B(n9402), .ZN(n9496)
         );
  MUX2_X1 U10629 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9496), .S(n9782), .Z(
        P1_U3551) );
  AOI22_X1 U10630 ( .A1(n9406), .A2(n9554), .B1(n9487), .B2(n9405), .ZN(n9407)
         );
  OAI211_X1 U10631 ( .C1(n9409), .C2(n9562), .A(n9408), .B(n9407), .ZN(n9497)
         );
  MUX2_X1 U10632 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9497), .S(n9782), .Z(
        P1_U3550) );
  AOI22_X1 U10633 ( .A1(n9411), .A2(n9554), .B1(n9487), .B2(n9410), .ZN(n9412)
         );
  OAI211_X1 U10634 ( .C1(n9414), .C2(n9562), .A(n9413), .B(n9412), .ZN(n9498)
         );
  MUX2_X1 U10635 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9498), .S(n9782), .Z(
        P1_U3549) );
  AOI22_X1 U10636 ( .A1(n9416), .A2(n9554), .B1(n9487), .B2(n9415), .ZN(n9417)
         );
  OAI211_X1 U10637 ( .C1(n9419), .C2(n9562), .A(n9418), .B(n9417), .ZN(n9499)
         );
  MUX2_X1 U10638 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9499), .S(n9782), .Z(
        P1_U3548) );
  AOI21_X1 U10639 ( .B1(n9487), .B2(n9421), .A(n9420), .ZN(n9422) );
  OAI211_X1 U10640 ( .C1(n9424), .C2(n9562), .A(n9423), .B(n9422), .ZN(n9500)
         );
  MUX2_X1 U10641 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9500), .S(n9782), .Z(
        P1_U3547) );
  AOI22_X1 U10642 ( .A1(n9426), .A2(n9554), .B1(n9487), .B2(n9425), .ZN(n9427)
         );
  OAI211_X1 U10643 ( .C1(n9429), .C2(n9562), .A(n9428), .B(n9427), .ZN(n9501)
         );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9501), .S(n9782), .Z(
        P1_U3546) );
  AOI22_X1 U10645 ( .A1(n9431), .A2(n9554), .B1(n9487), .B2(n9430), .ZN(n9432)
         );
  OAI211_X1 U10646 ( .C1(n9434), .C2(n9562), .A(n9433), .B(n9432), .ZN(n9502)
         );
  MUX2_X1 U10647 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9502), .S(n9782), .Z(
        P1_U3545) );
  AOI211_X1 U10648 ( .C1(n9487), .C2(n9437), .A(n9436), .B(n9435), .ZN(n9438)
         );
  OAI21_X1 U10649 ( .B1(n9562), .B2(n9439), .A(n9438), .ZN(n9503) );
  MUX2_X1 U10650 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9503), .S(n9782), .Z(
        P1_U3544) );
  AOI211_X1 U10651 ( .C1(n9487), .C2(n9442), .A(n9441), .B(n9440), .ZN(n9443)
         );
  OAI21_X1 U10652 ( .B1(n9444), .B2(n9562), .A(n9443), .ZN(n9504) );
  MUX2_X1 U10653 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9504), .S(n9782), .Z(
        P1_U3543) );
  AOI21_X1 U10654 ( .B1(n9487), .B2(n9446), .A(n9445), .ZN(n9447) );
  OAI211_X1 U10655 ( .C1(n9449), .C2(n9562), .A(n9448), .B(n9447), .ZN(n9505)
         );
  MUX2_X1 U10656 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9505), .S(n9782), .Z(
        P1_U3542) );
  AOI22_X1 U10657 ( .A1(n9451), .A2(n9554), .B1(n9487), .B2(n9450), .ZN(n9452)
         );
  OAI211_X1 U10658 ( .C1(n9454), .C2(n9562), .A(n9453), .B(n9452), .ZN(n9506)
         );
  MUX2_X1 U10659 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9506), .S(n9782), .Z(
        P1_U3541) );
  AOI22_X1 U10660 ( .A1(n9456), .A2(n9554), .B1(n9487), .B2(n9455), .ZN(n9457)
         );
  OAI211_X1 U10661 ( .C1(n9459), .C2(n9562), .A(n9458), .B(n9457), .ZN(n9507)
         );
  MUX2_X1 U10662 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9507), .S(n9782), .Z(
        P1_U3540) );
  AOI211_X1 U10663 ( .C1(n9487), .C2(n9462), .A(n9461), .B(n9460), .ZN(n9463)
         );
  OAI21_X1 U10664 ( .B1(n9562), .B2(n9464), .A(n9463), .ZN(n9508) );
  MUX2_X1 U10665 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9508), .S(n9782), .Z(
        P1_U3539) );
  AOI22_X1 U10666 ( .A1(n9466), .A2(n9554), .B1(n9487), .B2(n9465), .ZN(n9467)
         );
  OAI211_X1 U10667 ( .C1(n9469), .C2(n9491), .A(n9468), .B(n9467), .ZN(n9509)
         );
  MUX2_X1 U10668 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9509), .S(n9782), .Z(
        P1_U3538) );
  INV_X1 U10669 ( .A(n9470), .ZN(n9471) );
  OAI22_X1 U10670 ( .A1(n9472), .A2(n9767), .B1(n9471), .B2(n9765), .ZN(n9473)
         );
  AOI21_X1 U10671 ( .B1(n9474), .B2(n9772), .A(n9473), .ZN(n9475) );
  AND2_X1 U10672 ( .A1(n9476), .A2(n9475), .ZN(n9510) );
  MUX2_X1 U10673 ( .A(n7057), .B(n9510), .S(n9782), .Z(n9477) );
  INV_X1 U10674 ( .A(n9477), .ZN(P1_U3536) );
  AND2_X1 U10675 ( .A1(n9478), .A2(n9772), .ZN(n9483) );
  INV_X1 U10676 ( .A(n9479), .ZN(n9480) );
  OAI22_X1 U10677 ( .A1(n9481), .A2(n9767), .B1(n9480), .B2(n9765), .ZN(n9482)
         );
  MUX2_X1 U10678 ( .A(n9513), .B(P1_REG1_REG_11__SCAN_IN), .S(n9779), .Z(
        P1_U3534) );
  INV_X1 U10679 ( .A(n9485), .ZN(n9492) );
  AOI22_X1 U10680 ( .A1(n9488), .A2(n9554), .B1(n9487), .B2(n9486), .ZN(n9489)
         );
  OAI211_X1 U10681 ( .C1(n9492), .C2(n9491), .A(n9490), .B(n9489), .ZN(n9514)
         );
  MUX2_X1 U10682 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9514), .S(n9782), .Z(
        P1_U3532) );
  MUX2_X1 U10683 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9493), .S(n9774), .Z(
        P1_U3522) );
  MUX2_X1 U10684 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9494), .S(n9774), .Z(
        P1_U3521) );
  MUX2_X1 U10685 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9495), .S(n9774), .Z(
        P1_U3520) );
  MUX2_X1 U10686 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9496), .S(n9774), .Z(
        P1_U3519) );
  MUX2_X1 U10687 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9497), .S(n9774), .Z(
        P1_U3518) );
  MUX2_X1 U10688 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9498), .S(n9774), .Z(
        P1_U3517) );
  MUX2_X1 U10689 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9499), .S(n9774), .Z(
        P1_U3516) );
  MUX2_X1 U10690 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9500), .S(n9774), .Z(
        P1_U3515) );
  MUX2_X1 U10691 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9501), .S(n9774), .Z(
        P1_U3514) );
  MUX2_X1 U10692 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9502), .S(n9774), .Z(
        P1_U3513) );
  MUX2_X1 U10693 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9503), .S(n9774), .Z(
        P1_U3512) );
  MUX2_X1 U10694 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9504), .S(n9774), .Z(
        P1_U3511) );
  MUX2_X1 U10695 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9505), .S(n9774), .Z(
        P1_U3510) );
  MUX2_X1 U10696 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9506), .S(n9774), .Z(
        P1_U3508) );
  MUX2_X1 U10697 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9507), .S(n9774), .Z(
        P1_U3505) );
  MUX2_X1 U10698 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9508), .S(n9774), .Z(
        P1_U3502) );
  MUX2_X1 U10699 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9509), .S(n9774), .Z(
        P1_U3499) );
  INV_X1 U10700 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9511) );
  MUX2_X1 U10701 ( .A(n9511), .B(n9510), .S(n9774), .Z(n9512) );
  INV_X1 U10702 ( .A(n9512), .ZN(P1_U3493) );
  MUX2_X1 U10703 ( .A(n9513), .B(P1_REG0_REG_11__SCAN_IN), .S(n9773), .Z(
        P1_U3487) );
  MUX2_X1 U10704 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n9514), .S(n9774), .Z(
        P1_U3481) );
  MUX2_X1 U10705 ( .A(P1_D_REG_1__SCAN_IN), .B(n9516), .S(n9515), .Z(P1_U3441)
         );
  NOR4_X1 U10706 ( .A1(n9518), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9517), .ZN(n9519) );
  AOI21_X1 U10707 ( .B1(n9520), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9519), .ZN(
        n9521) );
  OAI21_X1 U10708 ( .B1(n9523), .B2(n9522), .A(n9521), .ZN(P1_U3322) );
  OAI222_X1 U10709 ( .A1(n9527), .A2(n9526), .B1(n5899), .B2(P1_U3084), .C1(
        n9525), .C2(n9524), .ZN(P1_U3324) );
  MUX2_X1 U10710 ( .A(n9528), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10711 ( .A1(n9711), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(n9529), .B2(
        n9704), .ZN(n9539) );
  OAI211_X1 U10712 ( .C1(n9532), .C2(n9531), .A(n9702), .B(n9530), .ZN(n9537)
         );
  OAI211_X1 U10713 ( .C1(n9535), .C2(n9534), .A(n9712), .B(n9533), .ZN(n9536)
         );
  NAND4_X1 U10714 ( .A1(n9539), .A2(n9538), .A3(n9537), .A4(n9536), .ZN(
        P1_U3244) );
  XNOR2_X1 U10715 ( .A(n9540), .B(n9543), .ZN(n9567) );
  NAND2_X1 U10716 ( .A1(n9542), .A2(n9541), .ZN(n9544) );
  XNOR2_X1 U10717 ( .A(n9544), .B(n9543), .ZN(n9547) );
  AOI222_X1 U10718 ( .A1(n9725), .A2(n9547), .B1(n9546), .B2(n9720), .C1(n9545), .C2(n9721), .ZN(n9564) );
  INV_X1 U10719 ( .A(n9564), .ZN(n9548) );
  AOI21_X1 U10720 ( .B1(n9549), .B2(n9567), .A(n9548), .ZN(n9561) );
  AOI222_X1 U10721 ( .A1(n9552), .A2(n9551), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n9743), .C1(n9728), .C2(n9550), .ZN(n9560) );
  OAI211_X1 U10722 ( .C1(n9555), .C2(n9565), .A(n9554), .B(n9553), .ZN(n9563)
         );
  INV_X1 U10723 ( .A(n9563), .ZN(n9556) );
  AOI22_X1 U10724 ( .A1(n9567), .A2(n9558), .B1(n9557), .B2(n9556), .ZN(n9559)
         );
  OAI211_X1 U10725 ( .C1(n9743), .C2(n9561), .A(n9560), .B(n9559), .ZN(
        P1_U3281) );
  INV_X1 U10726 ( .A(n9562), .ZN(n9595) );
  OAI211_X1 U10727 ( .C1(n9565), .C2(n9765), .A(n9564), .B(n9563), .ZN(n9566)
         );
  AOI21_X1 U10728 ( .B1(n9595), .B2(n9567), .A(n9566), .ZN(n9569) );
  AOI22_X1 U10729 ( .A1(n9774), .A2(n9569), .B1(n6115), .B2(n9773), .ZN(
        P1_U3484) );
  AOI22_X1 U10730 ( .A1(n9782), .A2(n9569), .B1(n9568), .B2(n9779), .ZN(
        P1_U3533) );
  AOI21_X1 U10731 ( .B1(n9571), .B2(n9578), .A(n9570), .ZN(n9574) );
  AOI21_X1 U10732 ( .B1(n9574), .B2(n9573), .A(n9572), .ZN(n9585) );
  AOI222_X1 U10733 ( .A1(n9576), .A2(n9805), .B1(n9575), .B2(n9821), .C1(
        P2_REG2_REG_14__SCAN_IN), .C2(n9831), .ZN(n9583) );
  OAI21_X1 U10734 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9588) );
  OAI211_X1 U10735 ( .C1(n9586), .C2(n4347), .A(n4297), .B(n9905), .ZN(n9584)
         );
  INV_X1 U10736 ( .A(n9584), .ZN(n9580) );
  AOI22_X1 U10737 ( .A1(n9588), .A2(n9581), .B1(n9812), .B2(n9580), .ZN(n9582)
         );
  OAI211_X1 U10738 ( .C1(n9831), .C2(n9585), .A(n9583), .B(n9582), .ZN(
        P2_U3282) );
  OAI211_X1 U10739 ( .C1(n9586), .C2(n9941), .A(n9585), .B(n9584), .ZN(n9587)
         );
  AOI21_X1 U10740 ( .B1(n9588), .B2(n9947), .A(n9587), .ZN(n9590) );
  AOI22_X1 U10741 ( .A1(n9967), .A2(n9590), .B1(n7813), .B2(n9965), .ZN(
        P2_U3534) );
  INV_X1 U10742 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9589) );
  AOI22_X1 U10743 ( .A1(n9951), .A2(n9590), .B1(n9589), .B2(n9949), .ZN(
        P2_U3493) );
  OAI21_X1 U10744 ( .B1(n9592), .B2(n9765), .A(n9591), .ZN(n9593) );
  AOI211_X1 U10745 ( .C1(n9596), .C2(n9595), .A(n9594), .B(n9593), .ZN(n9605)
         );
  AOI22_X1 U10746 ( .A1(n9782), .A2(n9605), .B1(n7275), .B2(n9779), .ZN(
        P1_U3537) );
  INV_X1 U10747 ( .A(n9597), .ZN(n9599) );
  OAI21_X1 U10748 ( .B1(n9599), .B2(n9765), .A(n9598), .ZN(n9600) );
  AOI21_X1 U10749 ( .B1(n9601), .B2(n9772), .A(n9600), .ZN(n9602) );
  AND2_X1 U10750 ( .A1(n9603), .A2(n9602), .ZN(n9606) );
  AOI22_X1 U10751 ( .A1(n9782), .A2(n9606), .B1(n6851), .B2(n9779), .ZN(
        P1_U3535) );
  INV_X1 U10752 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9604) );
  AOI22_X1 U10753 ( .A1(n9774), .A2(n9605), .B1(n9604), .B2(n9773), .ZN(
        P1_U3496) );
  AOI22_X1 U10754 ( .A1(n9774), .A2(n9606), .B1(n6192), .B2(n9773), .ZN(
        P1_U3490) );
  XNOR2_X1 U10755 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U10756 ( .A(P2_RD_REG_SCAN_IN), .B(n9607), .Z(U126) );
  AOI22_X1 U10757 ( .A1(n9711), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(n9608), .B2(
        n9704), .ZN(n9618) );
  OAI211_X1 U10758 ( .C1(n9619), .C2(n9610), .A(n9702), .B(n9609), .ZN(n9617)
         );
  NOR2_X1 U10759 ( .A1(n4431), .A2(n9611), .ZN(n9614) );
  OAI211_X1 U10760 ( .C1(n9614), .C2(n9613), .A(n9712), .B(n9612), .ZN(n9616)
         );
  NAND2_X1 U10761 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n9615) );
  NAND4_X1 U10762 ( .A1(n9618), .A2(n9617), .A3(n9616), .A4(n9615), .ZN(
        P1_U3242) );
  INV_X1 U10763 ( .A(n9619), .ZN(n9622) );
  MUX2_X1 U10764 ( .A(n9622), .B(n9621), .S(n9620), .Z(n9625) );
  OAI211_X1 U10765 ( .C1(n9625), .C2(n9624), .A(P1_U4006), .B(n9623), .ZN(
        n9650) );
  OAI211_X1 U10766 ( .C1(n9628), .C2(n9627), .A(n9702), .B(n9626), .ZN(n9629)
         );
  OAI211_X1 U10767 ( .C1(n9641), .C2(n9630), .A(n9650), .B(n9629), .ZN(n9631)
         );
  AOI21_X1 U10768 ( .B1(n9711), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n9631), .ZN(
        n9636) );
  OAI211_X1 U10769 ( .C1(n9634), .C2(n9633), .A(n9712), .B(n9632), .ZN(n9635)
         );
  OAI211_X1 U10770 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6569), .A(n9636), .B(
        n9635), .ZN(P1_U3243) );
  AOI21_X1 U10771 ( .B1(n9639), .B2(n9638), .A(n9637), .ZN(n9642) );
  OAI22_X1 U10772 ( .A1(n9642), .A2(n9688), .B1(n9641), .B2(n9640), .ZN(n9643)
         );
  AOI21_X1 U10773 ( .B1(n9711), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9643), .ZN(
        n9652) );
  AOI21_X1 U10774 ( .B1(n9646), .B2(n9645), .A(n9644), .ZN(n9647) );
  OR2_X1 U10775 ( .A1(n9648), .A2(n9647), .ZN(n9649) );
  NAND4_X1 U10776 ( .A1(n9652), .A2(n9651), .A3(n9650), .A4(n9649), .ZN(
        P1_U3245) );
  AOI22_X1 U10777 ( .A1(n9711), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9653), .B2(
        n9704), .ZN(n9664) );
  AOI21_X1 U10778 ( .B1(n9656), .B2(n9655), .A(n9654), .ZN(n9657) );
  OR2_X1 U10779 ( .A1(n9688), .A2(n9657), .ZN(n9662) );
  OAI211_X1 U10780 ( .C1(n9660), .C2(n9659), .A(n9712), .B(n9658), .ZN(n9661)
         );
  NAND4_X1 U10781 ( .A1(n9664), .A2(n9663), .A3(n9662), .A4(n9661), .ZN(
        P1_U3246) );
  INV_X1 U10782 ( .A(n9680), .ZN(n9667) );
  INV_X1 U10783 ( .A(n9665), .ZN(n9675) );
  NAND3_X1 U10784 ( .A1(n9667), .A2(n9666), .A3(n9675), .ZN(n9668) );
  AND3_X1 U10785 ( .A1(n9669), .A2(n9712), .A3(n9668), .ZN(n9670) );
  AOI211_X1 U10786 ( .C1(n9711), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9671), .B(
        n9670), .ZN(n9684) );
  AOI21_X1 U10787 ( .B1(n9673), .B2(n9672), .A(n9704), .ZN(n9674) );
  OR2_X1 U10788 ( .A1(n9674), .A2(n9675), .ZN(n9683) );
  NAND3_X1 U10789 ( .A1(n9676), .A2(n7384), .A3(n9675), .ZN(n9677) );
  NAND3_X1 U10790 ( .A1(n9702), .A2(n9678), .A3(n9677), .ZN(n9682) );
  NAND3_X1 U10791 ( .A1(n9680), .A2(n9712), .A3(n9679), .ZN(n9681) );
  NAND4_X1 U10792 ( .A1(n9684), .A2(n9683), .A3(n9682), .A4(n9681), .ZN(
        P1_U3249) );
  OAI21_X1 U10793 ( .B1(n9687), .B2(n9686), .A(n9685), .ZN(n9694) );
  AOI211_X1 U10794 ( .C1(n9691), .C2(n9690), .A(n9689), .B(n9688), .ZN(n9692)
         );
  AOI211_X1 U10795 ( .C1(n9712), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9697)
         );
  AOI22_X1 U10796 ( .A1(n9711), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9695), .B2(
        n9704), .ZN(n9696) );
  NAND2_X1 U10797 ( .A1(n9697), .A2(n9696), .ZN(P1_U3251) );
  AOI21_X1 U10798 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9701) );
  NAND2_X1 U10799 ( .A1(n9702), .A2(n9701), .ZN(n9707) );
  NAND2_X1 U10800 ( .A1(n9704), .A2(n9703), .ZN(n9706) );
  AND3_X1 U10801 ( .A1(n9707), .A2(n9706), .A3(n9705), .ZN(n9715) );
  OAI21_X1 U10802 ( .B1(n9710), .B2(n9709), .A(n9708), .ZN(n9713) );
  AOI22_X1 U10803 ( .A1(n9713), .A2(n9712), .B1(n9711), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9714) );
  NAND2_X1 U10804 ( .A1(n9715), .A2(n9714), .ZN(P1_U3259) );
  OAI21_X1 U10805 ( .B1(n9718), .B2(n4837), .A(n9717), .ZN(n9734) );
  AOI22_X1 U10806 ( .A1(n6818), .A2(n9721), .B1(n9720), .B2(n9719), .ZN(n9722)
         );
  OAI21_X1 U10807 ( .B1(n9734), .B2(n9723), .A(n9722), .ZN(n9724) );
  AOI21_X1 U10808 ( .B1(n9726), .B2(n9725), .A(n9724), .ZN(n9753) );
  AOI22_X1 U10809 ( .A1(n9728), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9727), .B2(
        n9730), .ZN(n9739) );
  INV_X1 U10810 ( .A(n9729), .ZN(n9733) );
  AOI21_X1 U10811 ( .B1(n9731), .B2(n9730), .A(n9767), .ZN(n9732) );
  NAND2_X1 U10812 ( .A1(n9733), .A2(n9732), .ZN(n9751) );
  INV_X1 U10813 ( .A(n9734), .ZN(n9749) );
  NAND2_X1 U10814 ( .A1(n9749), .A2(n9735), .ZN(n9737) );
  MUX2_X1 U10815 ( .A(n9751), .B(n9737), .S(n9736), .Z(n9738) );
  AND3_X1 U10816 ( .A1(n9753), .A2(n9739), .A3(n9738), .ZN(n9741) );
  AOI22_X1 U10817 ( .A1(n9743), .A2(n9742), .B1(n9741), .B2(n9740), .ZN(
        P1_U3290) );
  AND2_X1 U10818 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9748), .ZN(P1_U3292) );
  AND2_X1 U10819 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9748), .ZN(P1_U3293) );
  AND2_X1 U10820 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9748), .ZN(P1_U3294) );
  AND2_X1 U10821 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9748), .ZN(P1_U3295) );
  AND2_X1 U10822 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9748), .ZN(P1_U3296) );
  AND2_X1 U10823 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9748), .ZN(P1_U3297) );
  AND2_X1 U10824 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9748), .ZN(P1_U3298) );
  AND2_X1 U10825 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9748), .ZN(P1_U3299) );
  AND2_X1 U10826 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9748), .ZN(P1_U3300) );
  AND2_X1 U10827 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9748), .ZN(P1_U3301) );
  AND2_X1 U10828 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9748), .ZN(P1_U3302) );
  AND2_X1 U10829 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9748), .ZN(P1_U3303) );
  NOR2_X1 U10830 ( .A1(n9747), .A2(n9744), .ZN(P1_U3304) );
  AND2_X1 U10831 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9748), .ZN(P1_U3305) );
  AND2_X1 U10832 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9748), .ZN(P1_U3306) );
  AND2_X1 U10833 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9748), .ZN(P1_U3307) );
  AND2_X1 U10834 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9748), .ZN(P1_U3308) );
  AND2_X1 U10835 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9748), .ZN(P1_U3309) );
  NOR2_X1 U10836 ( .A1(n9747), .A2(n9745), .ZN(P1_U3310) );
  AND2_X1 U10837 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9748), .ZN(P1_U3311) );
  AND2_X1 U10838 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9748), .ZN(P1_U3312) );
  AND2_X1 U10839 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9748), .ZN(P1_U3313) );
  AND2_X1 U10840 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9748), .ZN(P1_U3314) );
  AND2_X1 U10841 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9748), .ZN(P1_U3315) );
  NOR2_X1 U10842 ( .A1(n9747), .A2(n9746), .ZN(P1_U3316) );
  AND2_X1 U10843 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9748), .ZN(P1_U3317) );
  AND2_X1 U10844 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9748), .ZN(P1_U3318) );
  AND2_X1 U10845 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9748), .ZN(P1_U3319) );
  AND2_X1 U10846 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9748), .ZN(P1_U3320) );
  AND2_X1 U10847 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9748), .ZN(P1_U3321) );
  NAND2_X1 U10848 ( .A1(n9749), .A2(n9772), .ZN(n9750) );
  AND4_X1 U10849 ( .A1(n9753), .A2(n9752), .A3(n9751), .A4(n9750), .ZN(n9775)
         );
  INV_X1 U10850 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9754) );
  AOI22_X1 U10851 ( .A1(n9774), .A2(n9775), .B1(n9754), .B2(n9773), .ZN(
        P1_U3457) );
  OAI22_X1 U10852 ( .A1(n9756), .A2(n9767), .B1(n9755), .B2(n9765), .ZN(n9758)
         );
  AOI211_X1 U10853 ( .C1(n9772), .C2(n9759), .A(n9758), .B(n9757), .ZN(n9777)
         );
  AOI22_X1 U10854 ( .A1(n9774), .A2(n9777), .B1(n5961), .B2(n9773), .ZN(
        P1_U3460) );
  OAI22_X1 U10855 ( .A1(n9761), .A2(n9767), .B1(n9760), .B2(n9765), .ZN(n9763)
         );
  AOI211_X1 U10856 ( .C1(n9772), .C2(n9764), .A(n9763), .B(n9762), .ZN(n9778)
         );
  AOI22_X1 U10857 ( .A1(n9774), .A2(n9778), .B1(n5992), .B2(n9773), .ZN(
        P1_U3466) );
  OAI22_X1 U10858 ( .A1(n9768), .A2(n9767), .B1(n9766), .B2(n9765), .ZN(n9770)
         );
  AOI211_X1 U10859 ( .C1(n9772), .C2(n9771), .A(n9770), .B(n9769), .ZN(n9781)
         );
  AOI22_X1 U10860 ( .A1(n9774), .A2(n9781), .B1(n6027), .B2(n9773), .ZN(
        P1_U3472) );
  AOI22_X1 U10861 ( .A1(n9782), .A2(n9775), .B1(n6528), .B2(n9779), .ZN(
        P1_U3524) );
  AOI22_X1 U10862 ( .A1(n9782), .A2(n9777), .B1(n9776), .B2(n9779), .ZN(
        P1_U3525) );
  AOI22_X1 U10863 ( .A1(n9782), .A2(n9778), .B1(n5990), .B2(n9779), .ZN(
        P1_U3527) );
  AOI22_X1 U10864 ( .A1(n9782), .A2(n9781), .B1(n9780), .B2(n9779), .ZN(
        P1_U3529) );
  AOI22_X1 U10865 ( .A1(n9784), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9783), .ZN(n9793) );
  AOI22_X1 U10866 ( .A1(n9785), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9792) );
  OAI21_X1 U10867 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n9787), .A(n9786), .ZN(
        n9790) );
  NOR2_X1 U10868 ( .A1(n9788), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9789) );
  OAI21_X1 U10869 ( .B1(n9790), .B2(n9789), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9791) );
  OAI211_X1 U10870 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9793), .A(n9792), .B(
        n9791), .ZN(P2_U3245) );
  OAI21_X1 U10871 ( .B1(n9796), .B2(n9794), .A(n9795), .ZN(n9802) );
  OAI21_X1 U10872 ( .B1(n9798), .B2(n7556), .A(n9797), .ZN(n9807) );
  NOR2_X1 U10873 ( .A1(n9807), .A2(n9799), .ZN(n9800) );
  AOI211_X1 U10874 ( .C1(n9803), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9915)
         );
  AOI222_X1 U10875 ( .A1(n9806), .A2(n9805), .B1(P2_REG2_REG_8__SCAN_IN), .B2(
        n9831), .C1(n9821), .C2(n9804), .ZN(n9815) );
  INV_X1 U10876 ( .A(n9807), .ZN(n9918) );
  INV_X1 U10877 ( .A(n9808), .ZN(n9813) );
  OAI211_X1 U10878 ( .C1(n9810), .C2(n9914), .A(n9809), .B(n9905), .ZN(n9913)
         );
  INV_X1 U10879 ( .A(n9913), .ZN(n9811) );
  AOI22_X1 U10880 ( .A1(n9918), .A2(n9813), .B1(n9812), .B2(n9811), .ZN(n9814)
         );
  OAI211_X1 U10881 ( .C1(n9831), .C2(n9915), .A(n9815), .B(n9814), .ZN(
        P2_U3288) );
  INV_X1 U10882 ( .A(n9816), .ZN(n9827) );
  INV_X1 U10883 ( .A(n9817), .ZN(n9824) );
  AOI22_X1 U10884 ( .A1(n9821), .A2(n9820), .B1(n9819), .B2(n9818), .ZN(n9822)
         );
  OAI21_X1 U10885 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9826) );
  AOI211_X1 U10886 ( .C1(n9828), .C2(n9827), .A(n9826), .B(n9825), .ZN(n9830)
         );
  AOI22_X1 U10887 ( .A1(n9831), .A2(n6891), .B1(n9830), .B2(n9829), .ZN(
        P2_U3291) );
  INV_X1 U10888 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9834) );
  NOR2_X1 U10889 ( .A1(n9869), .A2(n9834), .ZN(P2_U3297) );
  INV_X1 U10890 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9835) );
  NOR2_X1 U10891 ( .A1(n9869), .A2(n9835), .ZN(P2_U3298) );
  INV_X1 U10892 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9836) );
  NOR2_X1 U10893 ( .A1(n9869), .A2(n9836), .ZN(P2_U3299) );
  INV_X1 U10894 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9837) );
  NOR2_X1 U10895 ( .A1(n9869), .A2(n9837), .ZN(P2_U3300) );
  INV_X1 U10896 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9838) );
  NOR2_X1 U10897 ( .A1(n9848), .A2(n9838), .ZN(P2_U3301) );
  INV_X1 U10898 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9839) );
  NOR2_X1 U10899 ( .A1(n9848), .A2(n9839), .ZN(P2_U3302) );
  NOR2_X1 U10900 ( .A1(n9848), .A2(n9840), .ZN(P2_U3303) );
  INV_X1 U10901 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9841) );
  NOR2_X1 U10902 ( .A1(n9848), .A2(n9841), .ZN(P2_U3304) );
  NOR2_X1 U10903 ( .A1(n9848), .A2(n9842), .ZN(P2_U3305) );
  INV_X1 U10904 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9843) );
  NOR2_X1 U10905 ( .A1(n9848), .A2(n9843), .ZN(P2_U3306) );
  INV_X1 U10906 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9844) );
  NOR2_X1 U10907 ( .A1(n9848), .A2(n9844), .ZN(P2_U3307) );
  INV_X1 U10908 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9845) );
  NOR2_X1 U10909 ( .A1(n9848), .A2(n9845), .ZN(P2_U3308) );
  INV_X1 U10910 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9846) );
  NOR2_X1 U10911 ( .A1(n9848), .A2(n9846), .ZN(P2_U3309) );
  INV_X1 U10912 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9847) );
  NOR2_X1 U10913 ( .A1(n9848), .A2(n9847), .ZN(P2_U3310) );
  INV_X1 U10914 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9849) );
  NOR2_X1 U10915 ( .A1(n9869), .A2(n9849), .ZN(P2_U3311) );
  INV_X1 U10916 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9850) );
  NOR2_X1 U10917 ( .A1(n9869), .A2(n9850), .ZN(P2_U3312) );
  INV_X1 U10918 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9851) );
  NOR2_X1 U10919 ( .A1(n9869), .A2(n9851), .ZN(P2_U3313) );
  INV_X1 U10920 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9852) );
  NOR2_X1 U10921 ( .A1(n9869), .A2(n9852), .ZN(P2_U3314) );
  INV_X1 U10922 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9853) );
  NOR2_X1 U10923 ( .A1(n9869), .A2(n9853), .ZN(P2_U3315) );
  INV_X1 U10924 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9854) );
  NOR2_X1 U10925 ( .A1(n9869), .A2(n9854), .ZN(P2_U3316) );
  INV_X1 U10926 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9855) );
  NOR2_X1 U10927 ( .A1(n9869), .A2(n9855), .ZN(P2_U3317) );
  INV_X1 U10928 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9856) );
  NOR2_X1 U10929 ( .A1(n9869), .A2(n9856), .ZN(P2_U3318) );
  INV_X1 U10930 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9857) );
  NOR2_X1 U10931 ( .A1(n9869), .A2(n9857), .ZN(P2_U3319) );
  INV_X1 U10932 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9858) );
  NOR2_X1 U10933 ( .A1(n9869), .A2(n9858), .ZN(P2_U3320) );
  INV_X1 U10934 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9859) );
  NOR2_X1 U10935 ( .A1(n9869), .A2(n9859), .ZN(P2_U3321) );
  INV_X1 U10936 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U10937 ( .A1(n9869), .A2(n9860), .ZN(P2_U3322) );
  NOR2_X1 U10938 ( .A1(n9869), .A2(n9861), .ZN(P2_U3323) );
  INV_X1 U10939 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9862) );
  NOR2_X1 U10940 ( .A1(n9869), .A2(n9862), .ZN(P2_U3324) );
  INV_X1 U10941 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9863) );
  NOR2_X1 U10942 ( .A1(n9869), .A2(n9863), .ZN(P2_U3325) );
  NOR2_X1 U10943 ( .A1(n9869), .A2(n9864), .ZN(P2_U3326) );
  OAI22_X1 U10944 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9869), .B1(n9868), .B2(
        n9865), .ZN(n9866) );
  INV_X1 U10945 ( .A(n9866), .ZN(P2_U3437) );
  OAI22_X1 U10946 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n9869), .B1(n9868), .B2(
        n9867), .ZN(n9870) );
  INV_X1 U10947 ( .A(n9870), .ZN(P2_U3438) );
  INV_X1 U10948 ( .A(n9871), .ZN(n9879) );
  OAI21_X1 U10949 ( .B1(n5561), .B2(n9873), .A(n9872), .ZN(n9876) );
  AOI21_X1 U10950 ( .B1(n9874), .B2(n5561), .A(n9947), .ZN(n9875) );
  AOI21_X1 U10951 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9878) );
  NOR2_X1 U10952 ( .A1(n9879), .A2(n9878), .ZN(n9953) );
  INV_X1 U10953 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9880) );
  AOI22_X1 U10954 ( .A1(n9951), .A2(n9953), .B1(n9880), .B2(n9949), .ZN(
        P2_U3451) );
  INV_X1 U10955 ( .A(n9881), .ZN(n9888) );
  NAND3_X1 U10956 ( .A1(n9883), .A2(n9905), .A3(n9882), .ZN(n9884) );
  OAI21_X1 U10957 ( .B1(n9885), .B2(n9941), .A(n9884), .ZN(n9887) );
  AOI211_X1 U10958 ( .C1(n9947), .C2(n9888), .A(n9887), .B(n9886), .ZN(n9954)
         );
  INV_X1 U10959 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U10960 ( .A1(n9951), .A2(n9954), .B1(n9889), .B2(n9949), .ZN(
        P2_U3454) );
  NAND3_X1 U10961 ( .A1(n9891), .A2(n9905), .A3(n9890), .ZN(n9892) );
  OAI211_X1 U10962 ( .C1(n4266), .C2(n9941), .A(n9893), .B(n9892), .ZN(n9894)
         );
  AOI21_X1 U10963 ( .B1(n9895), .B2(n9947), .A(n9894), .ZN(n9956) );
  INV_X1 U10964 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U10965 ( .A1(n9951), .A2(n9956), .B1(n9896), .B2(n9949), .ZN(
        P2_U3457) );
  NAND3_X1 U10966 ( .A1(n7751), .A2(n9897), .A3(n9947), .ZN(n9899) );
  OAI211_X1 U10967 ( .C1(n9900), .C2(n9941), .A(n9899), .B(n9898), .ZN(n9902)
         );
  NOR2_X1 U10968 ( .A1(n9902), .A2(n9901), .ZN(n9958) );
  INV_X1 U10969 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9903) );
  AOI22_X1 U10970 ( .A1(n9951), .A2(n9958), .B1(n9903), .B2(n9949), .ZN(
        P2_U3469) );
  AOI22_X1 U10971 ( .A1(n9906), .A2(n9905), .B1(n9929), .B2(n9904), .ZN(n9907)
         );
  OAI211_X1 U10972 ( .C1(n9910), .C2(n9909), .A(n9908), .B(n9907), .ZN(n9911)
         );
  INV_X1 U10973 ( .A(n9911), .ZN(n9960) );
  INV_X1 U10974 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9912) );
  AOI22_X1 U10975 ( .A1(n9951), .A2(n9960), .B1(n9912), .B2(n9949), .ZN(
        P2_U3472) );
  INV_X1 U10976 ( .A(n9931), .ZN(n9925) );
  OAI21_X1 U10977 ( .B1(n9914), .B2(n9941), .A(n9913), .ZN(n9917) );
  INV_X1 U10978 ( .A(n9915), .ZN(n9916) );
  AOI211_X1 U10979 ( .C1(n9925), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9961)
         );
  INV_X1 U10980 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U10981 ( .A1(n9951), .A2(n9961), .B1(n9919), .B2(n9949), .ZN(
        P2_U3475) );
  OAI22_X1 U10982 ( .A1(n9921), .A2(n9943), .B1(n9920), .B2(n9941), .ZN(n9923)
         );
  AOI211_X1 U10983 ( .C1(n9925), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9962)
         );
  INV_X1 U10984 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U10985 ( .A1(n9951), .A2(n9962), .B1(n9926), .B2(n9949), .ZN(
        P2_U3478) );
  AOI21_X1 U10986 ( .B1(n9929), .B2(n9928), .A(n9927), .ZN(n9930) );
  OAI21_X1 U10987 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(n9933) );
  NOR2_X1 U10988 ( .A1(n9934), .A2(n9933), .ZN(n9963) );
  INV_X1 U10989 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U10990 ( .A1(n9951), .A2(n9963), .B1(n9935), .B2(n9949), .ZN(
        P2_U3481) );
  OAI211_X1 U10991 ( .C1(n9938), .C2(n9941), .A(n9937), .B(n9936), .ZN(n9939)
         );
  AOI21_X1 U10992 ( .B1(n4359), .B2(n9947), .A(n9939), .ZN(n9964) );
  INV_X1 U10993 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U10994 ( .A1(n9951), .A2(n9964), .B1(n9940), .B2(n9949), .ZN(
        P2_U3484) );
  OAI22_X1 U10995 ( .A1(n9944), .A2(n9943), .B1(n9942), .B2(n9941), .ZN(n9946)
         );
  AOI211_X1 U10996 ( .C1(n9948), .C2(n9947), .A(n9946), .B(n9945), .ZN(n9966)
         );
  INV_X1 U10997 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U10998 ( .A1(n9951), .A2(n9966), .B1(n9950), .B2(n9949), .ZN(
        P2_U3487) );
  INV_X1 U10999 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9952) );
  AOI22_X1 U11000 ( .A1(n9967), .A2(n9953), .B1(n9952), .B2(n9965), .ZN(
        P2_U3520) );
  AOI22_X1 U11001 ( .A1(n9967), .A2(n9954), .B1(n4548), .B2(n9965), .ZN(
        P2_U3521) );
  AOI22_X1 U11002 ( .A1(n9967), .A2(n9956), .B1(n9955), .B2(n9965), .ZN(
        P2_U3522) );
  INV_X1 U11003 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9957) );
  AOI22_X1 U11004 ( .A1(n9967), .A2(n9958), .B1(n9957), .B2(n9965), .ZN(
        P2_U3526) );
  AOI22_X1 U11005 ( .A1(n9967), .A2(n9960), .B1(n9959), .B2(n9965), .ZN(
        P2_U3527) );
  AOI22_X1 U11006 ( .A1(n9967), .A2(n9961), .B1(n6916), .B2(n9965), .ZN(
        P2_U3528) );
  AOI22_X1 U11007 ( .A1(n9967), .A2(n9962), .B1(n7031), .B2(n9965), .ZN(
        P2_U3529) );
  AOI22_X1 U11008 ( .A1(n9967), .A2(n9963), .B1(n7123), .B2(n9965), .ZN(
        P2_U3530) );
  AOI22_X1 U11009 ( .A1(n9967), .A2(n9964), .B1(n7342), .B2(n9965), .ZN(
        P2_U3531) );
  AOI22_X1 U11010 ( .A1(n9967), .A2(n9966), .B1(n7474), .B2(n9965), .ZN(
        P2_U3532) );
  INV_X1 U11011 ( .A(n9968), .ZN(n9969) );
  NAND2_X1 U11012 ( .A1(n9970), .A2(n9969), .ZN(n9971) );
  XOR2_X1 U11013 ( .A(n9972), .B(n9971), .Z(ADD_1071_U5) );
  XOR2_X1 U11014 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11015 ( .B1(n9975), .B2(n9974), .A(n9973), .ZN(ADD_1071_U56) );
  OAI21_X1 U11016 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(ADD_1071_U57) );
  OAI21_X1 U11017 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(ADD_1071_U58) );
  OAI21_X1 U11018 ( .B1(n9984), .B2(n9983), .A(n9982), .ZN(ADD_1071_U59) );
  OAI21_X1 U11019 ( .B1(n9987), .B2(n9986), .A(n9985), .ZN(ADD_1071_U60) );
  OAI21_X1 U11020 ( .B1(n9990), .B2(n9989), .A(n9988), .ZN(ADD_1071_U61) );
  AOI21_X1 U11021 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(ADD_1071_U62) );
  AOI21_X1 U11022 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(ADD_1071_U63) );
  NOR2_X1 U11023 ( .A1(n9998), .A2(n9997), .ZN(n9999) );
  XOR2_X1 U11024 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9999), .Z(ADD_1071_U51) );
  XOR2_X1 U11025 ( .A(n10000), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  AOI21_X1 U11026 ( .B1(n10003), .B2(n10002), .A(n10001), .ZN(ADD_1071_U47) );
  OAI21_X1 U11027 ( .B1(n10006), .B2(n10005), .A(n10004), .ZN(n10007) );
  XNOR2_X1 U11028 ( .A(n10007), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11029 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10008), .Z(ADD_1071_U48) );
  XOR2_X1 U11030 ( .A(n10009), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11031 ( .A(n10011), .B(n10010), .Z(ADD_1071_U54) );
  XOR2_X1 U11032 ( .A(n10013), .B(n10012), .Z(ADD_1071_U53) );
  XNOR2_X1 U11033 ( .A(n10015), .B(n10014), .ZN(ADD_1071_U52) );
  INV_X1 U5859 ( .A(n5050), .ZN(n5087) );
  CLKBUF_X2 U4790 ( .A(n5935), .Z(n6406) );
  NAND2_X1 U4825 ( .A1(n8437), .A2(n5363), .ZN(n8311) );
  CLKBUF_X1 U6041 ( .A(n5113), .Z(n5489) );
endmodule

