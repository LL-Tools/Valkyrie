

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310;

  AND2_X1 U4817 ( .A1(n9354), .A2(n4991), .ZN(n8104) );
  NAND2_X1 U4818 ( .A1(n9575), .A2(n6625), .ZN(n9562) );
  NAND2_X1 U4819 ( .A1(n4848), .A2(n4846), .ZN(n9209) );
  NAND2_X1 U4820 ( .A1(n6611), .A2(n6610), .ZN(n9704) );
  NAND2_X1 U4821 ( .A1(n6521), .A2(n6520), .ZN(n9385) );
  NAND2_X1 U4822 ( .A1(n7569), .A2(n6057), .ZN(n7570) );
  AND2_X1 U4823 ( .A1(n9995), .A2(n6994), .ZN(n4975) );
  BUF_X2 U4824 ( .A(n7349), .Z(n7976) );
  INV_X1 U4826 ( .A(n6122), .ZN(n6100) );
  CLKBUF_X2 U4827 ( .A(n6394), .Z(n6551) );
  CLKBUF_X2 U4828 ( .A(n6363), .Z(n7271) );
  AND2_X1 U4829 ( .A1(n5994), .A2(n4980), .ZN(n5996) );
  NAND2_X2 U4830 ( .A1(n5993), .A2(n6840), .ZN(n6122) );
  INV_X2 U4831 ( .A(n5054), .ZN(n5582) );
  CLKBUF_X1 U4832 ( .A(n5982), .Z(n4319) );
  NAND2_X1 U4833 ( .A1(n9550), .A2(n8358), .ZN(n8369) );
  INV_X1 U4834 ( .A(n5015), .ZN(n4779) );
  OR2_X1 U4835 ( .A1(n6134), .A2(n6020), .ZN(n5970) );
  AND3_X1 U4836 ( .A1(n5992), .A2(n6003), .A3(n4825), .ZN(n6018) );
  NOR2_X1 U4837 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4825) );
  NAND2_X1 U4838 ( .A1(n8061), .A2(n8050), .ZN(n7349) );
  NOR2_X2 U4839 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6124) );
  NOR2_X1 U4840 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4933) );
  INV_X1 U4841 ( .A(n5585), .ZN(n5212) );
  INV_X1 U4842 ( .A(n8061), .ZN(n8048) );
  NAND3_X1 U4843 ( .A1(n9723), .A2(n9719), .A3(n4756), .ZN(n9678) );
  INV_X1 U4844 ( .A(n6017), .ZN(n6871) );
  NAND2_X1 U4845 ( .A1(n8325), .A2(n8114), .ZN(n8273) );
  AND2_X1 U4846 ( .A1(n6153), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6156) );
  CLKBUF_X2 U4849 ( .A(n5656), .Z(n6753) );
  OR2_X1 U4850 ( .A1(n8106), .A2(n6536), .ZN(n6542) );
  CLKBUF_X2 U4851 ( .A(n6382), .Z(n4316) );
  NAND2_X1 U4852 ( .A1(n9789), .A2(n9711), .ZN(n8310) );
  NAND2_X1 U4853 ( .A1(n4425), .A2(n10021), .ZN(n9970) );
  INV_X1 U4854 ( .A(n8277), .ZN(n8238) );
  NAND2_X1 U4855 ( .A1(n5996), .A2(n5995), .ZN(n7901) );
  AND2_X1 U4856 ( .A1(n6542), .A2(n6541), .ZN(n9360) );
  AND2_X1 U4857 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  INV_X1 U4858 ( .A(n6837), .ZN(n6840) );
  NAND2_X1 U4859 ( .A1(n6530), .A2(n6529), .ZN(n9384) );
  XNOR2_X1 U4860 ( .A(n5970), .B(n6133), .ZN(n5982) );
  OAI21_X1 U4861 ( .B1(n5093), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5051), .ZN(
        n5063) );
  NAND2_X2 U4864 ( .A1(n5195), .A2(n5194), .ZN(n5202) );
  OR2_X2 U4865 ( .A1(n6008), .A2(n6842), .ZN(n5994) );
  NOR2_X4 U4866 ( .A1(n9577), .A2(n9742), .ZN(n9576) );
  OAI21_X2 U4867 ( .B1(n8886), .B2(n8885), .A(n5879), .ZN(n8876) );
  NAND2_X2 U4868 ( .A1(n5345), .A2(n5869), .ZN(n8886) );
  NAND2_X1 U4869 ( .A1(n6593), .A2(n6592), .ZN(n7474) );
  INV_X1 U4870 ( .A(n4316), .ZN(n4311) );
  AOI21_X2 U4871 ( .B1(n9321), .B2(n9325), .A(n9202), .ZN(n9278) );
  BUF_X2 U4872 ( .A(n5993), .Z(n6017) );
  XNOR2_X1 U4873 ( .A(n5113), .B(n5123), .ZN(n6856) );
  OAI21_X2 U4874 ( .B1(n8141), .B2(n8246), .A(n6381), .ZN(n7297) );
  OR2_X1 U4875 ( .A1(n8375), .A2(n9550), .ZN(n8277) );
  OAI21_X1 U4876 ( .B1(n8103), .B2(n8104), .A(n9312), .ZN(n4444) );
  OAI21_X1 U4877 ( .B1(n7892), .B2(n8273), .A(n4920), .ZN(n9582) );
  CLKBUF_X1 U4878 ( .A(n8832), .Z(n8867) );
  CLKBUF_X1 U4879 ( .A(n8442), .Z(n4439) );
  CLKBUF_X1 U4880 ( .A(n9630), .Z(n9651) );
  NAND2_X1 U4881 ( .A1(n9705), .A2(n9706), .ZN(n6467) );
  CLKBUF_X1 U4882 ( .A(n7814), .Z(n4447) );
  NAND2_X1 U4883 ( .A1(n7475), .A2(n6403), .ZN(n7587) );
  NAND2_X1 U4884 ( .A1(n7488), .A2(n8142), .ZN(n7475) );
  OAI21_X2 U4885 ( .B1(n5397), .B2(n5396), .A(n5395), .ZN(n5435) );
  NAND2_X1 U4886 ( .A1(n6050), .A2(n6049), .ZN(n6597) );
  NAND2_X1 U4887 ( .A1(n5179), .A2(n5178), .ZN(n8502) );
  INV_X1 U4888 ( .A(n8602), .ZN(n8437) );
  INV_X1 U4889 ( .A(n8606), .ZN(n7370) );
  NAND2_X1 U4890 ( .A1(n6368), .A2(n6369), .ZN(n7055) );
  NAND4_X1 U4891 ( .A1(n5112), .A2(n5111), .A3(n5110), .A4(n5109), .ZN(n8606)
         );
  NAND2_X2 U4892 ( .A1(n6400), .A2(n8129), .ZN(n8142) );
  NAND2_X1 U4893 ( .A1(n5816), .A2(n5815), .ZN(n7112) );
  INV_X4 U4894 ( .A(n5108), .ZN(n5762) );
  XNOR2_X2 U4895 ( .A(n6573), .B(n7271), .ZN(n8249) );
  INV_X2 U4896 ( .A(n6380), .ZN(n7056) );
  INV_X4 U4897 ( .A(n4341), .ZN(n8058) );
  NAND2_X2 U4898 ( .A1(n6773), .A2(n6821), .ZN(n4341) );
  INV_X1 U4899 ( .A(n9001), .ZN(n6959) );
  NAND4_X1 U4900 ( .A1(n6338), .A2(n6337), .A3(n6336), .A4(n6335), .ZN(n9399)
         );
  INV_X1 U4901 ( .A(n6769), .ZN(n6773) );
  NAND2_X1 U4902 ( .A1(n8247), .A2(n8358), .ZN(n6769) );
  INV_X1 U4903 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5024) );
  NOR2_X1 U4904 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4999) );
  INV_X1 U4905 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6147) );
  AOI21_X1 U4906 ( .B1(n4927), .B2(n10064), .A(n4408), .ZN(n4926) );
  OR2_X1 U4907 ( .A1(n8367), .A2(n8366), .ZN(n4990) );
  NAND2_X1 U4908 ( .A1(n9239), .A2(n9240), .ZN(n9357) );
  NOR2_X1 U4909 ( .A1(n4928), .A2(n4758), .ZN(n4757) );
  AND2_X1 U4910 ( .A1(n4844), .A2(n4359), .ZN(n9219) );
  AOI211_X1 U4911 ( .C1(n9752), .C2(n9991), .A(n7896), .B(n7895), .ZN(n7897)
         );
  NOR2_X1 U4912 ( .A1(n8360), .A2(n8361), .ZN(n8367) );
  AND2_X1 U4913 ( .A1(n8776), .A2(n8775), .ZN(n9082) );
  NAND2_X1 U4914 ( .A1(n8083), .A2(n6308), .ZN(n6310) );
  NAND2_X1 U4915 ( .A1(n6572), .A2(n4368), .ZN(n4758) );
  AOI21_X1 U4916 ( .B1(n7882), .B2(n8317), .A(n4921), .ZN(n4920) );
  NOR2_X1 U4917 ( .A1(n6661), .A2(n4988), .ZN(n8721) );
  NAND2_X1 U4918 ( .A1(n9630), .A2(n6503), .ZN(n9607) );
  NAND2_X1 U4919 ( .A1(n6548), .A2(n6547), .ZN(n9383) );
  NAND2_X1 U4920 ( .A1(n4538), .A2(n8310), .ZN(n8342) );
  NAND3_X1 U4921 ( .A1(n4537), .A2(n4393), .A3(n4536), .ZN(n9630) );
  XNOR2_X1 U4922 ( .A(n5753), .B(n5752), .ZN(n9860) );
  OAI22_X1 U4923 ( .A1(n8514), .A2(n8515), .B1(n8938), .B2(n6233), .ZN(n8416)
         );
  NAND2_X1 U4924 ( .A1(n5570), .A2(n5569), .ZN(n5574) );
  CLKBUF_X1 U4925 ( .A(n7862), .Z(n4453) );
  NAND2_X1 U4926 ( .A1(n6118), .A2(n6117), .ZN(n9748) );
  NAND2_X1 U4927 ( .A1(n7831), .A2(n8178), .ZN(n6435) );
  CLKBUF_X1 U4928 ( .A(n7535), .Z(n4454) );
  AOI22_X1 U4929 ( .A1(n8646), .A2(P2_REG1_REG_11__SCAN_IN), .B1(n6692), .B2(
        n8648), .ZN(n7796) );
  XNOR2_X1 U4930 ( .A(n6691), .B(n8648), .ZN(n8646) );
  OR2_X1 U4931 ( .A1(n6487), .A2(n9327), .ZN(n6496) );
  NAND2_X1 U4932 ( .A1(n5442), .A2(n5441), .ZN(n9118) );
  NAND2_X1 U4933 ( .A1(n5423), .A2(n5422), .ZN(n9113) );
  NAND2_X1 U4934 ( .A1(n6108), .A2(n6107), .ZN(n9773) );
  NAND2_X1 U4935 ( .A1(n6404), .A2(n7587), .ZN(n7607) );
  NAND2_X1 U4936 ( .A1(n6595), .A2(n6594), .ZN(n7541) );
  AND2_X1 U4937 ( .A1(n8294), .A2(n8256), .ZN(n6404) );
  NAND2_X1 U4938 ( .A1(n6468), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U4939 ( .A1(n5401), .A2(n5400), .ZN(n9124) );
  NAND2_X1 U4940 ( .A1(n6104), .A2(n6103), .ZN(n9782) );
  INV_X1 U4941 ( .A(n6470), .ZN(n6468) );
  OR2_X1 U4942 ( .A1(n5612), .A2(n7713), .ZN(n5615) );
  NAND2_X1 U4943 ( .A1(n6102), .A2(n6101), .ZN(n9789) );
  NAND2_X1 U4944 ( .A1(n6082), .A2(n6081), .ZN(n9798) );
  NAND2_X1 U4945 ( .A1(n6074), .A2(n6073), .ZN(n9811) );
  NAND2_X1 U4946 ( .A1(n5299), .A2(n5298), .ZN(n9154) );
  NAND2_X2 U4947 ( .A1(n6078), .A2(n6077), .ZN(n9803) );
  NAND2_X1 U4948 ( .A1(n6293), .A2(n6292), .ZN(n8593) );
  OR2_X1 U4949 ( .A1(n8502), .A2(n8437), .ZN(n5841) );
  NAND2_X1 U4950 ( .A1(n5211), .A2(n5210), .ZN(n7690) );
  NAND2_X1 U4951 ( .A1(n6056), .A2(n6055), .ZN(n9826) );
  INV_X2 U4952 ( .A(n9073), .ZN(n4313) );
  NAND2_X1 U4953 ( .A1(n4751), .A2(n4752), .ZN(n5376) );
  NAND2_X1 U4954 ( .A1(n4596), .A2(n4363), .ZN(n4751) );
  AND2_X1 U4955 ( .A1(n7455), .A2(n5824), .ZN(n7385) );
  NAND2_X1 U4956 ( .A1(n4542), .A2(n6029), .ZN(n10039) );
  INV_X1 U4957 ( .A(n9967), .ZN(n10021) );
  NOR2_X2 U4958 ( .A1(n8743), .A2(n6750), .ZN(n6751) );
  XNOR2_X1 U4959 ( .A(n5172), .B(n5200), .ZN(n6869) );
  INV_X2 U4960 ( .A(n8383), .ZN(n6935) );
  OR2_X1 U4961 ( .A1(n5260), .A2(n4599), .ZN(n4596) );
  NAND2_X1 U4962 ( .A1(n7053), .A2(n7051), .ZN(n7052) );
  AOI21_X1 U4963 ( .B1(n5202), .B2(n4744), .A(n4745), .ZN(n5260) );
  XNOR2_X1 U4964 ( .A(n5166), .B(n5165), .ZN(n6863) );
  NAND2_X1 U4965 ( .A1(n6023), .A2(n6022), .ZN(n9967) );
  NAND2_X2 U4966 ( .A1(n6589), .A2(n8142), .ZN(n8253) );
  NAND2_X1 U4967 ( .A1(n6002), .A2(n7257), .ZN(n7300) );
  BUF_X1 U4968 ( .A(n6584), .Z(n8246) );
  NAND2_X1 U4969 ( .A1(n6196), .A2(n4669), .ZN(n4859) );
  INV_X1 U4970 ( .A(n10004), .ZN(n7302) );
  AND2_X1 U4971 ( .A1(n4608), .A2(n4603), .ZN(n4602) );
  OAI211_X2 U4973 ( .C1(n5759), .C2(n5059), .A(n5058), .B(n5057), .ZN(n8607)
         );
  OR2_X1 U4974 ( .A1(n8608), .A2(n6959), .ZN(n5816) );
  INV_X1 U4975 ( .A(n6400), .ZN(n8128) );
  NAND2_X1 U4976 ( .A1(n6398), .A2(n4968), .ZN(n6400) );
  OAI211_X1 U4977 ( .C1(n6856), .C2(n6008), .A(n6016), .B(n6015), .ZN(n10011)
         );
  NAND2_X1 U4978 ( .A1(n4888), .A2(n4886), .ZN(n7222) );
  NAND4_X2 U4979 ( .A1(n5042), .A2(n5041), .A3(n5040), .A4(n5039), .ZN(n8608)
         );
  NAND4_X1 U4980 ( .A1(n5035), .A2(n5034), .A3(n5033), .A4(n5032), .ZN(n8610)
         );
  AND3_X1 U4981 ( .A1(n5223), .A2(n5201), .A3(n5243), .ZN(n4744) );
  NAND2_X1 U4982 ( .A1(n5582), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5042) );
  AND4_X1 U4983 ( .A1(n6331), .A2(n6330), .A3(n6329), .A4(n6328), .ZN(n7790)
         );
  AND3_X2 U4984 ( .A1(n6001), .A2(n6000), .A3(n5999), .ZN(n7257) );
  AND4_X1 U4985 ( .A1(n6345), .A2(n6344), .A3(n6343), .A4(n6342), .ZN(n7753)
         );
  INV_X1 U4986 ( .A(n7320), .ZN(n6994) );
  CLKBUF_X1 U4987 ( .A(n5599), .Z(n7414) );
  NAND2_X1 U4988 ( .A1(n6382), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6575) );
  AND2_X1 U4989 ( .A1(n4747), .A2(n5243), .ZN(n4745) );
  NAND2_X1 U4990 ( .A1(n6354), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6414) );
  NAND2_X2 U4991 ( .A1(n4778), .A2(n4779), .ZN(n5236) );
  NAND2_X2 U4992 ( .A1(n6098), .A2(n6099), .ZN(n9550) );
  INV_X1 U4993 ( .A(n6356), .ZN(n6354) );
  NAND2_X1 U4994 ( .A1(n5598), .A2(n5597), .ZN(n5599) );
  XNOR2_X1 U4995 ( .A(n6127), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8247) );
  OR2_X1 U4996 ( .A1(n5596), .A2(n5589), .ZN(n5598) );
  AND2_X1 U4997 ( .A1(n4931), .A2(n8098), .ZN(n4315) );
  NAND2_X1 U4998 ( .A1(n4474), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6356) );
  INV_X1 U4999 ( .A(n6334), .ZN(n4474) );
  AND2_X1 U5000 ( .A1(n6139), .A2(n8098), .ZN(n6375) );
  NAND2_X1 U5001 ( .A1(n6131), .A2(n6130), .ZN(n8358) );
  AND2_X1 U5002 ( .A1(n5385), .A2(n5595), .ZN(n6697) );
  NAND2_X1 U5003 ( .A1(n6130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U5004 ( .A1(n5595), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U5005 ( .A1(n9175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5011) );
  OR2_X1 U5006 ( .A1(n5124), .A2(n5119), .ZN(n5126) );
  MUX2_X1 U5007 ( .A(n6129), .B(P1_IR_REG_31__SCAN_IN), .S(n6147), .Z(n6131)
         );
  NAND2_X1 U5008 ( .A1(n6136), .A2(n6138), .ZN(n8098) );
  NAND2_X1 U5009 ( .A1(n6128), .A2(n6147), .ZN(n6130) );
  XNOR2_X1 U5010 ( .A(n5020), .B(n5008), .ZN(n6754) );
  INV_X2 U5011 ( .A(n9859), .ZN(n9864) );
  OAI21_X1 U5012 ( .B1(n5670), .B2(n5590), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5591) );
  NAND2_X2 U5013 ( .A1(n6840), .A2(P1_U3086), .ZN(n9866) );
  NAND2_X1 U5014 ( .A1(n4532), .A2(n4530), .ZN(n6138) );
  NAND2_X1 U5015 ( .A1(n6136), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6135) );
  NOR2_X1 U5016 ( .A1(n6125), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4855) );
  AND2_X1 U5017 ( .A1(n5175), .A2(n5008), .ZN(n4430) );
  AND2_X2 U5018 ( .A1(n6667), .A2(n4912), .ZN(n5175) );
  NAND4_X1 U5019 ( .A1(n4999), .A2(n4998), .A3(n5132), .A4(n5075), .ZN(n5173)
         );
  NAND2_X1 U5020 ( .A1(n9869), .A2(n5024), .ZN(n4913) );
  NOR2_X1 U5021 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5964) );
  NOR2_X1 U5022 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6148) );
  NOR2_X2 U5023 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6667) );
  INV_X1 U5024 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5295) );
  NOR2_X1 U5025 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4821) );
  INV_X1 U5026 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6166) );
  INV_X1 U5027 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5132) );
  INV_X1 U5028 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5002) );
  AND2_X1 U5029 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9869) );
  INV_X4 U5030 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U5031 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5992) );
  INV_X1 U5032 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5075) );
  INV_X1 U5033 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6154) );
  OAI211_X1 U5034 ( .C1(n6636), .C2(n6641), .A(n5052), .B(n4348), .ZN(n9001)
         );
  AND2_X1 U5035 ( .A1(n4931), .A2(n8098), .ZN(n4314) );
  AND2_X1 U5036 ( .A1(n4931), .A2(n8098), .ZN(n6561) );
  AND2_X2 U5037 ( .A1(n7494), .A2(n8129), .ZN(n4425) );
  NAND3_X2 U5038 ( .A1(n6362), .A2(n6575), .A3(n6577), .ZN(n6573) );
  AND2_X1 U5039 ( .A1(n6578), .A2(n6576), .ZN(n6362) );
  NOR2_X4 U5040 ( .A1(n7570), .A2(n9820), .ZN(n7536) );
  NAND2_X2 U5041 ( .A1(n6374), .A2(n7130), .ZN(n8290) );
  INV_X2 U5042 ( .A(n7901), .ZN(n6374) );
  AND2_X2 U5043 ( .A1(n6139), .A2(n6321), .ZN(n6382) );
  AND3_X2 U5044 ( .A1(n4764), .A2(n4762), .A3(n6044), .ZN(n7569) );
  NAND2_X2 U5045 ( .A1(n6618), .A2(n6617), .ZN(n9606) );
  OR2_X2 U5046 ( .A1(n9622), .A2(n4401), .ZN(n6618) );
  NAND2_X2 U5047 ( .A1(n8290), .A2(n6581), .ZN(n7051) );
  AND2_X4 U5048 ( .A1(n9663), .A2(n9645), .ZN(n9641) );
  NOR2_X4 U5049 ( .A1(n4342), .A2(n9778), .ZN(n9663) );
  OR2_X2 U5050 ( .A1(n9678), .A2(n9782), .ZN(n4342) );
  OAI21_X2 U5051 ( .B1(n7541), .B2(n7544), .A(n7542), .ZN(n7648) );
  AND2_X1 U5052 ( .A1(n6139), .A2(n8098), .ZN(n4317) );
  INV_X4 U5053 ( .A(n6390), .ZN(n6498) );
  XNOR2_X2 U5054 ( .A(n6135), .B(n10193), .ZN(n6139) );
  INV_X4 U5055 ( .A(n4341), .ZN(n4318) );
  INV_X1 U5056 ( .A(n5600), .ZN(n4669) );
  OR2_X1 U5057 ( .A1(n9748), .A2(n9360), .ZN(n8325) );
  AND2_X1 U5058 ( .A1(n7806), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4807) );
  INV_X1 U5059 ( .A(n8653), .ZN(n4691) );
  NAND2_X1 U5060 ( .A1(n8937), .A2(n5622), .ZN(n4877) );
  NAND2_X1 U5061 ( .A1(n4586), .A2(n5550), .ZN(n5570) );
  NAND2_X1 U5062 ( .A1(n5549), .A2(n5548), .ZN(n4586) );
  OR2_X1 U5064 ( .A1(n5054), .A2(n5014), .ZN(n5018) );
  OR2_X1 U5065 ( .A1(n5236), .A2(n6964), .ZN(n5016) );
  NAND2_X1 U5066 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  NAND2_X1 U5067 ( .A1(n5643), .A2(n5642), .ZN(n8771) );
  INV_X1 U5068 ( .A(n4861), .ZN(n4860) );
  NOR2_X1 U5069 ( .A1(n6040), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6045) );
  OR2_X1 U5070 ( .A1(n4964), .A2(n4963), .ZN(n4961) );
  NAND2_X1 U5071 ( .A1(n4654), .A2(n4354), .ZN(n5860) );
  AND2_X1 U5072 ( .A1(n4643), .A2(n4635), .ZN(n4634) );
  AND2_X1 U5073 ( .A1(n4320), .A2(n4646), .ZN(n4635) );
  AND2_X1 U5074 ( .A1(n4643), .A2(n4320), .ZN(n4642) );
  NAND2_X1 U5075 ( .A1(n4629), .A2(n6495), .ZN(n4628) );
  INV_X1 U5076 ( .A(n8214), .ZN(n8212) );
  OR2_X1 U5077 ( .A1(n10039), .A2(n6353), .ZN(n8148) );
  NOR2_X1 U5078 ( .A1(n8784), .A2(n5639), .ZN(n4668) );
  NAND2_X1 U5079 ( .A1(n4742), .A2(n6634), .ZN(n4741) );
  NAND2_X1 U5080 ( .A1(n5687), .A2(n5685), .ZN(n6195) );
  NAND4_X1 U5081 ( .A1(n5001), .A2(n5000), .A3(n5295), .A4(n5317), .ZN(n5007)
         );
  INV_X1 U5082 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5000) );
  NOR2_X1 U5083 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5001) );
  NAND4_X1 U5084 ( .A1(n5005), .A2(n5004), .A3(n5003), .A4(n5002), .ZN(n5006)
         );
  INV_X1 U5085 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5005) );
  INV_X1 U5086 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5004) );
  INV_X1 U5087 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U5088 ( .A1(n8115), .A2(n8114), .ZN(n8345) );
  NAND2_X1 U5089 ( .A1(n4389), .A2(n5293), .ZN(n4754) );
  AOI21_X1 U5090 ( .B1(n5277), .B2(n4598), .A(n4382), .ZN(n4597) );
  INV_X1 U5091 ( .A(n5258), .ZN(n4598) );
  NAND2_X1 U5092 ( .A1(n5255), .A2(n5277), .ZN(n4599) );
  OAI21_X1 U5093 ( .B1(n6837), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n4452), .ZN(
        n5151) );
  NAND2_X1 U5094 ( .A1(n6837), .A2(n6866), .ZN(n4452) );
  NAND2_X1 U5095 ( .A1(n4562), .A2(n4563), .ZN(n6654) );
  AND2_X1 U5096 ( .A1(n4565), .A2(n4564), .ZN(n4563) );
  NAND2_X1 U5097 ( .A1(n4566), .A2(n6651), .ZN(n4564) );
  NAND2_X1 U5098 ( .A1(n4558), .A2(n4557), .ZN(n4556) );
  NAND2_X1 U5099 ( .A1(n8686), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4557) );
  OR2_X1 U5100 ( .A1(n5578), .A2(n6851), .ZN(n5029) );
  NOR2_X1 U5101 ( .A1(n6891), .A2(n5702), .ZN(n5725) );
  NAND2_X1 U5102 ( .A1(n5690), .A2(n5689), .ZN(n5722) );
  OR2_X1 U5103 ( .A1(n6891), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5690) );
  OR2_X1 U5104 ( .A1(n6300), .A2(n6315), .ZN(n5909) );
  OAI21_X1 U5105 ( .B1(n8897), .B2(n4862), .A(n5628), .ZN(n4861) );
  OAI211_X1 U5106 ( .C1(n4868), .C2(n4866), .A(n4865), .B(n5608), .ZN(n7386)
         );
  OR2_X1 U5107 ( .A1(n4867), .A2(n4866), .ZN(n4865) );
  NAND2_X1 U5108 ( .A1(n5607), .A2(n4355), .ZN(n4866) );
  OAI21_X1 U5109 ( .B1(n5280), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5316) );
  NOR2_X1 U5110 ( .A1(n7244), .A2(n4727), .ZN(n4726) );
  INV_X1 U5111 ( .A(n4729), .ZN(n4727) );
  INV_X1 U5112 ( .A(n8114), .ZN(n4921) );
  NOR2_X1 U5113 ( .A1(n9769), .A2(n9764), .ZN(n4761) );
  NAND2_X1 U5114 ( .A1(n4539), .A2(n4541), .ZN(n4536) );
  NAND2_X1 U5115 ( .A1(n6435), .A2(n4376), .ZN(n7814) );
  OR2_X1 U5116 ( .A1(n9826), .A2(n9336), .ZN(n8158) );
  OR2_X1 U5117 ( .A1(n6597), .A2(n7910), .ZN(n8157) );
  NAND2_X1 U5118 ( .A1(n5531), .A2(n5530), .ZN(n5549) );
  OR2_X1 U5119 ( .A1(n5369), .A2(n5371), .ZN(n5375) );
  NAND2_X1 U5120 ( .A1(n4596), .A2(n4597), .ZN(n5291) );
  NAND2_X1 U5121 ( .A1(n5195), .A2(n5190), .ZN(n5166) );
  OAI21_X1 U5122 ( .B1(n4446), .B2(n4386), .A(n5021), .ZN(n5656) );
  AOI21_X1 U5123 ( .B1(n5681), .B2(P2_IR_REG_31__SCAN_IN), .A(n4436), .ZN(
        n4446) );
  NAND2_X2 U5124 ( .A1(n6191), .A2(n5949), .ZN(n6634) );
  INV_X1 U5125 ( .A(n8803), .ZN(n8092) );
  NAND2_X1 U5126 ( .A1(n4324), .A2(n4375), .ZN(n4904) );
  INV_X1 U5127 ( .A(n8870), .ZN(n6255) );
  OAI21_X1 U5128 ( .B1(n8083), .B2(n8082), .A(n8081), .ZN(n8569) );
  AND2_X1 U5129 ( .A1(n8080), .A2(n8566), .ZN(n8081) );
  OR2_X1 U5130 ( .A1(n8390), .A2(n5581), .ZN(n5765) );
  INV_X1 U5131 ( .A(n5581), .ZN(n5562) );
  OR2_X1 U5132 ( .A1(n5762), .A2(n7202), .ZN(n5109) );
  NAND2_X1 U5133 ( .A1(n8384), .A2(n4779), .ZN(n5054) );
  INV_X1 U5134 ( .A(n8384), .ZN(n4778) );
  NAND2_X1 U5135 ( .A1(n6646), .A2(n6854), .ZN(n10085) );
  NAND2_X1 U5136 ( .A1(n4804), .A2(n6726), .ZN(n4808) );
  INV_X1 U5137 ( .A(n6652), .ZN(n4804) );
  NAND2_X1 U5138 ( .A1(n6652), .A2(n8648), .ZN(n4809) );
  AOI21_X1 U5139 ( .B1(n4689), .B2(n4694), .A(n4337), .ZN(n4688) );
  OR2_X1 U5140 ( .A1(n7466), .A2(n4690), .ZN(n4687) );
  NAND2_X1 U5141 ( .A1(n8683), .A2(n8682), .ZN(n8681) );
  AND2_X1 U5142 ( .A1(n10114), .A2(n4340), .ZN(n4769) );
  NAND2_X1 U5143 ( .A1(n8773), .A2(n5644), .ZN(n5954) );
  NAND2_X1 U5144 ( .A1(n5266), .A2(n4334), .ZN(n5320) );
  AOI21_X1 U5145 ( .B1(n5604), .B2(n7111), .A(n5603), .ZN(n5605) );
  OR2_X1 U5146 ( .A1(n6634), .A2(n5691), .ZN(n6986) );
  OR2_X1 U5147 ( .A1(n8771), .A2(n8770), .ZN(n8773) );
  AND2_X1 U5148 ( .A1(n4361), .A2(n5637), .ZN(n4870) );
  NAND2_X1 U5149 ( .A1(n5638), .A2(n5637), .ZN(n8793) );
  NOR2_X1 U5150 ( .A1(n8906), .A2(n8926), .ZN(n4876) );
  NAND2_X1 U5151 ( .A1(n4799), .A2(n5624), .ZN(n4798) );
  OR2_X1 U5152 ( .A1(n4321), .A2(n4800), .ZN(n4799) );
  XNOR2_X1 U5153 ( .A(n5154), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6720) );
  AND2_X1 U5154 ( .A1(n5116), .A2(n5131), .ZN(n6925) );
  INV_X1 U5155 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5043) );
  OAI21_X2 U5156 ( .B1(n6130), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6164) );
  NOR2_X1 U5157 ( .A1(n4448), .A2(n8276), .ZN(n8361) );
  NAND2_X1 U5158 ( .A1(n8239), .A2(n4449), .ZN(n4448) );
  AND2_X1 U5159 ( .A1(n8270), .A2(n4450), .ZN(n8274) );
  INV_X1 U5160 ( .A(n7290), .ZN(n8374) );
  NOR2_X1 U5161 ( .A1(n9468), .A2(n7020), .ZN(n7023) );
  AND2_X1 U5162 ( .A1(n9474), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7020) );
  NAND2_X1 U5163 ( .A1(n7249), .A2(n4500), .ZN(n4496) );
  OR2_X1 U5164 ( .A1(n9922), .A2(n4713), .ZN(n4711) );
  OR2_X1 U5165 ( .A1(n9498), .A2(n9940), .ZN(n4713) );
  OAI21_X1 U5166 ( .B1(n9606), .B2(n4955), .A(n4954), .ZN(n4953) );
  AOI21_X1 U5167 ( .B1(n4960), .B2(n8273), .A(n6624), .ZN(n4954) );
  NAND2_X1 U5168 ( .A1(n4957), .A2(n8273), .ZN(n4955) );
  NOR2_X1 U5169 ( .A1(n6621), .A2(n4965), .ZN(n4964) );
  INV_X1 U5170 ( .A(n4966), .ZN(n4965) );
  NAND2_X1 U5171 ( .A1(n6514), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6523) );
  INV_X1 U5172 ( .A(n6515), .ZN(n6514) );
  NAND2_X1 U5173 ( .A1(n4924), .A2(n4366), .ZN(n9598) );
  OR2_X1 U5174 ( .A1(n9764), .A2(n9386), .ZN(n4966) );
  OR2_X1 U5175 ( .A1(n9794), .A2(n9700), .ZN(n8200) );
  OR2_X1 U5176 ( .A1(n9815), .A2(n7818), .ZN(n8184) );
  NAND2_X1 U5177 ( .A1(n4935), .A2(n4937), .ZN(n4934) );
  INV_X1 U5178 ( .A(n4937), .ZN(n4936) );
  INV_X1 U5179 ( .A(n9962), .ZN(n9708) );
  NAND2_X1 U5180 ( .A1(n6062), .A2(n6061), .ZN(n9820) );
  OR2_X1 U5181 ( .A1(n8363), .A2(n7321), .ZN(n10020) );
  AND2_X1 U5182 ( .A1(n5474), .A2(n5462), .ZN(n5472) );
  AND2_X1 U5183 ( .A1(n5353), .A2(n5370), .ZN(n5355) );
  NOR2_X1 U5184 ( .A1(n7224), .A2(n4993), .ZN(n7232) );
  OR2_X2 U5185 ( .A1(n6758), .A2(P2_U3151), .ZN(n8743) );
  NAND2_X1 U5186 ( .A1(n8633), .A2(n8632), .ZN(n8631) );
  AOI21_X1 U5187 ( .B1(n8737), .B2(n8736), .A(n8735), .ZN(n8739) );
  OR2_X1 U5188 ( .A1(n7407), .A2(n6192), .ZN(n8817) );
  AND2_X1 U5189 ( .A1(n6048), .A2(n6052), .ZN(n7517) );
  NAND2_X1 U5190 ( .A1(n6132), .A2(n10012), .ZN(n9555) );
  NAND2_X1 U5191 ( .A1(n4323), .A2(n4659), .ZN(n4658) );
  OR2_X1 U5192 ( .A1(n5847), .A2(n5848), .ZN(n4656) );
  NAND2_X1 U5193 ( .A1(n4620), .A2(n4352), .ZN(n4619) );
  INV_X1 U5194 ( .A(n8943), .ZN(n4649) );
  INV_X1 U5195 ( .A(n5894), .ZN(n4645) );
  NAND2_X1 U5196 ( .A1(n4644), .A2(n5895), .ZN(n4636) );
  NAND2_X1 U5197 ( .A1(n5902), .A2(n4380), .ZN(n4643) );
  AND2_X1 U5198 ( .A1(n8203), .A2(n4440), .ZN(n8197) );
  INV_X1 U5199 ( .A(n8307), .ZN(n4440) );
  INV_X1 U5200 ( .A(n8784), .ZN(n4667) );
  NAND2_X1 U5201 ( .A1(n6657), .A2(n8707), .ZN(n4560) );
  NAND2_X1 U5202 ( .A1(n8330), .A2(n8329), .ZN(n8352) );
  AOI21_X1 U5203 ( .B1(n4627), .B2(n4358), .A(n4625), .ZN(n8224) );
  NAND2_X1 U5204 ( .A1(n8272), .A2(n4626), .ZN(n4625) );
  NOR2_X1 U5205 ( .A1(n8227), .A2(n8345), .ZN(n4469) );
  INV_X1 U5206 ( .A(n5241), .ZN(n4748) );
  NAND2_X1 U5207 ( .A1(n4592), .A2(SI_7_), .ZN(n5190) );
  NAND3_X1 U5208 ( .A1(n6195), .A2(n6194), .A3(n6193), .ZN(n6205) );
  INV_X1 U5209 ( .A(n8499), .ZN(n4911) );
  NAND2_X1 U5210 ( .A1(n4665), .A2(n4971), .ZN(n5930) );
  NAND2_X1 U5211 ( .A1(n8616), .A2(n6642), .ZN(n4792) );
  NAND2_X1 U5212 ( .A1(n8613), .A2(n6673), .ZN(n6674) );
  NOR2_X1 U5213 ( .A1(n6715), .A2(n7372), .ZN(n6647) );
  AND2_X1 U5214 ( .A1(n5336), .A2(n4678), .ZN(n4677) );
  INV_X1 U5215 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4678) );
  INV_X1 U5216 ( .A(n5338), .ZN(n5337) );
  NAND2_X1 U5217 ( .A1(n5615), .A2(n4442), .ZN(n5616) );
  NAND2_X1 U5218 ( .A1(n8462), .A2(n7711), .ZN(n4442) );
  AND2_X1 U5219 ( .A1(n4351), .A2(n4684), .ZN(n4683) );
  INV_X1 U5220 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n4684) );
  AND2_X1 U5221 ( .A1(n5189), .A2(n5825), .ZN(n4818) );
  INV_X1 U5222 ( .A(n5833), .ZN(n4781) );
  NAND2_X1 U5223 ( .A1(n5821), .A2(n5832), .ZN(n5604) );
  OR2_X1 U5224 ( .A1(n5723), .A2(n5722), .ZN(n6981) );
  INV_X1 U5225 ( .A(n8861), .ZN(n6258) );
  OR2_X1 U5226 ( .A1(n9124), .A2(n8455), .ZN(n5633) );
  OR2_X1 U5227 ( .A1(n9136), .A2(n8446), .ZN(n5879) );
  NAND2_X1 U5228 ( .A1(n9142), .A2(n8913), .ZN(n5869) );
  OR2_X1 U5229 ( .A1(n9142), .A2(n8913), .ZN(n5877) );
  OR2_X1 U5230 ( .A1(n7458), .A2(n5610), .ZN(n7580) );
  INV_X1 U5231 ( .A(n7677), .ZN(n5222) );
  AND2_X1 U5232 ( .A1(n4812), .A2(n4811), .ZN(n4810) );
  NOR2_X1 U5233 ( .A1(n5006), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4812) );
  NOR2_X1 U5234 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n4972) );
  NOR2_X1 U5235 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4977) );
  INV_X1 U5236 ( .A(n5682), .ZN(n4813) );
  INV_X1 U5237 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5673) );
  INV_X1 U5238 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5317) );
  OR2_X1 U5239 ( .A1(n5245), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5261) );
  OR2_X1 U5240 ( .A1(n5114), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U5241 ( .A1(n4842), .A2(n4841), .ZN(n4840) );
  INV_X1 U5242 ( .A(n8025), .ZN(n4841) );
  AOI21_X1 U5243 ( .B1(n4839), .B2(n4842), .A(n4388), .ZN(n4838) );
  NOR2_X1 U5244 ( .A1(n4346), .A2(n8025), .ZN(n4839) );
  NOR2_X1 U5245 ( .A1(n6784), .A2(n4981), .ZN(n6789) );
  OR2_X1 U5246 ( .A1(n4843), .A2(n8009), .ZN(n4842) );
  AND2_X1 U5247 ( .A1(n9220), .A2(n4359), .ZN(n4843) );
  NAND2_X1 U5248 ( .A1(n4853), .A2(n4852), .ZN(n7336) );
  AND2_X1 U5249 ( .A1(n6817), .A2(n6812), .ZN(n4852) );
  NAND2_X1 U5250 ( .A1(n8331), .A2(n8332), .ZN(n4590) );
  INV_X1 U5251 ( .A(n8352), .ZN(n4591) );
  NOR2_X1 U5252 ( .A1(n8241), .A2(n8240), .ZN(n8333) );
  NAND2_X1 U5253 ( .A1(n9448), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4721) );
  INV_X1 U5254 ( .A(n6620), .ZN(n4963) );
  AND2_X1 U5255 ( .A1(n8285), .A2(n4540), .ZN(n4539) );
  OR2_X1 U5256 ( .A1(n4326), .A2(n4541), .ZN(n4540) );
  INV_X1 U5257 ( .A(n8310), .ZN(n4541) );
  OR2_X1 U5258 ( .A1(n9778), .A2(n9648), .ZN(n8243) );
  NAND2_X1 U5259 ( .A1(n4514), .A2(n4512), .ZN(n6352) );
  INV_X1 U5260 ( .A(n8152), .ZN(n4514) );
  NOR2_X1 U5261 ( .A1(n6351), .A2(n6350), .ZN(n4512) );
  NAND2_X1 U5262 ( .A1(n6325), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6334) );
  OAI21_X1 U5263 ( .B1(n8398), .B2(n6008), .A(n5975), .ZN(n6569) );
  INV_X1 U5264 ( .A(n8265), .ZN(n6451) );
  NOR2_X1 U5265 ( .A1(n6860), .A2(n7289), .ZN(n6813) );
  AND2_X1 U5266 ( .A1(n5573), .A2(n5555), .ZN(n5569) );
  INV_X1 U5267 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5968) );
  AND2_X1 U5268 ( .A1(n5550), .A2(n5536), .ZN(n5548) );
  NAND2_X1 U5269 ( .A1(n4584), .A2(n5514), .ZN(n5529) );
  AND2_X1 U5270 ( .A1(n5530), .A2(n5518), .ZN(n5528) );
  AND2_X1 U5271 ( .A1(n4933), .A2(n4821), .ZN(n4820) );
  AND2_X1 U5272 ( .A1(n5495), .A2(n5479), .ZN(n5493) );
  INV_X1 U5273 ( .A(n5456), .ZN(n4615) );
  INV_X1 U5274 ( .A(n4754), .ZN(n4595) );
  AOI21_X1 U5275 ( .B1(n5200), .B2(n5199), .A(n5198), .ZN(n5201) );
  INV_X1 U5276 ( .A(n5193), .ZN(n5200) );
  NAND2_X1 U5277 ( .A1(n5126), .A2(n5125), .ZN(n5127) );
  XNOR2_X1 U5278 ( .A(n4592), .B(SI_7_), .ZN(n5148) );
  NAND2_X1 U5279 ( .A1(n5093), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U5280 ( .A1(n8558), .A2(n4369), .ZN(n7695) );
  XNOR2_X1 U5281 ( .A(n6196), .B(n6205), .ZN(n6197) );
  NOR2_X1 U5282 ( .A1(n6197), .A2(n8609), .ZN(n6199) );
  AND2_X1 U5283 ( .A1(n4324), .A2(n8443), .ZN(n4905) );
  INV_X1 U5284 ( .A(n8582), .ZN(n6237) );
  NAND2_X1 U5285 ( .A1(n5705), .A2(n5704), .ZN(n6749) );
  NAND2_X1 U5286 ( .A1(n5384), .A2(n5383), .ZN(n5595) );
  INV_X1 U5287 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5383) );
  INV_X1 U5288 ( .A(n5670), .ZN(n5384) );
  INV_X1 U5289 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5589) );
  AND4_X1 U5290 ( .A1(n5220), .A2(n5219), .A3(n5218), .A4(n5217), .ZN(n8537)
         );
  OR2_X1 U5291 ( .A1(n5585), .A2(n6701), .ZN(n5034) );
  XNOR2_X1 U5292 ( .A(n6700), .B(n6976), .ZN(n6970) );
  OAI21_X1 U5293 ( .B1(n6838), .B2(n6638), .A(n6639), .ZN(n6965) );
  OAI21_X1 U5294 ( .B1(n6753), .B2(n6964), .A(n4702), .ZN(n6700) );
  NAND2_X1 U5295 ( .A1(n6753), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4702) );
  NAND2_X1 U5296 ( .A1(n6969), .A2(n6970), .ZN(n6968) );
  XNOR2_X1 U5297 ( .A(n6641), .B(n6640), .ZN(n8618) );
  NAND2_X1 U5298 ( .A1(n4897), .A2(n4896), .ZN(n8615) );
  NAND2_X1 U5299 ( .A1(n6641), .A2(n6665), .ZN(n4896) );
  OR2_X1 U5300 ( .A1(n6641), .A2(n6665), .ZN(n4897) );
  AOI21_X1 U5301 ( .B1(n6922), .B2(n10085), .A(n10086), .ZN(n10088) );
  NAND2_X1 U5302 ( .A1(n10082), .A2(n6683), .ZN(n6684) );
  NAND2_X1 U5303 ( .A1(n4696), .A2(n4700), .ZN(n4695) );
  INV_X1 U5304 ( .A(n4698), .ZN(n4696) );
  AOI21_X1 U5305 ( .B1(n7467), .B2(n4407), .A(n4699), .ZN(n4698) );
  INV_X1 U5306 ( .A(n7441), .ZN(n4699) );
  AND2_X1 U5307 ( .A1(n4807), .A2(n8648), .ZN(n4805) );
  AND2_X1 U5308 ( .A1(n7806), .A2(n8648), .ZN(n4806) );
  NAND2_X1 U5309 ( .A1(n4568), .A2(n4567), .ZN(n6652) );
  AND2_X1 U5310 ( .A1(n4687), .A2(n4418), .ZN(n7799) );
  INV_X1 U5311 ( .A(n7801), .ZN(n4686) );
  AOI21_X1 U5312 ( .B1(n7463), .B2(n4576), .A(n4573), .ZN(n6691) );
  AND2_X1 U5313 ( .A1(n7440), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4576) );
  NAND2_X1 U5314 ( .A1(n6654), .A2(n8665), .ZN(n8677) );
  NOR2_X1 U5315 ( .A1(n4556), .A2(n4894), .ZN(n6656) );
  NAND2_X1 U5316 ( .A1(n8681), .A2(n4412), .ZN(n8697) );
  NAND2_X1 U5317 ( .A1(n4580), .A2(n4577), .ZN(n6694) );
  AND2_X1 U5318 ( .A1(n4890), .A2(n4895), .ZN(n4577) );
  OR2_X1 U5319 ( .A1(n6732), .A2(n10262), .ZN(n4895) );
  XNOR2_X1 U5320 ( .A(n6694), .B(n7033), .ZN(n4579) );
  XNOR2_X1 U5321 ( .A(n8774), .B(n8410), .ZN(n5953) );
  INV_X1 U5322 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n4679) );
  NAND2_X1 U5323 ( .A1(n5483), .A2(n5482), .ZN(n5504) );
  AND2_X1 U5324 ( .A1(n5599), .A2(n6697), .ZN(n6192) );
  OR2_X1 U5325 ( .A1(n5465), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5484) );
  OR2_X1 U5326 ( .A1(n5445), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U5327 ( .A1(n5425), .A2(n5424), .ZN(n5445) );
  INV_X1 U5328 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5424) );
  INV_X1 U5329 ( .A(n5443), .ZN(n5425) );
  OR2_X1 U5330 ( .A1(n5402), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5443) );
  AND2_X1 U5331 ( .A1(n4869), .A2(n4397), .ZN(n4867) );
  OR2_X1 U5332 ( .A1(n7312), .A2(n7235), .ZN(n4869) );
  INV_X1 U5333 ( .A(n5604), .ZN(n7113) );
  INV_X1 U5334 ( .A(n7112), .ZN(n4445) );
  NAND2_X1 U5335 ( .A1(n6191), .A2(n5599), .ZN(n7036) );
  NAND2_X1 U5336 ( .A1(n5602), .A2(n5601), .ZN(n6955) );
  OR2_X1 U5337 ( .A1(n8610), .A2(n7216), .ZN(n7038) );
  NOR2_X1 U5338 ( .A1(n8753), .A2(n8752), .ZN(n9076) );
  NAND2_X1 U5339 ( .A1(n5501), .A2(n5500), .ZN(n6300) );
  NAND2_X1 U5340 ( .A1(n8839), .A2(n4372), .ZN(n4815) );
  AND2_X1 U5341 ( .A1(n8839), .A2(n8810), .ZN(n8823) );
  OR2_X1 U5342 ( .A1(n9118), .A2(n6255), .ZN(n8835) );
  NAND2_X1 U5343 ( .A1(n8898), .A2(n8897), .ZN(n8896) );
  NAND2_X1 U5344 ( .A1(n5877), .A2(n5869), .ZN(n8897) );
  INV_X1 U5345 ( .A(n8939), .ZN(n8912) );
  OR2_X1 U5346 ( .A1(n6634), .A2(n6276), .ZN(n8969) );
  NOR2_X1 U5347 ( .A1(n5305), .A2(n4803), .ZN(n4802) );
  INV_X1 U5348 ( .A(n5274), .ZN(n4803) );
  NAND2_X1 U5349 ( .A1(n8959), .A2(n5273), .ZN(n5275) );
  AND2_X1 U5350 ( .A1(n5866), .A2(n5875), .ZN(n8926) );
  NAND2_X1 U5351 ( .A1(n5248), .A2(n5247), .ZN(n9058) );
  INV_X1 U5352 ( .A(n8969), .ZN(n8954) );
  XNOR2_X1 U5353 ( .A(n5706), .B(n5707), .ZN(n6748) );
  NOR2_X1 U5354 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4912) );
  NAND2_X1 U5355 ( .A1(n4554), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4553) );
  NAND2_X1 U5356 ( .A1(n4431), .A2(n5043), .ZN(n4554) );
  INV_X1 U5357 ( .A(n9233), .ZN(n4830) );
  NAND2_X1 U5358 ( .A1(n7255), .A2(n7256), .ZN(n4853) );
  CLKBUF_X1 U5359 ( .A(n7336), .Z(n7396) );
  INV_X1 U5360 ( .A(n7919), .ZN(n4831) );
  AOI21_X1 U5361 ( .B1(n4849), .B2(n4851), .A(n4847), .ZN(n4846) );
  INV_X1 U5362 ( .A(n9263), .ZN(n4847) );
  NAND2_X1 U5363 ( .A1(n8375), .A2(n8247), .ZN(n8354) );
  NOR2_X1 U5364 ( .A1(n7015), .A2(n7016), .ZN(n7017) );
  INV_X1 U5365 ( .A(n7017), .ZN(n4720) );
  AOI21_X1 U5366 ( .B1(n9431), .B2(n4720), .A(n9442), .ZN(n4719) );
  NOR2_X1 U5367 ( .A1(n9432), .A2(n9431), .ZN(n9430) );
  OR2_X1 U5368 ( .A1(n7242), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4729) );
  OR2_X1 U5369 ( .A1(n6047), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U5370 ( .A1(n4728), .A2(n7416), .ZN(n4723) );
  NAND2_X1 U5371 ( .A1(n7241), .A2(n4726), .ZN(n4724) );
  INV_X1 U5372 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10247) );
  OR2_X1 U5373 ( .A1(n9935), .A2(n9506), .ZN(n4485) );
  NAND2_X1 U5374 ( .A1(n4485), .A2(n4484), .ZN(n9524) );
  INV_X1 U5375 ( .A(n9509), .ZN(n4484) );
  NOR2_X1 U5376 ( .A1(n4710), .A2(n9932), .ZN(n4709) );
  INV_X1 U5377 ( .A(n4712), .ZN(n4710) );
  AOI21_X1 U5378 ( .B1(n4506), .B2(n4508), .A(n4428), .ZN(n4505) );
  AOI21_X1 U5379 ( .B1(n4734), .B2(n4732), .A(n4731), .ZN(n4730) );
  INV_X1 U5380 ( .A(n4734), .ZN(n4733) );
  NAND2_X1 U5381 ( .A1(n4919), .A2(n4917), .ZN(n9581) );
  AOI21_X1 U5382 ( .B1(n4920), .B2(n8273), .A(n4918), .ZN(n4917) );
  NAND2_X1 U5383 ( .A1(n7881), .A2(n7882), .ZN(n7880) );
  NAND2_X1 U5384 ( .A1(n7892), .A2(n8219), .ZN(n7881) );
  AND2_X1 U5385 ( .A1(n4327), .A2(n9367), .ZN(n4759) );
  NAND2_X1 U5386 ( .A1(n4479), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6515) );
  OAI21_X1 U5387 ( .B1(n6467), .B2(n4541), .A(n4539), .ZN(n4923) );
  INV_X1 U5388 ( .A(n4948), .ZN(n4947) );
  OAI22_X1 U5389 ( .A1(n6614), .A2(n4949), .B1(n9221), .B2(n9782), .ZN(n4948)
         );
  NAND2_X1 U5390 ( .A1(n4349), .A2(n6613), .ZN(n4949) );
  INV_X1 U5391 ( .A(n6613), .ZN(n4952) );
  NAND2_X1 U5392 ( .A1(n4520), .A2(n4521), .ZN(n9705) );
  AOI21_X1 U5393 ( .B1(n4524), .B2(n8180), .A(n4522), .ZN(n4521) );
  INV_X1 U5394 ( .A(n8199), .ZN(n4522) );
  AND2_X1 U5395 ( .A1(n8200), .A2(n8201), .ZN(n9706) );
  AND2_X1 U5396 ( .A1(n8265), .A2(n8181), .ZN(n4922) );
  AND2_X1 U5397 ( .A1(n8189), .A2(n8304), .ZN(n8265) );
  INV_X1 U5398 ( .A(n7832), .ZN(n8264) );
  NAND2_X1 U5399 ( .A1(n4454), .A2(n8261), .ZN(n7534) );
  NAND2_X1 U5400 ( .A1(n7530), .A2(n6426), .ZN(n7831) );
  NAND2_X1 U5401 ( .A1(n6353), .A2(n10039), .ZN(n8151) );
  NOR2_X1 U5402 ( .A1(n9970), .A2(n10029), .ZN(n7552) );
  OR2_X1 U5403 ( .A1(n8354), .A2(n7025), .ZN(n9712) );
  NAND2_X1 U5404 ( .A1(n6580), .A2(n6579), .ZN(n7053) );
  NAND2_X1 U5405 ( .A1(n9995), .A2(n4353), .ZN(n6579) );
  INV_X1 U5406 ( .A(n9712), .ZN(n9675) );
  OR2_X1 U5407 ( .A1(n7321), .A2(n8365), .ZN(n9724) );
  OR2_X1 U5408 ( .A1(n8363), .A2(n8354), .ZN(n7292) );
  AOI21_X1 U5409 ( .B1(n6185), .B2(n6184), .A(n6862), .ZN(n7295) );
  NOR2_X1 U5410 ( .A1(n6627), .A2(n10051), .ZN(n6628) );
  NAND2_X1 U5411 ( .A1(n4464), .A2(n4463), .ZN(n4462) );
  NAND2_X1 U5412 ( .A1(n6559), .A2(n8336), .ZN(n9962) );
  OAI21_X1 U5413 ( .B1(n5742), .B2(n5741), .A(n5740), .ZN(n5750) );
  XNOR2_X1 U5414 ( .A(n5750), .B(n5749), .ZN(n8379) );
  INV_X1 U5415 ( .A(n5574), .ZN(n5572) );
  NAND2_X1 U5416 ( .A1(n5574), .A2(n5573), .ZN(n5742) );
  INV_X1 U5417 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6133) );
  XNOR2_X1 U5418 ( .A(n5570), .B(n5569), .ZN(n8388) );
  OR2_X1 U5419 ( .A1(n6151), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U5420 ( .A1(n6071), .A2(n5967), .ZN(n6151) );
  OAI21_X1 U5421 ( .B1(n5260), .B2(n5259), .A(n5258), .ZN(n5278) );
  NAND2_X1 U5422 ( .A1(n5070), .A2(SI_3_), .ZN(n5071) );
  NAND2_X1 U5423 ( .A1(n4916), .A2(n5065), .ZN(n5068) );
  NAND2_X1 U5424 ( .A1(n4503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6005) );
  INV_X1 U5425 ( .A(n5992), .ZN(n4503) );
  NAND2_X1 U5426 ( .A1(n8089), .A2(n8088), .ZN(n8413) );
  AND4_X1 U5427 ( .A1(n5146), .A2(n5145), .A3(n5144), .A4(n5143), .ZN(n7700)
         );
  NAND2_X1 U5428 ( .A1(n6270), .A2(n6269), .ZN(n4435) );
  AOI21_X1 U5429 ( .B1(n8882), .B2(n5562), .A(n5393), .ZN(n8510) );
  AOI21_X1 U5430 ( .B1(n4901), .B2(n4903), .A(n4387), .ZN(n4899) );
  AND2_X1 U5431 ( .A1(n6278), .A2(n6277), .ZN(n8587) );
  INV_X1 U5432 ( .A(n8786), .ZN(n8576) );
  NAND2_X1 U5433 ( .A1(n6304), .A2(n8989), .ZN(n8578) );
  NAND2_X1 U5434 ( .A1(n5527), .A2(n5526), .ZN(n8803) );
  NAND2_X1 U5435 ( .A1(n5367), .A2(n5366), .ZN(n8899) );
  OAI211_X1 U5436 ( .C1(n5762), .C2(n8944), .A(n5288), .B(n5287), .ZN(n8953)
         );
  AND2_X1 U5437 ( .A1(n5056), .A2(n5055), .ZN(n5058) );
  NAND2_X1 U5438 ( .A1(n8631), .A2(n4706), .ZN(n6921) );
  OR2_X1 U5439 ( .A1(n6710), .A2(n8630), .ZN(n4706) );
  NAND2_X1 U5440 ( .A1(n6921), .A2(n6920), .ZN(n6919) );
  NAND2_X1 U5441 ( .A1(n4816), .A2(n10085), .ZN(n4552) );
  XNOR2_X1 U5442 ( .A(n6689), .B(n6721), .ZN(n7463) );
  NAND2_X1 U5443 ( .A1(n7463), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U5444 ( .A1(n4697), .A2(n4407), .ZN(n7442) );
  OR2_X1 U5445 ( .A1(n7466), .A2(n7467), .ZN(n4697) );
  AND2_X1 U5446 ( .A1(n6914), .A2(n6743), .ZN(n10114) );
  NAND2_X1 U5447 ( .A1(n4570), .A2(n10095), .ZN(n4569) );
  NAND2_X1 U5448 ( .A1(n4582), .A2(n4776), .ZN(n4581) );
  INV_X1 U5449 ( .A(n6761), .ZN(n4776) );
  AND2_X1 U5450 ( .A1(n10114), .A2(n4773), .ZN(n4771) );
  NAND2_X1 U5451 ( .A1(n4775), .A2(n4774), .ZN(n4773) );
  NAND2_X1 U5452 ( .A1(n6744), .A2(n6663), .ZN(n4775) );
  INV_X1 U5453 ( .A(n5665), .ZN(n5666) );
  NAND2_X1 U5454 ( .A1(n5959), .A2(n5958), .ZN(n8759) );
  NOR2_X1 U5455 ( .A1(n5957), .A2(n5956), .ZN(n5958) );
  OAI211_X1 U5456 ( .C1(n8771), .C2(n4881), .A(n4879), .B(n4878), .ZN(n5959)
         );
  NOR2_X1 U5457 ( .A1(n5955), .A2(n8969), .ZN(n5957) );
  INV_X1 U5458 ( .A(n8817), .ZN(n9002) );
  OR2_X1 U5459 ( .A1(n5578), .A2(n6842), .ZN(n5052) );
  NOR2_X1 U5460 ( .A1(n5727), .A2(n6980), .ZN(n5717) );
  NAND2_X1 U5461 ( .A1(n5755), .A2(n5754), .ZN(n9075) );
  NOR2_X1 U5462 ( .A1(n5732), .A2(n9095), .ZN(n5736) );
  AOI21_X1 U5463 ( .B1(n8765), .B2(n7501), .A(n8759), .ZN(n6763) );
  INV_X1 U5464 ( .A(n6300), .ZN(n9096) );
  NAND2_X1 U5465 ( .A1(n5464), .A2(n5463), .ZN(n9107) );
  OR2_X1 U5466 ( .A1(n6301), .A2(n5724), .ZN(n5730) );
  XNOR2_X1 U5467 ( .A(n6167), .B(n6166), .ZN(n6872) );
  NAND2_X1 U5468 ( .A1(n6068), .A2(n6067), .ZN(n9815) );
  NAND2_X1 U5469 ( .A1(n6110), .A2(n6109), .ZN(n9769) );
  INV_X1 U5470 ( .A(n9389), .ZN(n9700) );
  CLKBUF_X1 U5471 ( .A(n9294), .Z(n9295) );
  AND2_X1 U5472 ( .A1(n9269), .A2(n9675), .ZN(n9317) );
  NAND2_X1 U5473 ( .A1(n6089), .A2(n6088), .ZN(n9794) );
  AOI21_X2 U5474 ( .B1(n6832), .B2(n9975), .A(n9965), .ZN(n9366) );
  AND2_X1 U5475 ( .A1(n9355), .A2(n9356), .ZN(n8045) );
  AND4_X1 U5476 ( .A1(n6450), .A2(n6449), .A3(n6448), .A4(n6447), .ZN(n9376)
         );
  OR2_X1 U5477 ( .A1(n8370), .A2(n8369), .ZN(n4473) );
  INV_X1 U5478 ( .A(n9360), .ZN(n9586) );
  OR2_X1 U5479 ( .A1(n9595), .A2(n6536), .ZN(n6521) );
  NAND2_X1 U5480 ( .A1(n9476), .A2(n9477), .ZN(n9475) );
  NAND2_X1 U5481 ( .A1(n9462), .A2(n4486), .ZN(n9476) );
  NAND2_X1 U5482 ( .A1(n9461), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4486) );
  NOR2_X1 U5483 ( .A1(n6041), .A2(n6045), .ZN(n7415) );
  OR2_X1 U5484 ( .A1(n7247), .A2(n4496), .ZN(n7421) );
  INV_X1 U5485 ( .A(n4494), .ZN(n4493) );
  OAI21_X1 U5486 ( .B1(n4495), .B2(n4499), .A(n7424), .ZN(n4494) );
  NOR2_X1 U5487 ( .A1(n9500), .A2(n4487), .ZN(n9921) );
  AND2_X1 U5488 ( .A1(n9501), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4487) );
  NOR2_X1 U5489 ( .A1(n9937), .A2(n9936), .ZN(n9935) );
  NAND2_X1 U5490 ( .A1(n4736), .A2(n4734), .ZN(n9949) );
  NAND2_X1 U5491 ( .A1(n4736), .A2(n9541), .ZN(n9946) );
  NAND2_X1 U5492 ( .A1(n4483), .A2(n9546), .ZN(n4482) );
  AOI21_X1 U5493 ( .B1(n9548), .B2(n9545), .A(n9947), .ZN(n9546) );
  NAND2_X1 U5494 ( .A1(n9549), .A2(n9951), .ZN(n4483) );
  OAI22_X1 U5495 ( .A1(n9548), .A2(n9944), .B1(n9934), .B2(n9549), .ZN(n4738)
         );
  OAI21_X1 U5496 ( .B1(n9606), .B2(n4956), .A(n4959), .ZN(n7875) );
  NAND2_X1 U5497 ( .A1(n7886), .A2(n7885), .ZN(n4550) );
  AOI21_X1 U5498 ( .B1(n9383), .B2(n9675), .A(n7884), .ZN(n7885) );
  NAND2_X1 U5499 ( .A1(n7883), .A2(n9962), .ZN(n7886) );
  NOR2_X1 U5500 ( .A1(n9710), .A2(n6531), .ZN(n7884) );
  NAND2_X1 U5501 ( .A1(n4924), .A2(n8280), .ZN(n9601) );
  NAND2_X1 U5502 ( .A1(n4967), .A2(n4966), .ZN(n9592) );
  INV_X1 U5503 ( .A(n9987), .ZN(n9965) );
  OAI21_X1 U5504 ( .B1(n8234), .B2(n10020), .A(n9738), .ZN(n6145) );
  INV_X1 U5505 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10193) );
  NOR2_X1 U5506 ( .A1(n9895), .A2(n9894), .ZN(n10153) );
  NOR2_X1 U5507 ( .A1(n9906), .A2(n9905), .ZN(n10145) );
  NOR2_X1 U5508 ( .A1(n10147), .A2(n10146), .ZN(n9905) );
  OAI21_X1 U5509 ( .B1(n5820), .B2(n5819), .A(n7166), .ZN(n5835) );
  NOR2_X1 U5510 ( .A1(n5837), .A2(n5821), .ZN(n4659) );
  NOR2_X1 U5511 ( .A1(n4663), .A2(n4661), .ZN(n4660) );
  NAND2_X1 U5512 ( .A1(n5825), .A2(n5824), .ZN(n4663) );
  NAND2_X1 U5513 ( .A1(n4411), .A2(n4533), .ZN(n4620) );
  NAND2_X1 U5514 ( .A1(n4535), .A2(n4534), .ZN(n4533) );
  NOR2_X1 U5515 ( .A1(n8122), .A2(n8123), .ZN(n4534) );
  NAND2_X1 U5516 ( .A1(n7055), .A2(n8290), .ZN(n4535) );
  NOR2_X1 U5517 ( .A1(n5846), .A2(n6634), .ZN(n4657) );
  MUX2_X1 U5518 ( .A(n8153), .B(n8152), .S(n4312), .Z(n8154) );
  NAND2_X1 U5519 ( .A1(n4325), .A2(n8146), .ZN(n4441) );
  NAND2_X1 U5520 ( .A1(n4647), .A2(n8926), .ZN(n5876) );
  OR2_X1 U5521 ( .A1(n4800), .A2(n5925), .ZN(n5867) );
  INV_X1 U5522 ( .A(n8191), .ZN(n4517) );
  OR2_X1 U5523 ( .A1(n8190), .A2(n9811), .ZN(n4515) );
  NAND2_X1 U5524 ( .A1(n4457), .A2(n4456), .ZN(n4631) );
  NOR2_X1 U5525 ( .A1(n8305), .A2(n4383), .ZN(n4456) );
  NAND2_X1 U5526 ( .A1(n8179), .A2(n8178), .ZN(n4457) );
  NOR2_X1 U5527 ( .A1(n5880), .A2(n6634), .ZN(n5881) );
  AOI21_X1 U5528 ( .B1(n6573), .B2(n9995), .A(n8286), .ZN(n8289) );
  NAND2_X1 U5529 ( .A1(n4641), .A2(n4638), .ZN(n4742) );
  AOI21_X1 U5530 ( .B1(n4642), .B2(n4640), .A(n4639), .ZN(n4638) );
  INV_X1 U5531 ( .A(n5907), .ZN(n4639) );
  OAI21_X1 U5532 ( .B1(n4640), .B2(n4637), .A(n4385), .ZN(n5906) );
  NOR2_X1 U5533 ( .A1(n8211), .A2(n9600), .ZN(n4626) );
  NAND2_X1 U5534 ( .A1(n8198), .A2(n8238), .ZN(n4455) );
  NOR2_X1 U5535 ( .A1(n4930), .A2(n4929), .ZN(n8149) );
  INV_X1 U5536 ( .A(n8151), .ZN(n4930) );
  OAI21_X1 U5537 ( .B1(n6837), .B2(P1_DATAO_REG_9__SCAN_IN), .A(n5167), .ZN(
        n5170) );
  NAND2_X1 U5538 ( .A1(n6837), .A2(n6883), .ZN(n5167) );
  NAND2_X1 U5539 ( .A1(n4667), .A2(n5913), .ZN(n4666) );
  AOI21_X1 U5540 ( .B1(n4805), .B2(n4566), .A(n4416), .ZN(n4565) );
  INV_X1 U5541 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5381) );
  INV_X1 U5542 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4998) );
  AOI211_X1 U5543 ( .C1(n8320), .C2(n8319), .A(n8318), .B(n8317), .ZN(n8343)
         );
  INV_X1 U5544 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5963) );
  NOR2_X1 U5545 ( .A1(n4611), .A2(n4606), .ZN(n4605) );
  INV_X1 U5546 ( .A(n5395), .ZN(n4606) );
  AOI21_X1 U5547 ( .B1(n4614), .B2(n4610), .A(n4609), .ZN(n4608) );
  INV_X1 U5548 ( .A(n5472), .ZN(n4609) );
  OR2_X1 U5549 ( .A1(n4611), .A2(n4604), .ZN(n4603) );
  NAND2_X1 U5550 ( .A1(n5396), .A2(n5395), .ZN(n4604) );
  INV_X1 U5551 ( .A(SI_19_), .ZN(n10166) );
  INV_X1 U5552 ( .A(SI_21_), .ZN(n5410) );
  INV_X1 U5553 ( .A(n5432), .ZN(n5413) );
  INV_X1 U5554 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5354) );
  INV_X1 U5555 ( .A(SI_17_), .ZN(n5328) );
  NAND2_X1 U5556 ( .A1(n4545), .A2(n5123), .ZN(n5125) );
  INV_X1 U5557 ( .A(n5124), .ZN(n4545) );
  OAI21_X1 U5558 ( .B1(n6837), .B2(n4594), .A(n4593), .ZN(n4592) );
  NAND2_X1 U5559 ( .A1(n6837), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4593) );
  OAI21_X1 U5560 ( .B1(n5093), .B2(n5092), .A(n5091), .ZN(n5129) );
  NAND2_X1 U5561 ( .A1(n5093), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5091) );
  INV_X1 U5562 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5023) );
  INV_X1 U5563 ( .A(n5930), .ZN(n5924) );
  NAND2_X1 U5564 ( .A1(n4789), .A2(n8616), .ZN(n4788) );
  NOR2_X1 U5565 ( .A1(n4791), .A2(n4790), .ZN(n4789) );
  INV_X1 U5566 ( .A(n6642), .ZN(n4791) );
  INV_X1 U5567 ( .A(n7440), .ZN(n4574) );
  NOR2_X1 U5568 ( .A1(n8676), .A2(n10237), .ZN(n4889) );
  NAND2_X1 U5569 ( .A1(n4892), .A2(n4891), .ZN(n4890) );
  OAI21_X1 U5570 ( .B1(n8693), .B2(n4561), .A(n4559), .ZN(n6659) );
  INV_X1 U5571 ( .A(n8707), .ZN(n4561) );
  AND2_X1 U5572 ( .A1(n4560), .A2(n4421), .ZN(n4559) );
  AND2_X1 U5573 ( .A1(n6659), .A2(n8727), .ZN(n6661) );
  AND2_X1 U5574 ( .A1(n5953), .A2(n5644), .ZN(n4883) );
  AND2_X1 U5575 ( .A1(n5502), .A2(n4681), .ZN(n4680) );
  INV_X1 U5576 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n4681) );
  INV_X1 U5577 ( .A(n5504), .ZN(n5503) );
  INV_X1 U5578 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4675) );
  INV_X1 U5579 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5265) );
  INV_X1 U5580 ( .A(n5267), .ZN(n5266) );
  INV_X1 U5581 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n4685) );
  INV_X1 U5582 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5181) );
  INV_X1 U5583 ( .A(n5183), .ZN(n5182) );
  INV_X1 U5584 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5080) );
  AND2_X1 U5585 ( .A1(n5711), .A2(n6634), .ZN(n5713) );
  INV_X1 U5586 ( .A(n4874), .ZN(n4873) );
  AND2_X1 U5587 ( .A1(n4875), .A2(n5631), .ZN(n4874) );
  INV_X1 U5588 ( .A(n5627), .ZN(n4862) );
  OR2_X1 U5589 ( .A1(n9154), .A2(n8912), .ZN(n5866) );
  NOR2_X1 U5590 ( .A1(n4787), .A2(n5849), .ZN(n4785) );
  INV_X1 U5591 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5098) );
  AND2_X1 U5592 ( .A1(n5727), .A2(n5726), .ZN(n6283) );
  INV_X1 U5593 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U5594 ( .A1(n4322), .A2(n5357), .ZN(n5670) );
  OR2_X1 U5595 ( .A1(n5261), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5280) );
  INV_X1 U5596 ( .A(n7773), .ZN(n7764) );
  NOR2_X1 U5597 ( .A1(n6482), .A2(n10160), .ZN(n4480) );
  AND2_X1 U5598 ( .A1(n4850), .A2(n9264), .ZN(n4849) );
  OR2_X1 U5599 ( .A1(n7961), .A2(n4851), .ZN(n4850) );
  INV_X1 U5600 ( .A(n7966), .ZN(n4851) );
  NOR2_X1 U5601 ( .A1(n4451), .A2(n8273), .ZN(n4450) );
  NAND2_X1 U5602 ( .A1(n8272), .A2(n4378), .ZN(n4451) );
  OR3_X1 U5603 ( .A1(n9634), .A2(n9668), .A3(n8268), .ZN(n8269) );
  NOR2_X1 U5604 ( .A1(n8335), .A2(n8333), .ZN(n4449) );
  INV_X1 U5605 ( .A(n8222), .ZN(n4470) );
  NAND2_X1 U5606 ( .A1(n4469), .A2(n8331), .ZN(n4468) );
  AOI211_X1 U5607 ( .C1(n8348), .C2(n9382), .A(n8228), .B(n8335), .ZN(n8232)
         );
  INV_X1 U5608 ( .A(n7418), .ZN(n4728) );
  INV_X1 U5609 ( .A(n9953), .ZN(n4506) );
  INV_X1 U5610 ( .A(n9537), .ZN(n4507) );
  INV_X1 U5611 ( .A(n9538), .ZN(n4732) );
  INV_X1 U5612 ( .A(n9543), .ZN(n4731) );
  INV_X1 U5613 ( .A(n4525), .ZN(n4524) );
  OAI21_X1 U5614 ( .B1(n4922), .B2(n8180), .A(n8193), .ZN(n4525) );
  OAI21_X1 U5615 ( .B1(n6451), .B2(n4941), .A(n6609), .ZN(n4939) );
  NAND2_X1 U5616 ( .A1(n4475), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6454) );
  INV_X1 U5617 ( .A(n6445), .ZN(n4475) );
  NAND2_X1 U5618 ( .A1(n4476), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6445) );
  INV_X1 U5619 ( .A(n6437), .ZN(n4476) );
  NOR2_X1 U5620 ( .A1(n6605), .A2(n4938), .ZN(n4937) );
  INV_X1 U5621 ( .A(n6604), .ZN(n4938) );
  INV_X1 U5622 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6427) );
  OR2_X1 U5623 ( .A1(n6428), .A2(n6427), .ZN(n6437) );
  NOR2_X1 U5624 ( .A1(n6597), .A2(n4765), .ZN(n4762) );
  NOR2_X1 U5625 ( .A1(n10046), .A2(n9831), .ZN(n6044) );
  NOR2_X1 U5626 ( .A1(n6402), .A2(n6401), .ZN(n6403) );
  AND2_X1 U5627 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n6323) );
  AND2_X1 U5628 ( .A1(n7121), .A2(n7285), .ZN(n6583) );
  NAND2_X1 U5629 ( .A1(n9402), .A2(n7302), .ZN(n8137) );
  INV_X1 U5630 ( .A(n8358), .ZN(n8365) );
  INV_X1 U5631 ( .A(n6017), .ZN(n4464) );
  INV_X1 U5632 ( .A(n8369), .ZN(n8363) );
  NAND2_X1 U5633 ( .A1(n4585), .A2(n5495), .ZN(n5513) );
  AND2_X1 U5634 ( .A1(n5514), .A2(n5499), .ZN(n5512) );
  INV_X1 U5635 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6123) );
  OR2_X1 U5636 ( .A1(n5347), .A2(n5352), .ZN(n5369) );
  INV_X1 U5637 ( .A(n5347), .ZN(n4750) );
  INV_X1 U5638 ( .A(n4753), .ZN(n4752) );
  OAI21_X1 U5639 ( .B1(n5290), .B2(n4754), .A(n5311), .ZN(n4753) );
  NAND2_X1 U5640 ( .A1(n4748), .A2(n5225), .ZN(n4747) );
  NAND2_X1 U5641 ( .A1(n5093), .A2(n6857), .ZN(n4467) );
  INV_X1 U5642 ( .A(n5071), .ZN(n4623) );
  NAND2_X1 U5643 ( .A1(n4622), .A2(n4916), .ZN(n4621) );
  NAND2_X1 U5644 ( .A1(n4671), .A2(n5098), .ZN(n5107) );
  INV_X1 U5645 ( .A(n5105), .ZN(n4671) );
  NAND2_X1 U5646 ( .A1(n7229), .A2(n5080), .ZN(n5105) );
  NAND2_X1 U5647 ( .A1(n6217), .A2(n6216), .ZN(n7692) );
  AOI21_X1 U5648 ( .B1(n4909), .B2(n7693), .A(n4365), .ZN(n4908) );
  INV_X1 U5649 ( .A(n4904), .ZN(n4903) );
  INV_X1 U5650 ( .A(n4902), .ZN(n4901) );
  OAI21_X1 U5651 ( .B1(n4905), .B2(n4903), .A(n8452), .ZN(n4902) );
  CLKBUF_X1 U5652 ( .A(n8431), .Z(n8459) );
  NAND2_X1 U5653 ( .A1(n8476), .A2(n4907), .ZN(n8550) );
  AND2_X1 U5654 ( .A1(n4362), .A2(n6241), .ZN(n4907) );
  NAND2_X1 U5655 ( .A1(n8560), .A2(n8559), .ZN(n8558) );
  OR2_X1 U5656 ( .A1(n6270), .A2(n6269), .ZN(n8077) );
  NAND2_X1 U5657 ( .A1(n5926), .A2(n4672), .ZN(n5800) );
  NOR2_X1 U5658 ( .A1(n4673), .A2(n5796), .ZN(n4672) );
  OR2_X1 U5659 ( .A1(n4674), .A2(n5942), .ZN(n4673) );
  OR2_X1 U5660 ( .A1(n5943), .A2(n5942), .ZN(n4651) );
  AND2_X1 U5661 ( .A1(n5510), .A2(n5509), .ZN(n6315) );
  OR2_X1 U5662 ( .A1(n6965), .A2(n6964), .ZN(n6967) );
  XNOR2_X1 U5663 ( .A(n6674), .B(n6708), .ZN(n10066) );
  AND2_X1 U5664 ( .A1(n6643), .A2(n4788), .ZN(n10068) );
  NAND2_X1 U5665 ( .A1(n8634), .A2(n6678), .ZN(n6679) );
  XNOR2_X1 U5666 ( .A(n6679), .B(n6925), .ZN(n6923) );
  NAND2_X1 U5667 ( .A1(n8660), .A2(n4410), .ZN(n8683) );
  AND2_X1 U5668 ( .A1(n6693), .A2(n8665), .ZN(n4892) );
  NAND2_X1 U5669 ( .A1(n4797), .A2(n4336), .ZN(n8666) );
  OR2_X1 U5670 ( .A1(n8678), .A2(n8962), .ZN(n4796) );
  NAND2_X1 U5671 ( .A1(n8693), .A2(n6658), .ZN(n8708) );
  AOI21_X1 U5672 ( .B1(n8697), .B2(n8696), .A(n4703), .ZN(n8711) );
  AND2_X1 U5673 ( .A1(n7033), .A2(n6735), .ZN(n4703) );
  NAND2_X1 U5674 ( .A1(n4777), .A2(n6664), .ZN(n4774) );
  AND2_X1 U5675 ( .A1(n4880), .A2(n4884), .ZN(n4879) );
  INV_X1 U5676 ( .A(n4885), .ZN(n4884) );
  NAND2_X1 U5677 ( .A1(n4883), .A2(n8770), .ZN(n4880) );
  OAI21_X1 U5678 ( .B1(n5953), .B2(n5644), .A(n8949), .ZN(n4885) );
  NAND2_X1 U5679 ( .A1(n4882), .A2(n8768), .ZN(n4881) );
  INV_X1 U5680 ( .A(n5953), .ZN(n4882) );
  AND2_X1 U5681 ( .A1(n4677), .A2(n10154), .ZN(n4676) );
  NAND2_X1 U5682 ( .A1(n5337), .A2(n4677), .ZN(n5389) );
  NAND2_X1 U5683 ( .A1(n5337), .A2(n5336), .ZN(n5361) );
  OR2_X1 U5684 ( .A1(n5321), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U5685 ( .A1(n5266), .A2(n5265), .ZN(n5285) );
  NAND2_X1 U5686 ( .A1(n5182), .A2(n4682), .ZN(n5267) );
  AND2_X1 U5687 ( .A1(n4683), .A2(n5249), .ZN(n4682) );
  INV_X1 U5688 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U5689 ( .A1(n5182), .A2(n4351), .ZN(n5234) );
  OR2_X1 U5690 ( .A1(n5157), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U5691 ( .A1(n5182), .A2(n5181), .ZN(n5214) );
  NAND2_X1 U5692 ( .A1(n5164), .A2(n5825), .ZN(n7576) );
  NAND2_X1 U5693 ( .A1(n5139), .A2(n5138), .ZN(n5157) );
  INV_X1 U5694 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5138) );
  INV_X1 U5695 ( .A(n5140), .ZN(n5139) );
  NAND4_X1 U5696 ( .A1(n5098), .A2(n4670), .A3(n7229), .A4(n5080), .ZN(n5140)
         );
  INV_X1 U5697 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4670) );
  INV_X1 U5698 ( .A(n5822), .ZN(n4783) );
  CLKBUF_X1 U5699 ( .A(n7112), .Z(n4433) );
  INV_X1 U5700 ( .A(n6892), .ZN(n6303) );
  OR2_X1 U5701 ( .A1(n7407), .A2(n5712), .ZN(n6302) );
  AND2_X1 U5702 ( .A1(n5723), .A2(n5722), .ZN(n5727) );
  OR2_X1 U5703 ( .A1(n5915), .A2(n5777), .ZN(n8784) );
  AND2_X1 U5704 ( .A1(n8812), .A2(n5899), .ZN(n8825) );
  OR2_X1 U5705 ( .A1(n5452), .A2(n5451), .ZN(n5453) );
  NAND2_X1 U5706 ( .A1(n8877), .A2(n5630), .ZN(n5632) );
  NAND2_X1 U5707 ( .A1(n5632), .A2(n4874), .ZN(n8869) );
  INV_X1 U5708 ( .A(n5630), .ZN(n8878) );
  OR2_X1 U5709 ( .A1(n8921), .A2(n5778), .ZN(n8943) );
  NAND2_X1 U5710 ( .A1(n5614), .A2(n4466), .ZN(n7713) );
  OAI22_X1 U5711 ( .A1(n7386), .A2(n5609), .B1(n8604), .B2(n7631), .ZN(n7458)
         );
  NAND2_X1 U5712 ( .A1(n6283), .A2(n6892), .ZN(n6296) );
  NAND2_X1 U5713 ( .A1(n5687), .A2(n8110), .ZN(n6891) );
  AND2_X1 U5714 ( .A1(n6749), .A2(n5708), .ZN(n6892) );
  AND2_X1 U5715 ( .A1(n6748), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5708) );
  INV_X1 U5716 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5678) );
  INV_X1 U5717 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5207) );
  XNOR2_X1 U5718 ( .A(n5095), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6715) );
  AND2_X1 U5719 ( .A1(n8056), .A2(n8055), .ZN(n8099) );
  NAND2_X1 U5720 ( .A1(n4480), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U5721 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6391) );
  AOI21_X1 U5722 ( .B1(n4838), .B2(n4840), .A(n4835), .ZN(n4834) );
  INV_X1 U5723 ( .A(n9276), .ZN(n4835) );
  INV_X1 U5724 ( .A(n4480), .ZN(n6484) );
  NAND2_X1 U5725 ( .A1(n4837), .A2(n4842), .ZN(n9200) );
  NAND2_X1 U5726 ( .A1(n9304), .A2(n4346), .ZN(n4837) );
  AND2_X1 U5727 ( .A1(n8011), .A2(n8010), .ZN(n9322) );
  NOR2_X1 U5728 ( .A1(n6794), .A2(n4526), .ZN(n6796) );
  NOR2_X1 U5729 ( .A1(n4527), .A2(n7278), .ZN(n4526) );
  INV_X1 U5730 ( .A(n8063), .ZN(n4527) );
  INV_X1 U5731 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U5732 ( .A1(n7343), .A2(n7342), .ZN(n7667) );
  CLKBUF_X1 U5733 ( .A(n9248), .Z(n9249) );
  AND2_X1 U5734 ( .A1(n7952), .A2(n7951), .ZN(n7958) );
  AND2_X1 U5735 ( .A1(n4587), .A2(n8356), .ZN(n8370) );
  INV_X1 U5736 ( .A(n8333), .ZN(n4588) );
  NAND2_X1 U5737 ( .A1(n4591), .A2(n4590), .ZN(n4589) );
  INV_X1 U5738 ( .A(n6551), .ZN(n6536) );
  AND4_X1 U5739 ( .A1(n6408), .A2(n6407), .A3(n6406), .A4(n6405), .ZN(n7910)
         );
  OR2_X1 U5740 ( .A1(n4719), .A2(n4718), .ZN(n4717) );
  INV_X1 U5741 ( .A(n4721), .ZN(n4718) );
  OR2_X1 U5742 ( .A1(n6065), .A2(n6037), .ZN(n6040) );
  INV_X1 U5743 ( .A(n4496), .ZN(n4495) );
  OR2_X1 U5744 ( .A1(n7515), .A2(n7516), .ZN(n4489) );
  NAND2_X1 U5745 ( .A1(n9498), .A2(n9940), .ZN(n4712) );
  AND2_X1 U5746 ( .A1(n9524), .A2(n9523), .ZN(n9525) );
  NOR2_X1 U5747 ( .A1(n9945), .A2(n4735), .ZN(n4734) );
  INV_X1 U5748 ( .A(n9541), .ZN(n4735) );
  NAND2_X1 U5749 ( .A1(n9539), .A2(n9538), .ZN(n4736) );
  NAND2_X1 U5750 ( .A1(n4600), .A2(n6121), .ZN(n8241) );
  NAND2_X1 U5751 ( .A1(n8379), .A2(n6058), .ZN(n4600) );
  OR2_X1 U5752 ( .A1(n6569), .A2(n8067), .ZN(n8226) );
  INV_X1 U5753 ( .A(n6569), .ZN(n9569) );
  OR2_X1 U5754 ( .A1(n6623), .A2(n4963), .ZN(n4962) );
  NAND2_X1 U5755 ( .A1(n9598), .A2(n8316), .ZN(n7893) );
  NAND2_X1 U5756 ( .A1(n9641), .A2(n4761), .ZN(n9614) );
  AND2_X1 U5757 ( .A1(n9641), .A2(n4327), .ZN(n9593) );
  INV_X1 U5758 ( .A(n9600), .ZN(n6522) );
  INV_X1 U5759 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9204) );
  INV_X1 U5760 ( .A(n4479), .ZN(n6505) );
  NAND2_X1 U5761 ( .A1(n9641), .A2(n9625), .ZN(n9613) );
  AOI21_X1 U5762 ( .B1(n4944), .B2(n4951), .A(n4329), .ZN(n4943) );
  NOR2_X1 U5763 ( .A1(n9798), .A2(n9789), .ZN(n4756) );
  AND2_X1 U5764 ( .A1(n9713), .A2(n9719), .ZN(n9691) );
  AND2_X1 U5765 ( .A1(n9723), .A2(n9728), .ZN(n9713) );
  NAND2_X1 U5766 ( .A1(n4478), .A2(n4377), .ZN(n6420) );
  INV_X1 U5767 ( .A(n6414), .ZN(n4478) );
  NAND2_X1 U5768 ( .A1(n4477), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6428) );
  INV_X1 U5769 ( .A(n6420), .ZN(n4477) );
  NAND2_X1 U5770 ( .A1(n6599), .A2(n6598), .ZN(n6600) );
  AND2_X1 U5771 ( .A1(n8165), .A2(n8156), .ZN(n7650) );
  AND2_X1 U5772 ( .A1(n4764), .A2(n4763), .ZN(n7653) );
  AOI21_X1 U5773 ( .B1(n4316), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6349), .ZN(
        n8126) );
  NOR2_X2 U5774 ( .A1(n7300), .A2(n10004), .ZN(n7494) );
  NAND2_X1 U5775 ( .A1(n6773), .A2(n6772), .ZN(n7616) );
  NAND2_X1 U5776 ( .A1(n6116), .A2(n6115), .ZN(n9753) );
  INV_X1 U5777 ( .A(n4453), .ZN(n4942) );
  NAND2_X1 U5778 ( .A1(n6863), .A2(n6058), .ZN(n4542) );
  NAND2_X1 U5779 ( .A1(n6844), .A2(n6058), .ZN(n4630) );
  INV_X1 U5780 ( .A(n9724), .ZN(n10012) );
  OAI21_X1 U5781 ( .B1(n6860), .B2(P1_D_REG_0__SCAN_IN), .A(n9855), .ZN(n7293)
         );
  AND2_X1 U5782 ( .A1(n6187), .A2(n6186), .ZN(n6767) );
  NOR2_X1 U5783 ( .A1(n6183), .A2(n6813), .ZN(n6187) );
  OR2_X1 U5784 ( .A1(n6169), .A2(n6831), .ZN(n6183) );
  AND2_X1 U5785 ( .A1(n6168), .A2(n6872), .ZN(n7290) );
  XNOR2_X1 U5786 ( .A(n5457), .B(n5456), .ZN(n7638) );
  OAI21_X1 U5787 ( .B1(n5435), .B2(n5417), .A(n5416), .ZN(n5457) );
  XNOR2_X1 U5788 ( .A(n5440), .B(n5439), .ZN(n7527) );
  INV_X1 U5789 ( .A(n6149), .ZN(n6128) );
  NOR2_X1 U5790 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  AND2_X1 U5791 ( .A1(n6093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6094) );
  AND2_X1 U5792 ( .A1(n6020), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n6095) );
  CLKBUF_X1 U5793 ( .A(n6018), .Z(n6019) );
  INV_X1 U5794 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4932) );
  NAND2_X1 U5795 ( .A1(n4755), .A2(n5293), .ZN(n5312) );
  AND2_X1 U5796 ( .A1(n5201), .A2(n5223), .ZN(n4749) );
  XNOR2_X1 U5797 ( .A(n5226), .B(n5223), .ZN(n6858) );
  OAI21_X1 U5798 ( .B1(n5166), .B2(n5165), .A(n5196), .ZN(n5172) );
  OR2_X1 U5799 ( .A1(n6026), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6065) );
  XNOR2_X1 U5800 ( .A(n5088), .B(SI_5_), .ZN(n5123) );
  OAI21_X1 U5801 ( .B1(n6837), .B2(n6839), .A(n5045), .ZN(n5027) );
  NAND2_X1 U5802 ( .A1(n8558), .A2(n6213), .ZN(n7628) );
  AND2_X1 U5803 ( .A1(n5491), .A2(n5490), .ZN(n8427) );
  AND2_X1 U5804 ( .A1(n6197), .A2(n8609), .ZN(n6198) );
  NAND2_X1 U5805 ( .A1(n4439), .A2(n4905), .ZN(n4900) );
  AND4_X1 U5806 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n8970)
         );
  NAND2_X1 U5807 ( .A1(n8478), .A2(n8477), .ZN(n8476) );
  NAND2_X1 U5808 ( .A1(n8476), .A2(n6241), .ZN(n8484) );
  NAND2_X1 U5809 ( .A1(n7692), .A2(n6220), .ZN(n8498) );
  NAND2_X1 U5810 ( .A1(n4439), .A2(n8443), .ZN(n8505) );
  NAND2_X1 U5811 ( .A1(n4906), .A2(n6236), .ZN(n8583) );
  XNOR2_X1 U5812 ( .A(n5594), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5949) );
  OAI21_X1 U5813 ( .B1(n5595), .B2(n5593), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5594) );
  INV_X1 U5814 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5592) );
  AND2_X1 U5815 ( .A1(n5765), .A2(n5764), .ZN(n8753) );
  NAND2_X1 U5816 ( .A1(n5567), .A2(n5566), .ZN(n8774) );
  NAND2_X1 U5817 ( .A1(n5546), .A2(n5545), .ZN(n8786) );
  INV_X1 U5818 ( .A(n6315), .ZN(n8815) );
  INV_X1 U5819 ( .A(n8427), .ZN(n8826) );
  NAND2_X1 U5820 ( .A1(n5471), .A2(n5470), .ZN(n8846) );
  NAND2_X1 U5821 ( .A1(n5431), .A2(n5430), .ZN(n8861) );
  NAND2_X1 U5822 ( .A1(n5450), .A2(n5449), .ZN(n8870) );
  NAND2_X1 U5823 ( .A1(n5408), .A2(n5407), .ZN(n8879) );
  NAND2_X1 U5824 ( .A1(n5304), .A2(n5303), .ZN(n8939) );
  OR2_X1 U5825 ( .A1(n5054), .A2(n5031), .ZN(n5035) );
  OR2_X1 U5826 ( .A1(n5236), .A2(n10163), .ZN(n5032) );
  AND2_X1 U5827 ( .A1(n6755), .A2(n9182), .ZN(n6914) );
  NAND2_X1 U5828 ( .A1(n6968), .A2(n4701), .ZN(n8622) );
  OR2_X1 U5829 ( .A1(n6702), .A2(n6976), .ZN(n4701) );
  NOR2_X1 U5830 ( .A1(n10075), .A2(n4707), .ZN(n8633) );
  AND2_X1 U5831 ( .A1(n6707), .A2(n6708), .ZN(n4707) );
  NAND2_X1 U5832 ( .A1(n4809), .A2(n4808), .ZN(n8649) );
  NAND2_X1 U5833 ( .A1(n4692), .A2(n4695), .ZN(n8654) );
  NAND2_X1 U5834 ( .A1(n7466), .A2(n4693), .ZN(n4692) );
  INV_X1 U5835 ( .A(n4809), .ZN(n7807) );
  OAI21_X1 U5836 ( .B1(n6652), .B2(n4805), .A(n4566), .ZN(n7804) );
  NAND2_X1 U5837 ( .A1(n4687), .A2(n4688), .ZN(n7800) );
  AND2_X1 U5838 ( .A1(n6757), .A2(n6756), .ZN(n10111) );
  INV_X1 U5839 ( .A(n4558), .ZN(n8680) );
  INV_X1 U5840 ( .A(n4579), .ZN(n8692) );
  NAND2_X1 U5841 ( .A1(n4579), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4578) );
  AND2_X1 U5842 ( .A1(n9008), .A2(n7157), .ZN(n8764) );
  NAND2_X1 U5843 ( .A1(n4864), .A2(n5607), .ZN(n7368) );
  NAND2_X1 U5844 ( .A1(n4867), .A2(n4868), .ZN(n4864) );
  NAND2_X1 U5845 ( .A1(n4868), .A2(n4869), .ZN(n7152) );
  NAND2_X1 U5846 ( .A1(n5605), .A2(n5606), .ZN(n7165) );
  NAND2_X1 U5847 ( .A1(n5066), .A2(n5821), .ZN(n7164) );
  OR2_X1 U5848 ( .A1(n5060), .A2(n7874), .ZN(n4888) );
  INV_X1 U5849 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7229) );
  INV_X1 U5850 ( .A(n8989), .ZN(n9003) );
  INV_X2 U5851 ( .A(n8993), .ZN(n9008) );
  CLKBUF_X1 U5852 ( .A(n7041), .Z(n7145) );
  NAND2_X1 U5853 ( .A1(n6985), .A2(n9002), .ZN(n8991) );
  AND2_X1 U5854 ( .A1(n6988), .A2(n8989), .ZN(n8993) );
  AOI21_X1 U5855 ( .B1(n8379), .B2(n5537), .A(n5747), .ZN(n9081) );
  NAND2_X1 U5856 ( .A1(n5539), .A2(n5538), .ZN(n9084) );
  NAND2_X1 U5857 ( .A1(n5520), .A2(n5519), .ZN(n9090) );
  NAND2_X1 U5858 ( .A1(n5481), .A2(n5480), .ZN(n9102) );
  NAND2_X1 U5859 ( .A1(n5388), .A2(n5387), .ZN(n9130) );
  NAND2_X1 U5860 ( .A1(n5360), .A2(n5359), .ZN(n9136) );
  NAND2_X1 U5861 ( .A1(n8896), .A2(n5627), .ZN(n8888) );
  NAND2_X1 U5862 ( .A1(n4740), .A2(n5335), .ZN(n9142) );
  NAND2_X1 U5863 ( .A1(n7174), .A2(n5537), .ZN(n4740) );
  AND2_X1 U5864 ( .A1(n8901), .A2(n8900), .ZN(n9140) );
  NAND2_X1 U5865 ( .A1(n5319), .A2(n5318), .ZN(n9148) );
  AOI21_X1 U5866 ( .B1(n5275), .B2(n4802), .A(n4321), .ZN(n8907) );
  AND2_X1 U5867 ( .A1(n8932), .A2(n8931), .ZN(n9152) );
  NAND2_X1 U5868 ( .A1(n5282), .A2(n5281), .ZN(n9160) );
  NAND2_X1 U5869 ( .A1(n5264), .A2(n5263), .ZN(n9166) );
  INV_X1 U5870 ( .A(n4786), .ZN(n8973) );
  AOI21_X1 U5871 ( .B1(n7708), .B2(n5850), .A(n4787), .ZN(n4786) );
  INV_X1 U5872 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9176) );
  INV_X1 U5873 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5009) );
  INV_X1 U5874 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U5875 ( .A1(n5681), .A2(n5684), .ZN(n7849) );
  INV_X1 U5876 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7850) );
  INV_X1 U5877 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7826) );
  CLKBUF_X1 U5878 ( .A(n5686), .Z(n5703) );
  INV_X1 U5879 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7643) );
  INV_X1 U5880 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7528) );
  INV_X1 U5881 ( .A(n6191), .ZN(n7529) );
  INV_X1 U5882 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7330) );
  INV_X1 U5883 ( .A(n6697), .ZN(n7328) );
  INV_X1 U5884 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7253) );
  INV_X1 U5885 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7264) );
  INV_X1 U5886 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6906) );
  INV_X1 U5887 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6888) );
  NAND2_X1 U5888 ( .A1(n4432), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4766) );
  XNOR2_X1 U5889 ( .A(n5022), .B(n4555), .ZN(n6838) );
  INV_X1 U5890 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4555) );
  CLKBUF_X1 U5891 ( .A(n7766), .Z(n7348) );
  CLKBUF_X1 U5892 ( .A(n9188), .Z(n9189) );
  NAND2_X1 U5893 ( .A1(n6120), .A2(n6119), .ZN(n9742) );
  NAND2_X1 U5894 ( .A1(n9304), .A2(n8001), .ZN(n4844) );
  AOI21_X1 U5895 ( .B1(n4829), .B2(n4831), .A(n4335), .ZN(n4827) );
  AOI21_X1 U5896 ( .B1(n7919), .B2(n4833), .A(n4830), .ZN(n4829) );
  NAND2_X1 U5897 ( .A1(n9254), .A2(n7966), .ZN(n9266) );
  AND2_X1 U5898 ( .A1(n9269), .A2(n9673), .ZN(n9371) );
  NAND2_X1 U5899 ( .A1(n4853), .A2(n6812), .ZN(n6819) );
  AND4_X1 U5900 ( .A1(n6361), .A2(n6360), .A3(n6359), .A4(n6358), .ZN(n9289)
         );
  INV_X1 U5901 ( .A(n7656), .ZN(n10046) );
  AOI21_X1 U5902 ( .B1(n9295), .B2(n4832), .A(n4831), .ZN(n4828) );
  AND4_X1 U5903 ( .A1(n6419), .A2(n6418), .A3(n6417), .A4(n6416), .ZN(n9336)
         );
  NAND2_X1 U5904 ( .A1(n9673), .A2(n6573), .ZN(n7057) );
  AND2_X1 U5905 ( .A1(n6828), .A2(n6827), .ZN(n9349) );
  INV_X1 U5906 ( .A(n9371), .ZN(n9359) );
  NAND2_X1 U5907 ( .A1(n4858), .A2(n4857), .ZN(n4856) );
  INV_X1 U5908 ( .A(n9355), .ZN(n4857) );
  NAND2_X1 U5909 ( .A1(n9357), .A2(n9356), .ZN(n4858) );
  AND2_X1 U5910 ( .A1(n6534), .A2(n6524), .ZN(n9363) );
  INV_X1 U5911 ( .A(n9349), .ZN(n9372) );
  INV_X1 U5912 ( .A(n7958), .ZN(n9370) );
  INV_X1 U5913 ( .A(n9366), .ZN(n9378) );
  NAND2_X1 U5914 ( .A1(n6512), .A2(n6511), .ZN(n9386) );
  INV_X1 U5915 ( .A(n7790), .ZN(n9398) );
  NAND2_X1 U5916 ( .A1(n4316), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6337) );
  INV_X1 U5917 ( .A(P1_U3973), .ZN(n9403) );
  NAND2_X1 U5918 ( .A1(n9437), .A2(n9438), .ZN(n9436) );
  NAND2_X1 U5919 ( .A1(n7087), .A2(n4491), .ZN(n9437) );
  NAND2_X1 U5920 ( .A1(n4463), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4491) );
  NAND2_X1 U5921 ( .A1(n9436), .A2(n4490), .ZN(n9450) );
  NAND2_X1 U5922 ( .A1(n6014), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4490) );
  NAND2_X1 U5923 ( .A1(n9450), .A2(n9451), .ZN(n9449) );
  NOR2_X1 U5924 ( .A1(n9430), .A2(n7017), .ZN(n9443) );
  NAND2_X1 U5925 ( .A1(n9432), .A2(n4720), .ZN(n4716) );
  NAND2_X1 U5926 ( .A1(n9463), .A2(n9464), .ZN(n9462) );
  NAND2_X1 U5927 ( .A1(n9475), .A2(n4415), .ZN(n7005) );
  NAND2_X1 U5928 ( .A1(n7241), .A2(n4729), .ZN(n7243) );
  INV_X1 U5929 ( .A(n4724), .ZN(n7417) );
  INV_X1 U5930 ( .A(n4489), .ZN(n9481) );
  AND2_X1 U5931 ( .A1(n6059), .A2(n6054), .ZN(n9489) );
  AND2_X1 U5932 ( .A1(n4489), .A2(n4488), .ZN(n9485) );
  NAND2_X1 U5933 ( .A1(n9482), .A2(n7511), .ZN(n4488) );
  AND2_X1 U5934 ( .A1(n9485), .A2(n9484), .ZN(n9500) );
  INV_X1 U5935 ( .A(n4485), .ZN(n9510) );
  AND2_X1 U5936 ( .A1(n4714), .A2(n4357), .ZN(n9518) );
  NAND2_X1 U5937 ( .A1(n6874), .A2(n6876), .ZN(n9960) );
  INV_X1 U5938 ( .A(n8241), .ZN(n9740) );
  AOI22_X1 U5939 ( .A1(n9586), .A2(n9673), .B1(n9585), .B2(n9675), .ZN(n9587)
         );
  AOI21_X1 U5940 ( .B1(n9747), .B2(n9991), .A(n7887), .ZN(n4548) );
  INV_X1 U5941 ( .A(n9753), .ZN(n9367) );
  NAND2_X1 U5942 ( .A1(n4958), .A2(n6620), .ZN(n7888) );
  NAND2_X1 U5943 ( .A1(n4967), .A2(n4964), .ZN(n4958) );
  NAND2_X1 U5944 ( .A1(n6112), .A2(n6111), .ZN(n9764) );
  NAND2_X1 U5945 ( .A1(n4923), .A2(n8314), .ZN(n9647) );
  NAND2_X1 U5946 ( .A1(n4946), .A2(n4947), .ZN(n9669) );
  NAND2_X1 U5947 ( .A1(n9690), .A2(n4950), .ZN(n4946) );
  OAI21_X1 U5948 ( .B1(n9690), .B2(n4349), .A(n6613), .ZN(n9685) );
  NAND2_X1 U5949 ( .A1(n6467), .A2(n8200), .ZN(n9698) );
  NAND2_X1 U5950 ( .A1(n4447), .A2(n4922), .ZN(n4523) );
  NAND2_X1 U5951 ( .A1(n6435), .A2(n8184), .ZN(n7816) );
  NAND2_X1 U5952 ( .A1(n7534), .A2(n6604), .ZN(n7834) );
  INV_X1 U5953 ( .A(n9982), .ZN(n9991) );
  NAND2_X1 U5954 ( .A1(n6831), .A2(n7290), .ZN(n9987) );
  NAND2_X1 U5955 ( .A1(n9675), .A2(n6573), .ZN(n7322) );
  OAI21_X2 U5956 ( .B1(n6017), .B2(n7009), .A(n5991), .ZN(n7320) );
  INV_X1 U5957 ( .A(n4550), .ZN(n9750) );
  NAND2_X2 U5958 ( .A1(n7290), .A2(n6860), .ZN(n10003) );
  OAI21_X1 U5959 ( .B1(n5750), .B2(n5749), .A(n5748), .ZN(n5753) );
  NAND2_X1 U5960 ( .A1(n5577), .A2(n5576), .ZN(n8398) );
  OR2_X1 U5961 ( .A1(n5742), .A2(n5575), .ZN(n5576) );
  NAND2_X1 U5962 ( .A1(n4531), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4530) );
  OAI21_X1 U5963 ( .B1(n6137), .B2(n6020), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n4532) );
  INV_X1 U5964 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9865) );
  INV_X1 U5965 ( .A(n6153), .ZN(n5974) );
  INV_X1 U5966 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7853) );
  CLKBUF_X1 U5967 ( .A(n6171), .Z(n7855) );
  INV_X1 U5968 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7829) );
  INV_X1 U5969 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6159) );
  INV_X1 U5970 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7760) );
  INV_X1 U5971 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7646) );
  NAND2_X1 U5972 ( .A1(n4607), .A2(n4610), .ZN(n5473) );
  NAND2_X1 U5973 ( .A1(n5435), .A2(n4613), .ZN(n4607) );
  INV_X1 U5974 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7640) );
  INV_X1 U5975 ( .A(n8247), .ZN(n8286) );
  INV_X1 U5976 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7603) );
  AND2_X1 U5977 ( .A1(n6087), .A2(n6086), .ZN(n9948) );
  XNOR2_X1 U5978 ( .A(n6060), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9501) );
  INV_X1 U5979 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U5980 ( .A1(n5071), .A2(n4624), .ZN(n4461) );
  XNOR2_X1 U5981 ( .A(n4501), .B(n5998), .ZN(n7871) );
  NAND2_X1 U5982 ( .A1(n4502), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4501) );
  NAND2_X1 U5983 ( .A1(n6005), .A2(n5997), .ZN(n4502) );
  XNOR2_X1 U5984 ( .A(n6005), .B(n5997), .ZN(n7080) );
  XNOR2_X1 U5985 ( .A(n5977), .B(n5976), .ZN(n7007) );
  NOR2_X1 U5986 ( .A1(n9892), .A2(n9891), .ZN(n10300) );
  NOR2_X1 U5987 ( .A1(n9898), .A2(n9897), .ZN(n10151) );
  NOR2_X1 U5988 ( .A1(n10153), .A2(n10152), .ZN(n9897) );
  NOR2_X1 U5989 ( .A1(n9903), .A2(n9902), .ZN(n10147) );
  NOR2_X1 U5990 ( .A1(n10149), .A2(n10148), .ZN(n9902) );
  NOR2_X1 U5991 ( .A1(n9908), .A2(n9907), .ZN(n10143) );
  NAND2_X1 U5992 ( .A1(n4434), .A2(n8557), .ZN(n6306) );
  NAND2_X1 U5993 ( .A1(n6922), .A2(n4551), .ZN(n6930) );
  NAND2_X1 U5994 ( .A1(n6690), .A2(n4575), .ZN(n7439) );
  AOI21_X1 U5995 ( .B1(n8745), .B2(n4338), .A(n4704), .ZN(n4571) );
  NAND2_X1 U5996 ( .A1(n8749), .A2(n8750), .ZN(n4705) );
  OAI21_X1 U5997 ( .B1(n8739), .B2(n8738), .A(n10114), .ZN(n4572) );
  NAND2_X1 U5998 ( .A1(n6762), .A2(n6751), .ZN(n4767) );
  NAND2_X1 U5999 ( .A1(n4772), .A2(n4771), .ZN(n4770) );
  OR2_X1 U6000 ( .A1(n6763), .A2(n9073), .ZN(n6766) );
  OAI22_X1 U6001 ( .A1(n8762), .A2(n9065), .B1(n10259), .B2(n4313), .ZN(n6764)
         );
  NOR2_X1 U6002 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  AOI21_X1 U6003 ( .B1(n8410), .B2(n9167), .A(n5961), .ZN(n5962) );
  NOR2_X1 U6004 ( .A1(n5734), .A2(n5960), .ZN(n5961) );
  AND2_X1 U6005 ( .A1(n8108), .A2(n4417), .ZN(n4443) );
  OR2_X1 U6006 ( .A1(n8377), .A2(n8376), .ZN(n4437) );
  INV_X1 U6007 ( .A(n4528), .ZN(P1_U3555) );
  AOI21_X1 U6008 ( .B1(n9403), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n4529), .ZN(
        n4528) );
  NOR2_X1 U6009 ( .A1(n9403), .A2(n7278), .ZN(n4529) );
  NAND2_X1 U6010 ( .A1(n7421), .A2(n4498), .ZN(n7425) );
  AOI21_X1 U6011 ( .B1(n9552), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9551), .ZN(
        n4739) );
  NAND2_X1 U6012 ( .A1(n4738), .A2(n9550), .ZN(n4737) );
  NAND2_X1 U6013 ( .A1(n4482), .A2(n6772), .ZN(n4481) );
  NAND2_X1 U6014 ( .A1(n4549), .A2(n4546), .ZN(P1_U3266) );
  NAND2_X1 U6015 ( .A1(n4550), .A2(n9989), .ZN(n4549) );
  INV_X1 U6016 ( .A(n4547), .ZN(n4546) );
  OAI21_X1 U6017 ( .B1(n9751), .B2(n9736), .A(n4548), .ZN(n4547) );
  OAI21_X1 U6018 ( .B1(n9572), .B2(n4927), .A(n10055), .ZN(n6633) );
  AND2_X1 U6019 ( .A1(n5905), .A2(n8812), .ZN(n4320) );
  INV_X1 U6020 ( .A(n6573), .ZN(n7278) );
  INV_X1 U6021 ( .A(n7094), .ZN(n4463) );
  OAI22_X2 U6022 ( .A1(n9704), .A2(n6612), .B1(n9389), .B2(n9794), .ZN(n9690)
         );
  NOR2_X1 U6023 ( .A1(n5307), .A2(n5306), .ZN(n4321) );
  AND2_X1 U6024 ( .A1(n5356), .A2(n5381), .ZN(n4322) );
  AND2_X1 U6025 ( .A1(n5839), .A2(n5822), .ZN(n4323) );
  OR2_X1 U6026 ( .A1(n6253), .A2(n8507), .ZN(n4324) );
  AND3_X1 U6027 ( .A1(n6071), .A2(n5967), .A3(n4356), .ZN(n6134) );
  NOR2_X1 U6028 ( .A1(n5903), .A2(n4645), .ZN(n4644) );
  INV_X1 U6029 ( .A(n4644), .ZN(n4640) );
  AND4_X1 U6030 ( .A1(n4619), .A2(n4618), .A3(n4617), .A4(n4616), .ZN(n4325)
         );
  AND2_X1 U6031 ( .A1(n4367), .A2(n8200), .ZN(n4326) );
  AND2_X1 U6032 ( .A1(n4761), .A2(n4760), .ZN(n4327) );
  OAI211_X1 U6033 ( .C1(n9954), .C2(n4509), .A(n4505), .B(n4504), .ZN(n9547)
         );
  AND2_X1 U6034 ( .A1(n8972), .A2(n4373), .ZN(n4328) );
  AND2_X1 U6035 ( .A1(n9778), .A2(n9676), .ZN(n4329) );
  OR2_X1 U6036 ( .A1(n7842), .A2(n7818), .ZN(n4330) );
  OR2_X1 U6037 ( .A1(n9107), .A2(n8528), .ZN(n8812) );
  OR2_X1 U6038 ( .A1(n7153), .A2(n7170), .ZN(n4331) );
  AND2_X1 U6039 ( .A1(n4651), .A2(n5944), .ZN(n4332) );
  AND2_X1 U6040 ( .A1(n4808), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4333) );
  AND2_X1 U6041 ( .A1(n5265), .A2(n4675), .ZN(n4334) );
  NAND2_X1 U6042 ( .A1(n7927), .A2(n7926), .ZN(n4335) );
  AND2_X1 U6043 ( .A1(n8677), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4336) );
  NOR2_X1 U6044 ( .A1(n6727), .A2(n8648), .ZN(n4337) );
  AND2_X1 U6045 ( .A1(n6751), .A2(n8744), .ZN(n4338) );
  AND2_X1 U6046 ( .A1(n9953), .A2(n4510), .ZN(n4339) );
  NAND2_X1 U6047 ( .A1(n4774), .A2(n6744), .ZN(n4340) );
  NAND2_X1 U6048 ( .A1(n4792), .A2(n4790), .ZN(n6643) );
  NAND2_X1 U6049 ( .A1(n4877), .A2(n5623), .ZN(n8908) );
  AND2_X1 U6050 ( .A1(n4333), .A2(n4809), .ZN(n7805) );
  NOR2_X1 U6051 ( .A1(n8484), .A2(n8485), .ZN(n4343) );
  AND2_X1 U6052 ( .A1(n9295), .A2(n7782), .ZN(n4344) );
  NAND2_X1 U6053 ( .A1(n5357), .A2(n5356), .ZN(n4345) );
  XNOR2_X1 U6054 ( .A(n4553), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6708) );
  INV_X1 U6055 ( .A(n6708), .ZN(n4790) );
  OR2_X1 U6056 ( .A1(n9148), .A2(n8487), .ZN(n5624) );
  AND2_X1 U6057 ( .A1(n4845), .A2(n8001), .ZN(n4346) );
  NAND2_X1 U6058 ( .A1(n7906), .A2(n7915), .ZN(n4347) );
  OR2_X1 U6059 ( .A1(n5060), .A2(n6843), .ZN(n4348) );
  NOR2_X1 U6060 ( .A1(n9789), .A2(n9674), .ZN(n4349) );
  AND2_X1 U6061 ( .A1(n5175), .A2(n5174), .ZN(n5357) );
  NAND2_X1 U6062 ( .A1(n5182), .A2(n4683), .ZN(n4350) );
  NAND2_X1 U6063 ( .A1(n4900), .A2(n4904), .ZN(n8451) );
  INV_X1 U6064 ( .A(n4611), .ZN(n4610) );
  NAND2_X1 U6065 ( .A1(n4612), .A2(n5455), .ZN(n4611) );
  AND2_X1 U6066 ( .A1(n5181), .A2(n4685), .ZN(n4351) );
  NAND2_X1 U6067 ( .A1(n4523), .A2(n8189), .ZN(n9729) );
  NAND2_X1 U6068 ( .A1(n4863), .A2(n5629), .ZN(n8877) );
  NAND2_X1 U6069 ( .A1(n7861), .A2(n6608), .ZN(n9722) );
  NAND4_X1 U6070 ( .A1(n6379), .A2(n6378), .A3(n6377), .A4(n6376), .ZN(n6380)
         );
  NAND2_X1 U6071 ( .A1(n6028), .A2(n4630), .ZN(n10029) );
  AND4_X1 U6072 ( .A1(n8124), .A2(n8139), .A3(n6589), .A4(n4312), .ZN(n4352)
         );
  AND4_X1 U6073 ( .A1(n6575), .A2(n6577), .A3(n6576), .A4(n6578), .ZN(n4353)
         );
  AND2_X1 U6074 ( .A1(n5854), .A2(n8972), .ZN(n4354) );
  OR2_X1 U6075 ( .A1(n9068), .A2(n8605), .ZN(n4355) );
  NOR2_X1 U6076 ( .A1(n5969), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4356) );
  OR2_X2 U6077 ( .A1(n8538), .A2(n8970), .ZN(n6223) );
  INV_X1 U6078 ( .A(n6223), .ZN(n4787) );
  OR2_X1 U6079 ( .A1(n9499), .A2(n9505), .ZN(n4357) );
  NOR3_X1 U6080 ( .A1(n8209), .A2(n8281), .A3(n4312), .ZN(n4358) );
  NAND2_X1 U6081 ( .A1(n9302), .A2(n8000), .ZN(n4359) );
  AND2_X1 U6082 ( .A1(n8234), .A2(n8348), .ZN(n8335) );
  AND3_X1 U6083 ( .A1(n6148), .A2(n6147), .A3(n6166), .ZN(n4360) );
  NAND2_X1 U6084 ( .A1(n8226), .A2(n8329), .ZN(n9564) );
  NOR2_X1 U6085 ( .A1(n8794), .A2(n4987), .ZN(n4361) );
  NOR2_X1 U6086 ( .A1(n8485), .A2(n6244), .ZN(n4362) );
  AND2_X1 U6087 ( .A1(n4597), .A2(n4595), .ZN(n4363) );
  OR2_X1 U6088 ( .A1(n9778), .A2(n9676), .ZN(n4364) );
  AND2_X1 U6089 ( .A1(n6221), .A2(n8602), .ZN(n4365) );
  OR2_X1 U6090 ( .A1(n9803), .A2(n9376), .ZN(n8189) );
  AND2_X1 U6091 ( .A1(n6522), .A2(n8280), .ZN(n4366) );
  AND2_X1 U6092 ( .A1(n8195), .A2(n8310), .ZN(n4367) );
  OR2_X1 U6093 ( .A1(n9569), .A2(n10020), .ZN(n4368) );
  AND2_X1 U6094 ( .A1(n6213), .A2(n6215), .ZN(n4369) );
  AND2_X1 U6095 ( .A1(n5632), .A2(n5631), .ZN(n4370) );
  OR2_X1 U6096 ( .A1(n8233), .A2(n9740), .ZN(n4371) );
  AND2_X1 U6097 ( .A1(n5901), .A2(n5905), .ZN(n4372) );
  OR2_X1 U6098 ( .A1(n5850), .A2(n4787), .ZN(n4373) );
  NAND2_X1 U6099 ( .A1(n9250), .A2(n7958), .ZN(n4374) );
  NAND2_X1 U6100 ( .A1(n8504), .A2(n6251), .ZN(n4375) );
  AND2_X1 U6101 ( .A1(n6443), .A2(n8184), .ZN(n4376) );
  AND2_X1 U6102 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n4377) );
  INV_X1 U6103 ( .A(n4833), .ZN(n4832) );
  NAND2_X1 U6104 ( .A1(n7782), .A2(n4347), .ZN(n4833) );
  AND2_X1 U6105 ( .A1(n6522), .A2(n8271), .ZN(n4378) );
  INV_X1 U6106 ( .A(n4951), .ZN(n4950) );
  OR2_X1 U6107 ( .A1(n6614), .A2(n4952), .ZN(n4951) );
  AND2_X1 U6108 ( .A1(n6010), .A2(n4462), .ZN(n4379) );
  OR2_X1 U6109 ( .A1(n9130), .A2(n8510), .ZN(n5889) );
  INV_X1 U6110 ( .A(n5895), .ZN(n4646) );
  OR2_X1 U6111 ( .A1(n5898), .A2(n8836), .ZN(n4380) );
  OR2_X1 U6112 ( .A1(n8607), .A2(n7116), .ZN(n5821) );
  INV_X1 U6113 ( .A(n5821), .ZN(n4782) );
  INV_X1 U6114 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5672) );
  INV_X1 U6115 ( .A(n4500), .ZN(n4497) );
  NAND2_X1 U6116 ( .A1(n7248), .A2(n6996), .ZN(n4500) );
  INV_X1 U6117 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6326) );
  AND2_X1 U6118 ( .A1(n8206), .A2(n8205), .ZN(n4381) );
  INV_X1 U6119 ( .A(n4499), .ZN(n4498) );
  NOR2_X1 U6120 ( .A1(n7422), .A2(n7423), .ZN(n4499) );
  INV_X1 U6121 ( .A(n4765), .ZN(n4763) );
  NAND2_X1 U6122 ( .A1(n7758), .A2(n7483), .ZN(n4765) );
  AND2_X1 U6123 ( .A1(n5279), .A2(SI_13_), .ZN(n4382) );
  OR2_X1 U6124 ( .A1(n8177), .A2(n8238), .ZN(n4383) );
  INV_X1 U6125 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6079) );
  INV_X1 U6126 ( .A(n4960), .ZN(n4959) );
  OAI21_X1 U6127 ( .B1(n6623), .B2(n4961), .A(n6622), .ZN(n4960) );
  NAND2_X1 U6128 ( .A1(n8550), .A2(n8549), .ZN(n4384) );
  AND2_X1 U6129 ( .A1(n4636), .A2(n4643), .ZN(n4385) );
  NAND2_X1 U6130 ( .A1(n7962), .A2(n7961), .ZN(n9254) );
  AND2_X1 U6131 ( .A1(n8225), .A2(n8115), .ZN(n9583) );
  INV_X1 U6132 ( .A(n9583), .ZN(n4918) );
  AND2_X1 U6133 ( .A1(n4436), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4386) );
  AND2_X1 U6134 ( .A1(n6256), .A2(n6255), .ZN(n4387) );
  INV_X1 U6135 ( .A(n5870), .ZN(n4800) );
  NAND2_X1 U6136 ( .A1(n8024), .A2(n9275), .ZN(n4388) );
  INV_X1 U6137 ( .A(n4945), .ZN(n4944) );
  NAND2_X1 U6138 ( .A1(n4947), .A2(n4364), .ZN(n4945) );
  AND2_X1 U6139 ( .A1(n8324), .A2(n8219), .ZN(n8272) );
  INV_X1 U6140 ( .A(n4614), .ZN(n4613) );
  NAND2_X1 U6141 ( .A1(n5416), .A2(n4615), .ZN(n4614) );
  NAND2_X1 U6142 ( .A1(n5308), .A2(SI_15_), .ZN(n4389) );
  NAND2_X1 U6143 ( .A1(n8237), .A2(n8235), .ZN(n8239) );
  INV_X1 U6144 ( .A(n4957), .ZN(n4956) );
  NOR2_X1 U6145 ( .A1(n4962), .A2(n6619), .ZN(n4957) );
  OR2_X1 U6146 ( .A1(n9102), .A2(n8427), .ZN(n5905) );
  AND2_X1 U6147 ( .A1(n8708), .A2(n8707), .ZN(n4390) );
  INV_X1 U6148 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U6149 ( .A1(n4815), .A2(n5492), .ZN(n8792) );
  NAND2_X1 U6150 ( .A1(n8157), .A2(n8170), .ZN(n8245) );
  AND2_X1 U6151 ( .A1(n8906), .A2(n5866), .ZN(n4391) );
  AND2_X1 U6152 ( .A1(n5909), .A2(n5910), .ZN(n8798) );
  AND2_X1 U6153 ( .A1(n8216), .A2(n9631), .ZN(n4392) );
  AND2_X1 U6154 ( .A1(n8314), .A2(n6495), .ZN(n4393) );
  AND2_X1 U6155 ( .A1(n4802), .A2(n5624), .ZN(n4394) );
  AND2_X1 U6156 ( .A1(n5492), .A2(n5910), .ZN(n4395) );
  AND2_X1 U6157 ( .A1(n4855), .A2(n4360), .ZN(n4396) );
  INV_X1 U6158 ( .A(n8156), .ZN(n4513) );
  NAND2_X1 U6159 ( .A1(n7204), .A2(n8606), .ZN(n4397) );
  INV_X1 U6160 ( .A(n6608), .ZN(n4941) );
  AND2_X1 U6161 ( .A1(n4720), .A2(n4721), .ZN(n4398) );
  AND2_X1 U6162 ( .A1(n6237), .A2(n6236), .ZN(n4399) );
  AND2_X1 U6163 ( .A1(n4992), .A2(n4666), .ZN(n4400) );
  INV_X1 U6164 ( .A(n5942), .ZN(n4653) );
  NOR2_X1 U6165 ( .A1(n9769), .A2(n9387), .ZN(n4401) );
  AND2_X1 U6166 ( .A1(n4752), .A2(n4750), .ZN(n4402) );
  AND2_X1 U6167 ( .A1(n8339), .A2(n8340), .ZN(n4403) );
  AND2_X1 U6168 ( .A1(n5863), .A2(n5862), .ZN(n4404) );
  INV_X1 U6169 ( .A(n8009), .ZN(n4845) );
  AND2_X1 U6170 ( .A1(n4972), .A2(n4977), .ZN(n4405) );
  INV_X1 U6171 ( .A(n4690), .ZN(n4689) );
  NAND2_X1 U6172 ( .A1(n4695), .A2(n4691), .ZN(n4690) );
  OR2_X1 U6173 ( .A1(n8858), .A2(n4873), .ZN(n4406) );
  INV_X1 U6174 ( .A(n4910), .ZN(n4909) );
  NAND2_X1 U6175 ( .A1(n4911), .A2(n6220), .ZN(n4910) );
  INV_X1 U6176 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4531) );
  NAND2_X2 U6177 ( .A1(n7296), .A2(n9987), .ZN(n9989) );
  OR2_X1 U6178 ( .A1(n6722), .A2(n7465), .ZN(n4407) );
  OR2_X1 U6179 ( .A1(n6650), .A2(n6721), .ZN(n7447) );
  NAND2_X1 U6180 ( .A1(n5671), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U6181 ( .A1(n6114), .A2(n6113), .ZN(n9759) );
  INV_X1 U6182 ( .A(n9759), .ZN(n4760) );
  INV_X1 U6183 ( .A(n9970), .ZN(n4764) );
  NAND2_X1 U6184 ( .A1(n4942), .A2(n6451), .ZN(n7861) );
  NAND2_X1 U6185 ( .A1(n8375), .A2(n9550), .ZN(n6770) );
  AND2_X1 U6186 ( .A1(n10062), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4408) );
  INV_X1 U6187 ( .A(n7546), .ZN(n4929) );
  OR2_X1 U6188 ( .A1(n9096), .A2(n8596), .ZN(n4409) );
  AOI21_X1 U6189 ( .B1(n7446), .B2(n7447), .A(n7448), .ZN(n7445) );
  INV_X1 U6190 ( .A(n7445), .ZN(n4568) );
  NAND2_X1 U6191 ( .A1(n5275), .A2(n5274), .ZN(n8920) );
  INV_X1 U6192 ( .A(n8676), .ZN(n4891) );
  OR2_X1 U6193 ( .A1(n8665), .A2(n6731), .ZN(n4410) );
  NAND2_X1 U6194 ( .A1(n5222), .A2(n5221), .ZN(n7708) );
  AND2_X1 U6195 ( .A1(n8137), .A2(n8138), .ZN(n4411) );
  OR2_X1 U6196 ( .A1(n8686), .A2(n6733), .ZN(n4412) );
  AND2_X1 U6197 ( .A1(n4724), .A2(n4725), .ZN(n4413) );
  AND2_X1 U6198 ( .A1(n7692), .A2(n4909), .ZN(n4414) );
  INV_X1 U6199 ( .A(n4694), .ZN(n4693) );
  NAND2_X1 U6200 ( .A1(n4407), .A2(n4700), .ZN(n4694) );
  OR2_X1 U6201 ( .A1(n7004), .A2(n7551), .ZN(n4415) );
  INV_X1 U6202 ( .A(n7416), .ZN(n4725) );
  NOR2_X1 U6203 ( .A1(n6728), .A2(n6653), .ZN(n4416) );
  INV_X1 U6204 ( .A(n6651), .ZN(n4567) );
  AND2_X1 U6205 ( .A1(n7444), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6651) );
  INV_X1 U6206 ( .A(n8410), .ZN(n8762) );
  NAND2_X1 U6207 ( .A1(n5557), .A2(n5556), .ZN(n8410) );
  AND2_X1 U6208 ( .A1(n5633), .A2(n8852), .ZN(n8868) );
  INV_X1 U6209 ( .A(n8868), .ZN(n4875) );
  INV_X1 U6210 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6436) );
  AND2_X1 U6211 ( .A1(n8567), .A2(n6266), .ZN(n6268) );
  OR2_X1 U6212 ( .A1(n8109), .A2(n9366), .ZN(n4417) );
  AND2_X1 U6213 ( .A1(n4688), .A2(n4686), .ZN(n4418) );
  NOR2_X1 U6214 ( .A1(n8678), .A2(n6730), .ZN(n4419) );
  AND2_X1 U6215 ( .A1(n4728), .A2(n4726), .ZN(n4420) );
  OR2_X1 U6216 ( .A1(n6736), .A2(n8916), .ZN(n4421) );
  AND2_X1 U6217 ( .A1(n7447), .A2(n4819), .ZN(n4422) );
  INV_X1 U6218 ( .A(n4828), .ZN(n9232) );
  AND2_X1 U6219 ( .A1(n4334), .A2(n10221), .ZN(n4423) );
  INV_X1 U6220 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10154) );
  OR2_X1 U6221 ( .A1(n4807), .A2(n4806), .ZN(n4566) );
  NAND2_X1 U6222 ( .A1(n7444), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4424) );
  INV_X1 U6223 ( .A(n7033), .ZN(n4894) );
  INV_X1 U6224 ( .A(n5779), .ZN(n7037) );
  INV_X1 U6225 ( .A(n9934), .ZN(n9951) );
  INV_X1 U6226 ( .A(n9312), .ZN(n9380) );
  NOR2_X2 U6227 ( .A1(n6830), .A2(n6816), .ZN(n9312) );
  NAND2_X1 U6228 ( .A1(n8147), .A2(n7546), .ZN(n8135) );
  INV_X1 U6229 ( .A(n8135), .ZN(n4618) );
  NOR2_X1 U6230 ( .A1(n6122), .A2(n9856), .ZN(n4426) );
  OAI21_X1 U6231 ( .B1(n8748), .B2(n8747), .A(n8746), .ZN(n4704) );
  AND2_X1 U6232 ( .A1(n4716), .A2(n4719), .ZN(n4427) );
  AND2_X1 U6233 ( .A1(n4507), .A2(n4510), .ZN(n4428) );
  INV_X1 U6234 ( .A(n4509), .ZN(n4508) );
  NAND2_X1 U6235 ( .A1(n9537), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n4509) );
  AND2_X1 U6236 ( .A1(n4680), .A2(n4679), .ZN(n4429) );
  OR2_X1 U6237 ( .A1(n6872), .A2(P1_U3086), .ZN(n8378) );
  INV_X1 U6238 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4510) );
  INV_X1 U6239 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4594) );
  OAI21_X1 U6240 ( .B1(n4465), .B2(n5951), .A(n5950), .ZN(P2_U3296) );
  NAND2_X1 U6241 ( .A1(n5876), .A2(n4391), .ZN(n5868) );
  NAND2_X1 U6242 ( .A1(n4743), .A2(n4741), .ZN(n5914) );
  AOI22_X1 U6243 ( .A1(n5873), .A2(n5872), .B1(n5925), .B2(n5871), .ZN(n5885)
         );
  NAND2_X1 U6244 ( .A1(n4648), .A2(n5865), .ZN(n4647) );
  NAND2_X2 U6245 ( .A1(n8384), .A2(n5015), .ZN(n5585) );
  OAI21_X1 U6246 ( .B1(n4657), .B2(n4655), .A(n5852), .ZN(n4654) );
  NAND4_X1 U6247 ( .A1(n4810), .A2(n4430), .A3(n4813), .A4(n4814), .ZN(n5012)
         );
  NAND2_X1 U6248 ( .A1(n5212), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5019) );
  CLKBUF_X1 U6249 ( .A(n6667), .Z(n4431) );
  NAND2_X1 U6250 ( .A1(n7383), .A2(n5848), .ZN(n5164) );
  OAI21_X2 U6251 ( .B1(n5066), .B2(n4783), .A(n4780), .ZN(n7150) );
  NAND2_X1 U6252 ( .A1(n8975), .A2(n5856), .ZN(n8959) );
  NAND2_X1 U6253 ( .A1(n5394), .A2(n5889), .ZN(n8832) );
  OAI21_X2 U6254 ( .B1(n8781), .B2(n5915), .A(n5916), .ZN(n8769) );
  OAI21_X1 U6255 ( .B1(n5772), .B2(n5796), .A(n5771), .ZN(n5774) );
  NOR2_X1 U6256 ( .A1(n8422), .A2(n8846), .ZN(n8423) );
  NAND2_X1 U6257 ( .A1(n7143), .A2(n7142), .ZN(n7141) );
  INV_X1 U6258 ( .A(n6667), .ZN(n4432) );
  OAI21_X1 U6259 ( .B1(n6312), .B2(n4435), .A(n8571), .ZN(n4434) );
  NAND2_X4 U6260 ( .A1(n6754), .A2(n5656), .ZN(n6636) );
  INV_X1 U6261 ( .A(n4556), .ZN(n6655) );
  INV_X1 U6262 ( .A(n6659), .ZN(n6660) );
  NAND2_X1 U6263 ( .A1(n4795), .A2(n4797), .ZN(n4558) );
  NAND2_X1 U6264 ( .A1(n8739), .A2(n4769), .ZN(n4582) );
  NOR2_X1 U6265 ( .A1(n10088), .A2(n6647), .ZN(n6648) );
  AOI21_X1 U6266 ( .B1(n4583), .B2(n10095), .A(n4581), .ZN(n4768) );
  AOI21_X1 U6267 ( .B1(n7181), .B2(n7182), .A(n7183), .ZN(n7180) );
  NAND2_X2 U6268 ( .A1(n6636), .A2(n6837), .ZN(n5060) );
  NAND2_X1 U6269 ( .A1(n8522), .A2(n8523), .ZN(n6260) );
  NAND2_X1 U6270 ( .A1(n8416), .A2(n8415), .ZN(n4906) );
  OAI21_X1 U6271 ( .B1(n6217), .B2(n4910), .A(n4908), .ZN(n8431) );
  OAI21_X1 U6272 ( .B1(n6313), .B2(n6312), .A(n8557), .ZN(n6320) );
  NAND2_X1 U6273 ( .A1(n8550), .A2(n6247), .ZN(n8442) );
  AOI21_X1 U6274 ( .B1(n7308), .B2(n7307), .A(n7306), .ZN(n7310) );
  NAND2_X1 U6275 ( .A1(n5021), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U6276 ( .A1(n7232), .A2(n7231), .ZN(n7308) );
  NAND2_X1 U6277 ( .A1(n8584), .A2(n6239), .ZN(n8478) );
  NOR2_X1 U6278 ( .A1(n7225), .A2(n7226), .ZN(n7224) );
  NAND2_X1 U6279 ( .A1(n6232), .A2(n8464), .ZN(n8514) );
  NAND2_X1 U6280 ( .A1(n4438), .A2(n4437), .ZN(P1_U3242) );
  OAI21_X1 U6281 ( .B1(n8371), .B2(n4472), .A(n6824), .ZN(n4438) );
  NAND2_X1 U6282 ( .A1(n8341), .A2(n4403), .ZN(n8368) );
  NAND2_X1 U6283 ( .A1(n8236), .A2(n8239), .ZN(n8341) );
  MUX2_X1 U6284 ( .A(n8175), .B(n8174), .S(n8238), .Z(n8188) );
  AOI21_X1 U6285 ( .B1(n4441), .B2(n8155), .A(n8154), .ZN(n8168) );
  NAND2_X1 U6286 ( .A1(n4518), .A2(n4517), .ZN(n4516) );
  NAND2_X1 U6287 ( .A1(n4628), .A2(n4392), .ZN(n4627) );
  NAND2_X1 U6288 ( .A1(n8136), .A2(n9967), .ZN(n4616) );
  OAI21_X1 U6289 ( .B1(n8212), .B2(n8207), .A(n8243), .ZN(n4629) );
  AND2_X1 U6290 ( .A1(n7579), .A2(n5615), .ZN(n5613) );
  AOI21_X2 U6291 ( .B1(n7580), .B2(n5618), .A(n4969), .ZN(n8965) );
  NAND2_X1 U6292 ( .A1(n8844), .A2(n5635), .ZN(n8824) );
  AOI21_X1 U6293 ( .B1(n5954), .B2(n5651), .A(n5650), .ZN(n5668) );
  NAND2_X1 U6294 ( .A1(n5626), .A2(n5625), .ZN(n8898) );
  OAI21_X2 U6295 ( .B1(n8832), .B2(n5454), .A(n5453), .ZN(n8839) );
  NAND2_X1 U6296 ( .A1(n7578), .A2(n5841), .ZN(n7677) );
  INV_X2 U6298 ( .A(n8050), .ZN(n8063) );
  NAND2_X4 U6299 ( .A1(n6775), .A2(n7616), .ZN(n8050) );
  NAND2_X1 U6300 ( .A1(n7266), .A2(n7265), .ZN(n7267) );
  XNOR2_X1 U6301 ( .A(n6796), .B(n6795), .ZN(n7265) );
  NAND2_X1 U6302 ( .A1(n4444), .A2(n4443), .ZN(P1_U3214) );
  NAND2_X1 U6303 ( .A1(n6954), .A2(n4445), .ZN(n5053) );
  NAND2_X1 U6304 ( .A1(n5568), .A2(n5928), .ZN(n5757) );
  NAND4_X1 U6305 ( .A1(n4810), .A2(n4813), .A3(n4814), .A4(n5175), .ZN(n5021)
         );
  NAND2_X1 U6306 ( .A1(n4784), .A2(n4328), .ZN(n8975) );
  AND2_X1 U6307 ( .A1(n5613), .A2(n6222), .ZN(n5618) );
  NAND2_X1 U6308 ( .A1(n9607), .A2(n6513), .ZN(n4924) );
  NAND2_X1 U6309 ( .A1(n8258), .A2(n6352), .ZN(n8294) );
  AND4_X2 U6310 ( .A1(n6071), .A2(n5967), .A3(n4356), .A4(n6133), .ZN(n6137)
         );
  NAND2_X1 U6311 ( .A1(n5638), .A2(n4870), .ZN(n8783) );
  OAI21_X1 U6312 ( .B1(n8149), .B2(n8152), .A(n8156), .ZN(n6401) );
  OAI21_X2 U6313 ( .B1(n7055), .B2(n8123), .A(n8290), .ZN(n8141) );
  XNOR2_X1 U6314 ( .A(n6698), .B(n6745), .ZN(n4583) );
  XNOR2_X1 U6315 ( .A(n8734), .B(n8733), .ZN(n4570) );
  NAND3_X1 U6316 ( .A1(n6587), .A2(n6586), .A3(n7287), .ZN(n4459) );
  OR2_X1 U6317 ( .A1(n8359), .A2(n8358), .ZN(n8360) );
  NAND2_X1 U6318 ( .A1(n9565), .A2(n4757), .ZN(n4927) );
  NAND2_X1 U6319 ( .A1(n6631), .A2(n6630), .ZN(n4928) );
  INV_X1 U6320 ( .A(n4953), .ZN(n9575) );
  NAND2_X1 U6321 ( .A1(n5038), .A2(n5779), .ZN(n7040) );
  OAI21_X1 U6322 ( .B1(n8769), .B2(n8768), .A(n5547), .ZN(n5952) );
  NAND2_X1 U6323 ( .A1(n4801), .A2(n4798), .ZN(n8895) );
  NAND2_X1 U6324 ( .A1(n7150), .A2(n5839), .ZN(n5147) );
  NAND3_X1 U6325 ( .A1(n4543), .A2(n4381), .A3(n4455), .ZN(n8214) );
  AOI21_X1 U6326 ( .B1(n4471), .B2(n4470), .A(n4468), .ZN(n8230) );
  OAI21_X1 U6327 ( .B1(n4633), .B2(n4632), .A(n8193), .ZN(n8203) );
  NAND2_X1 U6328 ( .A1(n9357), .A2(n8045), .ZN(n9354) );
  NAND2_X1 U6329 ( .A1(n4836), .A2(n4834), .ZN(n9279) );
  NAND2_X1 U6330 ( .A1(n9188), .A2(n7947), .ZN(n9248) );
  NAND2_X1 U6331 ( .A1(n4458), .A2(n4371), .ZN(n8236) );
  OAI22_X1 U6332 ( .A1(n8230), .A2(n8231), .B1(n8229), .B2(n8232), .ZN(n4458)
         );
  NAND3_X1 U6333 ( .A1(n8368), .A2(n4990), .A3(n4473), .ZN(n4472) );
  AOI21_X1 U6334 ( .B1(n4516), .B2(n4515), .A(n4312), .ZN(n4633) );
  NOR2_X1 U6335 ( .A1(n8128), .A2(n8238), .ZN(n8130) );
  INV_X1 U6336 ( .A(n8134), .ZN(n4617) );
  NAND2_X1 U6337 ( .A1(n8224), .A2(n8223), .ZN(n4471) );
  NAND2_X1 U6338 ( .A1(n4519), .A2(n8189), .ZN(n4518) );
  OAI211_X1 U6339 ( .C1(n8197), .C2(n8311), .A(n8196), .B(n8310), .ZN(n4544)
         );
  NAND2_X1 U6340 ( .A1(n4544), .A2(n4312), .ZN(n4543) );
  OAI211_X2 U6341 ( .C1(n5632), .C2(n4872), .A(n4871), .B(n8836), .ZN(n8844)
         );
  NAND2_X1 U6342 ( .A1(n8783), .A2(n5641), .ZN(n5643) );
  NAND2_X1 U6343 ( .A1(n4749), .A2(n5202), .ZN(n4746) );
  NAND2_X1 U6344 ( .A1(n4746), .A2(n5225), .ZN(n5242) );
  NAND2_X1 U6345 ( .A1(n4459), .A2(n6588), .ZN(n7487) );
  NAND2_X1 U6346 ( .A1(n4460), .A2(n4940), .ZN(n6611) );
  NAND2_X1 U6347 ( .A1(n7862), .A2(n6608), .ZN(n4460) );
  XNOR2_X1 U6348 ( .A(n4461), .B(n5086), .ZN(n6007) );
  OR2_X2 U6349 ( .A1(n9606), .A2(n6619), .ZN(n4967) );
  XOR2_X2 U6350 ( .A(n8272), .B(n7888), .Z(n9756) );
  NAND2_X1 U6352 ( .A1(n5946), .A2(n4650), .ZN(n4465) );
  NAND2_X1 U6353 ( .A1(n5908), .A2(n5925), .ZN(n4743) );
  OAI21_X1 U6354 ( .B1(n5861), .B2(n4404), .A(n4649), .ZN(n4648) );
  OAI21_X1 U6355 ( .B1(n5845), .B2(n5925), .A(n4656), .ZN(n4655) );
  NAND3_X1 U6356 ( .A1(n5932), .A2(n5931), .A3(n4653), .ZN(n4652) );
  NAND2_X1 U6357 ( .A1(n5611), .A2(n7680), .ZN(n4466) );
  NAND2_X1 U6358 ( .A1(n4511), .A2(n5149), .ZN(n5195) );
  OAI21_X1 U6359 ( .B1(n8965), .B2(n5620), .A(n5619), .ZN(n8948) );
  NAND2_X1 U6360 ( .A1(n5202), .A2(n5201), .ZN(n5226) );
  OAI21_X1 U6361 ( .B1(n8898), .B2(n4862), .A(n4860), .ZN(n4863) );
  OAI21_X1 U6362 ( .B1(n5093), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4467), .ZN(
        n5088) );
  NAND2_X1 U6363 ( .A1(n4631), .A2(n8192), .ZN(n4632) );
  NAND2_X1 U6364 ( .A1(n4915), .A2(n5130), .ZN(n4511) );
  INV_X1 U6365 ( .A(n8204), .ZN(n8206) );
  NOR2_X2 U6366 ( .A1(n6496), .A2(n9204), .ZN(n4479) );
  NAND3_X1 U6367 ( .A1(n4481), .A2(n4737), .A3(n4739), .ZN(P1_U3262) );
  NAND2_X1 U6368 ( .A1(n4492), .A2(n4493), .ZN(n7512) );
  NAND2_X1 U6369 ( .A1(n7247), .A2(n4498), .ZN(n4492) );
  NOR2_X1 U6370 ( .A1(n7247), .A2(n4497), .ZN(n7250) );
  NAND2_X1 U6371 ( .A1(n9954), .A2(n4339), .ZN(n4504) );
  INV_X1 U6372 ( .A(n9547), .ZN(n9549) );
  NAND2_X1 U6373 ( .A1(n9954), .A2(n9953), .ZN(n9952) );
  XNOR2_X1 U6374 ( .A(n4511), .B(n5148), .ZN(n6844) );
  NAND2_X2 U6375 ( .A1(n7893), .A2(n8272), .ZN(n7892) );
  NAND2_X1 U6376 ( .A1(n8148), .A2(n8165), .ZN(n8152) );
  INV_X1 U6377 ( .A(n6401), .ZN(n8258) );
  OAI21_X1 U6378 ( .B1(n8188), .B2(n8297), .A(n8300), .ZN(n4519) );
  NAND2_X1 U6379 ( .A1(n7814), .A2(n4524), .ZN(n4520) );
  NAND2_X1 U6380 ( .A1(n8058), .A2(n6573), .ZN(n6792) );
  NAND2_X1 U6381 ( .A1(n6467), .A2(n4539), .ZN(n4537) );
  NAND2_X1 U6382 ( .A1(n6467), .A2(n4326), .ZN(n4538) );
  NAND3_X1 U6383 ( .A1(n4816), .A2(n10085), .A3(P2_REG2_REG_5__SCAN_IN), .ZN(
        n6922) );
  NAND2_X1 U6384 ( .A1(n4552), .A2(n7202), .ZN(n4551) );
  NAND2_X1 U6385 ( .A1(n7445), .A2(n4566), .ZN(n4562) );
  INV_X1 U6386 ( .A(n6654), .ZN(n4793) );
  NAND4_X1 U6387 ( .A1(n4572), .A2(n4705), .A3(n4571), .A4(n4569), .ZN(
        P2_U3200) );
  OAI21_X1 U6388 ( .B1(n6690), .B2(n4574), .A(n4424), .ZN(n4573) );
  NAND2_X1 U6389 ( .A1(n4893), .A2(n4578), .ZN(n8705) );
  NAND2_X1 U6390 ( .A1(n8659), .A2(n4889), .ZN(n4580) );
  NAND2_X1 U6391 ( .A1(n5513), .A2(n5512), .ZN(n4584) );
  NAND2_X1 U6392 ( .A1(n5494), .A2(n5493), .ZN(n4585) );
  NAND3_X1 U6393 ( .A1(n8239), .A2(n4589), .A3(n4588), .ZN(n4587) );
  NAND2_X1 U6394 ( .A1(n4601), .A2(n4602), .ZN(n5475) );
  NAND2_X1 U6395 ( .A1(n5397), .A2(n4605), .ZN(n4601) );
  NAND3_X1 U6396 ( .A1(n5416), .A2(n5417), .A3(n4615), .ZN(n4612) );
  OAI21_X1 U6397 ( .B1(n8168), .B2(n8167), .A(n8166), .ZN(n8173) );
  OAI211_X1 U6398 ( .C1(n4623), .C2(n5067), .A(n4621), .B(n5086), .ZN(n5122)
         );
  AND2_X1 U6399 ( .A1(n5071), .A2(n5065), .ZN(n4622) );
  NAND2_X1 U6400 ( .A1(n5068), .A2(n5067), .ZN(n4624) );
  NAND2_X1 U6401 ( .A1(n4637), .A2(n4634), .ZN(n4641) );
  NAND3_X1 U6402 ( .A1(n5887), .A2(n5888), .A3(n5886), .ZN(n4637) );
  NAND2_X1 U6403 ( .A1(n4652), .A2(n4651), .ZN(n5945) );
  NAND2_X1 U6404 ( .A1(n4652), .A2(n4332), .ZN(n4650) );
  NOR2_X1 U6405 ( .A1(n5823), .A2(n5837), .ZN(n4661) );
  NAND3_X1 U6406 ( .A1(n4662), .A2(n4660), .A3(n4658), .ZN(n5831) );
  NAND3_X1 U6407 ( .A1(n5835), .A2(n4323), .A3(n7385), .ZN(n4662) );
  NAND2_X1 U6408 ( .A1(n5914), .A2(n4668), .ZN(n4664) );
  NAND2_X1 U6409 ( .A1(n4664), .A2(n4400), .ZN(n4665) );
  INV_X1 U6410 ( .A(n6196), .ZN(n7041) );
  INV_X1 U6411 ( .A(n4859), .ZN(n5810) );
  OAI211_X1 U6412 ( .C1(n6636), .C2(n6838), .A(n5030), .B(n5029), .ZN(n6196)
         );
  NOR2_X2 U6413 ( .A1(n5173), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4814) );
  NAND3_X1 U6414 ( .A1(n5795), .A2(n5953), .A3(n8770), .ZN(n4674) );
  NAND2_X1 U6415 ( .A1(n5266), .A2(n4423), .ZN(n5321) );
  NAND2_X1 U6416 ( .A1(n5337), .A2(n4676), .ZN(n5402) );
  NAND2_X1 U6417 ( .A1(n5503), .A2(n4680), .ZN(n5540) );
  NAND2_X1 U6418 ( .A1(n5503), .A2(n4429), .ZN(n5560) );
  NAND2_X1 U6419 ( .A1(n5503), .A2(n5502), .ZN(n5521) );
  NAND2_X1 U6420 ( .A1(n6724), .A2(n6725), .ZN(n4700) );
  NAND4_X1 U6421 ( .A1(n5356), .A2(n4813), .A3(n5175), .A4(n4814), .ZN(n5681)
         );
  NAND4_X1 U6422 ( .A1(n4977), .A2(n4972), .A3(n4996), .A4(n4997), .ZN(n5682)
         );
  NAND3_X1 U6423 ( .A1(n4711), .A2(n4709), .A3(n4708), .ZN(n4714) );
  NAND2_X1 U6424 ( .A1(n9922), .A2(n9940), .ZN(n4708) );
  NAND3_X1 U6425 ( .A1(n4711), .A2(n4712), .A3(n4708), .ZN(n9933) );
  NOR2_X1 U6426 ( .A1(n9922), .A2(n9498), .ZN(n9499) );
  INV_X1 U6427 ( .A(n4714), .ZN(n9931) );
  NAND2_X1 U6428 ( .A1(n4715), .A2(n4717), .ZN(n9457) );
  NAND2_X1 U6429 ( .A1(n9432), .A2(n4398), .ZN(n4715) );
  NAND2_X1 U6430 ( .A1(n7241), .A2(n4420), .ZN(n4722) );
  NAND2_X1 U6431 ( .A1(n4722), .A2(n4723), .ZN(n7518) );
  OAI21_X1 U6432 ( .B1(n9539), .B2(n4733), .A(n4730), .ZN(n9544) );
  NOR2_X1 U6433 ( .A1(n7076), .A2(n4979), .ZN(n9419) );
  NOR2_X1 U6434 ( .A1(n9457), .A2(n9456), .ZN(n9455) );
  NOR2_X1 U6435 ( .A1(n7086), .A2(n7085), .ZN(n7084) );
  NOR2_X1 U6436 ( .A1(n7518), .A2(n4973), .ZN(n7519) );
  NOR3_X1 U6437 ( .A1(n9405), .A2(n7010), .A3(n7009), .ZN(n9404) );
  NOR2_X1 U6438 ( .A1(n9470), .A2(n9469), .ZN(n9468) );
  NOR2_X1 U6439 ( .A1(n9490), .A2(n9491), .ZN(n9497) );
  NOR2_X1 U6440 ( .A1(n9455), .A2(n4982), .ZN(n9470) );
  AOI21_X1 U6441 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n4463), .A(n7084), .ZN(
        n9432) );
  NAND2_X1 U6442 ( .A1(n7023), .A2(n7022), .ZN(n7241) );
  NOR2_X1 U6443 ( .A1(n9924), .A2(n9923), .ZN(n9922) );
  AOI21_X1 U6444 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n9423), .A(n9417), .ZN(
        n7086) );
  NAND2_X1 U6445 ( .A1(n7519), .A2(n7520), .ZN(n9488) );
  NOR2_X1 U6446 ( .A1(n9419), .A2(n9418), .ZN(n9417) );
  NOR2_X1 U6447 ( .A1(n7078), .A2(n7077), .ZN(n7076) );
  NOR2_X2 U6448 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9868) );
  NAND2_X1 U6449 ( .A1(n4751), .A2(n4402), .ZN(n5326) );
  NAND2_X1 U6450 ( .A1(n5291), .A2(n5290), .ZN(n4755) );
  NAND2_X1 U6451 ( .A1(n9641), .A2(n4759), .ZN(n7876) );
  NAND3_X1 U6452 ( .A1(n4764), .A2(n4763), .A3(n6044), .ZN(n7618) );
  XNOR2_X2 U6453 ( .A(n4766), .B(n5043), .ZN(n6641) );
  INV_X1 U6454 ( .A(n8739), .ZN(n4772) );
  NAND3_X1 U6455 ( .A1(n4770), .A2(n4768), .A3(n4767), .ZN(P2_U3201) );
  INV_X1 U6456 ( .A(n6744), .ZN(n4777) );
  OR2_X1 U6457 ( .A1(n8384), .A2(n4779), .ZN(n5079) );
  AOI21_X1 U6458 ( .B1(n5822), .B2(n4782), .A(n4781), .ZN(n4780) );
  NAND2_X1 U6459 ( .A1(n5222), .A2(n4785), .ZN(n4784) );
  NAND3_X1 U6460 ( .A1(n6643), .A2(P2_REG2_REG_3__SCAN_IN), .A3(n4788), .ZN(
        n10067) );
  NAND2_X1 U6461 ( .A1(n4793), .A2(n6730), .ZN(n4797) );
  NAND2_X1 U6462 ( .A1(n4794), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U6463 ( .A1(n6654), .A2(n4419), .ZN(n4794) );
  NAND2_X1 U6464 ( .A1(n4797), .A2(n8677), .ZN(n8667) );
  NAND2_X1 U6465 ( .A1(n4394), .A2(n5275), .ZN(n4801) );
  AND2_X1 U6466 ( .A1(n5807), .A2(n4859), .ZN(n5779) );
  INV_X1 U6467 ( .A(n5007), .ZN(n4811) );
  NOR2_X2 U6468 ( .A1(n5007), .A2(n5006), .ZN(n5356) );
  NAND2_X1 U6469 ( .A1(n4815), .A2(n4395), .ZN(n5511) );
  NAND2_X1 U6470 ( .A1(n4817), .A2(n6925), .ZN(n4816) );
  INV_X1 U6471 ( .A(n6646), .ZN(n4817) );
  NAND2_X1 U6472 ( .A1(n5164), .A2(n4818), .ZN(n7578) );
  NAND2_X1 U6473 ( .A1(n8694), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8693) );
  NAND3_X1 U6474 ( .A1(n7447), .A2(n4819), .A3(P2_REG2_REG_9__SCAN_IN), .ZN(
        n7446) );
  NAND2_X1 U6475 ( .A1(n6650), .A2(n6721), .ZN(n4819) );
  NOR2_X2 U6476 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6003) );
  AND3_X2 U6477 ( .A1(n6018), .A2(n6063), .A3(n4820), .ZN(n6071) );
  AND3_X2 U6478 ( .A1(n4824), .A2(n4823), .A3(n4822), .ZN(n6063) );
  NOR2_X2 U6479 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4822) );
  NOR2_X2 U6480 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4823) );
  NOR2_X2 U6481 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4824) );
  NAND2_X1 U6482 ( .A1(n9294), .A2(n4829), .ZN(n4826) );
  NAND2_X1 U6483 ( .A1(n4827), .A2(n4826), .ZN(n9235) );
  NAND2_X1 U6484 ( .A1(n9304), .A2(n4838), .ZN(n4836) );
  NAND2_X1 U6485 ( .A1(n7962), .A2(n4849), .ZN(n4848) );
  NAND3_X1 U6486 ( .A1(n7943), .A2(n7946), .A3(n7947), .ZN(n9188) );
  NAND2_X1 U6487 ( .A1(n7943), .A2(n7947), .ZN(n9191) );
  NAND2_X1 U6488 ( .A1(n6080), .A2(n4396), .ZN(n4854) );
  NAND2_X1 U6489 ( .A1(n6080), .A2(n4855), .ZN(n6149) );
  NAND2_X1 U6490 ( .A1(n4854), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U6491 ( .A1(n6080), .A2(n6079), .ZN(n6126) );
  NAND3_X1 U6492 ( .A1(n4856), .A2(n9354), .A3(n9312), .ZN(n9365) );
  NAND2_X1 U6493 ( .A1(n5806), .A2(n4859), .ZN(n5808) );
  NAND2_X1 U6494 ( .A1(n7040), .A2(n4859), .ZN(n6954) );
  NAND3_X1 U6495 ( .A1(n5606), .A2(n5605), .A3(n4331), .ZN(n4868) );
  NAND2_X1 U6496 ( .A1(n4406), .A2(n5634), .ZN(n4871) );
  INV_X1 U6497 ( .A(n5634), .ZN(n4872) );
  NAND3_X1 U6498 ( .A1(n4877), .A2(n5623), .A3(n4876), .ZN(n5626) );
  AND2_X1 U6499 ( .A1(n5624), .A2(n5870), .ZN(n8906) );
  NAND2_X1 U6500 ( .A1(n8771), .A2(n4883), .ZN(n4878) );
  INV_X2 U6501 ( .A(n6636), .ZN(n5386) );
  INV_X1 U6502 ( .A(n4887), .ZN(n4886) );
  OAI22_X1 U6503 ( .A1(n7873), .A2(n5578), .B1(n6636), .B2(n4790), .ZN(n4887)
         );
  NAND2_X2 U6504 ( .A1(n6636), .A2(n6840), .ZN(n5578) );
  NAND2_X1 U6505 ( .A1(n6923), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6681) );
  NAND2_X1 U6506 ( .A1(n8635), .A2(n8636), .ZN(n8634) );
  AOI21_X1 U6507 ( .B1(n8659), .B2(P2_REG1_REG_13__SCAN_IN), .A(n4892), .ZN(
        n8675) );
  OR2_X1 U6508 ( .A1(n6695), .A2(n7033), .ZN(n4893) );
  NAND2_X1 U6509 ( .A1(n8615), .A2(n8614), .ZN(n8613) );
  NAND2_X1 U6510 ( .A1(n8442), .A2(n4901), .ZN(n4898) );
  NAND2_X1 U6511 ( .A1(n4898), .A2(n4899), .ZN(n8522) );
  NAND2_X1 U6512 ( .A1(n4906), .A2(n4399), .ZN(n8584) );
  NAND3_X1 U6513 ( .A1(n5357), .A2(n4322), .A3(n4405), .ZN(n5671) );
  NAND2_X4 U6514 ( .A1(n4914), .A2(n4913), .ZN(n5093) );
  NAND2_X1 U6515 ( .A1(n9868), .A2(n5023), .ZN(n4914) );
  NAND2_X1 U6516 ( .A1(n5128), .A2(n5127), .ZN(n4915) );
  NAND2_X1 U6517 ( .A1(n5061), .A2(n5062), .ZN(n4916) );
  NAND2_X1 U6518 ( .A1(n7892), .A2(n4920), .ZN(n4919) );
  NAND2_X1 U6519 ( .A1(n9572), .A2(n10064), .ZN(n4925) );
  NAND2_X1 U6520 ( .A1(n4926), .A2(n4925), .ZN(P1_U3551) );
  INV_X1 U6521 ( .A(n6139), .ZN(n4931) );
  AND2_X2 U6522 ( .A1(n6321), .A2(n4931), .ZN(n6394) );
  NAND4_X1 U6523 ( .A1(n6019), .A2(n6063), .A3(n4933), .A4(n4932), .ZN(n6069)
         );
  OAI211_X2 U6524 ( .C1(n7535), .C2(n4936), .A(n4330), .B(n4934), .ZN(n7813)
         );
  INV_X1 U6525 ( .A(n8261), .ZN(n4935) );
  OAI21_X2 U6526 ( .B1(n7559), .B2(n7562), .A(n6603), .ZN(n7535) );
  INV_X1 U6527 ( .A(n4939), .ZN(n4940) );
  OAI21_X2 U6528 ( .B1(n9690), .B2(n4945), .A(n4943), .ZN(n9640) );
  INV_X2 U6529 ( .A(n5578), .ZN(n5537) );
  NAND2_X1 U6530 ( .A1(n9737), .A2(n10055), .ZN(n6190) );
  NAND2_X1 U6531 ( .A1(n5669), .A2(n8396), .ZN(n5731) );
  AND2_X1 U6532 ( .A1(n6636), .A2(n5657), .ZN(n6276) );
  NAND2_X1 U6533 ( .A1(n9584), .A2(n9962), .ZN(n9588) );
  NAND2_X1 U6534 ( .A1(n6394), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6578) );
  AOI21_X1 U6535 ( .B1(n5706), .B2(n5707), .A(n5672), .ZN(n5675) );
  INV_X1 U6536 ( .A(n7054), .ZN(n6002) );
  NAND2_X1 U6537 ( .A1(n4975), .A2(n6374), .ZN(n7054) );
  NAND2_X1 U6538 ( .A1(n6156), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n6157) );
  INV_X1 U6539 ( .A(n6080), .ZN(n6075) );
  INV_X2 U6540 ( .A(n5060), .ZN(n5244) );
  CLKBUF_X1 U6541 ( .A(n8584), .Z(n8585) );
  NOR2_X1 U6542 ( .A1(n6092), .A2(n6091), .ZN(n6097) );
  AOI211_X2 U6543 ( .C1(n9991), .C2(n9741), .A(n9590), .B(n9589), .ZN(n9591)
         );
  NAND2_X1 U6544 ( .A1(n7056), .A2(n7257), .ZN(n7285) );
  OR2_X1 U6545 ( .A1(n6122), .A2(n7872), .ZN(n6001) );
  OR2_X1 U6546 ( .A1(n6122), .A2(n6841), .ZN(n5995) );
  NAND2_X1 U6547 ( .A1(n5774), .A2(n4994), .ZN(n5803) );
  INV_X1 U6548 ( .A(n9576), .ZN(n6568) );
  AOI21_X1 U6549 ( .B1(n6272), .B2(n8079), .A(n6271), .ZN(n8571) );
  AND2_X1 U6550 ( .A1(n6272), .A2(n6267), .ZN(n6312) );
  CLKBUF_X1 U6551 ( .A(n7559), .Z(n7596) );
  XNOR2_X1 U6552 ( .A(n9556), .B(n8234), .ZN(n6132) );
  NAND2_X1 U6553 ( .A1(n7940), .A2(n7939), .ZN(n7943) );
  NAND2_X2 U6554 ( .A1(n6223), .A2(n5853), .ZN(n8462) );
  NAND2_X1 U6555 ( .A1(n6310), .A2(n6309), .ZN(n6311) );
  AND2_X1 U6556 ( .A1(n6821), .A2(n6769), .ZN(n6771) );
  AND2_X1 U6557 ( .A1(n6821), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6168) );
  INV_X1 U6558 ( .A(n7692), .ZN(n7697) );
  NAND2_X1 U6559 ( .A1(n4314), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6577) );
  CLKBUF_X1 U6560 ( .A(n5688), .Z(n8112) );
  AND2_X1 U6561 ( .A1(n8422), .A2(n8846), .ZN(n8424) );
  AND3_X1 U6562 ( .A1(n6397), .A2(n6396), .A3(n6395), .ZN(n4968) );
  NOR2_X1 U6563 ( .A1(n5617), .A2(n5616), .ZN(n4969) );
  NOR2_X1 U6564 ( .A1(n5371), .A2(n5370), .ZN(n4970) );
  AND2_X1 U6565 ( .A1(n5653), .A2(n5921), .ZN(n4971) );
  AND2_X1 U6566 ( .A1(n7517), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4973) );
  INV_X1 U6567 ( .A(n8193), .ZN(n9730) );
  AND2_X1 U6568 ( .A1(n5373), .A2(SI_18_), .ZN(n4974) );
  NAND2_X1 U6569 ( .A1(n5717), .A2(n5716), .ZN(n9073) );
  INV_X1 U6570 ( .A(n9646), .ZN(n6495) );
  INV_X1 U6571 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n5377) );
  AND2_X1 U6572 ( .A1(n8568), .A2(n8567), .ZN(n4976) );
  AND2_X1 U6573 ( .A1(n7187), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4978) );
  AND2_X1 U6574 ( .A1(n7012), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4979) );
  OR2_X1 U6575 ( .A1(n5993), .A2(n7080), .ZN(n4980) );
  AND2_X1 U6576 ( .A1(n4318), .A2(n7131), .ZN(n4981) );
  INV_X1 U6577 ( .A(n6375), .ZN(n6390) );
  AND2_X1 U6578 ( .A1(n9461), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4982) );
  INV_X1 U6579 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5336) );
  INV_X1 U6580 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n5399) );
  INV_X1 U6581 ( .A(n8387), .ZN(n9183) );
  NAND2_X1 U6582 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n4983) );
  INV_X1 U6583 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5092) );
  AND3_X1 U6584 ( .A1(n8406), .A2(n8402), .A3(n8557), .ZN(n4984) );
  AND2_X1 U6585 ( .A1(n5823), .A2(n7385), .ZN(n4985) );
  NAND2_X1 U6586 ( .A1(n8567), .A2(n8077), .ZN(n4986) );
  NOR2_X1 U6587 ( .A1(n6300), .A2(n8815), .ZN(n4987) );
  INV_X1 U6588 ( .A(n9826), .ZN(n6057) );
  AND2_X1 U6589 ( .A1(n6660), .A2(n6740), .ZN(n4988) );
  AND3_X1 U6590 ( .A1(n5802), .A2(n5801), .A3(n7604), .ZN(n4989) );
  OR2_X1 U6591 ( .A1(n8354), .A2(n4319), .ZN(n9710) );
  INV_X1 U6592 ( .A(n8124), .ZN(n6402) );
  NOR2_X1 U6593 ( .A1(n8100), .A2(n8099), .ZN(n4991) );
  AND2_X1 U6594 ( .A1(n8770), .A2(n5918), .ZN(n4992) );
  AND2_X1 U6595 ( .A1(n6206), .A2(n8607), .ZN(n4993) );
  INV_X1 U6596 ( .A(n7257), .ZN(n7430) );
  AND2_X1 U6597 ( .A1(n6191), .A2(n5799), .ZN(n4994) );
  AND2_X1 U6598 ( .A1(n6191), .A2(n5797), .ZN(n4995) );
  AND2_X1 U6599 ( .A1(n5647), .A2(n5646), .ZN(n8967) );
  AOI21_X1 U6600 ( .B1(n8304), .B2(n8181), .A(n8180), .ZN(n8191) );
  NAND2_X1 U6601 ( .A1(n5882), .A2(n6634), .ZN(n5883) );
  OAI21_X1 U6602 ( .B1(n5885), .B2(n5884), .A(n5883), .ZN(n5886) );
  INV_X1 U6603 ( .A(n5902), .ZN(n5903) );
  NOR2_X1 U6604 ( .A1(n7764), .A2(n7763), .ZN(n7765) );
  OR4_X1 U6605 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6179) );
  OR2_X1 U6606 ( .A1(n9058), .A2(n8951), .ZN(n5619) );
  INV_X1 U6607 ( .A(n8244), .ZN(n6443) );
  INV_X1 U6608 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5458) );
  INV_X1 U6609 ( .A(n8608), .ZN(n6202) );
  NAND2_X1 U6610 ( .A1(n5924), .A2(n5923), .ZN(n5932) );
  OR2_X1 U6611 ( .A1(n6634), .A2(n5944), .ZN(n6282) );
  INV_X1 U6612 ( .A(n7581), .ZN(n5189) );
  INV_X1 U6613 ( .A(n6820), .ZN(n6817) );
  OAI21_X1 U6614 ( .B1(n8370), .B2(n8365), .A(n8364), .ZN(n8366) );
  INV_X1 U6615 ( .A(n8098), .ZN(n6321) );
  INV_X1 U6616 ( .A(n7015), .ZN(n6014) );
  NAND2_X1 U6617 ( .A1(n7491), .A2(n10004), .ZN(n8139) );
  INV_X1 U6618 ( .A(SI_24_), .ZN(n5476) );
  INV_X1 U6619 ( .A(SI_22_), .ZN(n5418) );
  INV_X1 U6620 ( .A(n5368), .ZN(n5371) );
  INV_X1 U6621 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6035) );
  INV_X1 U6622 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6024) );
  INV_X1 U6623 ( .A(n7627), .ZN(n6215) );
  NOR2_X1 U6624 ( .A1(n5732), .A2(n9065), .ZN(n5718) );
  NOR2_X1 U6625 ( .A1(n8576), .A2(n8971), .ZN(n5956) );
  INV_X1 U6626 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10221) );
  OR2_X1 U6627 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5590) );
  INV_X1 U6628 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U6629 ( .A1(n5980), .A2(n5979), .ZN(n5985) );
  NAND2_X1 U6630 ( .A1(n6532), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U6631 ( .A1(n6452), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6462) );
  AND2_X1 U6632 ( .A1(n7415), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7416) );
  AOI21_X1 U6633 ( .B1(n9860), .B2(n6058), .A(n4426), .ZN(n8234) );
  NAND2_X1 U6634 ( .A1(n6871), .A2(n6014), .ZN(n6015) );
  NOR2_X1 U6635 ( .A1(n4970), .A2(n4974), .ZN(n5374) );
  OR2_X1 U6636 ( .A1(n5352), .A2(n5351), .ZN(n5370) );
  NAND2_X1 U6637 ( .A1(n5171), .A2(n5197), .ZN(n5193) );
  NAND2_X1 U6638 ( .A1(n5093), .A2(n6841), .ZN(n5051) );
  NAND2_X1 U6639 ( .A1(n6211), .A2(n8605), .ZN(n6213) );
  INV_X1 U6640 ( .A(n8899), .ZN(n8446) );
  INV_X1 U6641 ( .A(n8879), .ZN(n8455) );
  INV_X1 U6642 ( .A(n8889), .ZN(n8913) );
  INV_X1 U6643 ( .A(n8587), .ZN(n8575) );
  OR2_X1 U6644 ( .A1(n6296), .A2(n6295), .ZN(n8590) );
  INV_X1 U6645 ( .A(n10114), .ZN(n8668) );
  OR3_X1 U6646 ( .A1(n5709), .A2(n5725), .A3(n6303), .ZN(n6980) );
  INV_X1 U6647 ( .A(n8971), .ZN(n8952) );
  INV_X1 U6648 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10160) );
  INV_X1 U6649 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9327) );
  OR2_X1 U6650 ( .A1(n6826), .A2(n8374), .ZN(n6830) );
  NAND2_X1 U6651 ( .A1(n9518), .A2(n9517), .ZN(n9520) );
  OR2_X1 U6652 ( .A1(n9773), .A2(n9388), .ZN(n6615) );
  AND2_X1 U6653 ( .A1(n8199), .A2(n8194), .ZN(n8193) );
  INV_X1 U6654 ( .A(n7569), .ZN(n7619) );
  INV_X1 U6655 ( .A(n6363), .ZN(n9995) );
  NOR2_X1 U6656 ( .A1(n9724), .A2(n9550), .ZN(n6831) );
  NAND2_X1 U6657 ( .A1(n9562), .A2(n6629), .ZN(n6630) );
  INV_X1 U6658 ( .A(n10020), .ZN(n10047) );
  NAND2_X1 U6659 ( .A1(n7639), .A2(n8286), .ZN(n7321) );
  XNOR2_X1 U6660 ( .A(n5260), .B(n5255), .ZN(n6051) );
  OAI21_X1 U6661 ( .B1(n8818), .B2(n8596), .A(n6317), .ZN(n6318) );
  NAND2_X1 U6662 ( .A1(n7038), .A2(n5805), .ZN(n7218) );
  INV_X1 U6663 ( .A(n8590), .ZN(n8572) );
  NAND2_X1 U6664 ( .A1(n6275), .A2(n6274), .ZN(n8557) );
  OR2_X1 U6665 ( .A1(n6749), .A2(n8111), .ZN(n6758) );
  INV_X1 U6666 ( .A(n8748), .ZN(n10118) );
  OR2_X1 U6667 ( .A1(n6303), .A2(n6302), .ZN(n8989) );
  INV_X1 U6668 ( .A(n8991), .ZN(n8977) );
  INV_X1 U6669 ( .A(n9065), .ZN(n9054) );
  OAI21_X1 U6670 ( .B1(n6982), .B2(n5715), .A(n6983), .ZN(n5716) );
  NAND2_X1 U6671 ( .A1(n7529), .A2(n7641), .ZN(n7407) );
  INV_X1 U6672 ( .A(n9095), .ZN(n9167) );
  NAND2_X1 U6673 ( .A1(n7687), .A2(n7103), .ZN(n7501) );
  OR2_X1 U6674 ( .A1(n6296), .A2(n5728), .ZN(n5729) );
  INV_X1 U6675 ( .A(n7849), .ZN(n8110) );
  XNOR2_X1 U6676 ( .A(n5246), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6728) );
  AND2_X1 U6677 ( .A1(n6557), .A2(n6556), .ZN(n8067) );
  INV_X1 U6678 ( .A(n6561), .ZN(n6554) );
  AND4_X1 U6679 ( .A1(n6425), .A2(n6424), .A3(n6423), .A4(n6422), .ZN(n9231)
         );
  INV_X1 U6680 ( .A(n7095), .ZN(n9947) );
  INV_X1 U6681 ( .A(n9710), .ZN(n9673) );
  INV_X1 U6682 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6188) );
  AND2_X1 U6683 ( .A1(n7835), .A2(n10031), .ZN(n10051) );
  INV_X1 U6684 ( .A(n10051), .ZN(n10026) );
  NAND2_X1 U6685 ( .A1(n6173), .A2(n6172), .ZN(n6860) );
  AND2_X1 U6686 ( .A1(n6027), .A2(n6065), .ZN(n9461) );
  INV_X1 U6687 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9878) );
  INV_X1 U6688 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9884) );
  INV_X1 U6689 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9893) );
  NOR2_X1 U6690 ( .A1(n10151), .A2(n10150), .ZN(n9900) );
  NOR2_X1 U6691 ( .A1(n10145), .A2(n10144), .ZN(n9907) );
  NAND2_X1 U6692 ( .A1(n8413), .A2(n4984), .ZN(n8412) );
  INV_X1 U6693 ( .A(n8557), .ZN(n8581) );
  INV_X1 U6694 ( .A(n8578), .ZN(n8596) );
  INV_X1 U6695 ( .A(n8537), .ZN(n8601) );
  OR2_X1 U6696 ( .A1(P2_U3150), .A2(n6759), .ZN(n8748) );
  OR2_X1 U6697 ( .A1(n6699), .A2(n6743), .ZN(n10106) );
  INV_X1 U6698 ( .A(n8764), .ZN(n8980) );
  NOR2_X1 U6699 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  OR2_X1 U6700 ( .A1(n9073), .A2(n7407), .ZN(n9065) );
  OR2_X1 U6701 ( .A1(n9073), .A2(n9072), .ZN(n9061) );
  NAND2_X1 U6702 ( .A1(n5734), .A2(n9069), .ZN(n9095) );
  NAND2_X1 U6703 ( .A1(n5734), .A2(n7501), .ZN(n9173) );
  AND2_X1 U6704 ( .A1(n5730), .A2(n5729), .ZN(n10292) );
  INV_X1 U6705 ( .A(n5949), .ZN(n7641) );
  INV_X1 U6706 ( .A(n6730), .ZN(n8665) );
  INV_X1 U6707 ( .A(n6925), .ZN(n6854) );
  INV_X1 U6708 ( .A(n9789), .ZN(n9694) );
  INV_X1 U6709 ( .A(n9317), .ZN(n9375) );
  INV_X1 U6710 ( .A(n8067), .ZN(n9585) );
  OR2_X1 U6711 ( .A1(n6466), .A2(n6465), .ZN(n9389) );
  INV_X1 U6712 ( .A(n7910), .ZN(n9396) );
  OR2_X1 U6713 ( .A1(n7026), .A2(n8372), .ZN(n9934) );
  OR2_X1 U6714 ( .A1(n7026), .A2(n7067), .ZN(n9944) );
  NAND2_X1 U6715 ( .A1(n9989), .A2(n9981), .ZN(n9736) );
  INV_X2 U6716 ( .A(n9989), .ZN(n10001) );
  INV_X1 U6717 ( .A(n10064), .ZN(n10062) );
  AND2_X2 U6718 ( .A1(n6767), .A2(n6815), .ZN(n10064) );
  INV_X1 U6719 ( .A(n10055), .ZN(n10053) );
  AND2_X2 U6720 ( .A1(n6767), .A2(n7293), .ZN(n10055) );
  AND2_X1 U6721 ( .A1(n7855), .A2(n7830), .ZN(n6862) );
  XNOR2_X1 U6722 ( .A(n6160), .B(n6159), .ZN(n7830) );
  INV_X1 U6723 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7438) );
  INV_X1 U6724 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6908) );
  NOR2_X1 U6725 ( .A1(n9889), .A2(n9888), .ZN(n10304) );
  NOR2_X1 U6726 ( .A1(n9901), .A2(n9900), .ZN(n10149) );
  INV_X1 U6727 ( .A(n8743), .ZN(P2_U3893) );
  OAI21_X1 U6728 ( .B1(n6763), .B2(n10292), .A(n5962), .ZN(P2_U3455) );
  AND2_X2 U6729 ( .A1(n6768), .A2(n6872), .ZN(P1_U3973) );
  NAND2_X1 U6730 ( .A1(n6190), .A2(n6189), .ZN(P1_U3521) );
  NOR2_X1 U6731 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4997) );
  NOR2_X1 U6732 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n4996) );
  INV_X1 U6733 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5008) );
  INV_X1 U6734 ( .A(n5012), .ZN(n5010) );
  NAND2_X1 U6735 ( .A1(n5010), .A2(n5009), .ZN(n9175) );
  XNOR2_X2 U6736 ( .A(n5011), .B(n9176), .ZN(n8384) );
  NAND2_X1 U6737 ( .A1(n5012), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5013) );
  INV_X1 U6738 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5014) );
  INV_X1 U6739 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7149) );
  OR2_X1 U6740 ( .A1(n5079), .A2(n7149), .ZN(n5017) );
  INV_X1 U6741 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6964) );
  NAND4_X1 U6742 ( .A1(n5019), .A2(n5018), .A3(n5017), .A4(n5016), .ZN(n5600)
         );
  NAND2_X1 U6743 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5022) );
  BUF_X8 U6744 ( .A(n5093), .Z(n6837) );
  INV_X1 U6745 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6839) );
  OR2_X1 U6746 ( .A1(n5060), .A2(n6839), .ZN(n5030) );
  NAND2_X1 U6747 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5026) );
  AND2_X1 U6748 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6749 ( .A1(n5093), .A2(n5025), .ZN(n5989) );
  OAI21_X1 U6750 ( .B1(n5093), .B2(n5026), .A(n5989), .ZN(n5047) );
  XNOR2_X1 U6751 ( .A(n5047), .B(SI_1_), .ZN(n5028) );
  XNOR2_X1 U6752 ( .A(n5027), .B(n5028), .ZN(n5981) );
  INV_X1 U6753 ( .A(n5981), .ZN(n6851) );
  NAND2_X1 U6754 ( .A1(n5600), .A2(n7041), .ZN(n5807) );
  INV_X1 U6755 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5031) );
  INV_X1 U6756 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6701) );
  INV_X1 U6757 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7220) );
  OR2_X1 U6758 ( .A1(n5079), .A2(n7220), .ZN(n5033) );
  INV_X1 U6759 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10163) );
  INV_X1 U6760 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U6761 ( .A1(n6840), .A2(SI_0_), .ZN(n5037) );
  INV_X1 U6762 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5036) );
  XNOR2_X1 U6763 ( .A(n5037), .B(n5036), .ZN(n9186) );
  MUX2_X1 U6764 ( .A(n6666), .B(n9186), .S(n6636), .Z(n7216) );
  INV_X1 U6765 ( .A(n7038), .ZN(n5038) );
  INV_X1 U6766 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8611) );
  OR2_X1 U6767 ( .A1(n5079), .A2(n8611), .ZN(n5041) );
  INV_X1 U6768 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6640) );
  OR2_X1 U6769 ( .A1(n5236), .A2(n6640), .ZN(n5040) );
  INV_X1 U6770 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6665) );
  OR2_X1 U6771 ( .A1(n5585), .A2(n6665), .ZN(n5039) );
  INV_X1 U6772 ( .A(SI_1_), .ZN(n5044) );
  OAI211_X1 U6773 ( .C1(n5093), .C2(n6839), .A(n5045), .B(n5044), .ZN(n5046)
         );
  NAND2_X1 U6774 ( .A1(n5047), .A2(n5046), .ZN(n5050) );
  INV_X1 U6775 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U6776 ( .A1(n5093), .A2(n6850), .ZN(n5048) );
  OAI211_X1 U6777 ( .C1(n5093), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n5048), .B(
        SI_1_), .ZN(n5049) );
  NAND2_X1 U6778 ( .A1(n5050), .A2(n5049), .ZN(n5062) );
  INV_X1 U6779 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6843) );
  INV_X1 U6780 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6841) );
  XNOR2_X1 U6781 ( .A(n5063), .B(SI_2_), .ZN(n5061) );
  XNOR2_X1 U6782 ( .A(n5062), .B(n5061), .ZN(n6842) );
  NAND2_X1 U6783 ( .A1(n8608), .A2(n6959), .ZN(n5815) );
  NAND2_X1 U6784 ( .A1(n5053), .A2(n5816), .ZN(n7110) );
  INV_X1 U6785 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5059) );
  INV_X1 U6786 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7160) );
  OR2_X1 U6787 ( .A1(n5236), .A2(n7160), .ZN(n5056) );
  OR2_X1 U6788 ( .A1(n5079), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5055) );
  INV_X1 U6789 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10065) );
  OR2_X1 U6790 ( .A1(n5585), .A2(n10065), .ZN(n5057) );
  INV_X1 U6791 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7874) );
  INV_X1 U6792 ( .A(n5063), .ZN(n5064) );
  NAND2_X1 U6793 ( .A1(n5064), .A2(SI_2_), .ZN(n5065) );
  INV_X1 U6794 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7872) );
  MUX2_X1 U6795 ( .A(n7874), .B(n7872), .S(n5093), .Z(n5069) );
  XNOR2_X1 U6796 ( .A(n5069), .B(SI_3_), .ZN(n5067) );
  XNOR2_X1 U6797 ( .A(n5067), .B(n5068), .ZN(n7873) );
  INV_X1 U6798 ( .A(n7222), .ZN(n7116) );
  NAND2_X1 U6799 ( .A1(n8607), .A2(n7116), .ZN(n5832) );
  NAND2_X1 U6800 ( .A1(n7110), .A2(n7113), .ZN(n5066) );
  INV_X1 U6801 ( .A(n5069), .ZN(n5070) );
  MUX2_X1 U6802 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5093), .Z(n5087) );
  INV_X1 U6803 ( .A(SI_4_), .ZN(n5072) );
  XNOR2_X1 U6804 ( .A(n5087), .B(n5072), .ZN(n5086) );
  OR2_X1 U6805 ( .A1(n6007), .A2(n5578), .ZN(n5078) );
  INV_X1 U6806 ( .A(n5175), .ZN(n5073) );
  NAND2_X1 U6807 ( .A1(n5073), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5074) );
  MUX2_X1 U6808 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5074), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5076) );
  NAND2_X1 U6809 ( .A1(n5175), .A2(n5075), .ZN(n5114) );
  NAND2_X1 U6810 ( .A1(n5076), .A2(n5114), .ZN(n6852) );
  INV_X1 U6811 ( .A(n6852), .ZN(n8630) );
  AOI22_X1 U6812 ( .A1(n5244), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8630), .B2(
        n5386), .ZN(n5077) );
  NAND2_X1 U6813 ( .A1(n5078), .A2(n5077), .ZN(n7170) );
  INV_X2 U6814 ( .A(n7170), .ZN(n7235) );
  NAND2_X1 U6815 ( .A1(n5582), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5085) );
  INV_X1 U6816 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6677) );
  OR2_X1 U6817 ( .A1(n5585), .A2(n6677), .ZN(n5084) );
  NAND2_X1 U6818 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5081) );
  AND2_X1 U6819 ( .A1(n5105), .A2(n5081), .ZN(n7239) );
  OR2_X1 U6820 ( .A1(n5079), .A2(n7239), .ZN(n5083) );
  INV_X1 U6821 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7168) );
  OR2_X1 U6822 ( .A1(n5236), .A2(n7168), .ZN(n5082) );
  NAND4_X1 U6823 ( .A1(n5085), .A2(n5084), .A3(n5083), .A4(n5082), .ZN(n7153)
         );
  NAND2_X1 U6824 ( .A1(n7235), .A2(n7153), .ZN(n5822) );
  OR2_X1 U6825 ( .A1(n7153), .A2(n7235), .ZN(n5833) );
  NAND2_X1 U6826 ( .A1(n5087), .A2(SI_4_), .ZN(n5120) );
  NAND2_X1 U6827 ( .A1(n5122), .A2(n5120), .ZN(n5113) );
  INV_X1 U6828 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6855) );
  INV_X1 U6829 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U6830 ( .A1(n5113), .A2(n5123), .ZN(n5090) );
  INV_X1 U6831 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6832 ( .A1(n5089), .A2(SI_5_), .ZN(n5119) );
  NAND2_X1 U6833 ( .A1(n5090), .A2(n5119), .ZN(n5094) );
  XNOR2_X1 U6834 ( .A(n5129), .B(SI_6_), .ZN(n5124) );
  XNOR2_X1 U6835 ( .A(n5094), .B(n5124), .ZN(n6847) );
  NAND2_X1 U6836 ( .A1(n6847), .A2(n5537), .ZN(n5097) );
  NAND2_X1 U6837 ( .A1(n5131), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5095) );
  AOI22_X1 U6838 ( .A1(n5244), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6715), .B2(
        n5386), .ZN(n5096) );
  NAND2_X1 U6839 ( .A1(n5097), .A2(n5096), .ZN(n9068) );
  NAND2_X1 U6840 ( .A1(n5582), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5103) );
  INV_X1 U6841 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7372) );
  OR2_X1 U6842 ( .A1(n5236), .A2(n7372), .ZN(n5102) );
  NAND2_X1 U6843 ( .A1(n5107), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5099) );
  AND2_X1 U6844 ( .A1(n5140), .A2(n5099), .ZN(n7373) );
  OR2_X1 U6845 ( .A1(n5581), .A2(n7373), .ZN(n5101) );
  INV_X1 U6846 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6682) );
  OR2_X1 U6847 ( .A1(n5585), .A2(n6682), .ZN(n5100) );
  NAND4_X1 U6848 ( .A1(n5103), .A2(n5102), .A3(n5101), .A4(n5100), .ZN(n8605)
         );
  INV_X1 U6849 ( .A(n8605), .ZN(n6212) );
  OR2_X1 U6850 ( .A1(n9068), .A2(n6212), .ZN(n7379) );
  NAND2_X1 U6851 ( .A1(n5582), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5112) );
  INV_X1 U6852 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5104) );
  OR2_X1 U6853 ( .A1(n5585), .A2(n5104), .ZN(n5111) );
  NAND2_X1 U6854 ( .A1(n5105), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5106) );
  AND2_X1 U6855 ( .A1(n5107), .A2(n5106), .ZN(n7319) );
  OR2_X1 U6856 ( .A1(n5581), .A2(n7319), .ZN(n5110) );
  INV_X2 U6857 ( .A(n5236), .ZN(n5108) );
  INV_X1 U6858 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7202) );
  OR2_X1 U6859 ( .A1(n6856), .A2(n5578), .ZN(n5118) );
  NAND2_X1 U6860 ( .A1(n5114), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5115) );
  MUX2_X1 U6861 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5115), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5116) );
  AOI22_X1 U6862 ( .A1(n5244), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6925), .B2(
        n5386), .ZN(n5117) );
  NAND2_X1 U6863 ( .A1(n5118), .A2(n5117), .ZN(n7204) );
  OR2_X1 U6864 ( .A1(n7370), .A2(n7204), .ZN(n7364) );
  AND2_X1 U6865 ( .A1(n7379), .A2(n7364), .ZN(n5839) );
  NAND2_X1 U6866 ( .A1(n9068), .A2(n6212), .ZN(n5836) );
  NAND2_X1 U6867 ( .A1(n7370), .A2(n7204), .ZN(n7365) );
  NAND2_X1 U6868 ( .A1(n5836), .A2(n7365), .ZN(n7376) );
  NAND2_X1 U6869 ( .A1(n7376), .A2(n7379), .ZN(n5823) );
  AND2_X1 U6870 ( .A1(n5120), .A2(n5126), .ZN(n5121) );
  NAND2_X1 U6871 ( .A1(n5122), .A2(n5121), .ZN(n5128) );
  NAND2_X1 U6872 ( .A1(n5129), .A2(SI_6_), .ZN(n5130) );
  NAND2_X1 U6873 ( .A1(n6844), .A2(n5537), .ZN(n5136) );
  INV_X1 U6874 ( .A(n5131), .ZN(n5133) );
  NAND2_X1 U6875 ( .A1(n5133), .A2(n5132), .ZN(n5153) );
  NAND2_X1 U6876 ( .A1(n5153), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5134) );
  XNOR2_X1 U6877 ( .A(n5134), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6716) );
  AOI22_X1 U6878 ( .A1(n5244), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6716), .B2(
        n5386), .ZN(n5135) );
  NAND2_X1 U6879 ( .A1(n5136), .A2(n5135), .ZN(n7631) );
  NAND2_X1 U6880 ( .A1(n5582), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5146) );
  INV_X1 U6881 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5137) );
  OR2_X1 U6882 ( .A1(n5236), .A2(n5137), .ZN(n5145) );
  NAND2_X1 U6883 ( .A1(n5140), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5141) );
  AND2_X1 U6884 ( .A1(n5157), .A2(n5141), .ZN(n7629) );
  OR2_X1 U6885 ( .A1(n5581), .A2(n7629), .ZN(n5144) );
  INV_X1 U6886 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5142) );
  OR2_X1 U6887 ( .A1(n5585), .A2(n5142), .ZN(n5143) );
  OR2_X1 U6888 ( .A1(n7631), .A2(n7700), .ZN(n7455) );
  NAND2_X1 U6889 ( .A1(n7631), .A2(n7700), .ZN(n5824) );
  NAND2_X1 U6890 ( .A1(n5147), .A2(n4985), .ZN(n7383) );
  INV_X1 U6891 ( .A(n5148), .ZN(n5149) );
  INV_X1 U6892 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6864) );
  INV_X1 U6893 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6866) );
  INV_X1 U6894 ( .A(SI_8_), .ZN(n5150) );
  NAND2_X1 U6895 ( .A1(n5151), .A2(n5150), .ZN(n5196) );
  INV_X1 U6896 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6897 ( .A1(n5152), .A2(SI_8_), .ZN(n5191) );
  NAND2_X1 U6898 ( .A1(n5196), .A2(n5191), .ZN(n5165) );
  NAND2_X1 U6899 ( .A1(n6863), .A2(n5537), .ZN(n5156) );
  OAI21_X1 U6900 ( .B1(n5153), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5154) );
  AOI22_X1 U6901 ( .A1(n5244), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6720), .B2(
        n5386), .ZN(n5155) );
  NAND2_X1 U6902 ( .A1(n5156), .A2(n5155), .ZN(n7701) );
  NAND2_X1 U6903 ( .A1(n5582), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5162) );
  INV_X1 U6904 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7506) );
  OR2_X1 U6905 ( .A1(n5236), .A2(n7506), .ZN(n5161) );
  NAND2_X1 U6906 ( .A1(n5157), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5158) );
  AND2_X1 U6907 ( .A1(n5183), .A2(n5158), .ZN(n7507) );
  OR2_X1 U6908 ( .A1(n5581), .A2(n7507), .ZN(n5160) );
  INV_X1 U6909 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7502) );
  OR2_X1 U6910 ( .A1(n5585), .A2(n7502), .ZN(n5159) );
  NAND4_X1 U6911 ( .A1(n5162), .A2(n5161), .A3(n5160), .A4(n5159), .ZN(n8603)
         );
  INV_X1 U6912 ( .A(n8603), .ZN(n5163) );
  OR2_X1 U6913 ( .A1(n7701), .A2(n5163), .ZN(n5826) );
  AND2_X1 U6914 ( .A1(n5826), .A2(n7455), .ZN(n5848) );
  NAND2_X1 U6915 ( .A1(n7701), .A2(n5163), .ZN(n5825) );
  INV_X1 U6916 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6870) );
  INV_X1 U6917 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6883) );
  INV_X1 U6918 ( .A(n5170), .ZN(n5168) );
  NAND2_X1 U6919 ( .A1(n5168), .A2(SI_9_), .ZN(n5171) );
  INV_X1 U6920 ( .A(SI_9_), .ZN(n5169) );
  NAND2_X1 U6921 ( .A1(n5170), .A2(n5169), .ZN(n5197) );
  NAND2_X1 U6922 ( .A1(n6869), .A2(n5537), .ZN(n5179) );
  INV_X1 U6923 ( .A(n5173), .ZN(n5174) );
  INV_X1 U6924 ( .A(n5357), .ZN(n5176) );
  NAND2_X1 U6925 ( .A1(n5176), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5177) );
  XNOR2_X1 U6926 ( .A(n5177), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6721) );
  AOI22_X1 U6927 ( .A1(n5244), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6721), .B2(
        n5386), .ZN(n5178) );
  NAND2_X1 U6928 ( .A1(n5582), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5188) );
  INV_X1 U6929 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5180) );
  OR2_X1 U6930 ( .A1(n5762), .A2(n5180), .ZN(n5187) );
  NAND2_X1 U6931 ( .A1(n5183), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5184) );
  AND2_X1 U6932 ( .A1(n5214), .A2(n5184), .ZN(n8990) );
  OR2_X1 U6933 ( .A1(n5581), .A2(n8990), .ZN(n5186) );
  INV_X1 U6934 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7728) );
  OR2_X1 U6935 ( .A1(n5585), .A2(n7728), .ZN(n5185) );
  NAND4_X1 U6936 ( .A1(n5188), .A2(n5187), .A3(n5186), .A4(n5185), .ZN(n8602)
         );
  NAND2_X1 U6937 ( .A1(n8502), .A2(n8437), .ZN(n5828) );
  NAND2_X1 U6938 ( .A1(n5841), .A2(n5828), .ZN(n7581) );
  NAND2_X1 U6939 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  NOR2_X1 U6940 ( .A1(n5193), .A2(n5192), .ZN(n5194) );
  INV_X1 U6941 ( .A(n5196), .ZN(n5199) );
  INV_X1 U6942 ( .A(n5197), .ZN(n5198) );
  MUX2_X1 U6943 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6837), .Z(n5224) );
  INV_X1 U6944 ( .A(SI_10_), .ZN(n5203) );
  XNOR2_X1 U6945 ( .A(n5224), .B(n5203), .ZN(n5223) );
  NAND2_X1 U6946 ( .A1(n6858), .A2(n5537), .ZN(n5211) );
  INV_X1 U6947 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5204) );
  AND2_X1 U6948 ( .A1(n5357), .A2(n5204), .ZN(n5208) );
  INV_X1 U6949 ( .A(n5208), .ZN(n5205) );
  NAND2_X1 U6950 ( .A1(n5205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5206) );
  MUX2_X1 U6951 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5206), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n5209) );
  NAND2_X1 U6952 ( .A1(n5208), .A2(n5207), .ZN(n5245) );
  NAND2_X1 U6953 ( .A1(n5209), .A2(n5245), .ZN(n7444) );
  INV_X1 U6954 ( .A(n7444), .ZN(n6725) );
  AOI22_X1 U6955 ( .A1(n5244), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6725), .B2(
        n5386), .ZN(n5210) );
  NAND2_X1 U6956 ( .A1(n5758), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5220) );
  INV_X1 U6957 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5213) );
  OR2_X1 U6958 ( .A1(n5759), .A2(n5213), .ZN(n5219) );
  NAND2_X1 U6959 ( .A1(n5214), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5215) );
  AND2_X1 U6960 ( .A1(n5234), .A2(n5215), .ZN(n8983) );
  OR2_X1 U6961 ( .A1(n5581), .A2(n8983), .ZN(n5218) );
  INV_X1 U6962 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5216) );
  OR2_X1 U6963 ( .A1(n5236), .A2(n5216), .ZN(n5217) );
  NOR2_X1 U6964 ( .A1(n7690), .A2(n8537), .ZN(n5849) );
  INV_X1 U6965 ( .A(n5849), .ZN(n5221) );
  NAND2_X1 U6966 ( .A1(n5224), .A2(SI_10_), .ZN(n5225) );
  MUX2_X1 U6967 ( .A(n6888), .B(n6890), .S(n6837), .Z(n5228) );
  INV_X1 U6968 ( .A(SI_11_), .ZN(n5227) );
  NAND2_X1 U6969 ( .A1(n5228), .A2(n5227), .ZN(n5243) );
  INV_X1 U6970 ( .A(n5228), .ZN(n5229) );
  NAND2_X1 U6971 ( .A1(n5229), .A2(SI_11_), .ZN(n5230) );
  NAND2_X1 U6972 ( .A1(n5243), .A2(n5230), .ZN(n5241) );
  XNOR2_X1 U6973 ( .A(n5242), .B(n5241), .ZN(n6887) );
  NAND2_X1 U6974 ( .A1(n6887), .A2(n5537), .ZN(n5233) );
  NAND2_X1 U6975 ( .A1(n5245), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5231) );
  XNOR2_X1 U6976 ( .A(n5231), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6726) );
  AOI22_X1 U6977 ( .A1(n5244), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6726), .B2(
        n5386), .ZN(n5232) );
  NAND2_X2 U6978 ( .A1(n5233), .A2(n5232), .ZN(n8538) );
  NAND2_X1 U6979 ( .A1(n5758), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5240) );
  INV_X1 U6980 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7717) );
  OR2_X1 U6981 ( .A1(n5759), .A2(n7717), .ZN(n5239) );
  NAND2_X1 U6982 ( .A1(n5234), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5235) );
  AND2_X1 U6983 ( .A1(n4350), .A2(n5235), .ZN(n7723) );
  OR2_X1 U6984 ( .A1(n5581), .A2(n7723), .ZN(n5238) );
  INV_X1 U6985 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10261) );
  OR2_X1 U6986 ( .A1(n5236), .A2(n10261), .ZN(n5237) );
  NAND2_X1 U6987 ( .A1(n8538), .A2(n8970), .ZN(n5853) );
  NAND2_X1 U6988 ( .A1(n7690), .A2(n8537), .ZN(n7709) );
  AND2_X1 U6989 ( .A1(n5853), .A2(n7709), .ZN(n5850) );
  MUX2_X1 U6990 ( .A(n6906), .B(n6908), .S(n6837), .Z(n5256) );
  XNOR2_X1 U6991 ( .A(n5256), .B(SI_12_), .ZN(n5255) );
  NAND2_X1 U6992 ( .A1(n6051), .A2(n5537), .ZN(n5248) );
  NAND2_X1 U6993 ( .A1(n5261), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U6994 ( .A1(n5244), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6728), .B2(
        n5386), .ZN(n5247) );
  NAND2_X1 U6995 ( .A1(n4350), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6996 ( .A1(n5267), .A2(n5250), .ZN(n8976) );
  NAND2_X1 U6997 ( .A1(n5562), .A2(n8976), .ZN(n5254) );
  INV_X1 U6998 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9059) );
  OR2_X1 U6999 ( .A1(n5585), .A2(n9059), .ZN(n5253) );
  INV_X1 U7000 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10170) );
  OR2_X1 U7001 ( .A1(n5759), .A2(n10170), .ZN(n5252) );
  INV_X1 U7002 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6653) );
  OR2_X1 U7003 ( .A1(n5762), .A2(n6653), .ZN(n5251) );
  NAND4_X1 U7004 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n8951)
         );
  XNOR2_X1 U7005 ( .A(n9058), .B(n8951), .ZN(n8972) );
  INV_X1 U7006 ( .A(n8951), .ZN(n8517) );
  OR2_X1 U7007 ( .A1(n9058), .A2(n8517), .ZN(n5856) );
  INV_X1 U7008 ( .A(n5255), .ZN(n5259) );
  INV_X1 U7009 ( .A(n5256), .ZN(n5257) );
  NAND2_X1 U7010 ( .A1(n5257), .A2(SI_12_), .ZN(n5258) );
  MUX2_X1 U7011 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6837), .Z(n5279) );
  XNOR2_X1 U7012 ( .A(n5279), .B(SI_13_), .ZN(n5276) );
  XNOR2_X1 U7013 ( .A(n5278), .B(n5276), .ZN(n6909) );
  NAND2_X1 U7014 ( .A1(n6909), .A2(n5537), .ZN(n5264) );
  NAND2_X1 U7015 ( .A1(n5280), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5262) );
  XNOR2_X1 U7016 ( .A(n5262), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6730) );
  AOI22_X1 U7017 ( .A1(n6730), .A2(n5386), .B1(n5244), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U7018 ( .A1(n5267), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U7019 ( .A1(n5285), .A2(n5268), .ZN(n8957) );
  NAND2_X1 U7020 ( .A1(n5562), .A2(n8957), .ZN(n5272) );
  INV_X1 U7021 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9165) );
  OR2_X1 U7022 ( .A1(n5759), .A2(n9165), .ZN(n5271) );
  INV_X1 U7023 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8962) );
  OR2_X1 U7024 ( .A1(n5762), .A2(n8962), .ZN(n5270) );
  INV_X1 U7025 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10237) );
  OR2_X1 U7026 ( .A1(n5585), .A2(n10237), .ZN(n5269) );
  NAND4_X1 U7027 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n8938)
         );
  INV_X1 U7028 ( .A(n8938), .ZN(n8968) );
  NAND2_X1 U7029 ( .A1(n9166), .A2(n8968), .ZN(n5273) );
  OR2_X1 U7030 ( .A1(n9166), .A2(n8968), .ZN(n5274) );
  INV_X1 U7031 ( .A(n5276), .ZN(n5277) );
  MUX2_X1 U7032 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6837), .Z(n5292) );
  XNOR2_X1 U7033 ( .A(n5292), .B(SI_14_), .ZN(n5289) );
  XNOR2_X1 U7034 ( .A(n5291), .B(n5289), .ZN(n6933) );
  NAND2_X1 U7035 ( .A1(n6933), .A2(n5537), .ZN(n5282) );
  XNOR2_X1 U7036 ( .A(n5316), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6732) );
  AOI22_X1 U7037 ( .A1(n6732), .A2(n5386), .B1(n5244), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5281) );
  INV_X1 U7038 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8944) );
  INV_X1 U7039 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9159) );
  OR2_X1 U7040 ( .A1(n5759), .A2(n9159), .ZN(n5284) );
  INV_X1 U7041 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10262) );
  OR2_X1 U7042 ( .A1(n5585), .A2(n10262), .ZN(n5283) );
  AND2_X1 U7043 ( .A1(n5284), .A2(n5283), .ZN(n5288) );
  NAND2_X1 U7044 ( .A1(n5285), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U7045 ( .A1(n5320), .A2(n5286), .ZN(n8941) );
  NAND2_X1 U7046 ( .A1(n8941), .A2(n5562), .ZN(n5287) );
  INV_X1 U7047 ( .A(n8953), .ZN(n8591) );
  NOR2_X1 U7048 ( .A1(n9160), .A2(n8591), .ZN(n8921) );
  INV_X1 U7049 ( .A(n5289), .ZN(n5290) );
  NAND2_X1 U7050 ( .A1(n5292), .A2(SI_14_), .ZN(n5293) );
  MUX2_X1 U7051 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6837), .Z(n5308) );
  XNOR2_X1 U7052 ( .A(n5308), .B(SI_15_), .ZN(n5294) );
  XNOR2_X1 U7053 ( .A(n5312), .B(n5294), .ZN(n7031) );
  NAND2_X1 U7054 ( .A1(n7031), .A2(n5537), .ZN(n5299) );
  NAND2_X1 U7055 ( .A1(n5316), .A2(n5295), .ZN(n5296) );
  NAND2_X1 U7056 ( .A1(n5296), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5297) );
  XNOR2_X1 U7057 ( .A(n5297), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7033) );
  AOI22_X1 U7058 ( .A1(n7033), .A2(n5386), .B1(n5244), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5298) );
  XNOR2_X1 U7059 ( .A(n5320), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U7060 ( .A1(n8934), .A2(n5562), .ZN(n5304) );
  INV_X1 U7061 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U7062 ( .A1(n5108), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U7063 ( .A1(n5582), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5300) );
  OAI211_X1 U7064 ( .C1(n5585), .C2(n9049), .A(n5301), .B(n5300), .ZN(n5302)
         );
  INV_X1 U7065 ( .A(n5302), .ZN(n5303) );
  INV_X1 U7066 ( .A(n5866), .ZN(n5307) );
  OR2_X1 U7067 ( .A1(n8921), .A2(n5307), .ZN(n5305) );
  NAND2_X1 U7068 ( .A1(n9154), .A2(n8912), .ZN(n5875) );
  NAND2_X1 U7069 ( .A1(n9160), .A2(n8591), .ZN(n8922) );
  AND2_X1 U7070 ( .A1(n5875), .A2(n8922), .ZN(n5306) );
  INV_X1 U7071 ( .A(n5308), .ZN(n5310) );
  INV_X1 U7072 ( .A(SI_15_), .ZN(n5309) );
  NAND2_X1 U7073 ( .A1(n5310), .A2(n5309), .ZN(n5311) );
  MUX2_X1 U7074 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6837), .Z(n5325) );
  INV_X1 U7075 ( .A(SI_16_), .ZN(n5313) );
  XNOR2_X1 U7076 ( .A(n5325), .B(n5313), .ZN(n5314) );
  XNOR2_X1 U7077 ( .A(n5376), .B(n5314), .ZN(n7119) );
  NAND2_X1 U7078 ( .A1(n7119), .A2(n5537), .ZN(n5319) );
  OAI21_X1 U7079 ( .B1(P2_IR_REG_15__SCAN_IN), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U7080 ( .A1(n5316), .A2(n5315), .ZN(n5333) );
  XNOR2_X1 U7081 ( .A(n5333), .B(n5317), .ZN(n6736) );
  AOI22_X1 U7082 ( .A1(n6736), .A2(n5386), .B1(P1_DATAO_REG_16__SCAN_IN), .B2(
        n5244), .ZN(n5318) );
  INV_X1 U7083 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U7084 ( .A1(n5321), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U7085 ( .A1(n5338), .A2(n5322), .ZN(n8917) );
  NAND2_X1 U7086 ( .A1(n8917), .A2(n5562), .ZN(n5324) );
  AOI22_X1 U7087 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n5758), .B1(n5582), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n5323) );
  OAI211_X1 U7088 ( .C1(n5762), .C2(n8916), .A(n5324), .B(n5323), .ZN(n8930)
         );
  INV_X1 U7089 ( .A(n8930), .ZN(n8487) );
  NAND2_X1 U7090 ( .A1(n9148), .A2(n8487), .ZN(n5870) );
  INV_X1 U7091 ( .A(n5624), .ZN(n5874) );
  NOR2_X1 U7092 ( .A1(n5325), .A2(SI_16_), .ZN(n5347) );
  NAND2_X1 U7093 ( .A1(n5325), .A2(SI_16_), .ZN(n5348) );
  NAND2_X1 U7094 ( .A1(n5326), .A2(n5348), .ZN(n5332) );
  INV_X1 U7095 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5327) );
  MUX2_X1 U7096 ( .A(n7264), .B(n5327), .S(n6837), .Z(n5329) );
  NAND2_X1 U7097 ( .A1(n5329), .A2(n5328), .ZN(n5346) );
  INV_X1 U7098 ( .A(n5329), .ZN(n5330) );
  NAND2_X1 U7099 ( .A1(n5330), .A2(SI_17_), .ZN(n5331) );
  NAND2_X1 U7100 ( .A1(n5346), .A2(n5331), .ZN(n5350) );
  XNOR2_X1 U7101 ( .A(n5332), .B(n5350), .ZN(n7174) );
  OAI21_X1 U7102 ( .B1(n5333), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5334) );
  XNOR2_X1 U7103 ( .A(n5334), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6740) );
  AOI22_X1 U7104 ( .A1(n6740), .A2(n5386), .B1(n5244), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U7105 ( .A1(n5338), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U7106 ( .A1(n5361), .A2(n5339), .ZN(n8903) );
  NAND2_X1 U7107 ( .A1(n8903), .A2(n5562), .ZN(n5344) );
  INV_X1 U7108 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U7109 ( .A1(n5108), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U7110 ( .A1(n5582), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5340) );
  OAI211_X1 U7111 ( .C1(n5585), .C2(n9043), .A(n5341), .B(n5340), .ZN(n5342)
         );
  INV_X1 U7112 ( .A(n5342), .ZN(n5343) );
  NAND2_X1 U7113 ( .A1(n5344), .A2(n5343), .ZN(n8889) );
  NAND2_X1 U7114 ( .A1(n8895), .A2(n5877), .ZN(n5345) );
  INV_X1 U7115 ( .A(n5346), .ZN(n5352) );
  OR2_X1 U7116 ( .A1(n5376), .A2(n5369), .ZN(n5353) );
  INV_X1 U7117 ( .A(n5348), .ZN(n5349) );
  NOR2_X1 U7118 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  MUX2_X1 U7119 ( .A(n7253), .B(n5354), .S(n6837), .Z(n5372) );
  XNOR2_X1 U7120 ( .A(n5372), .B(SI_18_), .ZN(n5368) );
  XNOR2_X1 U7121 ( .A(n5355), .B(n5368), .ZN(n7197) );
  NAND2_X1 U7122 ( .A1(n7197), .A2(n5537), .ZN(n5360) );
  NAND2_X1 U7123 ( .A1(n4345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5358) );
  XNOR2_X1 U7124 ( .A(n5358), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8750) );
  AOI22_X1 U7125 ( .A1(n5244), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8750), .B2(
        n5386), .ZN(n5359) );
  NAND2_X1 U7126 ( .A1(n5361), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U7127 ( .A1(n5389), .A2(n5362), .ZN(n8892) );
  NAND2_X1 U7128 ( .A1(n8892), .A2(n5562), .ZN(n5367) );
  INV_X1 U7129 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n10246) );
  NAND2_X1 U7130 ( .A1(n5758), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U7131 ( .A1(n5582), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5363) );
  OAI211_X1 U7132 ( .C1(n5762), .C2(n10246), .A(n5364), .B(n5363), .ZN(n5365)
         );
  INV_X1 U7133 ( .A(n5365), .ZN(n5366) );
  NAND2_X1 U7134 ( .A1(n9136), .A2(n8446), .ZN(n5882) );
  NAND2_X1 U7135 ( .A1(n5879), .A2(n5882), .ZN(n8885) );
  INV_X1 U7136 ( .A(n5372), .ZN(n5373) );
  OAI21_X2 U7137 ( .B1(n5376), .B2(n5375), .A(n5374), .ZN(n5397) );
  MUX2_X1 U7138 ( .A(n7330), .B(n5377), .S(n6837), .Z(n5378) );
  NAND2_X1 U7139 ( .A1(n5378), .A2(n10166), .ZN(n5395) );
  INV_X1 U7140 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U7141 ( .A1(n5379), .A2(SI_19_), .ZN(n5380) );
  NAND2_X1 U7142 ( .A1(n5395), .A2(n5380), .ZN(n5396) );
  XNOR2_X1 U7143 ( .A(n5397), .B(n5396), .ZN(n7327) );
  NAND2_X1 U7144 ( .A1(n7327), .A2(n5537), .ZN(n5388) );
  NAND2_X1 U7145 ( .A1(n5670), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5382) );
  MUX2_X1 U7146 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5382), .S(
        P2_IR_REG_19__SCAN_IN), .Z(n5385) );
  AOI22_X1 U7147 ( .A1(n5244), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6697), .B2(
        n5386), .ZN(n5387) );
  NAND2_X1 U7148 ( .A1(n5389), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U7149 ( .A1(n5402), .A2(n5390), .ZN(n8882) );
  INV_X1 U7150 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U7151 ( .A1(n5108), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U7152 ( .A1(n5582), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5391) );
  OAI211_X1 U7153 ( .C1(n5585), .C2(n9037), .A(n5392), .B(n5391), .ZN(n5393)
         );
  NAND2_X1 U7154 ( .A1(n9130), .A2(n8510), .ZN(n5888) );
  NAND2_X1 U7155 ( .A1(n5889), .A2(n5888), .ZN(n5630) );
  NAND2_X1 U7156 ( .A1(n8876), .A2(n8878), .ZN(n5394) );
  MUX2_X1 U7157 ( .A(n5399), .B(n7438), .S(n6837), .Z(n5432) );
  XNOR2_X1 U7158 ( .A(n5432), .B(SI_20_), .ZN(n5398) );
  XNOR2_X1 U7159 ( .A(n5435), .B(n5398), .ZN(n7413) );
  NAND2_X1 U7160 ( .A1(n7413), .A2(n5537), .ZN(n5401) );
  OR2_X1 U7161 ( .A1(n5060), .A2(n5399), .ZN(n5400) );
  NAND2_X1 U7162 ( .A1(n5402), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U7163 ( .A1(n5443), .A2(n5403), .ZN(n8873) );
  NAND2_X1 U7164 ( .A1(n8873), .A2(n5562), .ZN(n5408) );
  INV_X1 U7165 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U7166 ( .A1(n5582), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U7167 ( .A1(n5758), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5404) );
  OAI211_X1 U7168 ( .C1(n8872), .C2(n5762), .A(n5405), .B(n5404), .ZN(n5406)
         );
  INV_X1 U7169 ( .A(n5406), .ZN(n5407) );
  INV_X1 U7170 ( .A(n5633), .ZN(n8833) );
  MUX2_X1 U7171 ( .A(n7528), .B(n7603), .S(n6837), .Z(n5438) );
  NAND2_X1 U7172 ( .A1(n5438), .A2(n5410), .ZN(n5409) );
  OAI21_X1 U7173 ( .B1(n5413), .B2(SI_20_), .A(n5409), .ZN(n5417) );
  NAND2_X1 U7174 ( .A1(n5413), .A2(SI_20_), .ZN(n5411) );
  NAND2_X1 U7175 ( .A1(n5411), .A2(n5410), .ZN(n5415) );
  INV_X1 U7176 ( .A(n5438), .ZN(n5414) );
  AND2_X1 U7177 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5412) );
  AOI22_X1 U7178 ( .A1(n5415), .A2(n5414), .B1(n5413), .B2(n5412), .ZN(n5416)
         );
  MUX2_X1 U7179 ( .A(n7643), .B(n7640), .S(n6837), .Z(n5419) );
  NAND2_X1 U7180 ( .A1(n5419), .A2(n5418), .ZN(n5455) );
  INV_X1 U7181 ( .A(n5419), .ZN(n5420) );
  NAND2_X1 U7182 ( .A1(n5420), .A2(SI_22_), .ZN(n5421) );
  NAND2_X1 U7183 ( .A1(n5455), .A2(n5421), .ZN(n5456) );
  NAND2_X1 U7184 ( .A1(n7638), .A2(n5537), .ZN(n5423) );
  NAND2_X1 U7185 ( .A1(n5244), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U7186 ( .A1(n5445), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U7187 ( .A1(n5465), .A2(n5426), .ZN(n8849) );
  NAND2_X1 U7188 ( .A1(n8849), .A2(n5562), .ZN(n5431) );
  INV_X1 U7189 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U7190 ( .A1(n5758), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U7191 ( .A1(n5582), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5427) );
  OAI211_X1 U7192 ( .C1(n8848), .C2(n5762), .A(n5428), .B(n5427), .ZN(n5429)
         );
  INV_X1 U7193 ( .A(n5429), .ZN(n5430) );
  XNOR2_X1 U7194 ( .A(n9113), .B(n6258), .ZN(n8836) );
  INV_X1 U7195 ( .A(SI_20_), .ZN(n5434) );
  OR2_X1 U7196 ( .A1(n5435), .A2(n5434), .ZN(n5433) );
  NAND2_X1 U7197 ( .A1(n5433), .A2(n5432), .ZN(n5437) );
  NAND2_X1 U7198 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  NAND2_X1 U7199 ( .A1(n5437), .A2(n5436), .ZN(n5440) );
  XNOR2_X1 U7200 ( .A(n5438), .B(SI_21_), .ZN(n5439) );
  NAND2_X1 U7201 ( .A1(n7527), .A2(n5537), .ZN(n5442) );
  NAND2_X1 U7202 ( .A1(n5244), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U7203 ( .A1(n5443), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U7204 ( .A1(n5445), .A2(n5444), .ZN(n8864) );
  NAND2_X1 U7205 ( .A1(n8864), .A2(n5562), .ZN(n5450) );
  INV_X1 U7206 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U7207 ( .A1(n5758), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U7208 ( .A1(n5108), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5446) );
  OAI211_X1 U7209 ( .C1(n5759), .C2(n10218), .A(n5447), .B(n5446), .ZN(n5448)
         );
  INV_X1 U7210 ( .A(n5448), .ZN(n5449) );
  NOR2_X1 U7211 ( .A1(n8836), .A2(n8835), .ZN(n5452) );
  OR2_X1 U7212 ( .A1(n8833), .A2(n5452), .ZN(n5454) );
  NAND2_X1 U7213 ( .A1(n9118), .A2(n6255), .ZN(n5896) );
  NAND2_X1 U7214 ( .A1(n9124), .A2(n8455), .ZN(n8852) );
  AND2_X1 U7215 ( .A1(n5896), .A2(n8852), .ZN(n8834) );
  INV_X1 U7216 ( .A(n8836), .ZN(n8843) );
  AND2_X1 U7217 ( .A1(n8834), .A2(n8843), .ZN(n5451) );
  MUX2_X1 U7218 ( .A(n5458), .B(n7646), .S(n6837), .Z(n5460) );
  INV_X1 U7219 ( .A(SI_23_), .ZN(n5459) );
  NAND2_X1 U7220 ( .A1(n5460), .A2(n5459), .ZN(n5474) );
  INV_X1 U7221 ( .A(n5460), .ZN(n5461) );
  NAND2_X1 U7222 ( .A1(n5461), .A2(SI_23_), .ZN(n5462) );
  XNOR2_X1 U7223 ( .A(n5473), .B(n5472), .ZN(n7644) );
  NAND2_X1 U7224 ( .A1(n7644), .A2(n5537), .ZN(n5464) );
  NAND2_X1 U7225 ( .A1(n5244), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U7226 ( .A1(n5465), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7227 ( .A1(n5484), .A2(n5466), .ZN(n8829) );
  NAND2_X1 U7228 ( .A1(n8829), .A2(n5562), .ZN(n5471) );
  INV_X1 U7229 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10206) );
  NAND2_X1 U7230 ( .A1(n5758), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U7231 ( .A1(n5108), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5467) );
  OAI211_X1 U7232 ( .C1(n5759), .C2(n10206), .A(n5468), .B(n5467), .ZN(n5469)
         );
  INV_X1 U7233 ( .A(n5469), .ZN(n5470) );
  INV_X1 U7234 ( .A(n8846), .ZN(n8528) );
  OR2_X1 U7235 ( .A1(n9113), .A2(n6258), .ZN(n8810) );
  AND2_X1 U7236 ( .A1(n8812), .A2(n8810), .ZN(n5901) );
  NAND2_X1 U7237 ( .A1(n5475), .A2(n5474), .ZN(n5494) );
  MUX2_X1 U7238 ( .A(n7826), .B(n7760), .S(n6837), .Z(n5477) );
  NAND2_X1 U7239 ( .A1(n5477), .A2(n5476), .ZN(n5495) );
  INV_X1 U7240 ( .A(n5477), .ZN(n5478) );
  NAND2_X1 U7241 ( .A1(n5478), .A2(SI_24_), .ZN(n5479) );
  XNOR2_X1 U7242 ( .A(n5494), .B(n5493), .ZN(n7759) );
  NAND2_X1 U7243 ( .A1(n7759), .A2(n5537), .ZN(n5481) );
  NAND2_X1 U7244 ( .A1(n5244), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5480) );
  INV_X1 U7245 ( .A(n5484), .ZN(n5483) );
  INV_X1 U7246 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U7247 ( .A1(n5484), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U7248 ( .A1(n5504), .A2(n5485), .ZN(n8820) );
  NAND2_X1 U7249 ( .A1(n8820), .A2(n5562), .ZN(n5491) );
  INV_X1 U7250 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7251 ( .A1(n5582), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7252 ( .A1(n5758), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5486) );
  OAI211_X1 U7253 ( .C1(n5488), .C2(n5762), .A(n5487), .B(n5486), .ZN(n5489)
         );
  INV_X1 U7254 ( .A(n5489), .ZN(n5490) );
  NAND2_X1 U7255 ( .A1(n9102), .A2(n8427), .ZN(n5907) );
  NAND2_X1 U7256 ( .A1(n9107), .A2(n8528), .ZN(n5899) );
  NAND2_X1 U7257 ( .A1(n5907), .A2(n5899), .ZN(n5904) );
  NAND2_X1 U7258 ( .A1(n5904), .A2(n5905), .ZN(n5492) );
  MUX2_X1 U7259 ( .A(n7850), .B(n7829), .S(n6837), .Z(n5497) );
  INV_X1 U7260 ( .A(SI_25_), .ZN(n5496) );
  NAND2_X1 U7261 ( .A1(n5497), .A2(n5496), .ZN(n5514) );
  INV_X1 U7262 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U7263 ( .A1(n5498), .A2(SI_25_), .ZN(n5499) );
  XNOR2_X1 U7264 ( .A(n5513), .B(n5512), .ZN(n7828) );
  NAND2_X1 U7265 ( .A1(n7828), .A2(n5537), .ZN(n5501) );
  NAND2_X1 U7266 ( .A1(n5244), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5500) );
  INV_X1 U7267 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7268 ( .A1(n5504), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7269 ( .A1(n5521), .A2(n5505), .ZN(n8807) );
  NAND2_X1 U7270 ( .A1(n8807), .A2(n5562), .ZN(n5510) );
  INV_X1 U7271 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10167) );
  NAND2_X1 U7272 ( .A1(n5758), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7273 ( .A1(n5108), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5506) );
  OAI211_X1 U7274 ( .C1(n5759), .C2(n10167), .A(n5507), .B(n5506), .ZN(n5508)
         );
  INV_X1 U7275 ( .A(n5508), .ZN(n5509) );
  NAND2_X1 U7276 ( .A1(n6300), .A2(n6315), .ZN(n5910) );
  NAND2_X1 U7277 ( .A1(n5511), .A2(n5909), .ZN(n8781) );
  MUX2_X1 U7278 ( .A(n7848), .B(n7853), .S(n6837), .Z(n5516) );
  INV_X1 U7279 ( .A(SI_26_), .ZN(n5515) );
  NAND2_X1 U7280 ( .A1(n5516), .A2(n5515), .ZN(n5530) );
  INV_X1 U7281 ( .A(n5516), .ZN(n5517) );
  NAND2_X1 U7282 ( .A1(n5517), .A2(SI_26_), .ZN(n5518) );
  XNOR2_X1 U7283 ( .A(n5529), .B(n5528), .ZN(n7847) );
  NAND2_X1 U7284 ( .A1(n7847), .A2(n5537), .ZN(n5520) );
  NAND2_X1 U7285 ( .A1(n5244), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7286 ( .A1(n5521), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7287 ( .A1(n5540), .A2(n5522), .ZN(n8789) );
  NAND2_X1 U7288 ( .A1(n8789), .A2(n5562), .ZN(n5527) );
  INV_X1 U7289 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8788) );
  NAND2_X1 U7290 ( .A1(n5758), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7291 ( .A1(n5582), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5523) );
  OAI211_X1 U7292 ( .C1(n8788), .C2(n5762), .A(n5524), .B(n5523), .ZN(n5525)
         );
  INV_X1 U7293 ( .A(n5525), .ZN(n5526) );
  NOR2_X1 U7294 ( .A1(n9090), .A2(n8092), .ZN(n5915) );
  NAND2_X1 U7295 ( .A1(n9090), .A2(n8092), .ZN(n5916) );
  NAND2_X1 U7296 ( .A1(n5529), .A2(n5528), .ZN(n5531) );
  INV_X1 U7297 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5532) );
  MUX2_X1 U7298 ( .A(n5532), .B(n9865), .S(n6837), .Z(n5534) );
  INV_X1 U7299 ( .A(SI_27_), .ZN(n5533) );
  NAND2_X1 U7300 ( .A1(n5534), .A2(n5533), .ZN(n5550) );
  INV_X1 U7301 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U7302 ( .A1(n5535), .A2(SI_27_), .ZN(n5536) );
  XNOR2_X1 U7303 ( .A(n5549), .B(n5548), .ZN(n7856) );
  NAND2_X1 U7304 ( .A1(n7856), .A2(n5537), .ZN(n5539) );
  NAND2_X1 U7305 ( .A1(n5244), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7306 ( .A1(n5540), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7307 ( .A1(n5560), .A2(n5541), .ZN(n8778) );
  NAND2_X1 U7308 ( .A1(n8778), .A2(n5562), .ZN(n5546) );
  INV_X1 U7309 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U7310 ( .A1(n5758), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7311 ( .A1(n5582), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5542) );
  OAI211_X1 U7312 ( .C1(n8777), .C2(n5762), .A(n5543), .B(n5542), .ZN(n5544)
         );
  INV_X1 U7313 ( .A(n5544), .ZN(n5545) );
  XNOR2_X1 U7314 ( .A(n9084), .B(n8786), .ZN(n8770) );
  INV_X1 U7315 ( .A(n8770), .ZN(n8768) );
  OR2_X1 U7316 ( .A1(n9084), .A2(n8576), .ZN(n5547) );
  INV_X1 U7317 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5551) );
  INV_X1 U7318 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8389) );
  MUX2_X1 U7319 ( .A(n5551), .B(n8389), .S(n6837), .Z(n5553) );
  INV_X1 U7320 ( .A(SI_28_), .ZN(n5552) );
  NAND2_X1 U7321 ( .A1(n5553), .A2(n5552), .ZN(n5573) );
  INV_X1 U7322 ( .A(n5553), .ZN(n5554) );
  NAND2_X1 U7323 ( .A1(n5554), .A2(SI_28_), .ZN(n5555) );
  NAND2_X1 U7324 ( .A1(n8388), .A2(n5537), .ZN(n5557) );
  NAND2_X1 U7325 ( .A1(n5244), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5556) );
  INV_X1 U7326 ( .A(n5560), .ZN(n5559) );
  INV_X1 U7327 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7328 ( .A1(n5559), .A2(n5558), .ZN(n8390) );
  NAND2_X1 U7329 ( .A1(n5560), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7330 ( .A1(n8390), .A2(n5561), .ZN(n8760) );
  NAND2_X1 U7331 ( .A1(n8760), .A2(n5562), .ZN(n5567) );
  INV_X1 U7332 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U7333 ( .A1(n5108), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7334 ( .A1(n5582), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5563) );
  OAI211_X1 U7335 ( .C1(n5585), .C2(n10259), .A(n5564), .B(n5563), .ZN(n5565)
         );
  INV_X1 U7336 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7337 ( .A1(n5952), .A2(n5953), .ZN(n5568) );
  INV_X1 U7338 ( .A(n8774), .ZN(n5933) );
  OR2_X1 U7339 ( .A1(n8410), .A2(n5933), .ZN(n5928) );
  INV_X1 U7340 ( .A(n5573), .ZN(n5571) );
  MUX2_X1 U7341 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6837), .Z(n5739) );
  XNOR2_X1 U7342 ( .A(n5739), .B(SI_29_), .ZN(n5575) );
  OAI21_X1 U7343 ( .B1(n5572), .B2(n5571), .A(n5575), .ZN(n5577) );
  OR2_X1 U7344 ( .A1(n8398), .A2(n5578), .ZN(n5580) );
  INV_X1 U7345 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8397) );
  OR2_X1 U7346 ( .A1(n5060), .A2(n8397), .ZN(n5579) );
  NAND2_X1 U7347 ( .A1(n5580), .A2(n5579), .ZN(n8391) );
  INV_X1 U7348 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7349 ( .A1(n5108), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7350 ( .A1(n5582), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5583) );
  OAI211_X1 U7351 ( .C1(n5586), .C2(n5585), .A(n5584), .B(n5583), .ZN(n5587)
         );
  INV_X1 U7352 ( .A(n5587), .ZN(n5588) );
  NAND2_X1 U7353 ( .A1(n5765), .A2(n5588), .ZN(n8599) );
  INV_X1 U7354 ( .A(n8599), .ZN(n5955) );
  OR2_X1 U7355 ( .A1(n8391), .A2(n5955), .ZN(n5775) );
  NAND2_X1 U7356 ( .A1(n8391), .A2(n5955), .ZN(n5935) );
  NAND2_X1 U7357 ( .A1(n5775), .A2(n5935), .ZN(n5927) );
  XNOR2_X1 U7358 ( .A(n5757), .B(n5927), .ZN(n8393) );
  XNOR2_X2 U7359 ( .A(n5591), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7360 ( .A1(n5589), .A2(n5592), .ZN(n5593) );
  NAND2_X1 U7361 ( .A1(n5596), .A2(n5589), .ZN(n5597) );
  NAND2_X1 U7362 ( .A1(n7414), .A2(n7328), .ZN(n5691) );
  NAND2_X1 U7363 ( .A1(n7036), .A2(n7641), .ZN(n5710) );
  NAND3_X1 U7364 ( .A1(n6986), .A2(n7328), .A3(n5710), .ZN(n7687) );
  NAND2_X1 U7365 ( .A1(n7641), .A2(n6192), .ZN(n7103) );
  NAND2_X1 U7366 ( .A1(n8393), .A2(n7501), .ZN(n5669) );
  INV_X1 U7367 ( .A(n7216), .ZN(n6991) );
  NAND2_X1 U7368 ( .A1(n8610), .A2(n6991), .ZN(n7042) );
  NAND2_X1 U7369 ( .A1(n7037), .A2(n7042), .ZN(n5602) );
  OR2_X1 U7370 ( .A1(n8609), .A2(n6196), .ZN(n5601) );
  NAND3_X1 U7371 ( .A1(n5604), .A2(n6955), .A3(n7112), .ZN(n5606) );
  NOR2_X1 U7372 ( .A1(n8608), .A2(n9001), .ZN(n7111) );
  NOR2_X1 U7373 ( .A1(n8607), .A2(n7222), .ZN(n5603) );
  INV_X1 U7374 ( .A(n7153), .ZN(n7312) );
  OR2_X1 U7375 ( .A1(n7204), .A2(n8606), .ZN(n5607) );
  NAND2_X1 U7376 ( .A1(n9068), .A2(n8605), .ZN(n5608) );
  INV_X1 U7377 ( .A(n7700), .ZN(n8604) );
  AND2_X1 U7378 ( .A1(n7631), .A2(n8604), .ZN(n5609) );
  NOR2_X1 U7379 ( .A1(n7701), .A2(n8603), .ZN(n5610) );
  NAND2_X1 U7380 ( .A1(n7701), .A2(n8603), .ZN(n7579) );
  INV_X1 U7381 ( .A(n8462), .ZN(n5612) );
  OR2_X1 U7382 ( .A1(n7690), .A2(n8601), .ZN(n5614) );
  NAND2_X1 U7383 ( .A1(n8502), .A2(n8602), .ZN(n7680) );
  NAND2_X1 U7384 ( .A1(n7690), .A2(n8601), .ZN(n5611) );
  INV_X1 U7385 ( .A(n8970), .ZN(n8600) );
  NAND2_X1 U7386 ( .A1(n8538), .A2(n8600), .ZN(n6222) );
  INV_X1 U7387 ( .A(n6222), .ZN(n5617) );
  OR2_X1 U7388 ( .A1(n8502), .A2(n8602), .ZN(n7679) );
  AND2_X1 U7389 ( .A1(n7679), .A2(n5614), .ZN(n7711) );
  AND2_X1 U7390 ( .A1(n9058), .A2(n8951), .ZN(n5620) );
  NAND2_X1 U7391 ( .A1(n9166), .A2(n8938), .ZN(n5858) );
  NAND2_X1 U7392 ( .A1(n8948), .A2(n5858), .ZN(n5621) );
  OR2_X1 U7393 ( .A1(n9166), .A2(n8938), .ZN(n5862) );
  NAND2_X1 U7394 ( .A1(n5621), .A2(n5862), .ZN(n8937) );
  NAND2_X1 U7395 ( .A1(n9160), .A2(n8953), .ZN(n5622) );
  OR2_X1 U7396 ( .A1(n9160), .A2(n8953), .ZN(n5623) );
  INV_X1 U7397 ( .A(n8906), .ZN(n8910) );
  AND2_X1 U7398 ( .A1(n9154), .A2(n8939), .ZN(n8909) );
  AOI22_X1 U7399 ( .A1(n8910), .A2(n8909), .B1(n9148), .B2(n8930), .ZN(n5625)
         );
  NAND2_X1 U7400 ( .A1(n9142), .A2(n8889), .ZN(n5627) );
  OR2_X1 U7401 ( .A1(n9136), .A2(n8899), .ZN(n5628) );
  NAND2_X1 U7402 ( .A1(n9136), .A2(n8899), .ZN(n5629) );
  INV_X1 U7403 ( .A(n8510), .ZN(n8890) );
  NAND2_X1 U7404 ( .A1(n9130), .A2(n8890), .ZN(n5631) );
  NAND2_X1 U7405 ( .A1(n8835), .A2(n5896), .ZN(n8854) );
  INV_X1 U7406 ( .A(n8854), .ZN(n8858) );
  NOR2_X1 U7407 ( .A1(n9124), .A2(n8879), .ZN(n8856) );
  NOR2_X1 U7408 ( .A1(n9118), .A2(n8870), .ZN(n8841) );
  AOI21_X1 U7409 ( .B1(n8856), .B2(n8854), .A(n8841), .ZN(n5634) );
  OR2_X1 U7410 ( .A1(n9113), .A2(n8861), .ZN(n5635) );
  NAND2_X1 U7411 ( .A1(n9107), .A2(n8846), .ZN(n5636) );
  NAND2_X1 U7412 ( .A1(n8824), .A2(n5636), .ZN(n5638) );
  OR2_X1 U7413 ( .A1(n9107), .A2(n8846), .ZN(n5637) );
  NOR2_X1 U7414 ( .A1(n9102), .A2(n8826), .ZN(n8794) );
  NAND2_X1 U7415 ( .A1(n9090), .A2(n8803), .ZN(n5640) );
  INV_X1 U7416 ( .A(n8798), .ZN(n5639) );
  NAND2_X1 U7417 ( .A1(n9102), .A2(n8826), .ZN(n8796) );
  AND2_X1 U7418 ( .A1(n5639), .A2(n8796), .ZN(n8795) );
  OR2_X1 U7419 ( .A1(n4987), .A2(n8795), .ZN(n8782) );
  AND2_X1 U7420 ( .A1(n5640), .A2(n8782), .ZN(n5641) );
  OR2_X1 U7421 ( .A1(n9090), .A2(n8803), .ZN(n5642) );
  NAND2_X1 U7422 ( .A1(n9084), .A2(n8786), .ZN(n5644) );
  OR2_X1 U7423 ( .A1(n8410), .A2(n8774), .ZN(n5649) );
  AND2_X1 U7424 ( .A1(n5927), .A2(n5649), .ZN(n5651) );
  AND2_X1 U7425 ( .A1(n8410), .A2(n8774), .ZN(n5652) );
  NAND2_X1 U7426 ( .A1(n5927), .A2(n5652), .ZN(n5648) );
  INV_X1 U7427 ( .A(n7414), .ZN(n5645) );
  NAND2_X1 U7428 ( .A1(n6191), .A2(n5645), .ZN(n5647) );
  NAND2_X1 U7429 ( .A1(n5949), .A2(n6697), .ZN(n5646) );
  INV_X2 U7430 ( .A(n8967), .ZN(n8949) );
  OAI211_X1 U7431 ( .C1(n5927), .C2(n5649), .A(n5648), .B(n8949), .ZN(n5650)
         );
  INV_X1 U7432 ( .A(n5954), .ZN(n5655) );
  INV_X1 U7433 ( .A(n5652), .ZN(n5654) );
  INV_X1 U7434 ( .A(n5927), .ZN(n5653) );
  NAND3_X1 U7435 ( .A1(n5655), .A2(n5654), .A3(n5653), .ZN(n5667) );
  INV_X1 U7436 ( .A(n6754), .ZN(n6750) );
  INV_X1 U7437 ( .A(n6753), .ZN(n6743) );
  NAND2_X1 U7438 ( .A1(n6750), .A2(n6743), .ZN(n5657) );
  INV_X1 U7439 ( .A(n6276), .ZN(n6294) );
  OR2_X1 U7440 ( .A1(n6634), .A2(n6294), .ZN(n8971) );
  INV_X1 U7441 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7442 ( .A1(n5758), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5660) );
  INV_X1 U7443 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n5658) );
  OR2_X1 U7444 ( .A1(n5759), .A2(n5658), .ZN(n5659) );
  OAI211_X1 U7445 ( .C1(n5661), .C2(n5762), .A(n5660), .B(n5659), .ZN(n5662)
         );
  INV_X1 U7446 ( .A(n5662), .ZN(n5663) );
  NAND2_X1 U7447 ( .A1(n5765), .A2(n5663), .ZN(n8598) );
  AND2_X1 U7448 ( .A1(n6636), .A2(P2_B_REG_SCAN_IN), .ZN(n5664) );
  NOR2_X1 U7449 ( .A1(n8969), .A2(n5664), .ZN(n8751) );
  AOI22_X1 U7450 ( .A1(n8774), .A2(n8952), .B1(n8598), .B2(n8751), .ZN(n5665)
         );
  AOI21_X2 U7451 ( .B1(n5667), .B2(n5668), .A(n5666), .ZN(n8396) );
  INV_X1 U7452 ( .A(n5675), .ZN(n5674) );
  NAND2_X1 U7453 ( .A1(n5674), .A2(n5673), .ZN(n5677) );
  NAND2_X1 U7454 ( .A1(n5675), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7455 ( .A1(n5677), .A2(n5676), .ZN(n5686) );
  XNOR2_X1 U7456 ( .A(n5686), .B(P2_B_REG_SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7457 ( .A1(n5677), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5679) );
  XNOR2_X1 U7458 ( .A(n5679), .B(n5678), .ZN(n5688) );
  NAND2_X1 U7459 ( .A1(n5680), .A2(n5688), .ZN(n5687) );
  OAI21_X1 U7460 ( .B1(n4345), .B2(n5682), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5683) );
  MUX2_X1 U7461 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5683), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5684) );
  NOR2_X1 U7462 ( .A1(n7849), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7463 ( .A1(n5703), .A2(n7849), .ZN(n6193) );
  NAND2_X1 U7464 ( .A1(n6195), .A2(n6193), .ZN(n5723) );
  NAND2_X1 U7465 ( .A1(n8112), .A2(n7849), .ZN(n5689) );
  INV_X1 U7466 ( .A(n5691), .ZN(n5944) );
  INV_X1 U7467 ( .A(n6282), .ZN(n5709) );
  NOR2_X1 U7468 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5695) );
  NOR4_X1 U7469 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5694) );
  NOR4_X1 U7470 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5693) );
  NOR4_X1 U7471 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5692) );
  NAND4_X1 U7472 ( .A1(n5695), .A2(n5694), .A3(n5693), .A4(n5692), .ZN(n5701)
         );
  NOR4_X1 U7473 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5699) );
  NOR4_X1 U7474 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5698) );
  NOR4_X1 U7475 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5697) );
  NOR4_X1 U7476 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5696) );
  NAND4_X1 U7477 ( .A1(n5699), .A2(n5698), .A3(n5697), .A4(n5696), .ZN(n5700)
         );
  NOR2_X1 U7478 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  INV_X1 U7479 ( .A(n8112), .ZN(n5705) );
  NOR2_X1 U7480 ( .A1(n5703), .A2(n7849), .ZN(n5704) );
  NOR2_X1 U7481 ( .A1(n7414), .A2(n6697), .ZN(n5799) );
  NAND2_X1 U7482 ( .A1(n5710), .A2(n5799), .ZN(n5711) );
  NAND2_X1 U7483 ( .A1(n5722), .A2(n5713), .ZN(n6982) );
  INV_X1 U7484 ( .A(n6192), .ZN(n5712) );
  INV_X1 U7485 ( .A(n6302), .ZN(n5715) );
  INV_X1 U7486 ( .A(n5713), .ZN(n5714) );
  NAND2_X1 U7487 ( .A1(n5723), .A2(n5714), .ZN(n6983) );
  NAND2_X1 U7488 ( .A1(n5731), .A2(n4313), .ZN(n5721) );
  NOR2_X1 U7489 ( .A1(n4313), .A2(n5586), .ZN(n5719) );
  NAND2_X1 U7490 ( .A1(n5721), .A2(n5720), .ZN(P2_U3488) );
  NOR2_X1 U7491 ( .A1(n6981), .A2(n5725), .ZN(n6279) );
  NAND2_X1 U7492 ( .A1(n6279), .A2(n6892), .ZN(n6301) );
  NOR2_X1 U7493 ( .A1(n7414), .A2(n7328), .ZN(n5797) );
  NAND3_X1 U7494 ( .A1(n7529), .A2(n5797), .A3(n5949), .ZN(n6284) );
  AND2_X1 U7495 ( .A1(n6986), .A2(n6284), .ZN(n5724) );
  INV_X1 U7496 ( .A(n5725), .ZN(n5726) );
  NAND3_X1 U7497 ( .A1(n6284), .A2(n6634), .A3(n7407), .ZN(n6273) );
  NAND2_X1 U7498 ( .A1(n6273), .A2(n8817), .ZN(n6280) );
  INV_X1 U7499 ( .A(n6280), .ZN(n5728) );
  INV_X2 U7500 ( .A(n10292), .ZN(n5734) );
  NAND2_X1 U7501 ( .A1(n5731), .A2(n5734), .ZN(n5738) );
  INV_X1 U7502 ( .A(n8391), .ZN(n5732) );
  INV_X1 U7503 ( .A(n7407), .ZN(n9069) );
  INV_X1 U7504 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5733) );
  NOR2_X1 U7505 ( .A1(n5734), .A2(n5733), .ZN(n5735) );
  NAND2_X1 U7506 ( .A1(n5738), .A2(n5737), .ZN(P2_U3456) );
  INV_X1 U7507 ( .A(n5775), .ZN(n5756) );
  NOR2_X1 U7508 ( .A1(n5739), .A2(SI_29_), .ZN(n5741) );
  NAND2_X1 U7509 ( .A1(n5739), .A2(SI_29_), .ZN(n5740) );
  INV_X1 U7510 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8380) );
  INV_X1 U7511 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8386) );
  MUX2_X1 U7512 ( .A(n8380), .B(n8386), .S(n6840), .Z(n5744) );
  INV_X1 U7513 ( .A(SI_30_), .ZN(n5743) );
  NAND2_X1 U7514 ( .A1(n5744), .A2(n5743), .ZN(n5748) );
  INV_X1 U7515 ( .A(n5744), .ZN(n5745) );
  NAND2_X1 U7516 ( .A1(n5745), .A2(SI_30_), .ZN(n5746) );
  NAND2_X1 U7517 ( .A1(n5748), .A2(n5746), .ZN(n5749) );
  NOR2_X1 U7518 ( .A1(n5060), .A2(n8386), .ZN(n5747) );
  INV_X1 U7519 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9856) );
  INV_X1 U7520 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9177) );
  MUX2_X1 U7521 ( .A(n9856), .B(n9177), .S(n6840), .Z(n5751) );
  XNOR2_X1 U7522 ( .A(n5751), .B(SI_31_), .ZN(n5752) );
  NAND2_X1 U7523 ( .A1(n9860), .A2(n5537), .ZN(n5755) );
  OR2_X1 U7524 ( .A1(n5060), .A2(n9177), .ZN(n5754) );
  OAI22_X1 U7525 ( .A1(n5757), .A2(n5756), .B1(n9081), .B2(n9075), .ZN(n5772)
         );
  INV_X1 U7526 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U7527 ( .A1(n5758), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5761) );
  INV_X1 U7528 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9078) );
  OR2_X1 U7529 ( .A1(n5759), .A2(n9078), .ZN(n5760) );
  OAI211_X1 U7530 ( .C1(n8756), .C2(n5762), .A(n5761), .B(n5760), .ZN(n5763)
         );
  INV_X1 U7531 ( .A(n5763), .ZN(n5764) );
  NOR2_X1 U7532 ( .A1(n9075), .A2(n8753), .ZN(n5940) );
  INV_X1 U7533 ( .A(n5940), .ZN(n5770) );
  INV_X1 U7534 ( .A(n9081), .ZN(n5767) );
  INV_X1 U7535 ( .A(n8598), .ZN(n5766) );
  AND2_X1 U7536 ( .A1(n5767), .A2(n5766), .ZN(n5939) );
  INV_X1 U7537 ( .A(n5939), .ZN(n5768) );
  AND2_X1 U7538 ( .A1(n5768), .A2(n5935), .ZN(n5769) );
  NAND2_X1 U7539 ( .A1(n5770), .A2(n5769), .ZN(n5796) );
  AND2_X1 U7540 ( .A1(n9081), .A2(n8598), .ZN(n5922) );
  OAI21_X1 U7541 ( .B1(n5922), .B2(n8753), .A(n9075), .ZN(n5771) );
  INV_X1 U7542 ( .A(n5774), .ZN(n5773) );
  NAND2_X1 U7543 ( .A1(n5773), .A2(n4995), .ZN(n5804) );
  AND2_X1 U7544 ( .A1(n8753), .A2(n9075), .ZN(n5942) );
  INV_X1 U7545 ( .A(n5922), .ZN(n5776) );
  AND2_X1 U7546 ( .A1(n5776), .A2(n5775), .ZN(n5926) );
  INV_X1 U7547 ( .A(n5926), .ZN(n5938) );
  INV_X1 U7548 ( .A(n5916), .ZN(n5777) );
  NAND2_X1 U7549 ( .A1(n5905), .A2(n5907), .ZN(n8814) );
  INV_X1 U7550 ( .A(n8885), .ZN(n8887) );
  INV_X1 U7551 ( .A(n8922), .ZN(n5778) );
  NAND2_X1 U7552 ( .A1(n5862), .A2(n5858), .ZN(n8960) );
  NAND2_X1 U7553 ( .A1(n8610), .A2(n7216), .ZN(n5805) );
  NOR2_X1 U7554 ( .A1(n4433), .A2(n7218), .ZN(n5780) );
  AND2_X1 U7555 ( .A1(n5833), .A2(n5822), .ZN(n7166) );
  NAND4_X1 U7556 ( .A1(n5779), .A2(n7113), .A3(n5780), .A4(n7166), .ZN(n5781)
         );
  NAND2_X1 U7557 ( .A1(n7379), .A2(n5836), .ZN(n7367) );
  NOR2_X1 U7558 ( .A1(n5781), .A2(n7367), .ZN(n5782) );
  XNOR2_X1 U7559 ( .A(n7204), .B(n8606), .ZN(n7151) );
  NAND3_X1 U7560 ( .A1(n7385), .A2(n5782), .A3(n7151), .ZN(n5783) );
  INV_X1 U7561 ( .A(n7709), .ZN(n5830) );
  OR2_X1 U7562 ( .A1(n5849), .A2(n5830), .ZN(n7678) );
  NAND2_X1 U7563 ( .A1(n5826), .A2(n5825), .ZN(n7457) );
  OR4_X1 U7564 ( .A1(n5783), .A2(n7678), .A3(n7581), .A4(n7457), .ZN(n5784) );
  NOR2_X1 U7565 ( .A1(n5784), .A2(n8462), .ZN(n5785) );
  NAND3_X1 U7566 ( .A1(n8960), .A2(n5785), .A3(n8972), .ZN(n5786) );
  NOR2_X1 U7567 ( .A1(n8943), .A2(n5786), .ZN(n5787) );
  NAND3_X1 U7568 ( .A1(n8906), .A2(n8926), .A3(n5787), .ZN(n5788) );
  NOR2_X1 U7569 ( .A1(n8897), .A2(n5788), .ZN(n5789) );
  NAND4_X1 U7570 ( .A1(n8868), .A2(n8878), .A3(n8887), .A4(n5789), .ZN(n5790)
         );
  NOR2_X1 U7571 ( .A1(n8854), .A2(n5790), .ZN(n5791) );
  NAND3_X1 U7572 ( .A1(n8825), .A2(n5791), .A3(n8843), .ZN(n5792) );
  NOR2_X1 U7573 ( .A1(n8814), .A2(n5792), .ZN(n5793) );
  NAND2_X1 U7574 ( .A1(n8798), .A2(n5793), .ZN(n5794) );
  NOR2_X1 U7575 ( .A1(n8784), .A2(n5794), .ZN(n5795) );
  INV_X1 U7576 ( .A(n5800), .ZN(n5798) );
  NAND3_X1 U7577 ( .A1(n5798), .A2(n5797), .A3(n7529), .ZN(n5802) );
  NAND3_X1 U7578 ( .A1(n5800), .A2(n5799), .A3(n7529), .ZN(n5801) );
  INV_X4 U7579 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U7580 ( .A1(n6748), .A2(P2_U3151), .ZN(n7604) );
  NAND3_X1 U7581 ( .A1(n5804), .A2(n5803), .A3(n4989), .ZN(n5951) );
  INV_X1 U7582 ( .A(n6634), .ZN(n5925) );
  MUX2_X1 U7583 ( .A(n8938), .B(n9166), .S(n5925), .Z(n5857) );
  INV_X1 U7584 ( .A(n5857), .ZN(n5863) );
  NAND3_X1 U7585 ( .A1(n5828), .A2(n6634), .A3(n5825), .ZN(n5847) );
  INV_X1 U7586 ( .A(n5805), .ZN(n5806) );
  NAND2_X1 U7587 ( .A1(n5808), .A2(n5807), .ZN(n5811) );
  INV_X1 U7588 ( .A(n5811), .ZN(n5809) );
  NOR2_X1 U7589 ( .A1(n5809), .A2(n7112), .ZN(n5814) );
  NOR3_X1 U7590 ( .A1(n7218), .A2(n5810), .A3(n6191), .ZN(n5812) );
  NOR3_X1 U7591 ( .A1(n5812), .A2(n7112), .A3(n5811), .ZN(n5813) );
  MUX2_X1 U7592 ( .A(n5814), .B(n5813), .S(n6634), .Z(n5820) );
  NAND2_X1 U7593 ( .A1(n5832), .A2(n5815), .ZN(n5818) );
  NAND2_X1 U7594 ( .A1(n5821), .A2(n5816), .ZN(n5817) );
  MUX2_X1 U7595 ( .A(n5818), .B(n5817), .S(n6634), .Z(n5819) );
  INV_X1 U7596 ( .A(n7385), .ZN(n5837) );
  NAND3_X1 U7597 ( .A1(n5841), .A2(n5925), .A3(n5826), .ZN(n5827) );
  NAND2_X1 U7598 ( .A1(n5847), .A2(n5827), .ZN(n5843) );
  INV_X1 U7599 ( .A(n5828), .ZN(n5829) );
  AOI211_X1 U7600 ( .C1(n5831), .C2(n5843), .A(n5830), .B(n5829), .ZN(n5846)
         );
  INV_X1 U7601 ( .A(n5832), .ZN(n5834) );
  OAI211_X1 U7602 ( .C1(n5835), .C2(n5834), .A(n7365), .B(n5833), .ZN(n5840)
         );
  INV_X1 U7603 ( .A(n5836), .ZN(n5838) );
  AOI211_X1 U7604 ( .C1(n5840), .C2(n5839), .A(n5838), .B(n5837), .ZN(n5844)
         );
  INV_X1 U7605 ( .A(n5841), .ZN(n5842) );
  AOI211_X1 U7606 ( .C1(n5844), .C2(n5843), .A(n5849), .B(n5842), .ZN(n5845)
         );
  NOR2_X1 U7607 ( .A1(n4787), .A2(n5849), .ZN(n5851) );
  MUX2_X1 U7608 ( .A(n5851), .B(n5850), .S(n6634), .Z(n5852) );
  MUX2_X1 U7609 ( .A(n5853), .B(n6223), .S(n6634), .Z(n5854) );
  NAND2_X1 U7610 ( .A1(n9058), .A2(n8517), .ZN(n5855) );
  MUX2_X1 U7611 ( .A(n5856), .B(n5855), .S(n6634), .Z(n5859) );
  AOI22_X1 U7612 ( .A1(n5860), .A2(n5859), .B1(n5858), .B2(n5857), .ZN(n5861)
         );
  INV_X1 U7613 ( .A(n8921), .ZN(n5864) );
  MUX2_X1 U7614 ( .A(n5864), .B(n8922), .S(n6634), .Z(n5865) );
  NAND2_X1 U7615 ( .A1(n5868), .A2(n5867), .ZN(n5873) );
  INV_X1 U7616 ( .A(n8897), .ZN(n5872) );
  OAI211_X1 U7617 ( .C1(n8897), .C2(n5870), .A(n5882), .B(n5869), .ZN(n5871)
         );
  AOI211_X1 U7618 ( .C1(n5876), .C2(n5875), .A(n5925), .B(n5874), .ZN(n5878)
         );
  OAI211_X1 U7619 ( .C1(n5885), .C2(n5878), .A(n5879), .B(n5877), .ZN(n5887)
         );
  INV_X1 U7620 ( .A(n5879), .ZN(n5880) );
  NAND2_X1 U7621 ( .A1(n5881), .A2(n5889), .ZN(n5884) );
  NAND2_X1 U7622 ( .A1(n8852), .A2(n5888), .ZN(n5891) );
  NAND2_X1 U7623 ( .A1(n8868), .A2(n5889), .ZN(n5890) );
  MUX2_X1 U7624 ( .A(n5891), .B(n5890), .S(n6634), .Z(n5895) );
  INV_X1 U7625 ( .A(n8835), .ZN(n5892) );
  NOR2_X1 U7626 ( .A1(n5892), .A2(n8833), .ZN(n5893) );
  MUX2_X1 U7627 ( .A(n5893), .B(n8834), .S(n6634), .Z(n5894) );
  MUX2_X1 U7628 ( .A(n5896), .B(n8835), .S(n6634), .Z(n5897) );
  INV_X1 U7629 ( .A(n5897), .ZN(n5898) );
  INV_X1 U7630 ( .A(n5899), .ZN(n8811) );
  AOI21_X1 U7631 ( .B1(n6258), .B2(n9113), .A(n8811), .ZN(n5900) );
  MUX2_X1 U7632 ( .A(n5901), .B(n5900), .S(n6634), .Z(n5902) );
  OAI21_X1 U7633 ( .B1(n5906), .B2(n5904), .A(n5905), .ZN(n5908) );
  INV_X1 U7634 ( .A(n5909), .ZN(n5912) );
  INV_X1 U7635 ( .A(n5910), .ZN(n5911) );
  MUX2_X1 U7636 ( .A(n5912), .B(n5911), .S(n6634), .Z(n5913) );
  INV_X1 U7637 ( .A(n5915), .ZN(n5917) );
  MUX2_X1 U7638 ( .A(n5917), .B(n5916), .S(n6634), .Z(n5918) );
  NAND2_X1 U7639 ( .A1(n8786), .A2(n6634), .ZN(n5920) );
  NAND2_X1 U7640 ( .A1(n8576), .A2(n5925), .ZN(n5919) );
  MUX2_X1 U7641 ( .A(n5920), .B(n5919), .S(n9084), .Z(n5921) );
  NOR2_X1 U7642 ( .A1(n5922), .A2(n5925), .ZN(n5934) );
  NAND2_X1 U7643 ( .A1(n5934), .A2(n5928), .ZN(n5923) );
  OAI211_X1 U7644 ( .C1(n5928), .C2(n5927), .A(n5926), .B(n5925), .ZN(n5929)
         );
  NAND2_X1 U7645 ( .A1(n5930), .A2(n5929), .ZN(n5931) );
  NAND2_X1 U7646 ( .A1(n8410), .A2(n5933), .ZN(n5937) );
  INV_X1 U7647 ( .A(n5934), .ZN(n5936) );
  OAI22_X1 U7648 ( .A1(n5938), .A2(n5937), .B1(n5936), .B2(n5935), .ZN(n5941)
         );
  NOR3_X1 U7649 ( .A1(n5941), .A2(n5940), .A3(n5939), .ZN(n5943) );
  NAND2_X1 U7650 ( .A1(n5945), .A2(n6192), .ZN(n5946) );
  INV_X1 U7651 ( .A(n7604), .ZN(n5948) );
  NOR2_X1 U7652 ( .A1(n6303), .A2(n6986), .ZN(n6290) );
  NAND3_X1 U7653 ( .A1(n6290), .A2(n6750), .A3(n6753), .ZN(n5947) );
  OAI211_X1 U7654 ( .C1(n5949), .C2(n5948), .A(n5947), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5950) );
  XOR2_X1 U7655 ( .A(n5952), .B(n5953), .Z(n8765) );
  INV_X1 U7656 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5960) );
  NAND4_X1 U7657 ( .A1(n6124), .A2(n5963), .A3(n6147), .A4(n6166), .ZN(n5966)
         );
  NAND2_X1 U7658 ( .A1(n6148), .A2(n5964), .ZN(n5965) );
  NOR2_X2 U7659 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  NAND2_X1 U7660 ( .A1(n6154), .A2(n5968), .ZN(n5969) );
  NAND2_X1 U7661 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5971) );
  AOI22_X1 U7662 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(n6020), .B1(n5971), .B2(
        P1_IR_REG_31__SCAN_IN), .ZN(n5972) );
  NOR2_X1 U7663 ( .A1(n6134), .A2(n5972), .ZN(n5973) );
  OAI21_X2 U7664 ( .B1(n5974), .B2(n4983), .A(n5973), .ZN(n9862) );
  NAND2_X2 U7665 ( .A1(n5982), .A2(n9862), .ZN(n5993) );
  NAND2_X2 U7666 ( .A1(n5993), .A2(n6837), .ZN(n6008) );
  INV_X1 U7667 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8097) );
  OR2_X1 U7668 ( .A1(n6122), .A2(n8097), .ZN(n5975) );
  INV_X1 U7669 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7670 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5976) );
  OR2_X1 U7671 ( .A1(n6017), .A2(n7007), .ZN(n5986) );
  NAND2_X1 U7672 ( .A1(n6851), .A2(n6837), .ZN(n5980) );
  NOR2_X1 U7673 ( .A1(n6837), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5978) );
  NOR2_X1 U7674 ( .A1(n9862), .A2(n5978), .ZN(n5979) );
  MUX2_X1 U7675 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n5981), .S(n6837), .Z(n5983)
         );
  INV_X1 U7676 ( .A(n4319), .ZN(n7025) );
  NAND2_X1 U7677 ( .A1(n5983), .A2(n7025), .ZN(n5984) );
  NAND3_X1 U7678 ( .A1(n5986), .A2(n5985), .A3(n5984), .ZN(n6363) );
  NAND2_X1 U7679 ( .A1(n6837), .A2(SI_0_), .ZN(n5988) );
  INV_X1 U7680 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7681 ( .A1(n5988), .A2(n5987), .ZN(n5990) );
  AND2_X1 U7682 ( .A1(n5990), .A2(n5989), .ZN(n9867) );
  NAND2_X1 U7683 ( .A1(n6017), .A2(n9867), .ZN(n5991) );
  INV_X1 U7684 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5997) );
  INV_X1 U7685 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5998) );
  OR2_X1 U7686 ( .A1(n6017), .A2(n7871), .ZN(n6000) );
  OR2_X1 U7687 ( .A1(n6008), .A2(n7873), .ZN(n5999) );
  OR2_X1 U7688 ( .A1(n6003), .A2(n6020), .ZN(n6004) );
  NAND2_X1 U7689 ( .A1(n6005), .A2(n6004), .ZN(n6011) );
  XNOR2_X1 U7690 ( .A(n6011), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7094) );
  INV_X1 U7691 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7692 ( .A1(n6122), .A2(n6006), .ZN(n6010) );
  OR2_X1 U7693 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  OR2_X1 U7694 ( .A1(n6122), .A2(n6857), .ZN(n6016) );
  OAI21_X1 U7695 ( .B1(n6011), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6013) );
  INV_X1 U7696 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6012) );
  XNOR2_X1 U7697 ( .A(n6013), .B(n6012), .ZN(n7015) );
  INV_X2 U7698 ( .A(n10011), .ZN(n8129) );
  INV_X2 U7699 ( .A(n6008), .ZN(n6058) );
  NAND2_X1 U7700 ( .A1(n6847), .A2(n6058), .ZN(n6023) );
  INV_X1 U7701 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6020) );
  OR2_X1 U7702 ( .A1(n6019), .A2(n6020), .ZN(n6021) );
  XNOR2_X1 U7703 ( .A(n6021), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9448) );
  AOI22_X1 U7704 ( .A1(n6100), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6871), .B2(
        n9448), .ZN(n6022) );
  NAND2_X1 U7705 ( .A1(n6019), .A2(n6024), .ZN(n6026) );
  NAND2_X1 U7706 ( .A1(n6026), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6025) );
  MUX2_X1 U7707 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6025), .S(
        P1_IR_REG_7__SCAN_IN), .Z(n6027) );
  AOI22_X1 U7708 ( .A1(n6100), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6871), .B2(
        n9461), .ZN(n6028) );
  NAND2_X1 U7709 ( .A1(n6065), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6030) );
  XNOR2_X1 U7710 ( .A(n6030), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9474) );
  AOI22_X1 U7711 ( .A1(n6100), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6871), .B2(
        n9474), .ZN(n6029) );
  INV_X1 U7712 ( .A(n10039), .ZN(n7758) );
  NAND2_X1 U7713 ( .A1(n6869), .A2(n6058), .ZN(n6034) );
  NAND2_X1 U7714 ( .A1(n6030), .A2(n6035), .ZN(n6031) );
  NAND2_X1 U7715 ( .A1(n6031), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6032) );
  XNOR2_X1 U7716 ( .A(n6032), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7242) );
  AOI22_X1 U7717 ( .A1(n6100), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6871), .B2(
        n7242), .ZN(n6033) );
  NAND2_X1 U7718 ( .A1(n6034), .A2(n6033), .ZN(n9299) );
  INV_X1 U7719 ( .A(n9299), .ZN(n7656) );
  NAND2_X1 U7720 ( .A1(n6858), .A2(n6058), .ZN(n6043) );
  INV_X1 U7721 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7722 ( .A1(n6036), .A2(n6035), .ZN(n6037) );
  NAND2_X1 U7723 ( .A1(n6040), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6038) );
  MUX2_X1 U7724 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6038), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n6039) );
  INV_X1 U7725 ( .A(n6039), .ZN(n6041) );
  AOI22_X1 U7726 ( .A1(n6100), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6871), .B2(
        n7415), .ZN(n6042) );
  NAND2_X1 U7727 ( .A1(n6043), .A2(n6042), .ZN(n9831) );
  INV_X1 U7728 ( .A(n9831), .ZN(n7795) );
  NAND2_X1 U7729 ( .A1(n6887), .A2(n6058), .ZN(n6050) );
  INV_X1 U7730 ( .A(n6045), .ZN(n6047) );
  NAND2_X1 U7731 ( .A1(n6047), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6046) );
  MUX2_X1 U7732 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6046), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n6048) );
  AOI22_X1 U7733 ( .A1(n6100), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6871), .B2(
        n7517), .ZN(n6049) );
  NAND2_X1 U7734 ( .A1(n6051), .A2(n6058), .ZN(n6056) );
  NAND2_X1 U7735 ( .A1(n6052), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7736 ( .A1(n6053), .A2(n10247), .ZN(n6059) );
  OR2_X1 U7737 ( .A1(n6053), .A2(n10247), .ZN(n6054) );
  AOI22_X1 U7738 ( .A1(n6100), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6871), .B2(
        n9489), .ZN(n6055) );
  NAND2_X1 U7739 ( .A1(n6909), .A2(n6058), .ZN(n6062) );
  NAND2_X1 U7740 ( .A1(n6059), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6060) );
  AOI22_X1 U7741 ( .A1(n6100), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6871), .B2(
        n9501), .ZN(n6061) );
  NAND2_X1 U7742 ( .A1(n6933), .A2(n6058), .ZN(n6068) );
  INV_X1 U7743 ( .A(n6063), .ZN(n6064) );
  OAI21_X1 U7744 ( .B1(n6065), .B2(n6064), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6066) );
  XNOR2_X1 U7745 ( .A(n6066), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9927) );
  AOI22_X1 U7746 ( .A1(n6100), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4464), .B2(
        n9927), .ZN(n6067) );
  INV_X1 U7747 ( .A(n9815), .ZN(n7842) );
  NAND2_X1 U7748 ( .A1(n7536), .A2(n7842), .ZN(n7819) );
  NAND2_X1 U7749 ( .A1(n7031), .A2(n6058), .ZN(n6074) );
  NAND2_X1 U7750 ( .A1(n6069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6070) );
  MUX2_X1 U7751 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6070), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6072) );
  NAND2_X1 U7752 ( .A1(n6072), .A2(n6075), .ZN(n9505) );
  INV_X1 U7753 ( .A(n9505), .ZN(n9940) );
  AOI22_X1 U7754 ( .A1(n6100), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6871), .B2(
        n9940), .ZN(n6073) );
  OR2_X2 U7755 ( .A1(n7819), .A2(n9811), .ZN(n7865) );
  NAND2_X1 U7756 ( .A1(n7119), .A2(n6058), .ZN(n6078) );
  NAND2_X1 U7757 ( .A1(n6075), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6076) );
  XNOR2_X1 U7758 ( .A(n6076), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9522) );
  AOI22_X1 U7759 ( .A1(n6100), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4464), .B2(
        n9522), .ZN(n6077) );
  NOR2_X4 U7760 ( .A1(n7865), .A2(n9803), .ZN(n9723) );
  NAND2_X1 U7761 ( .A1(n7174), .A2(n6058), .ZN(n6082) );
  NAND2_X1 U7762 ( .A1(n6126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6083) );
  XNOR2_X1 U7763 ( .A(n6083), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9540) );
  AOI22_X1 U7764 ( .A1(n6100), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4464), .B2(
        n9540), .ZN(n6081) );
  INV_X1 U7765 ( .A(n9798), .ZN(n9728) );
  NAND2_X1 U7766 ( .A1(n7197), .A2(n6058), .ZN(n6089) );
  NAND2_X1 U7767 ( .A1(n6083), .A2(n6123), .ZN(n6092) );
  NAND2_X1 U7768 ( .A1(n6092), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6085) );
  INV_X1 U7769 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6084) );
  OR2_X1 U7770 ( .A1(n6085), .A2(n6084), .ZN(n6087) );
  NAND2_X1 U7771 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  AOI22_X1 U7772 ( .A1(n6100), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6871), .B2(
        n9948), .ZN(n6088) );
  INV_X1 U7773 ( .A(n9794), .ZN(n9719) );
  NAND2_X1 U7774 ( .A1(n7327), .A2(n6058), .ZN(n6102) );
  AND2_X1 U7775 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6090) );
  NAND2_X1 U7776 ( .A1(n6092), .A2(n6090), .ZN(n6099) );
  INV_X1 U7777 ( .A(n6124), .ZN(n6091) );
  NAND2_X1 U7778 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n6093) );
  NOR2_X1 U7779 ( .A1(n6097), .A2(n6096), .ZN(n6098) );
  INV_X1 U7780 ( .A(n9550), .ZN(n6772) );
  AOI22_X1 U7781 ( .A1(n6100), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6772), .B2(
        n4464), .ZN(n6101) );
  NAND2_X1 U7782 ( .A1(n7413), .A2(n6058), .ZN(n6104) );
  OR2_X1 U7783 ( .A1(n6122), .A2(n7438), .ZN(n6103) );
  NAND2_X1 U7784 ( .A1(n7527), .A2(n6058), .ZN(n6106) );
  OR2_X1 U7785 ( .A1(n6122), .A2(n7603), .ZN(n6105) );
  NAND2_X2 U7786 ( .A1(n6106), .A2(n6105), .ZN(n9778) );
  NAND2_X1 U7787 ( .A1(n7638), .A2(n6058), .ZN(n6108) );
  OR2_X1 U7788 ( .A1(n6122), .A2(n7640), .ZN(n6107) );
  INV_X1 U7789 ( .A(n9773), .ZN(n9645) );
  NAND2_X1 U7790 ( .A1(n7644), .A2(n6058), .ZN(n6110) );
  OR2_X1 U7791 ( .A1(n6122), .A2(n7646), .ZN(n6109) );
  INV_X1 U7792 ( .A(n9769), .ZN(n9625) );
  NAND2_X1 U7793 ( .A1(n7759), .A2(n6058), .ZN(n6112) );
  OR2_X1 U7794 ( .A1(n6122), .A2(n7760), .ZN(n6111) );
  NAND2_X1 U7795 ( .A1(n7828), .A2(n6058), .ZN(n6114) );
  OR2_X1 U7796 ( .A1(n6122), .A2(n7829), .ZN(n6113) );
  NAND2_X1 U7797 ( .A1(n7847), .A2(n6058), .ZN(n6116) );
  OR2_X1 U7798 ( .A1(n6122), .A2(n7853), .ZN(n6115) );
  NAND2_X1 U7799 ( .A1(n7856), .A2(n6058), .ZN(n6118) );
  OR2_X1 U7800 ( .A1(n6122), .A2(n9865), .ZN(n6117) );
  OR2_X2 U7801 ( .A1(n7876), .A2(n9748), .ZN(n9577) );
  NAND2_X1 U7802 ( .A1(n8388), .A2(n6058), .ZN(n6120) );
  OR2_X1 U7803 ( .A1(n6122), .A2(n8389), .ZN(n6119) );
  NAND2_X1 U7804 ( .A1(n9569), .A2(n9576), .ZN(n6570) );
  INV_X1 U7805 ( .A(n6570), .ZN(n9557) );
  OR2_X1 U7806 ( .A1(n6122), .A2(n8380), .ZN(n6121) );
  NAND2_X1 U7807 ( .A1(n9557), .A2(n9740), .ZN(n9556) );
  NAND2_X1 U7808 ( .A1(n6124), .A2(n6123), .ZN(n6125) );
  XNOR2_X2 U7809 ( .A(n6164), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8375) );
  INV_X1 U7810 ( .A(n8375), .ZN(n7639) );
  NAND2_X1 U7811 ( .A1(n6149), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7812 ( .A1(n6137), .A2(n4531), .ZN(n6136) );
  NAND2_X1 U7813 ( .A1(n4316), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7814 ( .A1(n6561), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7815 ( .A1(n6498), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6140) );
  NAND3_X1 U7816 ( .A1(n6142), .A2(n6141), .A3(n6140), .ZN(n8348) );
  INV_X1 U7817 ( .A(P1_B_REG_SCAN_IN), .ZN(n6143) );
  NOR2_X1 U7818 ( .A1(n9862), .A2(n6143), .ZN(n6144) );
  NOR2_X1 U7819 ( .A1(n9712), .A2(n6144), .ZN(n6564) );
  NAND2_X1 U7820 ( .A1(n8348), .A2(n6564), .ZN(n9738) );
  INV_X1 U7821 ( .A(n6145), .ZN(n6146) );
  NAND2_X1 U7822 ( .A1(n9555), .A2(n6146), .ZN(n9737) );
  MUX2_X1 U7823 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6150), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6152) );
  NAND2_X1 U7824 ( .A1(n6152), .A2(n6151), .ZN(n7761) );
  INV_X1 U7825 ( .A(n7761), .ZN(n6162) );
  INV_X1 U7826 ( .A(n6156), .ZN(n6155) );
  NAND2_X1 U7827 ( .A1(n6155), .A2(n6154), .ZN(n6158) );
  NAND2_X1 U7828 ( .A1(n6158), .A2(n6157), .ZN(n6171) );
  NAND2_X1 U7829 ( .A1(n6151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6160) );
  NOR2_X1 U7830 ( .A1(n6171), .A2(n7830), .ZN(n6161) );
  NAND2_X2 U7831 ( .A1(n6162), .A2(n6161), .ZN(n6821) );
  NAND2_X1 U7832 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7833 ( .A1(n6165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7834 ( .A1(n7290), .A2(n7292), .ZN(n6169) );
  NAND2_X1 U7835 ( .A1(n7830), .A2(P1_B_REG_SCAN_IN), .ZN(n6170) );
  MUX2_X1 U7836 ( .A(P1_B_REG_SCAN_IN), .B(n6170), .S(n7761), .Z(n6173) );
  INV_X1 U7837 ( .A(n7855), .ZN(n6172) );
  NOR4_X1 U7838 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6182) );
  NOR4_X1 U7839 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6181) );
  NOR4_X1 U7840 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6177) );
  NOR4_X1 U7841 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6176) );
  NOR4_X1 U7842 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6175) );
  NOR4_X1 U7843 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6174) );
  NAND4_X1 U7844 ( .A1(n6177), .A2(n6176), .A3(n6175), .A4(n6174), .ZN(n6178)
         );
  NOR4_X1 U7845 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6179), .A4(n6178), .ZN(n6180) );
  AND3_X1 U7846 ( .A1(n6182), .A2(n6181), .A3(n6180), .ZN(n7289) );
  INV_X1 U7847 ( .A(n6860), .ZN(n6185) );
  INV_X1 U7848 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6184) );
  INV_X1 U7849 ( .A(n7295), .ZN(n6186) );
  NAND2_X1 U7850 ( .A1(n7761), .A2(n7855), .ZN(n9855) );
  OR2_X1 U7851 ( .A1(n10055), .A2(n6188), .ZN(n6189) );
  OAI21_X1 U7852 ( .B1(n6192), .B2(n6191), .A(n7036), .ZN(n6194) );
  INV_X2 U7853 ( .A(n6205), .ZN(n8399) );
  INV_X4 U7854 ( .A(n8399), .ZN(n8461) );
  XNOR2_X1 U7855 ( .A(n8461), .B(n7204), .ZN(n6209) );
  INV_X1 U7856 ( .A(n6209), .ZN(n6210) );
  NOR2_X1 U7857 ( .A1(n6199), .A2(n6198), .ZN(n7143) );
  OAI21_X1 U7858 ( .B1(n8399), .B2(n6991), .A(n7038), .ZN(n7142) );
  INV_X1 U7859 ( .A(n6199), .ZN(n6200) );
  NAND2_X1 U7860 ( .A1(n7141), .A2(n6200), .ZN(n7209) );
  XNOR2_X1 U7861 ( .A(n9001), .B(n6205), .ZN(n6201) );
  XOR2_X1 U7862 ( .A(n8608), .B(n6201), .Z(n7210) );
  NAND2_X1 U7863 ( .A1(n7209), .A2(n7210), .ZN(n7208) );
  INV_X1 U7864 ( .A(n6201), .ZN(n6203) );
  NAND2_X1 U7865 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  NAND2_X1 U7866 ( .A1(n7208), .A2(n6204), .ZN(n7225) );
  XNOR2_X1 U7867 ( .A(n6205), .B(n7222), .ZN(n6206) );
  XNOR2_X1 U7868 ( .A(n6206), .B(n8607), .ZN(n7226) );
  XNOR2_X1 U7869 ( .A(n8461), .B(n7170), .ZN(n6207) );
  NOR2_X1 U7870 ( .A1(n6207), .A2(n7153), .ZN(n6208) );
  AOI21_X1 U7871 ( .B1(n7153), .B2(n6207), .A(n6208), .ZN(n7231) );
  INV_X1 U7872 ( .A(n6208), .ZN(n7307) );
  XNOR2_X1 U7873 ( .A(n6209), .B(n8606), .ZN(n7306) );
  AOI21_X1 U7874 ( .B1(n6210), .B2(n7370), .A(n7310), .ZN(n8560) );
  XNOR2_X1 U7875 ( .A(n9068), .B(n8461), .ZN(n6211) );
  XOR2_X1 U7876 ( .A(n8605), .B(n6211), .Z(n8559) );
  XNOR2_X1 U7877 ( .A(n7631), .B(n8399), .ZN(n6214) );
  NAND2_X1 U7878 ( .A1(n6214), .A2(n7700), .ZN(n7694) );
  OAI21_X1 U7879 ( .B1(n6214), .B2(n7700), .A(n7694), .ZN(n7627) );
  NAND2_X1 U7880 ( .A1(n7695), .A2(n7694), .ZN(n6217) );
  XNOR2_X1 U7881 ( .A(n7701), .B(n8461), .ZN(n6218) );
  XNOR2_X1 U7882 ( .A(n6218), .B(n8603), .ZN(n7693) );
  INV_X1 U7883 ( .A(n7693), .ZN(n6216) );
  INV_X1 U7884 ( .A(n6218), .ZN(n6219) );
  NAND2_X1 U7885 ( .A1(n6219), .A2(n5163), .ZN(n6220) );
  XNOR2_X1 U7886 ( .A(n8502), .B(n8461), .ZN(n6221) );
  XNOR2_X1 U7887 ( .A(n6221), .B(n8602), .ZN(n8499) );
  XNOR2_X1 U7888 ( .A(n7690), .B(n8399), .ZN(n8433) );
  MUX2_X1 U7889 ( .A(n6223), .B(n6222), .S(n8461), .Z(n8463) );
  OAI21_X1 U7890 ( .B1(n8537), .B2(n8433), .A(n8463), .ZN(n6230) );
  AND2_X1 U7891 ( .A1(n6222), .A2(n8461), .ZN(n6228) );
  NAND3_X1 U7892 ( .A1(n8462), .A2(n8399), .A3(n6223), .ZN(n6226) );
  INV_X1 U7893 ( .A(n7690), .ZN(n9066) );
  NAND4_X1 U7894 ( .A1(n6222), .A2(n8537), .A3(n9066), .A4(n8461), .ZN(n6225)
         );
  NAND4_X1 U7895 ( .A1(n6223), .A2(n8537), .A3(n8399), .A4(n7690), .ZN(n6224)
         );
  NAND3_X1 U7896 ( .A1(n6226), .A2(n6225), .A3(n6224), .ZN(n6227) );
  XNOR2_X1 U7897 ( .A(n9058), .B(n8461), .ZN(n6231) );
  NOR2_X1 U7898 ( .A1(n6231), .A2(n8951), .ZN(n8466) );
  AOI211_X1 U7899 ( .C1(n5612), .C2(n6228), .A(n6227), .B(n8466), .ZN(n6229)
         );
  OAI21_X1 U7900 ( .B1(n8431), .B2(n6230), .A(n6229), .ZN(n6232) );
  NAND2_X1 U7901 ( .A1(n6231), .A2(n8951), .ZN(n8464) );
  XNOR2_X1 U7902 ( .A(n9166), .B(n8461), .ZN(n6233) );
  XNOR2_X1 U7903 ( .A(n6233), .B(n8938), .ZN(n8515) );
  XNOR2_X1 U7904 ( .A(n9160), .B(n8461), .ZN(n6234) );
  XOR2_X1 U7905 ( .A(n8953), .B(n6234), .Z(n8415) );
  INV_X1 U7906 ( .A(n6234), .ZN(n6235) );
  NAND2_X1 U7907 ( .A1(n6235), .A2(n8591), .ZN(n6236) );
  XNOR2_X1 U7908 ( .A(n9154), .B(n8461), .ZN(n6238) );
  XNOR2_X1 U7909 ( .A(n6238), .B(n8939), .ZN(n8582) );
  NAND2_X1 U7910 ( .A1(n6238), .A2(n8939), .ZN(n6239) );
  XNOR2_X1 U7911 ( .A(n9148), .B(n8461), .ZN(n6240) );
  XOR2_X1 U7912 ( .A(n8930), .B(n6240), .Z(n8477) );
  NAND2_X1 U7913 ( .A1(n6240), .A2(n8930), .ZN(n6241) );
  XNOR2_X1 U7914 ( .A(n9142), .B(n8461), .ZN(n6242) );
  XNOR2_X1 U7915 ( .A(n6242), .B(n8889), .ZN(n8485) );
  XNOR2_X1 U7916 ( .A(n9136), .B(n8399), .ZN(n6245) );
  XNOR2_X1 U7917 ( .A(n6245), .B(n8899), .ZN(n8547) );
  INV_X1 U7918 ( .A(n8547), .ZN(n6244) );
  INV_X1 U7919 ( .A(n6242), .ZN(n6243) );
  NAND2_X1 U7920 ( .A1(n6243), .A2(n8913), .ZN(n8546) );
  OR2_X1 U7921 ( .A1(n6244), .A2(n8546), .ZN(n8549) );
  NAND2_X1 U7922 ( .A1(n6245), .A2(n8446), .ZN(n6246) );
  AND2_X1 U7923 ( .A1(n8549), .A2(n6246), .ZN(n6247) );
  XNOR2_X1 U7924 ( .A(n9130), .B(n8461), .ZN(n6248) );
  XNOR2_X1 U7925 ( .A(n6248), .B(n8510), .ZN(n8443) );
  INV_X1 U7926 ( .A(n6248), .ZN(n6249) );
  NAND2_X1 U7927 ( .A1(n6249), .A2(n8510), .ZN(n8504) );
  XNOR2_X1 U7928 ( .A(n9124), .B(n8461), .ZN(n6252) );
  INV_X1 U7929 ( .A(n6252), .ZN(n6250) );
  NAND2_X1 U7930 ( .A1(n6250), .A2(n8455), .ZN(n6251) );
  INV_X1 U7931 ( .A(n6251), .ZN(n6253) );
  XOR2_X1 U7932 ( .A(n8879), .B(n6252), .Z(n8507) );
  XNOR2_X1 U7933 ( .A(n9118), .B(n8461), .ZN(n6254) );
  XOR2_X1 U7934 ( .A(n8870), .B(n6254), .Z(n8452) );
  INV_X1 U7935 ( .A(n6254), .ZN(n6256) );
  XNOR2_X1 U7936 ( .A(n9113), .B(n8461), .ZN(n6257) );
  NAND2_X1 U7937 ( .A1(n6257), .A2(n8861), .ZN(n8523) );
  INV_X1 U7938 ( .A(n6257), .ZN(n6259) );
  NAND2_X1 U7939 ( .A1(n6259), .A2(n6258), .ZN(n8524) );
  NAND2_X2 U7940 ( .A1(n6260), .A2(n8524), .ZN(n8083) );
  INV_X1 U7941 ( .A(n8083), .ZN(n6262) );
  XNOR2_X1 U7942 ( .A(n9107), .B(n8461), .ZN(n6307) );
  NOR2_X1 U7943 ( .A1(n6307), .A2(n8846), .ZN(n8078) );
  INV_X1 U7944 ( .A(n8078), .ZN(n6261) );
  NAND2_X1 U7945 ( .A1(n6262), .A2(n6261), .ZN(n6272) );
  XNOR2_X1 U7946 ( .A(n9102), .B(n8399), .ZN(n6263) );
  NAND2_X1 U7947 ( .A1(n6263), .A2(n8427), .ZN(n6269) );
  OAI21_X1 U7948 ( .B1(n6263), .B2(n8427), .A(n6269), .ZN(n6309) );
  AOI21_X1 U7949 ( .B1(n8846), .B2(n6307), .A(n6309), .ZN(n6267) );
  XNOR2_X1 U7950 ( .A(n6300), .B(n8399), .ZN(n6264) );
  NAND2_X1 U7951 ( .A1(n6264), .A2(n6315), .ZN(n8567) );
  INV_X1 U7952 ( .A(n6264), .ZN(n6265) );
  NAND2_X1 U7953 ( .A1(n6265), .A2(n8815), .ZN(n6266) );
  AND2_X1 U7954 ( .A1(n6267), .A2(n6268), .ZN(n8079) );
  INV_X1 U7955 ( .A(n6268), .ZN(n6270) );
  INV_X1 U7956 ( .A(n8077), .ZN(n6271) );
  OR2_X1 U7957 ( .A1(n6301), .A2(n6273), .ZN(n6275) );
  OR2_X1 U7958 ( .A1(n6296), .A2(n6284), .ZN(n6274) );
  INV_X1 U7959 ( .A(n6296), .ZN(n6278) );
  NOR2_X1 U7960 ( .A1(n6986), .A2(n6276), .ZN(n6277) );
  INV_X1 U7961 ( .A(n8807), .ZN(n6298) );
  INV_X1 U7962 ( .A(n6279), .ZN(n6281) );
  NAND2_X1 U7963 ( .A1(n6281), .A2(n6280), .ZN(n6288) );
  AND2_X1 U7964 ( .A1(n6282), .A2(n6748), .ZN(n6287) );
  INV_X1 U7965 ( .A(n6283), .ZN(n6291) );
  INV_X1 U7966 ( .A(n6284), .ZN(n6285) );
  NAND2_X1 U7967 ( .A1(n6291), .A2(n6285), .ZN(n6286) );
  NAND4_X1 U7968 ( .A1(n6288), .A2(n6287), .A3(n6749), .A4(n6286), .ZN(n6289)
         );
  NAND2_X1 U7969 ( .A1(n6289), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7970 ( .A1(n6291), .A2(n6290), .ZN(n6292) );
  INV_X1 U7971 ( .A(n8593), .ZN(n7318) );
  OR2_X1 U7972 ( .A1(n6986), .A2(n6294), .ZN(n6295) );
  AOI22_X1 U7973 ( .A1(n8826), .A2(n8572), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n6297) );
  OAI21_X1 U7974 ( .B1(n6298), .B2(n7318), .A(n6297), .ZN(n6299) );
  AOI21_X1 U7975 ( .B1(n8587), .B2(n8803), .A(n6299), .ZN(n6305) );
  OR2_X1 U7976 ( .A1(n6301), .A2(n7407), .ZN(n6304) );
  NAND3_X1 U7977 ( .A1(n6306), .A2(n6305), .A3(n4409), .ZN(P2_U3165) );
  INV_X1 U7978 ( .A(n6307), .ZN(n6308) );
  OAI21_X1 U7979 ( .B1(n8083), .B2(n6308), .A(n6310), .ZN(n8422) );
  NOR2_X1 U7980 ( .A1(n8423), .A2(n6311), .ZN(n6313) );
  INV_X1 U7981 ( .A(n9102), .ZN(n8818) );
  AOI22_X1 U7982 ( .A1(n8846), .A2(n8572), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n6314) );
  OAI21_X1 U7983 ( .B1(n6315), .B2(n8575), .A(n6314), .ZN(n6316) );
  AOI21_X1 U7984 ( .B1(n8820), .B2(n8593), .A(n6316), .ZN(n6317) );
  INV_X1 U7985 ( .A(n6318), .ZN(n6319) );
  NAND2_X1 U7986 ( .A1(n6320), .A2(n6319), .ZN(P2_U3169) );
  NAND2_X1 U7987 ( .A1(n6498), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7988 ( .A1(n4316), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6330) );
  INV_X1 U7989 ( .A(n6391), .ZN(n6322) );
  NAND2_X1 U7990 ( .A1(n6322), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6393) );
  INV_X1 U7991 ( .A(n6393), .ZN(n6324) );
  NAND2_X1 U7992 ( .A1(n6324), .A2(n6323), .ZN(n6341) );
  INV_X1 U7993 ( .A(n6341), .ZN(n6325) );
  NAND2_X1 U7994 ( .A1(n6334), .A2(n6326), .ZN(n6327) );
  AND2_X1 U7995 ( .A1(n6356), .A2(n6327), .ZN(n9286) );
  NAND2_X1 U7996 ( .A1(n6551), .A2(n9286), .ZN(n6329) );
  NAND2_X1 U7997 ( .A1(n4315), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6328) );
  OR2_X1 U7998 ( .A1(n9299), .A2(n7790), .ZN(n8165) );
  NAND2_X1 U7999 ( .A1(n6498), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6338) );
  INV_X1 U8000 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U8001 ( .A1(n6341), .A2(n6332), .ZN(n6333) );
  AND2_X1 U8002 ( .A1(n6334), .A2(n6333), .ZN(n7554) );
  NAND2_X1 U8003 ( .A1(n6551), .A2(n7554), .ZN(n6336) );
  NAND2_X1 U8004 ( .A1(n4315), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6335) );
  INV_X1 U8005 ( .A(n9399), .ZN(n6353) );
  NAND2_X1 U8006 ( .A1(n4316), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U8007 ( .A1(n6498), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6344) );
  INV_X1 U8008 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7662) );
  INV_X1 U8009 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6339) );
  OAI21_X1 U8010 ( .B1(n6393), .B2(n7662), .A(n6339), .ZN(n6340) );
  AND2_X1 U8011 ( .A1(n6341), .A2(n6340), .ZN(n7481) );
  NAND2_X1 U8012 ( .A1(n6551), .A2(n7481), .ZN(n6343) );
  NAND2_X1 U8013 ( .A1(n4314), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6342) );
  OR2_X1 U8014 ( .A1(n7753), .A2(n10029), .ZN(n8147) );
  INV_X1 U8015 ( .A(n8147), .ZN(n6351) );
  NAND2_X1 U8016 ( .A1(n4317), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8017 ( .A1(n4314), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6347) );
  XNOR2_X1 U8018 ( .A(n6393), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U8019 ( .A1(n6394), .A2(n9964), .ZN(n6346) );
  NAND3_X1 U8020 ( .A1(n6348), .A2(n6347), .A3(n6346), .ZN(n6349) );
  INV_X1 U8021 ( .A(n8126), .ZN(n9401) );
  NAND2_X1 U8022 ( .A1(n9401), .A2(n10021), .ZN(n8145) );
  INV_X1 U8023 ( .A(n8145), .ZN(n6350) );
  INV_X1 U8024 ( .A(n6352), .ZN(n8257) );
  NAND2_X1 U8025 ( .A1(n7753), .A2(n10029), .ZN(n7546) );
  NAND2_X1 U8026 ( .A1(n9299), .A2(n7790), .ZN(n8156) );
  NAND2_X1 U8027 ( .A1(n4316), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U8028 ( .A1(n4314), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6360) );
  INV_X1 U8029 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8030 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  AND2_X1 U8031 ( .A1(n6414), .A2(n6357), .ZN(n7788) );
  NAND2_X1 U8032 ( .A1(n6551), .A2(n7788), .ZN(n6359) );
  NAND2_X1 U8033 ( .A1(n6498), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6358) );
  OR2_X1 U8034 ( .A1(n9831), .A2(n9289), .ZN(n8159) );
  NAND2_X1 U8035 ( .A1(n9831), .A2(n9289), .ZN(n8166) );
  NAND2_X1 U8036 ( .A1(n8159), .A2(n8166), .ZN(n7588) );
  INV_X1 U8037 ( .A(n7588), .ZN(n8256) );
  NAND2_X1 U8038 ( .A1(n6375), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U8039 ( .A1(n4315), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6367) );
  NAND2_X1 U8040 ( .A1(n4317), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U8041 ( .A1(n6382), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U8042 ( .A1(n6394), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6364) );
  NOR2_X1 U8043 ( .A1(n7131), .A2(n6994), .ZN(n7129) );
  NAND2_X1 U8044 ( .A1(n8249), .A2(n7129), .ZN(n6369) );
  NAND2_X1 U8045 ( .A1(n7278), .A2(n7271), .ZN(n6368) );
  NAND2_X1 U8046 ( .A1(n4315), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8047 ( .A1(n6382), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U8048 ( .A1(n6375), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U8049 ( .A1(n6394), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6370) );
  AND4_X2 U8050 ( .A1(n6373), .A2(n6372), .A3(n6371), .A4(n6370), .ZN(n6582)
         );
  NAND2_X1 U8051 ( .A1(n6582), .A2(n7901), .ZN(n6581) );
  INV_X1 U8052 ( .A(n6581), .ZN(n8123) );
  INV_X1 U8053 ( .A(n6582), .ZN(n7130) );
  NAND2_X1 U8054 ( .A1(n4315), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6379) );
  INV_X1 U8055 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7260) );
  NAND2_X1 U8056 ( .A1(n6394), .A2(n7260), .ZN(n6378) );
  NAND2_X1 U8057 ( .A1(n4317), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U8058 ( .A1(n6382), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U8059 ( .A1(n6380), .A2(n7257), .ZN(n8138) );
  NAND2_X1 U8060 ( .A1(n7056), .A2(n7430), .ZN(n6381) );
  NAND2_X1 U8061 ( .A1(n8138), .A2(n6381), .ZN(n6584) );
  INV_X1 U8062 ( .A(n6381), .ZN(n8122) );
  NAND2_X1 U8063 ( .A1(n6498), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U8064 ( .A1(n6382), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6387) );
  INV_X1 U8065 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U8066 ( .A1(n7260), .A2(n6383), .ZN(n6384) );
  AND2_X1 U8067 ( .A1(n6384), .A2(n6391), .ZN(n6829) );
  NAND2_X1 U8068 ( .A1(n6394), .A2(n6829), .ZN(n6386) );
  NAND2_X1 U8069 ( .A1(n4315), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6385) );
  AND4_X2 U8070 ( .A1(n6388), .A2(n6387), .A3(n6386), .A4(n6385), .ZN(n7491)
         );
  INV_X1 U8071 ( .A(n7491), .ZN(n9402) );
  NAND2_X1 U8072 ( .A1(n7297), .A2(n8137), .ZN(n6389) );
  NAND2_X1 U8073 ( .A1(n6389), .A2(n8139), .ZN(n7490) );
  INV_X1 U8074 ( .A(n7490), .ZN(n6399) );
  NAND2_X1 U8075 ( .A1(n6382), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U8076 ( .A1(n6498), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U8077 ( .A1(n4314), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6396) );
  INV_X1 U8078 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7402) );
  NAND2_X1 U8079 ( .A1(n6391), .A2(n7402), .ZN(n6392) );
  AND2_X1 U8080 ( .A1(n6393), .A2(n6392), .ZN(n7496) );
  NAND2_X1 U8081 ( .A1(n6394), .A2(n7496), .ZN(n6395) );
  NAND2_X1 U8082 ( .A1(n8128), .A2(n10011), .ZN(n6589) );
  NAND2_X1 U8083 ( .A1(n6399), .A2(n6589), .ZN(n7488) );
  NAND2_X1 U8084 ( .A1(n8126), .A2(n9967), .ZN(n8124) );
  NAND2_X1 U8085 ( .A1(n4316), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U8086 ( .A1(n6498), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6407) );
  XNOR2_X1 U8087 ( .A(n6414), .B(P1_REG3_REG_11__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U8088 ( .A1(n6551), .A2(n9333), .ZN(n6406) );
  NAND2_X1 U8089 ( .A1(n6561), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U8090 ( .A1(n6597), .A2(n7910), .ZN(n8170) );
  INV_X1 U8091 ( .A(n8166), .ZN(n6409) );
  NOR2_X1 U8092 ( .A1(n8245), .A2(n6409), .ZN(n6410) );
  NAND2_X1 U8093 ( .A1(n7607), .A2(n6410), .ZN(n6411) );
  NAND2_X1 U8094 ( .A1(n6411), .A2(n8157), .ZN(n7566) );
  NAND2_X1 U8095 ( .A1(n4317), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8096 ( .A1(n4316), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6418) );
  INV_X1 U8097 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6413) );
  INV_X1 U8098 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6412) );
  OAI21_X1 U8099 ( .B1(n6414), .B2(n6413), .A(n6412), .ZN(n6415) );
  AND2_X1 U8100 ( .A1(n6415), .A2(n6420), .ZN(n9228) );
  NAND2_X1 U8101 ( .A1(n6551), .A2(n9228), .ZN(n6417) );
  NAND2_X1 U8102 ( .A1(n6561), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8103 ( .A1(n9826), .A2(n9336), .ZN(n8171) );
  NAND2_X1 U8104 ( .A1(n8158), .A2(n8171), .ZN(n7567) );
  INV_X1 U8105 ( .A(n7567), .ZN(n8260) );
  NAND2_X1 U8106 ( .A1(n7566), .A2(n8260), .ZN(n7530) );
  NAND2_X1 U8107 ( .A1(n6498), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U8108 ( .A1(n4316), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6424) );
  INV_X1 U8109 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10235) );
  NAND2_X1 U8110 ( .A1(n6420), .A2(n10235), .ZN(n6421) );
  AND2_X1 U8111 ( .A1(n6428), .A2(n6421), .ZN(n9314) );
  NAND2_X1 U8112 ( .A1(n6551), .A2(n9314), .ZN(n6423) );
  NAND2_X1 U8113 ( .A1(n6561), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6422) );
  OR2_X1 U8114 ( .A1(n9820), .A2(n9231), .ZN(n8183) );
  NAND2_X1 U8115 ( .A1(n9820), .A2(n9231), .ZN(n8185) );
  NAND2_X1 U8116 ( .A1(n8183), .A2(n8185), .ZN(n8261) );
  INV_X1 U8117 ( .A(n8158), .ZN(n8169) );
  NOR2_X1 U8118 ( .A1(n8261), .A2(n8169), .ZN(n6426) );
  NAND2_X1 U8119 ( .A1(n6498), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U8120 ( .A1(n4316), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U8121 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  AND2_X1 U8122 ( .A1(n6437), .A2(n6429), .ZN(n9193) );
  NAND2_X1 U8123 ( .A1(n6551), .A2(n9193), .ZN(n6431) );
  NAND2_X1 U8124 ( .A1(n6561), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6430) );
  NAND4_X1 U8125 ( .A1(n6433), .A2(n6432), .A3(n6431), .A4(n6430), .ZN(n9393)
         );
  INV_X1 U8126 ( .A(n9393), .ZN(n7818) );
  NAND2_X1 U8127 ( .A1(n9815), .A2(n7818), .ZN(n8186) );
  NAND2_X1 U8128 ( .A1(n8184), .A2(n8186), .ZN(n7832) );
  INV_X1 U8129 ( .A(n8185), .ZN(n6434) );
  NOR2_X1 U8130 ( .A1(n7832), .A2(n6434), .ZN(n8178) );
  NAND2_X1 U8131 ( .A1(n6498), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8132 ( .A1(n4316), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U8133 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  AND2_X1 U8134 ( .A1(n6445), .A2(n6438), .ZN(n9373) );
  NAND2_X1 U8135 ( .A1(n6551), .A2(n9373), .ZN(n6440) );
  NAND2_X1 U8136 ( .A1(n6561), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6439) );
  NAND4_X1 U8137 ( .A1(n6442), .A2(n6441), .A3(n6440), .A4(n6439), .ZN(n9392)
         );
  INV_X1 U8138 ( .A(n9392), .ZN(n9258) );
  OR2_X1 U8139 ( .A1(n9811), .A2(n9258), .ZN(n8176) );
  NAND2_X1 U8140 ( .A1(n9811), .A2(n9258), .ZN(n8181) );
  NAND2_X1 U8141 ( .A1(n8176), .A2(n8181), .ZN(n8244) );
  NAND2_X1 U8142 ( .A1(n6498), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8143 ( .A1(n4316), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6449) );
  INV_X1 U8144 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8145 ( .A1(n6445), .A2(n6444), .ZN(n6446) );
  AND2_X1 U8146 ( .A1(n6454), .A2(n6446), .ZN(n7863) );
  NAND2_X1 U8147 ( .A1(n6551), .A2(n7863), .ZN(n6448) );
  NAND2_X1 U8148 ( .A1(n6561), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8149 ( .A1(n9803), .A2(n9376), .ZN(n8304) );
  INV_X1 U8150 ( .A(n8181), .ZN(n8302) );
  NAND2_X1 U8151 ( .A1(n4317), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U8152 ( .A1(n4316), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6458) );
  INV_X1 U8153 ( .A(n6454), .ZN(n6452) );
  INV_X1 U8154 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U8155 ( .A1(n6454), .A2(n6453), .ZN(n6455) );
  AND2_X1 U8156 ( .A1(n6462), .A2(n6455), .ZN(n9726) );
  NAND2_X1 U8157 ( .A1(n6551), .A2(n9726), .ZN(n6457) );
  NAND2_X1 U8158 ( .A1(n6561), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6456) );
  NAND4_X1 U8159 ( .A1(n6459), .A2(n6458), .A3(n6457), .A4(n6456), .ZN(n9390)
         );
  INV_X1 U8160 ( .A(n9390), .ZN(n9709) );
  OR2_X1 U8161 ( .A1(n9798), .A2(n9709), .ZN(n8199) );
  NAND2_X1 U8162 ( .A1(n9798), .A2(n9709), .ZN(n8194) );
  NAND2_X1 U8163 ( .A1(n4316), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U8164 ( .A1(n6498), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8165 ( .A1(n6461), .A2(n6460), .ZN(n6466) );
  OR2_X2 U8166 ( .A1(n6462), .A2(n9348), .ZN(n6470) );
  NAND2_X1 U8167 ( .A1(n6462), .A2(n9348), .ZN(n6463) );
  NAND2_X1 U8168 ( .A1(n6470), .A2(n6463), .ZN(n9715) );
  INV_X1 U8169 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n6464) );
  OAI22_X1 U8170 ( .A1(n9715), .A2(n6536), .B1(n6554), .B2(n6464), .ZN(n6465)
         );
  NAND2_X1 U8171 ( .A1(n9794), .A2(n9700), .ZN(n8201) );
  INV_X1 U8172 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U8173 ( .A1(n6470), .A2(n6469), .ZN(n6471) );
  NAND2_X1 U8174 ( .A1(n6482), .A2(n6471), .ZN(n9695) );
  OR2_X1 U8175 ( .A1(n9695), .A2(n6536), .ZN(n6473) );
  AOI22_X1 U8176 ( .A1(n4317), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n4316), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n6472) );
  OAI211_X1 U8177 ( .C1(n6554), .C2(n4510), .A(n6473), .B(n6472), .ZN(n9674)
         );
  NAND2_X1 U8178 ( .A1(n9694), .A2(n9674), .ZN(n8195) );
  INV_X1 U8179 ( .A(n9674), .ZN(n9711) );
  INV_X1 U8180 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U8181 ( .A1(n6484), .A2(n6474), .ZN(n6475) );
  NAND2_X1 U8182 ( .A1(n6487), .A2(n6475), .ZN(n9664) );
  OR2_X1 U8183 ( .A1(n9664), .A2(n6536), .ZN(n6481) );
  INV_X1 U8184 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8185 ( .A1(n6498), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8186 ( .A1(n4316), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6476) );
  OAI211_X1 U8187 ( .C1(n6478), .C2(n6554), .A(n6477), .B(n6476), .ZN(n6479)
         );
  INV_X1 U8188 ( .A(n6479), .ZN(n6480) );
  NAND2_X1 U8189 ( .A1(n6481), .A2(n6480), .ZN(n9676) );
  INV_X1 U8190 ( .A(n9676), .ZN(n9648) );
  NAND2_X1 U8191 ( .A1(n6482), .A2(n10160), .ZN(n6483) );
  NAND2_X1 U8192 ( .A1(n6484), .A2(n6483), .ZN(n9680) );
  AOI22_X1 U8193 ( .A1(n6561), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n4316), .B2(
        P1_REG1_REG_20__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U8194 ( .A1(n6498), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6485) );
  OAI211_X1 U8195 ( .C1(n9680), .C2(n6536), .A(n6486), .B(n6485), .ZN(n9221)
         );
  INV_X1 U8196 ( .A(n9221), .ZN(n9701) );
  OR2_X1 U8197 ( .A1(n9782), .A2(n9701), .ZN(n8205) );
  AND2_X1 U8198 ( .A1(n8243), .A2(n8205), .ZN(n8285) );
  NAND2_X1 U8199 ( .A1(n9778), .A2(n9648), .ZN(n8242) );
  NAND2_X1 U8200 ( .A1(n9782), .A2(n9701), .ZN(n8196) );
  NAND2_X1 U8201 ( .A1(n8242), .A2(n8196), .ZN(n8207) );
  NAND2_X1 U8202 ( .A1(n8207), .A2(n8243), .ZN(n8314) );
  NAND2_X1 U8203 ( .A1(n6487), .A2(n9327), .ZN(n6488) );
  AND2_X1 U8204 ( .A1(n6496), .A2(n6488), .ZN(n9643) );
  NAND2_X1 U8205 ( .A1(n9643), .A2(n6551), .ZN(n6494) );
  INV_X1 U8206 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U8207 ( .A1(n4317), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8208 ( .A1(n4316), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6489) );
  OAI211_X1 U8209 ( .C1(n6491), .C2(n6554), .A(n6490), .B(n6489), .ZN(n6492)
         );
  INV_X1 U8210 ( .A(n6492), .ZN(n6493) );
  NAND2_X1 U8211 ( .A1(n6494), .A2(n6493), .ZN(n9388) );
  INV_X1 U8212 ( .A(n9388), .ZN(n9636) );
  XNOR2_X1 U8213 ( .A(n9773), .B(n9636), .ZN(n9646) );
  NAND2_X1 U8214 ( .A1(n6496), .A2(n9204), .ZN(n6497) );
  NAND2_X1 U8215 ( .A1(n6505), .A2(n6497), .ZN(n9627) );
  INV_X1 U8216 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U8217 ( .A1(n6498), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U8218 ( .A1(n4316), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6499) );
  OAI211_X1 U8219 ( .C1(n9626), .C2(n6554), .A(n6500), .B(n6499), .ZN(n6501)
         );
  INV_X1 U8220 ( .A(n6501), .ZN(n6502) );
  OAI21_X2 U8221 ( .B1(n9627), .B2(n6536), .A(n6502), .ZN(n9387) );
  INV_X1 U8222 ( .A(n9387), .ZN(n9649) );
  OR2_X1 U8223 ( .A1(n9769), .A2(n9649), .ZN(n8216) );
  NAND2_X1 U8224 ( .A1(n9769), .A2(n9649), .ZN(n9608) );
  NAND2_X1 U8225 ( .A1(n8216), .A2(n9608), .ZN(n9634) );
  NOR2_X1 U8226 ( .A1(n9773), .A2(n9636), .ZN(n8208) );
  NOR2_X1 U8227 ( .A1(n9634), .A2(n8208), .ZN(n6503) );
  INV_X1 U8228 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U8229 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  AND2_X1 U8230 ( .A1(n6515), .A2(n6506), .ZN(n9616) );
  NAND2_X1 U8231 ( .A1(n9616), .A2(n6551), .ZN(n6512) );
  INV_X1 U8232 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U8233 ( .A1(n6498), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U8234 ( .A1(n4316), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6507) );
  OAI211_X1 U8235 ( .C1(n6509), .C2(n6554), .A(n6508), .B(n6507), .ZN(n6510)
         );
  INV_X1 U8236 ( .A(n6510), .ZN(n6511) );
  INV_X1 U8237 ( .A(n9386), .ZN(n9637) );
  OR2_X1 U8238 ( .A1(n9764), .A2(n9637), .ZN(n8280) );
  NAND2_X1 U8239 ( .A1(n9764), .A2(n9637), .ZN(n8313) );
  NAND2_X1 U8240 ( .A1(n8280), .A2(n8313), .ZN(n9609) );
  INV_X1 U8241 ( .A(n9608), .ZN(n8281) );
  NOR2_X1 U8242 ( .A1(n9609), .A2(n8281), .ZN(n6513) );
  INV_X1 U8243 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U8244 ( .A1(n6515), .A2(n9243), .ZN(n6516) );
  NAND2_X1 U8245 ( .A1(n6523), .A2(n6516), .ZN(n9595) );
  INV_X1 U8246 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9594) );
  NAND2_X1 U8247 ( .A1(n4317), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U8248 ( .A1(n4316), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6517) );
  OAI211_X1 U8249 ( .C1(n9594), .C2(n6554), .A(n6518), .B(n6517), .ZN(n6519)
         );
  INV_X1 U8250 ( .A(n6519), .ZN(n6520) );
  INV_X1 U8251 ( .A(n9385), .ZN(n9612) );
  OR2_X1 U8252 ( .A1(n9759), .A2(n9612), .ZN(n8282) );
  NAND2_X1 U8253 ( .A1(n9759), .A2(n9612), .ZN(n8316) );
  NAND2_X1 U8254 ( .A1(n8282), .A2(n8316), .ZN(n9600) );
  INV_X1 U8255 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9358) );
  OR2_X2 U8256 ( .A1(n6523), .A2(n9358), .ZN(n6534) );
  NAND2_X1 U8257 ( .A1(n6523), .A2(n9358), .ZN(n6524) );
  NAND2_X1 U8258 ( .A1(n9363), .A2(n6551), .ZN(n6530) );
  INV_X1 U8259 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U8260 ( .A1(n6498), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U8261 ( .A1(n4316), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6525) );
  OAI211_X1 U8262 ( .C1(n6527), .C2(n6554), .A(n6526), .B(n6525), .ZN(n6528)
         );
  INV_X1 U8263 ( .A(n6528), .ZN(n6529) );
  INV_X1 U8264 ( .A(n9384), .ZN(n6531) );
  OR2_X1 U8265 ( .A1(n9753), .A2(n6531), .ZN(n8324) );
  NAND2_X1 U8266 ( .A1(n9753), .A2(n6531), .ZN(n8219) );
  INV_X1 U8267 ( .A(n6534), .ZN(n6532) );
  INV_X1 U8268 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8269 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  NAND2_X1 U8270 ( .A1(n6550), .A2(n6535), .ZN(n8106) );
  INV_X1 U8271 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U8272 ( .A1(n6498), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U8273 ( .A1(n4316), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6537) );
  OAI211_X1 U8274 ( .C1(n6539), .C2(n6554), .A(n6538), .B(n6537), .ZN(n6540)
         );
  INV_X1 U8275 ( .A(n6540), .ZN(n6541) );
  NAND2_X1 U8276 ( .A1(n9748), .A2(n9360), .ZN(n8114) );
  INV_X1 U8277 ( .A(n8273), .ZN(n7882) );
  XNOR2_X1 U8278 ( .A(n6550), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U8279 ( .A1(n9578), .A2(n6551), .ZN(n6548) );
  INV_X1 U8280 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U8281 ( .A1(n6498), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U8282 ( .A1(n6561), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6543) );
  OAI211_X1 U8283 ( .C1(n6545), .C2(n4311), .A(n6544), .B(n6543), .ZN(n6546)
         );
  INV_X1 U8284 ( .A(n6546), .ZN(n6547) );
  INV_X1 U8285 ( .A(n9383), .ZN(n6549) );
  OR2_X1 U8286 ( .A1(n9742), .A2(n6549), .ZN(n8225) );
  NAND2_X1 U8287 ( .A1(n9742), .A2(n6549), .ZN(n8115) );
  NAND2_X1 U8288 ( .A1(n9581), .A2(n8115), .ZN(n6558) );
  INV_X1 U8289 ( .A(n6550), .ZN(n9566) );
  NAND3_X1 U8290 ( .A1(n9566), .A2(n6551), .A3(P1_REG3_REG_28__SCAN_IN), .ZN(
        n6557) );
  INV_X1 U8291 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n10238) );
  NAND2_X1 U8292 ( .A1(n4317), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U8293 ( .A1(n4316), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6552) );
  OAI211_X1 U8294 ( .C1(n10238), .C2(n6554), .A(n6553), .B(n6552), .ZN(n6555)
         );
  INV_X1 U8295 ( .A(n6555), .ZN(n6556) );
  NAND2_X1 U8296 ( .A1(n6569), .A2(n8067), .ZN(n8329) );
  INV_X1 U8297 ( .A(n9564), .ZN(n8275) );
  XNOR2_X1 U8298 ( .A(n6558), .B(n8275), .ZN(n6560) );
  NAND2_X1 U8299 ( .A1(n8375), .A2(n6772), .ZN(n6559) );
  NAND2_X1 U8300 ( .A1(n8247), .A2(n8365), .ZN(n8336) );
  NAND2_X1 U8301 ( .A1(n6560), .A2(n9962), .ZN(n6566) );
  INV_X1 U8302 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10220) );
  NAND2_X1 U8303 ( .A1(n4316), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U8304 ( .A1(n6561), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6562) );
  OAI211_X1 U8305 ( .C1(n6390), .C2(n10220), .A(n6563), .B(n6562), .ZN(n9382)
         );
  AOI22_X1 U8306 ( .A1(n9383), .A2(n9673), .B1(n6564), .B2(n9382), .ZN(n6565)
         );
  NAND2_X1 U8307 ( .A1(n6566), .A2(n6565), .ZN(n9572) );
  OR2_X1 U8308 ( .A1(n6770), .A2(n6769), .ZN(n8373) );
  NAND2_X1 U8309 ( .A1(n6770), .A2(n8369), .ZN(n6567) );
  NAND3_X1 U8310 ( .A1(n8373), .A2(n7321), .A3(n6567), .ZN(n7835) );
  NAND2_X1 U8311 ( .A1(n8238), .A2(n8358), .ZN(n10031) );
  NAND2_X1 U8312 ( .A1(n9742), .A2(n9383), .ZN(n9561) );
  OR3_X1 U8313 ( .A1(n9564), .A2(n10051), .A3(n9561), .ZN(n6572) );
  AOI21_X1 U8314 ( .B1(n6569), .B2(n6568), .A(n9724), .ZN(n6571) );
  NAND2_X1 U8315 ( .A1(n6571), .A2(n6570), .ZN(n9565) );
  NAND2_X1 U8316 ( .A1(n7131), .A2(n7320), .ZN(n7128) );
  NAND2_X1 U8317 ( .A1(n6573), .A2(n7271), .ZN(n6574) );
  NAND2_X1 U8318 ( .A1(n7128), .A2(n6574), .ZN(n6580) );
  NAND2_X1 U8319 ( .A1(n6582), .A2(n6374), .ZN(n7121) );
  NAND2_X1 U8320 ( .A1(n7052), .A2(n6583), .ZN(n6587) );
  INV_X1 U8321 ( .A(n6584), .ZN(n6585) );
  NAND2_X1 U8322 ( .A1(n6585), .A2(n7285), .ZN(n6586) );
  NAND2_X1 U8323 ( .A1(n8137), .A2(n8139), .ZN(n7287) );
  NAND2_X1 U8324 ( .A1(n7491), .A2(n7302), .ZN(n6588) );
  NAND2_X1 U8325 ( .A1(n7487), .A2(n8253), .ZN(n6591) );
  NAND2_X1 U8326 ( .A1(n8128), .A2(n8129), .ZN(n6590) );
  NAND2_X1 U8327 ( .A1(n6591), .A2(n6590), .ZN(n9968) );
  NAND2_X1 U8328 ( .A1(n8124), .A2(n8145), .ZN(n9969) );
  NAND2_X1 U8329 ( .A1(n9968), .A2(n9969), .ZN(n6593) );
  NAND2_X1 U8330 ( .A1(n8126), .A2(n10021), .ZN(n6592) );
  NAND2_X1 U8331 ( .A1(n7474), .A2(n8135), .ZN(n6595) );
  INV_X1 U8332 ( .A(n10029), .ZN(n7483) );
  NAND2_X1 U8333 ( .A1(n7483), .A2(n7753), .ZN(n6594) );
  NOR2_X1 U8334 ( .A1(n10039), .A2(n9399), .ZN(n7544) );
  NAND2_X1 U8335 ( .A1(n10039), .A2(n9399), .ZN(n7542) );
  OR2_X1 U8336 ( .A1(n9299), .A2(n9398), .ZN(n6596) );
  OAI21_X2 U8337 ( .B1(n7648), .B2(n7650), .A(n6596), .ZN(n7595) );
  NAND2_X1 U8338 ( .A1(n7595), .A2(n7588), .ZN(n7559) );
  INV_X1 U8339 ( .A(n8245), .ZN(n6599) );
  NOR2_X1 U8340 ( .A1(n6597), .A2(n9396), .ZN(n7558) );
  INV_X1 U8341 ( .A(n7558), .ZN(n6598) );
  NAND2_X1 U8342 ( .A1(n7567), .A2(n6600), .ZN(n7562) );
  INV_X1 U8343 ( .A(n7562), .ZN(n6602) );
  INV_X1 U8344 ( .A(n9289), .ZN(n9397) );
  OR2_X1 U8345 ( .A1(n9831), .A2(n9397), .ZN(n7560) );
  NAND2_X1 U8346 ( .A1(n6598), .A2(n7560), .ZN(n7561) );
  INV_X1 U8347 ( .A(n9336), .ZN(n9395) );
  NOR2_X1 U8348 ( .A1(n9826), .A2(n9395), .ZN(n6601) );
  AOI21_X1 U8349 ( .B1(n6602), .B2(n7561), .A(n6601), .ZN(n6603) );
  INV_X1 U8350 ( .A(n9231), .ZN(n9394) );
  OR2_X1 U8351 ( .A1(n9820), .A2(n9394), .ZN(n6604) );
  NOR2_X1 U8352 ( .A1(n9815), .A2(n9393), .ZN(n6605) );
  AND2_X1 U8353 ( .A1(n9811), .A2(n9392), .ZN(n6607) );
  OR2_X1 U8354 ( .A1(n9811), .A2(n9392), .ZN(n6606) );
  OAI21_X2 U8355 ( .B1(n7813), .B2(n6607), .A(n6606), .ZN(n7862) );
  INV_X1 U8356 ( .A(n9376), .ZN(n9391) );
  NAND2_X1 U8357 ( .A1(n9803), .A2(n9391), .ZN(n6608) );
  OR2_X1 U8358 ( .A1(n9798), .A2(n9390), .ZN(n6609) );
  NAND2_X1 U8359 ( .A1(n9798), .A2(n9390), .ZN(n6610) );
  AND2_X1 U8360 ( .A1(n9794), .A2(n9389), .ZN(n6612) );
  NAND2_X1 U8361 ( .A1(n9789), .A2(n9674), .ZN(n6613) );
  AND2_X1 U8362 ( .A1(n9782), .A2(n9221), .ZN(n6614) );
  AND2_X1 U8363 ( .A1(n9773), .A2(n9388), .ZN(n6616) );
  OAI21_X2 U8364 ( .B1(n9640), .B2(n6616), .A(n6615), .ZN(n9622) );
  NAND2_X1 U8365 ( .A1(n9769), .A2(n9387), .ZN(n6617) );
  AND2_X1 U8366 ( .A1(n9764), .A2(n9386), .ZN(n6619) );
  NOR2_X1 U8367 ( .A1(n9759), .A2(n9385), .ZN(n6621) );
  NAND2_X1 U8368 ( .A1(n9759), .A2(n9385), .ZN(n6620) );
  AND2_X1 U8369 ( .A1(n9753), .A2(n9384), .ZN(n6623) );
  OR2_X1 U8370 ( .A1(n9753), .A2(n9384), .ZN(n6622) );
  NOR2_X1 U8371 ( .A1(n9748), .A2(n9586), .ZN(n6624) );
  OR2_X1 U8372 ( .A1(n9742), .A2(n9383), .ZN(n6625) );
  INV_X1 U8373 ( .A(n9562), .ZN(n6626) );
  NAND3_X1 U8374 ( .A1(n6626), .A2(n10026), .A3(n8275), .ZN(n6631) );
  INV_X1 U8375 ( .A(n9561), .ZN(n6627) );
  AND2_X1 U8376 ( .A1(n9564), .A2(n6628), .ZN(n6629) );
  NAND2_X1 U8377 ( .A1(n10053), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U8378 ( .A1(n6633), .A2(n6632), .ZN(P1_U3519) );
  NAND2_X1 U8379 ( .A1(n6749), .A2(n6634), .ZN(n6635) );
  NAND2_X1 U8380 ( .A1(n6635), .A2(n6748), .ZN(n6755) );
  NAND2_X1 U8381 ( .A1(n6755), .A2(n6636), .ZN(n6637) );
  NAND2_X1 U8382 ( .A1(n6637), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8383 ( .A(n6732), .ZN(n8686) );
  AND2_X1 U8384 ( .A1(n6666), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U8385 ( .A1(n4431), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U8386 ( .A1(n6967), .A2(n6639), .ZN(n8617) );
  NAND2_X1 U8387 ( .A1(n8617), .A2(n8618), .ZN(n8616) );
  NAND2_X1 U8388 ( .A1(n6641), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U8389 ( .A1(n10067), .A2(n6643), .ZN(n8638) );
  NAND2_X1 U8390 ( .A1(n6852), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6645) );
  OAI21_X1 U8391 ( .B1(n6852), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6645), .ZN(
        n6644) );
  INV_X1 U8392 ( .A(n6644), .ZN(n8639) );
  NAND2_X1 U8393 ( .A1(n8638), .A2(n8639), .ZN(n8637) );
  NAND2_X1 U8394 ( .A1(n8637), .A2(n6645), .ZN(n6646) );
  XNOR2_X1 U8395 ( .A(n6715), .B(n7372), .ZN(n10086) );
  INV_X1 U8396 ( .A(n6715), .ZN(n10092) );
  NOR2_X1 U8397 ( .A1(n6648), .A2(n6716), .ZN(n6649) );
  AOI21_X1 U8398 ( .B1(n6648), .B2(n6716), .A(n6649), .ZN(n10104) );
  NAND2_X1 U8399 ( .A1(n10104), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7181) );
  INV_X1 U8400 ( .A(n6649), .ZN(n7182) );
  XNOR2_X1 U8401 ( .A(n6720), .B(n7506), .ZN(n7183) );
  INV_X1 U8402 ( .A(n6720), .ZN(n7187) );
  NOR2_X1 U8403 ( .A1(n7180), .A2(n4978), .ZN(n6650) );
  XNOR2_X1 U8404 ( .A(n7444), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7448) );
  INV_X1 U8405 ( .A(n6726), .ZN(n8648) );
  XNOR2_X1 U8406 ( .A(n6728), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7806) );
  XNOR2_X1 U8407 ( .A(n6732), .B(n8944), .ZN(n8678) );
  NOR2_X1 U8408 ( .A1(n6655), .A2(n7033), .ZN(n6657) );
  NOR2_X1 U8409 ( .A1(n6657), .A2(n6656), .ZN(n8694) );
  INV_X1 U8410 ( .A(n6657), .ZN(n6658) );
  XNOR2_X1 U8411 ( .A(n6736), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8707) );
  INV_X1 U8412 ( .A(n6736), .ZN(n8714) );
  INV_X1 U8413 ( .A(n6740), .ZN(n8727) );
  NAND2_X1 U8414 ( .A1(n8721), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8737) );
  INV_X1 U8415 ( .A(n6661), .ZN(n8736) );
  OR2_X1 U8416 ( .A1(n8750), .A2(n10246), .ZN(n6663) );
  NAND2_X1 U8417 ( .A1(n8750), .A2(n10246), .ZN(n6662) );
  NAND2_X1 U8418 ( .A1(n6663), .A2(n6662), .ZN(n8735) );
  INV_X1 U8419 ( .A(n6663), .ZN(n6664) );
  XNOR2_X1 U8420 ( .A(n7328), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6744) );
  NOR2_X1 U8421 ( .A1(n6754), .A2(P2_U3151), .ZN(n9182) );
  NAND2_X1 U8422 ( .A1(n4431), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8423 ( .A1(n6838), .A2(n6671), .ZN(n6670) );
  NAND2_X1 U8424 ( .A1(n6666), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6668) );
  OR2_X1 U8425 ( .A1(n6668), .A2(n4431), .ZN(n6669) );
  NAND2_X1 U8426 ( .A1(n6670), .A2(n6669), .ZN(n6974) );
  NAND2_X1 U8427 ( .A1(n6974), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U8428 ( .A1(n6672), .A2(n6671), .ZN(n8614) );
  NAND2_X1 U8429 ( .A1(n6641), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U8430 ( .A1(n10066), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6676) );
  NAND2_X1 U8431 ( .A1(n6674), .A2(n4790), .ZN(n6675) );
  NAND2_X1 U8432 ( .A1(n6676), .A2(n6675), .ZN(n8635) );
  MUX2_X1 U8433 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6677), .S(n6852), .Z(n8636)
         );
  NAND2_X1 U8434 ( .A1(n6852), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6678) );
  NAND2_X1 U8435 ( .A1(n6679), .A2(n6854), .ZN(n6680) );
  NAND2_X1 U8436 ( .A1(n6681), .A2(n6680), .ZN(n10083) );
  MUX2_X1 U8437 ( .A(n6682), .B(P2_REG1_REG_6__SCAN_IN), .S(n6715), .Z(n10084)
         );
  NAND2_X1 U8438 ( .A1(n10083), .A2(n10084), .ZN(n10082) );
  OR2_X1 U8439 ( .A1(n6715), .A2(n6682), .ZN(n6683) );
  XNOR2_X1 U8440 ( .A(n6684), .B(n6716), .ZN(n10105) );
  NAND2_X1 U8441 ( .A1(n10105), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6686) );
  INV_X1 U8442 ( .A(n6716), .ZN(n10110) );
  NAND2_X1 U8443 ( .A1(n6684), .A2(n10110), .ZN(n6685) );
  NAND2_X1 U8444 ( .A1(n6686), .A2(n6685), .ZN(n7176) );
  XNOR2_X1 U8445 ( .A(n6720), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7177) );
  NAND2_X1 U8446 ( .A1(n7176), .A2(n7177), .ZN(n6688) );
  OR2_X1 U8447 ( .A1(n6720), .A2(n7502), .ZN(n6687) );
  INV_X1 U8448 ( .A(n6721), .ZN(n7465) );
  NAND2_X1 U8449 ( .A1(n6689), .A2(n7465), .ZN(n6690) );
  INV_X1 U8450 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9063) );
  XNOR2_X1 U8451 ( .A(n7444), .B(n9063), .ZN(n7440) );
  INV_X1 U8452 ( .A(n6691), .ZN(n6692) );
  XOR2_X1 U8453 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6728), .Z(n7797) );
  OAI22_X1 U8454 ( .A1(n7796), .A2(n7797), .B1(n6728), .B2(n9059), .ZN(n6693)
         );
  XNOR2_X1 U8455 ( .A(n6693), .B(n6730), .ZN(n8659) );
  XOR2_X1 U8456 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n6732), .Z(n8676) );
  INV_X1 U8457 ( .A(n6694), .ZN(n6695) );
  XNOR2_X1 U8458 ( .A(n6736), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8706) );
  AOI22_X1 U8459 ( .A1(n8705), .A2(n8706), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n8714), .ZN(n6696) );
  XNOR2_X1 U8460 ( .A(n6696), .B(n6740), .ZN(n8720) );
  OAI22_X1 U8461 ( .A1(n8720), .A2(n9043), .B1(n6740), .B2(n6696), .ZN(n8733)
         );
  XNOR2_X1 U8462 ( .A(n8750), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8734) );
  INV_X1 U8463 ( .A(n8750), .ZN(n8744) );
  AOI22_X1 U8464 ( .A1(n8733), .A2(n8734), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8744), .ZN(n6698) );
  XNOR2_X1 U8465 ( .A(n6697), .B(n9037), .ZN(n6745) );
  INV_X1 U8466 ( .A(n6914), .ZN(n6699) );
  MUX2_X1 U8467 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6753), .Z(n6733) );
  MUX2_X1 U8468 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6753), .Z(n6731) );
  MUX2_X1 U8469 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6753), .Z(n6729) );
  INV_X1 U8470 ( .A(n6728), .ZN(n7798) );
  MUX2_X1 U8471 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n6753), .Z(n6713) );
  INV_X1 U8472 ( .A(n6713), .ZN(n6714) );
  MUX2_X1 U8473 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6753), .Z(n6711) );
  INV_X1 U8474 ( .A(n6711), .ZN(n6712) );
  MUX2_X1 U8475 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6753), .Z(n6709) );
  INV_X1 U8476 ( .A(n6709), .ZN(n6710) );
  MUX2_X1 U8477 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6753), .Z(n6706) );
  INV_X1 U8478 ( .A(n6706), .ZN(n6707) );
  INV_X1 U8479 ( .A(n6641), .ZN(n6705) );
  MUX2_X1 U8480 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6753), .Z(n6703) );
  INV_X1 U8481 ( .A(n6703), .ZN(n6704) );
  INV_X1 U8482 ( .A(n6838), .ZN(n6976) );
  INV_X1 U8483 ( .A(n6700), .ZN(n6702) );
  MUX2_X1 U8484 ( .A(n10163), .B(n6701), .S(n6753), .Z(n6912) );
  NAND2_X1 U8485 ( .A1(n6912), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6969) );
  XOR2_X1 U8486 ( .A(n6641), .B(n6703), .Z(n8623) );
  NAND2_X1 U8487 ( .A1(n8622), .A2(n8623), .ZN(n8621) );
  OAI21_X1 U8488 ( .B1(n6705), .B2(n6704), .A(n8621), .ZN(n10076) );
  XOR2_X1 U8489 ( .A(n6708), .B(n6706), .Z(n10077) );
  NOR2_X1 U8490 ( .A1(n10076), .A2(n10077), .ZN(n10075) );
  XNOR2_X1 U8491 ( .A(n6709), .B(n8630), .ZN(n8632) );
  XNOR2_X1 U8492 ( .A(n6711), .B(n6925), .ZN(n6920) );
  OAI21_X1 U8493 ( .B1(n6925), .B2(n6712), .A(n6919), .ZN(n10097) );
  XOR2_X1 U8494 ( .A(n6715), .B(n6713), .Z(n10098) );
  NOR2_X1 U8495 ( .A1(n10097), .A2(n10098), .ZN(n10096) );
  AOI21_X1 U8496 ( .B1(n6715), .B2(n6714), .A(n10096), .ZN(n10117) );
  MUX2_X1 U8497 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n6753), .Z(n6717) );
  XOR2_X1 U8498 ( .A(n6716), .B(n6717), .Z(n10116) );
  OAI22_X1 U8499 ( .A1(n10117), .A2(n10116), .B1(n6717), .B2(n10110), .ZN(
        n7179) );
  MUX2_X1 U8500 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6753), .Z(n6718) );
  XNOR2_X1 U8501 ( .A(n6718), .B(n6720), .ZN(n7178) );
  INV_X1 U8502 ( .A(n6718), .ZN(n6719) );
  AOI22_X1 U8503 ( .A1(n7179), .A2(n7178), .B1(n6720), .B2(n6719), .ZN(n7466)
         );
  MUX2_X1 U8504 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n6753), .Z(n6722) );
  XOR2_X1 U8505 ( .A(n6721), .B(n6722), .Z(n7467) );
  MUX2_X1 U8506 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n6753), .Z(n6723) );
  XNOR2_X1 U8507 ( .A(n6723), .B(n6725), .ZN(n7441) );
  INV_X1 U8508 ( .A(n6723), .ZN(n6724) );
  MUX2_X1 U8509 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n6753), .Z(n6727) );
  XOR2_X1 U8510 ( .A(n6726), .B(n6727), .Z(n8653) );
  XOR2_X1 U8511 ( .A(n6728), .B(n6729), .Z(n7801) );
  AOI21_X1 U8512 ( .B1(n6729), .B2(n7798), .A(n7799), .ZN(n8662) );
  XNOR2_X1 U8513 ( .A(n6730), .B(n6731), .ZN(n8661) );
  NAND2_X1 U8514 ( .A1(n8662), .A2(n8661), .ZN(n8660) );
  XNOR2_X1 U8515 ( .A(n6732), .B(n6733), .ZN(n8682) );
  MUX2_X1 U8516 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6753), .Z(n6734) );
  XNOR2_X1 U8517 ( .A(n7033), .B(n6734), .ZN(n8696) );
  INV_X1 U8518 ( .A(n6734), .ZN(n6735) );
  MUX2_X1 U8519 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6753), .Z(n6737) );
  XOR2_X1 U8520 ( .A(n6737), .B(n6736), .Z(n8710) );
  OAI22_X1 U8521 ( .A1(n8711), .A2(n8710), .B1(n8714), .B2(n6737), .ZN(n8724)
         );
  MUX2_X1 U8522 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n6753), .Z(n6738) );
  XNOR2_X1 U8523 ( .A(n6740), .B(n6738), .ZN(n8723) );
  INV_X1 U8524 ( .A(n6738), .ZN(n6739) );
  AOI22_X1 U8525 ( .A1(n8724), .A2(n8723), .B1(n6740), .B2(n6739), .ZN(n6742)
         );
  MUX2_X1 U8526 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6753), .Z(n6741) );
  NOR2_X1 U8527 ( .A1(n6742), .A2(n6741), .ZN(n8740) );
  NAND2_X1 U8528 ( .A1(n6742), .A2(n6741), .ZN(n8741) );
  OAI21_X1 U8529 ( .B1(n8740), .B2(n8750), .A(n8741), .ZN(n6747) );
  MUX2_X1 U8530 ( .A(n6745), .B(n6744), .S(n6743), .Z(n6746) );
  XNOR2_X1 U8531 ( .A(n6747), .B(n6746), .ZN(n6762) );
  INV_X1 U8532 ( .A(n6748), .ZN(n8111) );
  INV_X1 U8533 ( .A(n9182), .ZN(n6752) );
  OR2_X1 U8534 ( .A1(n6758), .A2(n6752), .ZN(n6757) );
  NOR2_X1 U8535 ( .A1(n6753), .A2(P2_U3151), .ZN(n7857) );
  NAND3_X1 U8536 ( .A1(n6755), .A2(n7857), .A3(n6754), .ZN(n6756) );
  INV_X1 U8537 ( .A(n6758), .ZN(n6759) );
  NAND2_X1 U8538 ( .A1(n10118), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U8539 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8444) );
  OAI211_X1 U8540 ( .C1(n10111), .C2(n7328), .A(n6760), .B(n8444), .ZN(n6761)
         );
  INV_X1 U8541 ( .A(n6764), .ZN(n6765) );
  NAND2_X1 U8542 ( .A1(n6766), .A2(n6765), .ZN(P2_U3487) );
  INV_X1 U8543 ( .A(n7293), .ZN(n6815) );
  NOR2_X1 U8544 ( .A1(n6821), .A2(P1_U3086), .ZN(n6768) );
  NAND2_X4 U8545 ( .A1(n6771), .A2(n6770), .ZN(n8061) );
  OAI21_X1 U8546 ( .B1(n8375), .B2(n8369), .A(n6821), .ZN(n6774) );
  INV_X1 U8547 ( .A(n6774), .ZN(n6775) );
  INV_X1 U8548 ( .A(n7349), .ZN(n6799) );
  OAI22_X1 U8549 ( .A1(n7491), .A2(n4341), .B1(n7302), .B2(n6799), .ZN(n6776)
         );
  XNOR2_X1 U8550 ( .A(n6776), .B(n8061), .ZN(n6779) );
  OR2_X1 U8551 ( .A1(n7491), .A2(n8050), .ZN(n6778) );
  NAND2_X1 U8552 ( .A1(n10004), .A2(n8058), .ZN(n6777) );
  NAND2_X1 U8553 ( .A1(n6778), .A2(n6777), .ZN(n6780) );
  NAND2_X1 U8554 ( .A1(n6779), .A2(n6780), .ZN(n7395) );
  INV_X1 U8555 ( .A(n6779), .ZN(n6782) );
  INV_X1 U8556 ( .A(n6780), .ZN(n6781) );
  NAND2_X1 U8557 ( .A1(n6782), .A2(n6781), .ZN(n6783) );
  NAND2_X1 U8558 ( .A1(n7395), .A2(n6783), .ZN(n6820) );
  AND2_X1 U8559 ( .A1(n7349), .A2(n7320), .ZN(n6784) );
  INV_X1 U8560 ( .A(n6821), .ZN(n6786) );
  NAND2_X1 U8561 ( .A1(n6786), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U8562 ( .A1(n6789), .A2(n6785), .ZN(n7064) );
  NAND2_X1 U8563 ( .A1(n7131), .A2(n8063), .ZN(n6788) );
  AOI22_X1 U8564 ( .A1(n7320), .A2(n8058), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6786), .ZN(n6787) );
  NAND2_X1 U8565 ( .A1(n6788), .A2(n6787), .ZN(n7063) );
  NAND2_X1 U8566 ( .A1(n7064), .A2(n7063), .ZN(n7066) );
  NAND2_X1 U8567 ( .A1(n6789), .A2(n8048), .ZN(n6790) );
  AND2_X1 U8568 ( .A1(n7066), .A2(n6790), .ZN(n7266) );
  NAND2_X1 U8569 ( .A1(n7349), .A2(n7271), .ZN(n6791) );
  NAND2_X1 U8570 ( .A1(n6792), .A2(n6791), .ZN(n6793) );
  XNOR2_X1 U8571 ( .A(n6793), .B(n8061), .ZN(n6795) );
  AND2_X1 U8572 ( .A1(n8058), .A2(n7271), .ZN(n6794) );
  INV_X1 U8573 ( .A(n6795), .ZN(n6797) );
  NAND2_X1 U8574 ( .A1(n6797), .A2(n6796), .ZN(n6798) );
  NAND2_X1 U8575 ( .A1(n7267), .A2(n6798), .ZN(n7898) );
  OAI22_X1 U8576 ( .A1(n6582), .A2(n4341), .B1(n6374), .B2(n6799), .ZN(n6800)
         );
  XNOR2_X1 U8577 ( .A(n6800), .B(n8048), .ZN(n6805) );
  OR2_X1 U8578 ( .A1(n6582), .A2(n8050), .ZN(n6802) );
  NAND2_X1 U8579 ( .A1(n7901), .A2(n8058), .ZN(n6801) );
  NAND2_X1 U8580 ( .A1(n6802), .A2(n6801), .ZN(n6803) );
  XNOR2_X1 U8581 ( .A(n6805), .B(n6803), .ZN(n7899) );
  NAND2_X1 U8582 ( .A1(n7898), .A2(n7899), .ZN(n6807) );
  INV_X1 U8583 ( .A(n6803), .ZN(n6804) );
  NAND2_X1 U8584 ( .A1(n6805), .A2(n6804), .ZN(n6806) );
  NAND2_X1 U8585 ( .A1(n6807), .A2(n6806), .ZN(n7255) );
  OAI22_X1 U8586 ( .A1(n7056), .A2(n4341), .B1(n7257), .B2(n6799), .ZN(n6808)
         );
  XNOR2_X1 U8587 ( .A(n6808), .B(n8048), .ZN(n6809) );
  OAI22_X1 U8588 ( .A1(n7056), .A2(n8050), .B1(n7257), .B2(n4341), .ZN(n6810)
         );
  XNOR2_X1 U8589 ( .A(n6809), .B(n6810), .ZN(n7256) );
  INV_X1 U8590 ( .A(n6809), .ZN(n6811) );
  OR2_X1 U8591 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  INV_X1 U8592 ( .A(n6813), .ZN(n6814) );
  NAND3_X1 U8593 ( .A1(n6815), .A2(n7295), .A3(n6814), .ZN(n6826) );
  NAND2_X1 U8594 ( .A1(n10020), .A2(n8354), .ZN(n6816) );
  INV_X1 U8595 ( .A(n7396), .ZN(n6818) );
  AOI211_X1 U8596 ( .C1(n6820), .C2(n6819), .A(n9380), .B(n6818), .ZN(n6836)
         );
  NAND2_X1 U8597 ( .A1(n6826), .A2(n10020), .ZN(n6822) );
  NAND3_X1 U8598 ( .A1(n6822), .A2(n7292), .A3(n6821), .ZN(n6823) );
  NAND2_X1 U8599 ( .A1(n6823), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6828) );
  NOR2_X1 U8600 ( .A1(n7321), .A2(n8358), .ZN(n9975) );
  AND2_X1 U8601 ( .A1(n9975), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6825) );
  INV_X1 U8602 ( .A(n8378), .ZN(n6824) );
  AOI21_X1 U8603 ( .B1(n6826), .B2(n6825), .A(n6824), .ZN(n6827) );
  INV_X1 U8604 ( .A(n6829), .ZN(n7301) );
  NOR2_X1 U8605 ( .A1(n9349), .A2(n7301), .ZN(n6835) );
  NOR2_X1 U8606 ( .A1(n6830), .A2(n8369), .ZN(n9269) );
  OAI22_X1 U8607 ( .A1(n8128), .A2(n9375), .B1(n9359), .B2(n7056), .ZN(n6834)
         );
  INV_X1 U8608 ( .A(n6830), .ZN(n6832) );
  NAND2_X1 U8609 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7092) );
  OAI21_X1 U8610 ( .B1(n9366), .B2(n7302), .A(n7092), .ZN(n6833) );
  OR4_X1 U8611 ( .A1(n6836), .A2(n6835), .A3(n6834), .A4(n6833), .ZN(P1_U3230)
         );
  XNOR2_X1 U8612 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X2 U8613 ( .A1(n6837), .A2(P2_U3151), .ZN(n8387) );
  AND2_X1 U8614 ( .A1(n6840), .A2(P2_U3151), .ZN(n9180) );
  INV_X2 U8615 ( .A(n9180), .ZN(n7852) );
  OAI222_X1 U8616 ( .A1(n8387), .A2(n6839), .B1(n7852), .B2(n6851), .C1(
        P2_U3151), .C2(n6838), .ZN(P2_U3294) );
  NOR2_X1 U8617 ( .A1(n6840), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9859) );
  OAI222_X1 U8618 ( .A1(n9866), .A2(n6841), .B1(n9864), .B2(n6842), .C1(
        P1_U3086), .C2(n7080), .ZN(P1_U3353) );
  OAI222_X1 U8619 ( .A1(n8387), .A2(n6843), .B1(n7852), .B2(n6842), .C1(
        P2_U3151), .C2(n6641), .ZN(P2_U3293) );
  INV_X1 U8620 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6845) );
  INV_X1 U8621 ( .A(n6844), .ZN(n6846) );
  INV_X1 U8622 ( .A(n9461), .ZN(n7003) );
  OAI222_X1 U8623 ( .A1(n9866), .A2(n6845), .B1(n9864), .B2(n6846), .C1(
        P1_U3086), .C2(n7003), .ZN(P1_U3348) );
  OAI222_X1 U8624 ( .A1(n8387), .A2(n4594), .B1(n7852), .B2(n6846), .C1(
        P2_U3151), .C2(n10110), .ZN(P2_U3288) );
  INV_X1 U8625 ( .A(n6847), .ZN(n6848) );
  OAI222_X1 U8626 ( .A1(n8387), .A2(n5092), .B1(n7852), .B2(n6848), .C1(
        P2_U3151), .C2(n10092), .ZN(P2_U3289) );
  INV_X1 U8627 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6849) );
  INV_X1 U8628 ( .A(n9448), .ZN(n7001) );
  OAI222_X1 U8629 ( .A1(n9866), .A2(n6849), .B1(n9864), .B2(n6848), .C1(
        P1_U3086), .C2(n7001), .ZN(P1_U3349) );
  OAI222_X1 U8630 ( .A1(n7007), .A2(P1_U3086), .B1(n9864), .B2(n6851), .C1(
        n6850), .C2(n9866), .ZN(P1_U3354) );
  INV_X1 U8631 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6853) );
  OAI222_X1 U8632 ( .A1(n8387), .A2(n6853), .B1(n7852), .B2(n6007), .C1(
        P2_U3151), .C2(n6852), .ZN(P2_U3291) );
  OAI222_X1 U8633 ( .A1(n8387), .A2(n6855), .B1(n7852), .B2(n6856), .C1(
        P2_U3151), .C2(n6854), .ZN(P2_U3290) );
  OAI222_X1 U8634 ( .A1(n9866), .A2(n6857), .B1(n9864), .B2(n6856), .C1(
        P1_U3086), .C2(n7015), .ZN(P1_U3350) );
  INV_X1 U8635 ( .A(n6858), .ZN(n6867) );
  INV_X1 U8636 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6859) );
  OAI222_X1 U8637 ( .A1(n7852), .A2(n6867), .B1(n7444), .B2(P2_U3151), .C1(
        n6859), .C2(n8387), .ZN(P2_U3285) );
  NAND2_X1 U8638 ( .A1(n10003), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6861) );
  OAI21_X1 U8639 ( .B1(n10003), .B2(n6862), .A(n6861), .ZN(P1_U3440) );
  INV_X1 U8640 ( .A(n6863), .ZN(n6865) );
  OAI222_X1 U8641 ( .A1(n8387), .A2(n6864), .B1(n7852), .B2(n6865), .C1(
        P2_U3151), .C2(n7187), .ZN(P2_U3287) );
  INV_X1 U8642 ( .A(n9474), .ZN(n7004) );
  OAI222_X1 U8643 ( .A1(n9866), .A2(n6866), .B1(n9864), .B2(n6865), .C1(
        P1_U3086), .C2(n7004), .ZN(P1_U3347) );
  INV_X1 U8644 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6868) );
  INV_X1 U8645 ( .A(n7415), .ZN(n7422) );
  OAI222_X1 U8646 ( .A1(n9866), .A2(n6868), .B1(n9864), .B2(n6867), .C1(n7422), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  OAI222_X1 U8647 ( .A1(n9864), .A2(n6007), .B1(P1_U3086), .B2(n7094), .C1(
        n9866), .C2(n6006), .ZN(P1_U3351) );
  INV_X1 U8648 ( .A(n6869), .ZN(n6882) );
  OAI222_X1 U8649 ( .A1(n7852), .A2(n6882), .B1(n7465), .B2(P2_U3151), .C1(
        n6870), .C2(n8387), .ZN(P2_U3286) );
  INV_X1 U8650 ( .A(n8354), .ZN(n6873) );
  AOI21_X1 U8651 ( .B1(n6873), .B2(n6872), .A(n4464), .ZN(n6875) );
  INV_X1 U8652 ( .A(n6875), .ZN(n6874) );
  NAND2_X1 U8653 ( .A1(n8374), .A2(n8378), .ZN(n6876) );
  INV_X1 U8654 ( .A(n9960), .ZN(n9552) );
  NOR2_X1 U8655 ( .A1(n9552), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8656 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U8657 ( .A1(n6876), .A2(n6875), .ZN(n7026) );
  INV_X1 U8658 ( .A(n7026), .ZN(n6879) );
  INV_X1 U8659 ( .A(n9862), .ZN(n7067) );
  INV_X1 U8660 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10182) );
  AOI21_X1 U8661 ( .B1(n7067), .B2(n10182), .A(n4319), .ZN(n7069) );
  OAI21_X1 U8662 ( .B1(n7067), .B2(P1_REG1_REG_0__SCAN_IN), .A(n7069), .ZN(
        n6877) );
  XNOR2_X1 U8663 ( .A(n6877), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6878) );
  AOI22_X1 U8664 ( .A1(n6879), .A2(n6878), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6880) );
  OAI21_X1 U8665 ( .B1(n9960), .B2(n6881), .A(n6880), .ZN(P1_U3243) );
  INV_X1 U8666 ( .A(n7242), .ZN(n7248) );
  OAI222_X1 U8667 ( .A1(n9866), .A2(n6883), .B1(n9864), .B2(n6882), .C1(n7248), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  NAND2_X1 U8668 ( .A1(n8348), .A2(P1_U3973), .ZN(n6884) );
  OAI21_X1 U8669 ( .B1(P1_U3973), .B2(n9177), .A(n6884), .ZN(P1_U3585) );
  NAND2_X1 U8670 ( .A1(n7131), .A2(P1_U3973), .ZN(n6885) );
  OAI21_X1 U8671 ( .B1(P1_U3973), .B2(n5036), .A(n6885), .ZN(P1_U3554) );
  NAND2_X1 U8672 ( .A1(P2_U3893), .A2(n7153), .ZN(n6886) );
  OAI21_X1 U8673 ( .B1(P2_U3893), .B2(n6006), .A(n6886), .ZN(P2_U3495) );
  INV_X1 U8674 ( .A(n6887), .ZN(n6889) );
  OAI222_X1 U8675 ( .A1(n8387), .A2(n6888), .B1(n7852), .B2(n6889), .C1(
        P2_U3151), .C2(n8648), .ZN(P2_U3284) );
  INV_X1 U8676 ( .A(n7517), .ZN(n7514) );
  OAI222_X1 U8677 ( .A1(n9866), .A2(n6890), .B1(n9864), .B2(n6889), .C1(
        P1_U3086), .C2(n7514), .ZN(P1_U3344) );
  NAND2_X1 U8678 ( .A1(n6892), .A2(n6891), .ZN(n8383) );
  INV_X1 U8679 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6893) );
  NOR2_X1 U8680 ( .A1(n6935), .A2(n6893), .ZN(P2_U3246) );
  INV_X1 U8681 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6894) );
  NOR2_X1 U8682 ( .A1(n6935), .A2(n6894), .ZN(P2_U3257) );
  INV_X1 U8683 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6895) );
  NOR2_X1 U8684 ( .A1(n6935), .A2(n6895), .ZN(P2_U3249) );
  INV_X1 U8685 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6896) );
  NOR2_X1 U8686 ( .A1(n6935), .A2(n6896), .ZN(P2_U3248) );
  INV_X1 U8687 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6897) );
  NOR2_X1 U8688 ( .A1(n6935), .A2(n6897), .ZN(P2_U3250) );
  INV_X1 U8689 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6898) );
  NOR2_X1 U8690 ( .A1(n6935), .A2(n6898), .ZN(P2_U3251) );
  INV_X1 U8691 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6899) );
  NOR2_X1 U8692 ( .A1(n6935), .A2(n6899), .ZN(P2_U3254) );
  INV_X1 U8693 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6900) );
  NOR2_X1 U8694 ( .A1(n6935), .A2(n6900), .ZN(P2_U3247) );
  INV_X1 U8695 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6901) );
  NOR2_X1 U8696 ( .A1(n6935), .A2(n6901), .ZN(P2_U3255) );
  INV_X1 U8697 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6902) );
  NOR2_X1 U8698 ( .A1(n6935), .A2(n6902), .ZN(P2_U3253) );
  INV_X1 U8699 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6903) );
  NOR2_X1 U8700 ( .A1(n6935), .A2(n6903), .ZN(P2_U3256) );
  INV_X1 U8701 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6904) );
  NOR2_X1 U8702 ( .A1(n6935), .A2(n6904), .ZN(P2_U3252) );
  NAND2_X1 U8703 ( .A1(n9221), .A2(P1_U3973), .ZN(n6905) );
  OAI21_X1 U8704 ( .B1(n5399), .B2(P1_U3973), .A(n6905), .ZN(P1_U3574) );
  INV_X1 U8705 ( .A(n6051), .ZN(n6907) );
  OAI222_X1 U8706 ( .A1(n7852), .A2(n6907), .B1(n7798), .B2(P2_U3151), .C1(
        n6906), .C2(n8387), .ZN(P2_U3283) );
  INV_X1 U8707 ( .A(n9489), .ZN(n9482) );
  OAI222_X1 U8708 ( .A1(n9866), .A2(n6908), .B1(n9864), .B2(n6907), .C1(n9482), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8709 ( .A(n6909), .ZN(n6918) );
  INV_X1 U8710 ( .A(n9866), .ZN(n7198) );
  AOI22_X1 U8711 ( .A1(n9501), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7198), .ZN(n6910) );
  OAI21_X1 U8712 ( .B1(n6918), .B2(n9864), .A(n6910), .ZN(P1_U3342) );
  NAND2_X1 U8713 ( .A1(n8890), .A2(P2_U3893), .ZN(n6911) );
  OAI21_X1 U8714 ( .B1(P2_U3893), .B2(n5377), .A(n6911), .ZN(P2_U3510) );
  INV_X1 U8715 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6917) );
  INV_X1 U8716 ( .A(n10111), .ZN(n8629) );
  AOI22_X1 U8717 ( .A1(n8629), .A2(P2_IR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n6916) );
  OAI21_X1 U8718 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6912), .A(n6969), .ZN(n6913) );
  OAI21_X1 U8719 ( .B1(n6751), .B2(n6914), .A(n6913), .ZN(n6915) );
  OAI211_X1 U8720 ( .C1(n6917), .C2(n8748), .A(n6916), .B(n6915), .ZN(P2_U3182) );
  INV_X1 U8721 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10272) );
  OAI222_X1 U8722 ( .A1(n8387), .A2(n10272), .B1(n7852), .B2(n6918), .C1(
        P2_U3151), .C2(n8665), .ZN(P2_U3282) );
  OAI211_X1 U8723 ( .C1(n6921), .C2(n6920), .A(n6919), .B(n6751), .ZN(n6932)
         );
  XOR2_X1 U8724 ( .A(n6923), .B(P2_REG1_REG_5__SCAN_IN), .Z(n6924) );
  NOR2_X1 U8725 ( .A1(n10106), .A2(n6924), .ZN(n6929) );
  INV_X1 U8726 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U8727 ( .A1(n8629), .A2(n6925), .ZN(n6926) );
  NAND2_X1 U8728 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7311) );
  OAI211_X1 U8729 ( .C1(n6927), .C2(n8748), .A(n6926), .B(n7311), .ZN(n6928)
         );
  AOI211_X1 U8730 ( .C1(n10114), .C2(n6930), .A(n6929), .B(n6928), .ZN(n6931)
         );
  NAND2_X1 U8731 ( .A1(n6932), .A2(n6931), .ZN(P2_U3187) );
  INV_X1 U8732 ( .A(n6933), .ZN(n6962) );
  AOI22_X1 U8733 ( .A1(n9927), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7198), .ZN(n6934) );
  OAI21_X1 U8734 ( .B1(n6962), .B2(n9864), .A(n6934), .ZN(P1_U3341) );
  INV_X1 U8735 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6936) );
  NOR2_X1 U8736 ( .A1(n6935), .A2(n6936), .ZN(P2_U3238) );
  INV_X1 U8737 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6937) );
  NOR2_X1 U8738 ( .A1(n6935), .A2(n6937), .ZN(P2_U3235) );
  INV_X1 U8739 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6938) );
  NOR2_X1 U8740 ( .A1(n6935), .A2(n6938), .ZN(P2_U3239) );
  INV_X1 U8741 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6939) );
  NOR2_X1 U8742 ( .A1(n6935), .A2(n6939), .ZN(P2_U3240) );
  INV_X1 U8743 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6940) );
  NOR2_X1 U8744 ( .A1(n6935), .A2(n6940), .ZN(P2_U3263) );
  INV_X1 U8745 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6941) );
  NOR2_X1 U8746 ( .A1(n6935), .A2(n6941), .ZN(P2_U3262) );
  INV_X1 U8747 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6942) );
  NOR2_X1 U8748 ( .A1(n6935), .A2(n6942), .ZN(P2_U3261) );
  INV_X1 U8749 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6943) );
  NOR2_X1 U8750 ( .A1(n6935), .A2(n6943), .ZN(P2_U3260) );
  INV_X1 U8751 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6944) );
  NOR2_X1 U8752 ( .A1(n6935), .A2(n6944), .ZN(P2_U3259) );
  INV_X1 U8753 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6945) );
  NOR2_X1 U8754 ( .A1(n6935), .A2(n6945), .ZN(P2_U3258) );
  INV_X1 U8755 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6946) );
  NOR2_X1 U8756 ( .A1(n6935), .A2(n6946), .ZN(P2_U3241) );
  INV_X1 U8757 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6947) );
  NOR2_X1 U8758 ( .A1(n6935), .A2(n6947), .ZN(P2_U3234) );
  INV_X1 U8759 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6948) );
  NOR2_X1 U8760 ( .A1(n6935), .A2(n6948), .ZN(P2_U3244) );
  INV_X1 U8761 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6949) );
  NOR2_X1 U8762 ( .A1(n6935), .A2(n6949), .ZN(P2_U3236) );
  INV_X1 U8763 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6950) );
  NOR2_X1 U8764 ( .A1(n6935), .A2(n6950), .ZN(P2_U3245) );
  INV_X1 U8765 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6951) );
  NOR2_X1 U8766 ( .A1(n6935), .A2(n6951), .ZN(P2_U3243) );
  INV_X1 U8767 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6952) );
  NOR2_X1 U8768 ( .A1(n6935), .A2(n6952), .ZN(P2_U3242) );
  INV_X1 U8769 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6953) );
  NOR2_X1 U8770 ( .A1(n6935), .A2(n6953), .ZN(P2_U3237) );
  XNOR2_X1 U8771 ( .A(n6954), .B(n4433), .ZN(n9006) );
  XNOR2_X1 U8772 ( .A(n6955), .B(n4433), .ZN(n6957) );
  INV_X1 U8773 ( .A(n8609), .ZN(n7215) );
  INV_X1 U8774 ( .A(n8607), .ZN(n7234) );
  OAI22_X1 U8775 ( .A1(n7215), .A2(n8971), .B1(n7234), .B2(n8969), .ZN(n6956)
         );
  AOI21_X1 U8776 ( .B1(n6957), .B2(n8949), .A(n6956), .ZN(n6958) );
  OAI21_X1 U8777 ( .B1(n9006), .B2(n7687), .A(n6958), .ZN(n9000) );
  OAI22_X1 U8778 ( .A1(n9006), .A2(n7103), .B1(n6959), .B2(n7407), .ZN(n6960)
         );
  NOR2_X1 U8779 ( .A1(n9000), .A2(n6960), .ZN(n10123) );
  NAND2_X1 U8780 ( .A1(n9073), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6961) );
  OAI21_X1 U8781 ( .B1(n10123), .B2(n9073), .A(n6961), .ZN(P2_U3461) );
  INV_X1 U8782 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6963) );
  OAI222_X1 U8783 ( .A1(n8387), .A2(n6963), .B1(n7852), .B2(n6962), .C1(
        P2_U3151), .C2(n8686), .ZN(P2_U3281) );
  INV_X1 U8784 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6979) );
  NAND2_X1 U8785 ( .A1(n6965), .A2(n6964), .ZN(n6966) );
  AOI21_X1 U8786 ( .B1(n6967), .B2(n6966), .A(n8668), .ZN(n6973) );
  OAI211_X1 U8787 ( .C1(n6970), .C2(n6969), .A(n6751), .B(n6968), .ZN(n6971)
         );
  OAI21_X1 U8788 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7149), .A(n6971), .ZN(n6972) );
  NOR2_X1 U8789 ( .A1(n6973), .A2(n6972), .ZN(n6978) );
  INV_X1 U8790 ( .A(n10106), .ZN(n10095) );
  XNOR2_X1 U8791 ( .A(n6974), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6975) );
  AOI22_X1 U8792 ( .A1(n6976), .A2(n8629), .B1(n10095), .B2(n6975), .ZN(n6977)
         );
  OAI211_X1 U8793 ( .C1(n8748), .C2(n6979), .A(n6978), .B(n6977), .ZN(P2_U3183) );
  INV_X1 U8794 ( .A(n6980), .ZN(n6984) );
  NAND4_X1 U8795 ( .A1(n6984), .A2(n6983), .A3(n6982), .A4(n6981), .ZN(n6988)
         );
  INV_X1 U8796 ( .A(n6988), .ZN(n6985) );
  NAND3_X1 U8797 ( .A1(n7218), .A2(n6986), .A3(n7407), .ZN(n6987) );
  NAND2_X1 U8798 ( .A1(n8954), .A2(n8609), .ZN(n7100) );
  OAI211_X1 U8799 ( .C1(n8989), .C2(n7220), .A(n6987), .B(n7100), .ZN(n6989)
         );
  MUX2_X1 U8800 ( .A(n6989), .B(P2_REG2_REG_0__SCAN_IN), .S(n8993), .Z(n6990)
         );
  AOI21_X1 U8801 ( .B1(n8977), .B2(n6991), .A(n6990), .ZN(n6992) );
  INV_X1 U8802 ( .A(n6992), .ZN(P2_U3233) );
  INV_X1 U8803 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7010) );
  AND2_X1 U8804 ( .A1(n7131), .A2(n6994), .ZN(n8287) );
  OR2_X1 U8805 ( .A1(n8287), .A2(n7129), .ZN(n8248) );
  OAI21_X1 U8806 ( .B1(n9962), .B2(n10026), .A(n8248), .ZN(n6993) );
  OAI211_X1 U8807 ( .C1(n6994), .C2(n7321), .A(n6993), .B(n7322), .ZN(n7138)
         );
  NAND2_X1 U8808 ( .A1(n7138), .A2(n10064), .ZN(n6995) );
  OAI21_X1 U8809 ( .B1(n10064), .B2(n7010), .A(n6995), .ZN(P1_U3522) );
  INV_X1 U8810 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6996) );
  MUX2_X1 U8811 ( .A(n6996), .B(P1_REG2_REG_9__SCAN_IN), .S(n7242), .Z(n7006)
         );
  INV_X1 U8812 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7551) );
  INV_X1 U8813 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7002) );
  INV_X1 U8814 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7299) );
  INV_X1 U8815 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6999) );
  INV_X1 U8816 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6998) );
  INV_X1 U8817 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6997) );
  MUX2_X1 U8818 ( .A(n6997), .B(P1_REG2_REG_1__SCAN_IN), .S(n7007), .Z(n9413)
         );
  NAND2_X1 U8819 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7068) );
  INV_X1 U8820 ( .A(n7068), .ZN(n9412) );
  NAND2_X1 U8821 ( .A1(n9413), .A2(n9412), .ZN(n9411) );
  OAI21_X1 U8822 ( .B1(n7007), .B2(n6997), .A(n9411), .ZN(n7073) );
  MUX2_X1 U8823 ( .A(n6998), .B(P1_REG2_REG_2__SCAN_IN), .S(n7080), .Z(n7074)
         );
  NAND2_X1 U8824 ( .A1(n7073), .A2(n7074), .ZN(n7072) );
  OAI21_X1 U8825 ( .B1(n7080), .B2(n6998), .A(n7072), .ZN(n9425) );
  MUX2_X1 U8826 ( .A(n6999), .B(P1_REG2_REG_3__SCAN_IN), .S(n7871), .Z(n9426)
         );
  NAND2_X1 U8827 ( .A1(n9425), .A2(n9426), .ZN(n9424) );
  OAI21_X1 U8828 ( .B1(n6999), .B2(n7871), .A(n9424), .ZN(n7088) );
  MUX2_X1 U8829 ( .A(n7299), .B(P1_REG2_REG_4__SCAN_IN), .S(n7094), .Z(n7089)
         );
  NAND2_X1 U8830 ( .A1(n7088), .A2(n7089), .ZN(n7087) );
  INV_X1 U8831 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7000) );
  MUX2_X1 U8832 ( .A(n7000), .B(P1_REG2_REG_5__SCAN_IN), .S(n7015), .Z(n9438)
         );
  MUX2_X1 U8833 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7002), .S(n9448), .Z(n9451)
         );
  OAI21_X1 U8834 ( .B1(n7002), .B2(n7001), .A(n9449), .ZN(n9463) );
  XOR2_X1 U8835 ( .A(n9461), .B(P1_REG2_REG_7__SCAN_IN), .Z(n9464) );
  MUX2_X1 U8836 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7551), .S(n9474), .Z(n9477)
         );
  NOR2_X1 U8837 ( .A1(n7005), .A2(n7006), .ZN(n7247) );
  AOI21_X1 U8838 ( .B1(n7006), .B2(n7005), .A(n7247), .ZN(n7030) );
  OR2_X1 U8839 ( .A1(n4319), .A2(n9862), .ZN(n8372) );
  INV_X1 U8840 ( .A(n7871), .ZN(n9423) );
  INV_X1 U8841 ( .A(n7007), .ZN(n9410) );
  INV_X1 U8842 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7008) );
  MUX2_X1 U8843 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n7008), .S(n7007), .Z(n9405)
         );
  INV_X1 U8844 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7009) );
  AOI21_X1 U8845 ( .B1(n9410), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9404), .ZN(
        n7078) );
  INV_X1 U8846 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7011) );
  MUX2_X1 U8847 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n7011), .S(n7080), .Z(n7077)
         );
  INV_X1 U8848 ( .A(n7080), .ZN(n7012) );
  INV_X1 U8849 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7013) );
  MUX2_X1 U8850 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7013), .S(n7871), .Z(n9418)
         );
  INV_X1 U8851 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7014) );
  MUX2_X1 U8852 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7014), .S(n7094), .Z(n7085)
         );
  MUX2_X1 U8853 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7016), .S(n7015), .Z(n9431)
         );
  INV_X1 U8854 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7016) );
  INV_X1 U8855 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7018) );
  MUX2_X1 U8856 ( .A(n7018), .B(P1_REG1_REG_6__SCAN_IN), .S(n9448), .Z(n9442)
         );
  XNOR2_X1 U8857 ( .A(n9461), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n9456) );
  INV_X1 U8858 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7019) );
  MUX2_X1 U8859 ( .A(n7019), .B(P1_REG1_REG_8__SCAN_IN), .S(n9474), .Z(n9469)
         );
  INV_X1 U8860 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7021) );
  MUX2_X1 U8861 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7021), .S(n7242), .Z(n7022)
         );
  OAI21_X1 U8862 ( .B1(n7023), .B2(n7022), .A(n7241), .ZN(n7024) );
  INV_X1 U8863 ( .A(n9944), .ZN(n9545) );
  NAND2_X1 U8864 ( .A1(n7024), .A2(n9545), .ZN(n7029) );
  OR2_X1 U8865 ( .A1(n7026), .A2(n7025), .ZN(n7095) );
  NAND2_X1 U8866 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9287) );
  OAI21_X1 U8867 ( .B1(n9960), .B2(n9893), .A(n9287), .ZN(n7027) );
  AOI21_X1 U8868 ( .B1(n7242), .B2(n9947), .A(n7027), .ZN(n7028) );
  OAI211_X1 U8869 ( .C1(n7030), .C2(n9934), .A(n7029), .B(n7028), .ZN(P1_U3252) );
  INV_X1 U8870 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7032) );
  INV_X1 U8871 ( .A(n7031), .ZN(n7034) );
  OAI222_X1 U8872 ( .A1(n9866), .A2(n7032), .B1(n9864), .B2(n7034), .C1(
        P1_U3086), .C2(n9505), .ZN(P1_U3340) );
  INV_X1 U8873 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7035) );
  OAI222_X1 U8874 ( .A1(n8387), .A2(n7035), .B1(n7852), .B2(n7034), .C1(
        P2_U3151), .C2(n4894), .ZN(P2_U3280) );
  OR2_X1 U8875 ( .A1(n7036), .A2(n7328), .ZN(n9007) );
  NOR2_X1 U8876 ( .A1(n8993), .A2(n9007), .ZN(n8997) );
  NAND2_X1 U8877 ( .A1(n7037), .A2(n7038), .ZN(n7039) );
  NAND2_X1 U8878 ( .A1(n7040), .A2(n7039), .ZN(n7104) );
  OAI22_X1 U8879 ( .A1(n8991), .A2(n7145), .B1(n8989), .B2(n7149), .ZN(n7049)
         );
  INV_X1 U8880 ( .A(n7042), .ZN(n7043) );
  XNOR2_X1 U8881 ( .A(n7037), .B(n7043), .ZN(n7047) );
  INV_X1 U8882 ( .A(n7687), .ZN(n7044) );
  NAND2_X1 U8883 ( .A1(n7104), .A2(n7044), .ZN(n7046) );
  AOI22_X1 U8884 ( .A1(n8952), .A2(n8610), .B1(n8954), .B2(n8608), .ZN(n7045)
         );
  OAI211_X1 U8885 ( .C1(n8967), .C2(n7047), .A(n7046), .B(n7045), .ZN(n7107)
         );
  MUX2_X1 U8886 ( .A(n7107), .B(P2_REG2_REG_1__SCAN_IN), .S(n8993), .Z(n7048)
         );
  AOI211_X1 U8887 ( .C1(n8997), .C2(n7104), .A(n7049), .B(n7048), .ZN(n7050)
         );
  INV_X1 U8888 ( .A(n7050), .ZN(P2_U3232) );
  OAI21_X1 U8889 ( .B1(n7051), .B2(n7053), .A(n7052), .ZN(n9980) );
  OAI211_X1 U8890 ( .C1(n4975), .C2(n6374), .A(n10012), .B(n7054), .ZN(n9983)
         );
  OAI21_X1 U8891 ( .B1(n6374), .B2(n10020), .A(n9983), .ZN(n7061) );
  XNOR2_X1 U8892 ( .A(n7055), .B(n7051), .ZN(n7060) );
  OR2_X1 U8893 ( .A1(n7056), .A2(n9712), .ZN(n7058) );
  NAND2_X1 U8894 ( .A1(n7058), .A2(n7057), .ZN(n7900) );
  INV_X1 U8895 ( .A(n7900), .ZN(n7059) );
  OAI21_X1 U8896 ( .B1(n7060), .B2(n9708), .A(n7059), .ZN(n9978) );
  AOI211_X1 U8897 ( .C1(n10026), .C2(n9980), .A(n7061), .B(n9978), .ZN(n7282)
         );
  NAND2_X1 U8898 ( .A1(n10062), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7062) );
  OAI21_X1 U8899 ( .B1(n7282), .B2(n10062), .A(n7062), .ZN(P1_U3524) );
  OR2_X1 U8900 ( .A1(n7064), .A2(n7063), .ZN(n7065) );
  AND2_X1 U8901 ( .A1(n7066), .A2(n7065), .ZN(n7275) );
  NOR3_X1 U8902 ( .A1(n7275), .A2(n7067), .A3(n4319), .ZN(n7071) );
  OAI22_X1 U8903 ( .A1(n7069), .A2(P1_IR_REG_0__SCAN_IN), .B1(n7068), .B2(
        n8372), .ZN(n7070) );
  NOR3_X1 U8904 ( .A1(n7071), .A2(n9403), .A3(n7070), .ZN(n7099) );
  OAI211_X1 U8905 ( .C1(n7074), .C2(n7073), .A(n9951), .B(n7072), .ZN(n7075)
         );
  INV_X1 U8906 ( .A(n7075), .ZN(n7083) );
  AOI211_X1 U8907 ( .C1(n7078), .C2(n7077), .A(n7076), .B(n9944), .ZN(n7082)
         );
  AOI22_X1 U8908 ( .A1(n9552), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7079) );
  OAI21_X1 U8909 ( .B1(n7080), .B2(n7095), .A(n7079), .ZN(n7081) );
  OR4_X1 U8910 ( .A1(n7099), .A2(n7083), .A3(n7082), .A4(n7081), .ZN(P1_U3245)
         );
  AOI211_X1 U8911 ( .C1(n7086), .C2(n7085), .A(n9944), .B(n7084), .ZN(n7098)
         );
  OAI211_X1 U8912 ( .C1(n7089), .C2(n7088), .A(n9951), .B(n7087), .ZN(n7090)
         );
  INV_X1 U8913 ( .A(n7090), .ZN(n7097) );
  INV_X1 U8914 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7091) );
  OR2_X1 U8915 ( .A1(n9960), .A2(n7091), .ZN(n7093) );
  OAI211_X1 U8916 ( .C1(n7095), .C2(n7094), .A(n7093), .B(n7092), .ZN(n7096)
         );
  OR4_X1 U8917 ( .A1(n7099), .A2(n7098), .A3(n7097), .A4(n7096), .ZN(P1_U3247)
         );
  OAI21_X1 U8918 ( .B1(n7501), .B2(n8949), .A(n7218), .ZN(n7101) );
  OAI211_X1 U8919 ( .C1(n7407), .C2(n7216), .A(n7101), .B(n7100), .ZN(n9074)
         );
  NAND2_X1 U8920 ( .A1(n5734), .A2(n9074), .ZN(n7102) );
  OAI21_X1 U8921 ( .B1(n5734), .B2(n5031), .A(n7102), .ZN(P2_U3390) );
  INV_X1 U8922 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7108) );
  INV_X1 U8923 ( .A(n7103), .ZN(n7689) );
  NAND2_X1 U8924 ( .A1(n7104), .A2(n7689), .ZN(n7105) );
  OAI21_X1 U8925 ( .B1(n7145), .B2(n7407), .A(n7105), .ZN(n7106) );
  NOR2_X1 U8926 ( .A1(n7107), .A2(n7106), .ZN(n10122) );
  MUX2_X1 U8927 ( .A(n7108), .B(n10122), .S(n4313), .Z(n7109) );
  INV_X1 U8928 ( .A(n7109), .ZN(P2_U3460) );
  XNOR2_X1 U8929 ( .A(n7110), .B(n7113), .ZN(n7158) );
  AOI21_X1 U8930 ( .B1(n6955), .B2(n4433), .A(n7111), .ZN(n7114) );
  XNOR2_X1 U8931 ( .A(n7114), .B(n7113), .ZN(n7115) );
  AOI222_X1 U8932 ( .A1(n8949), .A2(n7115), .B1(n7153), .B2(n8954), .C1(n8608), 
        .C2(n8952), .ZN(n7159) );
  OAI21_X1 U8933 ( .B1(n7116), .B2(n7407), .A(n7159), .ZN(n7117) );
  AOI21_X1 U8934 ( .B1(n7158), .B2(n7501), .A(n7117), .ZN(n10125) );
  OR2_X1 U8935 ( .A1(n4313), .A2(n10065), .ZN(n7118) );
  OAI21_X1 U8936 ( .B1(n10125), .B2(n9073), .A(n7118), .ZN(P2_U3462) );
  INV_X1 U8937 ( .A(n7119), .ZN(n7127) );
  AOI22_X1 U8938 ( .A1(n9522), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7198), .ZN(n7120) );
  OAI21_X1 U8939 ( .B1(n7127), .B2(n9864), .A(n7120), .ZN(P1_U3339) );
  NAND2_X1 U8940 ( .A1(n7052), .A2(n7121), .ZN(n7122) );
  NAND2_X1 U8941 ( .A1(n7122), .A2(n8246), .ZN(n7286) );
  OAI21_X1 U8942 ( .B1(n7122), .B2(n8246), .A(n7286), .ZN(n7434) );
  OAI211_X1 U8943 ( .C1(n6002), .C2(n7257), .A(n10012), .B(n7300), .ZN(n7432)
         );
  OAI21_X1 U8944 ( .B1(n7257), .B2(n10020), .A(n7432), .ZN(n7124) );
  XOR2_X1 U8945 ( .A(n8141), .B(n8246), .Z(n7123) );
  OAI222_X1 U8946 ( .A1(n9710), .A2(n6582), .B1(n9712), .B2(n7491), .C1(n9708), 
        .C2(n7123), .ZN(n7428) );
  AOI211_X1 U8947 ( .C1(n10026), .C2(n7434), .A(n7124), .B(n7428), .ZN(n7279)
         );
  NAND2_X1 U8948 ( .A1(n10062), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7125) );
  OAI21_X1 U8949 ( .B1(n7279), .B2(n10062), .A(n7125), .ZN(P1_U3525) );
  INV_X1 U8950 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7126) );
  OAI222_X1 U8951 ( .A1(n7852), .A2(n7127), .B1(P2_U3151), .B2(n8714), .C1(
        n7126), .C2(n8387), .ZN(P2_U3279) );
  INV_X1 U8952 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7137) );
  XOR2_X1 U8953 ( .A(n8249), .B(n7128), .Z(n9997) );
  INV_X1 U8954 ( .A(n9997), .ZN(n7135) );
  INV_X1 U8955 ( .A(n7835), .ZN(n10036) );
  XOR2_X1 U8956 ( .A(n8249), .B(n7129), .Z(n7132) );
  AOI22_X1 U8957 ( .A1(n7130), .A2(n9675), .B1(n9673), .B2(n7131), .ZN(n7269)
         );
  OAI21_X1 U8958 ( .B1(n7132), .B2(n9708), .A(n7269), .ZN(n7133) );
  AOI21_X1 U8959 ( .B1(n10036), .B2(n9997), .A(n7133), .ZN(n10000) );
  AOI211_X1 U8960 ( .C1(n7320), .C2(n7271), .A(n9724), .B(n4975), .ZN(n9992)
         );
  AOI21_X1 U8961 ( .B1(n10047), .B2(n7271), .A(n9992), .ZN(n7134) );
  OAI211_X1 U8962 ( .C1(n10031), .C2(n7135), .A(n10000), .B(n7134), .ZN(n9835)
         );
  NAND2_X1 U8963 ( .A1(n9835), .A2(n10055), .ZN(n7136) );
  OAI21_X1 U8964 ( .B1(n10055), .B2(n7137), .A(n7136), .ZN(P1_U3456) );
  INV_X1 U8965 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7140) );
  NAND2_X1 U8966 ( .A1(n7138), .A2(n10055), .ZN(n7139) );
  OAI21_X1 U8967 ( .B1(n10055), .B2(n7140), .A(n7139), .ZN(P1_U3453) );
  NOR2_X1 U8968 ( .A1(n8593), .A2(P2_U3151), .ZN(n7221) );
  OAI21_X1 U8969 ( .B1(n7143), .B2(n7142), .A(n7141), .ZN(n7147) );
  AOI22_X1 U8970 ( .A1(n8572), .A2(n8610), .B1(n8587), .B2(n8608), .ZN(n7144)
         );
  OAI21_X1 U8971 ( .B1(n7145), .B2(n8596), .A(n7144), .ZN(n7146) );
  AOI21_X1 U8972 ( .B1(n8557), .B2(n7147), .A(n7146), .ZN(n7148) );
  OAI21_X1 U8973 ( .B1(n7221), .B2(n7149), .A(n7148), .ZN(P2_U3162) );
  XNOR2_X1 U8974 ( .A(n7150), .B(n7151), .ZN(n7200) );
  INV_X1 U8975 ( .A(n7204), .ZN(n7313) );
  XNOR2_X1 U8976 ( .A(n7152), .B(n7151), .ZN(n7154) );
  AOI222_X1 U8977 ( .A1(n8949), .A2(n7154), .B1(n8605), .B2(n8954), .C1(n7153), 
        .C2(n8952), .ZN(n7201) );
  OAI21_X1 U8978 ( .B1(n7313), .B2(n7407), .A(n7201), .ZN(n7155) );
  AOI21_X1 U8979 ( .B1(n7501), .B2(n7200), .A(n7155), .ZN(n10128) );
  OR2_X1 U8980 ( .A1(n4313), .A2(n5104), .ZN(n7156) );
  OAI21_X1 U8981 ( .B1(n10128), .B2(n9073), .A(n7156), .ZN(P2_U3464) );
  NAND2_X1 U8982 ( .A1(n7687), .A2(n9007), .ZN(n7157) );
  INV_X1 U8983 ( .A(n7158), .ZN(n7163) );
  MUX2_X1 U8984 ( .A(n7160), .B(n7159), .S(n9008), .Z(n7162) );
  AOI22_X1 U8985 ( .A1(n8977), .A2(n7222), .B1(n9003), .B2(n7229), .ZN(n7161)
         );
  OAI211_X1 U8986 ( .C1(n8980), .C2(n7163), .A(n7162), .B(n7161), .ZN(P2_U3230) );
  XNOR2_X1 U8987 ( .A(n7164), .B(n7166), .ZN(n7195) );
  INV_X1 U8988 ( .A(n7195), .ZN(n7173) );
  XOR2_X1 U8989 ( .A(n7166), .B(n7165), .Z(n7167) );
  AOI222_X1 U8990 ( .A1(n8949), .A2(n7167), .B1(n8606), .B2(n8954), .C1(n8607), 
        .C2(n8952), .ZN(n7193) );
  MUX2_X1 U8991 ( .A(n7168), .B(n7193), .S(n9008), .Z(n7172) );
  INV_X1 U8992 ( .A(n7239), .ZN(n7169) );
  AOI22_X1 U8993 ( .A1(n8977), .A2(n7170), .B1(n9003), .B2(n7169), .ZN(n7171)
         );
  OAI211_X1 U8994 ( .C1(n8980), .C2(n7173), .A(n7172), .B(n7171), .ZN(P2_U3229) );
  INV_X1 U8995 ( .A(n7174), .ZN(n7263) );
  AOI22_X1 U8996 ( .A1(n9540), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7198), .ZN(n7175) );
  OAI21_X1 U8997 ( .B1(n7263), .B2(n9864), .A(n7175), .ZN(P1_U3338) );
  XOR2_X1 U8998 ( .A(n7176), .B(n7177), .Z(n7192) );
  XNOR2_X1 U8999 ( .A(n7179), .B(n7178), .ZN(n7190) );
  INV_X1 U9000 ( .A(n7180), .ZN(n7185) );
  NAND3_X1 U9001 ( .A1(n7181), .A2(n7183), .A3(n7182), .ZN(n7184) );
  AOI21_X1 U9002 ( .B1(n7185), .B2(n7184), .A(n8668), .ZN(n7189) );
  NAND2_X1 U9003 ( .A1(n10118), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7186) );
  NAND2_X1 U9004 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7698) );
  OAI211_X1 U9005 ( .C1(n10111), .C2(n7187), .A(n7186), .B(n7698), .ZN(n7188)
         );
  AOI211_X1 U9006 ( .C1(n7190), .C2(n6751), .A(n7189), .B(n7188), .ZN(n7191)
         );
  OAI21_X1 U9007 ( .B1(n7192), .B2(n10106), .A(n7191), .ZN(P2_U3190) );
  OAI21_X1 U9008 ( .B1(n7235), .B2(n7407), .A(n7193), .ZN(n7194) );
  AOI21_X1 U9009 ( .B1(n7195), .B2(n7501), .A(n7194), .ZN(n10126) );
  NAND2_X1 U9010 ( .A1(n9073), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7196) );
  OAI21_X1 U9011 ( .B1(n10126), .B2(n9073), .A(n7196), .ZN(P2_U3463) );
  INV_X1 U9012 ( .A(n7197), .ZN(n7254) );
  AOI22_X1 U9013 ( .A1(n9948), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7198), .ZN(n7199) );
  OAI21_X1 U9014 ( .B1(n7254), .B2(n9864), .A(n7199), .ZN(P1_U3337) );
  INV_X1 U9015 ( .A(n7200), .ZN(n7207) );
  MUX2_X1 U9016 ( .A(n7202), .B(n7201), .S(n9008), .Z(n7206) );
  INV_X1 U9017 ( .A(n7319), .ZN(n7203) );
  AOI22_X1 U9018 ( .A1(n8977), .A2(n7204), .B1(n9003), .B2(n7203), .ZN(n7205)
         );
  OAI211_X1 U9019 ( .C1(n7207), .C2(n8980), .A(n7206), .B(n7205), .ZN(P2_U3228) );
  OAI21_X1 U9020 ( .B1(n7210), .B2(n7209), .A(n7208), .ZN(n7211) );
  NAND2_X1 U9021 ( .A1(n7211), .A2(n8557), .ZN(n7214) );
  OAI22_X1 U9022 ( .A1(n8575), .A2(n7234), .B1(n7215), .B2(n8590), .ZN(n7212)
         );
  AOI21_X1 U9023 ( .B1(n9001), .B2(n8578), .A(n7212), .ZN(n7213) );
  OAI211_X1 U9024 ( .C1(n7221), .C2(n8611), .A(n7214), .B(n7213), .ZN(P2_U3177) );
  OAI22_X1 U9025 ( .A1(n8596), .A2(n7216), .B1(n8575), .B2(n7215), .ZN(n7217)
         );
  AOI21_X1 U9026 ( .B1(n8557), .B2(n7218), .A(n7217), .ZN(n7219) );
  OAI21_X1 U9027 ( .B1(n7221), .B2(n7220), .A(n7219), .ZN(P2_U3172) );
  AOI22_X1 U9028 ( .A1(n8572), .A2(n8608), .B1(n8578), .B2(n7222), .ZN(n7223)
         );
  NAND2_X1 U9029 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10072) );
  OAI211_X1 U9030 ( .C1(n7312), .C2(n8575), .A(n7223), .B(n10072), .ZN(n7228)
         );
  AOI211_X1 U9031 ( .C1(n7226), .C2(n7225), .A(n8581), .B(n7224), .ZN(n7227)
         );
  AOI211_X1 U9032 ( .C1(n7229), .C2(n8593), .A(n7228), .B(n7227), .ZN(n7230)
         );
  INV_X1 U9033 ( .A(n7230), .ZN(P2_U3158) );
  OAI21_X1 U9034 ( .B1(n7232), .B2(n7231), .A(n7308), .ZN(n7233) );
  NAND2_X1 U9035 ( .A1(n7233), .A2(n8557), .ZN(n7238) );
  AND2_X1 U9036 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8628) );
  OAI22_X1 U9037 ( .A1(n8596), .A2(n7235), .B1(n7234), .B2(n8590), .ZN(n7236)
         );
  AOI211_X1 U9038 ( .C1(n8587), .C2(n8606), .A(n8628), .B(n7236), .ZN(n7237)
         );
  OAI211_X1 U9039 ( .C1(n7239), .C2(n7318), .A(n7238), .B(n7237), .ZN(P2_U3170) );
  INV_X1 U9040 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9896) );
  AND2_X1 U9041 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7792) );
  INV_X1 U9042 ( .A(n7792), .ZN(n7240) );
  OAI21_X1 U9043 ( .B1(n9960), .B2(n9896), .A(n7240), .ZN(n7246) );
  XNOR2_X1 U9044 ( .A(n7415), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7244) );
  AOI211_X1 U9045 ( .C1(n7244), .C2(n7243), .A(n9944), .B(n7417), .ZN(n7245)
         );
  AOI211_X1 U9046 ( .C1(n9947), .C2(n7415), .A(n7246), .B(n7245), .ZN(n7252)
         );
  XOR2_X1 U9047 ( .A(n7415), .B(P1_REG2_REG_10__SCAN_IN), .Z(n7249) );
  OAI211_X1 U9048 ( .C1(n7250), .C2(n7249), .A(n7421), .B(n9951), .ZN(n7251)
         );
  NAND2_X1 U9049 ( .A1(n7252), .A2(n7251), .ZN(P1_U3253) );
  OAI222_X1 U9050 ( .A1(n7852), .A2(n7254), .B1(n8744), .B2(P2_U3151), .C1(
        n7253), .C2(n8387), .ZN(P2_U3277) );
  XOR2_X1 U9051 ( .A(n7255), .B(n7256), .Z(n7262) );
  NAND2_X1 U9052 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9421) );
  OAI21_X1 U9053 ( .B1(n9366), .B2(n7257), .A(n9421), .ZN(n7259) );
  OAI22_X1 U9054 ( .A1(n7491), .A2(n9375), .B1(n9359), .B2(n6582), .ZN(n7258)
         );
  AOI211_X1 U9055 ( .C1(n7260), .C2(n9372), .A(n7259), .B(n7258), .ZN(n7261)
         );
  OAI21_X1 U9056 ( .B1(n7262), .B2(n9380), .A(n7261), .ZN(P1_U3218) );
  OAI222_X1 U9057 ( .A1(n8387), .A2(n7264), .B1(n7852), .B2(n7263), .C1(
        P2_U3151), .C2(n8727), .ZN(P2_U3278) );
  NAND2_X1 U9058 ( .A1(n9349), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7902) );
  INV_X1 U9059 ( .A(n7902), .ZN(n7274) );
  INV_X1 U9060 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9988) );
  OAI21_X1 U9061 ( .B1(n7265), .B2(n7266), .A(n7267), .ZN(n7268) );
  NAND2_X1 U9062 ( .A1(n7268), .A2(n9312), .ZN(n7273) );
  INV_X1 U9063 ( .A(n7269), .ZN(n7270) );
  AOI22_X1 U9064 ( .A1(n9378), .A2(n7271), .B1(n7270), .B2(n9269), .ZN(n7272)
         );
  OAI211_X1 U9065 ( .C1(n7274), .C2(n9988), .A(n7273), .B(n7272), .ZN(P1_U3222) );
  AOI22_X1 U9066 ( .A1(n9378), .A2(n7320), .B1(n7275), .B2(n9312), .ZN(n7277)
         );
  NAND2_X1 U9067 ( .A1(n7902), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7276) );
  OAI211_X1 U9068 ( .C1(n7278), .C2(n9375), .A(n7277), .B(n7276), .ZN(P1_U3232) );
  INV_X1 U9069 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7281) );
  OR2_X1 U9070 ( .A1(n7279), .A2(n10053), .ZN(n7280) );
  OAI21_X1 U9071 ( .B1(n10055), .B2(n7281), .A(n7280), .ZN(P1_U3462) );
  INV_X1 U9072 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7284) );
  OR2_X1 U9073 ( .A1(n7282), .A2(n10053), .ZN(n7283) );
  OAI21_X1 U9074 ( .B1(n10055), .B2(n7284), .A(n7283), .ZN(P1_U3459) );
  NAND2_X1 U9075 ( .A1(n7286), .A2(n7285), .ZN(n7288) );
  INV_X1 U9076 ( .A(n7287), .ZN(n8250) );
  XNOR2_X1 U9077 ( .A(n7288), .B(n8250), .ZN(n10008) );
  NAND2_X1 U9078 ( .A1(n7290), .A2(n7289), .ZN(n7291) );
  NAND2_X1 U9079 ( .A1(n10003), .A2(n7291), .ZN(n7294) );
  NAND4_X1 U9080 ( .A1(n7295), .A2(n7294), .A3(n7293), .A4(n7292), .ZN(n7296)
         );
  NAND2_X1 U9081 ( .A1(n7835), .A2(n7616), .ZN(n9981) );
  XNOR2_X1 U9082 ( .A(n7297), .B(n8250), .ZN(n7298) );
  AOI222_X1 U9083 ( .A1(n9962), .A2(n7298), .B1(n6380), .B2(n9673), .C1(n6400), 
        .C2(n9675), .ZN(n10007) );
  MUX2_X1 U9084 ( .A(n7299), .B(n10007), .S(n9989), .Z(n7305) );
  AOI21_X1 U9085 ( .B1(n10004), .B2(n7300), .A(n7494), .ZN(n10005) );
  NAND2_X1 U9086 ( .A1(n9989), .A2(n9550), .ZN(n9982) );
  NOR2_X1 U9087 ( .A1(n9982), .A2(n9724), .ZN(n9688) );
  NAND2_X2 U9088 ( .A1(n9989), .A2(n9975), .ZN(n9994) );
  OAI22_X1 U9089 ( .A1(n9994), .A2(n7302), .B1(n7301), .B2(n9987), .ZN(n7303)
         );
  AOI21_X1 U9090 ( .B1(n10005), .B2(n9688), .A(n7303), .ZN(n7304) );
  OAI211_X1 U9091 ( .C1(n10008), .C2(n9736), .A(n7305), .B(n7304), .ZN(
        P1_U3289) );
  AND3_X1 U9092 ( .A1(n7308), .A2(n7307), .A3(n7306), .ZN(n7309) );
  OAI21_X1 U9093 ( .B1(n7310), .B2(n7309), .A(n8557), .ZN(n7317) );
  INV_X1 U9094 ( .A(n7311), .ZN(n7315) );
  OAI22_X1 U9095 ( .A1(n8596), .A2(n7313), .B1(n7312), .B2(n8590), .ZN(n7314)
         );
  AOI211_X1 U9096 ( .C1(n8587), .C2(n8605), .A(n7315), .B(n7314), .ZN(n7316)
         );
  OAI211_X1 U9097 ( .C1(n7319), .C2(n7318), .A(n7317), .B(n7316), .ZN(P2_U3167) );
  INV_X1 U9098 ( .A(n9994), .ZN(n9966) );
  OAI21_X1 U9099 ( .B1(n9688), .B2(n9966), .A(n7320), .ZN(n7326) );
  INV_X1 U9100 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10248) );
  NAND3_X1 U9101 ( .A1(n8248), .A2(n8373), .A3(n7321), .ZN(n7323) );
  OAI211_X1 U9102 ( .C1(n10248), .C2(n9987), .A(n7323), .B(n7322), .ZN(n7324)
         );
  NAND2_X1 U9103 ( .A1(n7324), .A2(n9989), .ZN(n7325) );
  OAI211_X1 U9104 ( .C1(n10182), .C2(n9989), .A(n7326), .B(n7325), .ZN(
        P1_U3293) );
  INV_X1 U9105 ( .A(n7327), .ZN(n7329) );
  OAI222_X1 U9106 ( .A1(P1_U3086), .A2(n9550), .B1(n9864), .B2(n7329), .C1(
        n9866), .C2(n5377), .ZN(P1_U3336) );
  OAI222_X1 U9107 ( .A1(n8387), .A2(n7330), .B1(n7852), .B2(n7329), .C1(
        P2_U3151), .C2(n7328), .ZN(P2_U3276) );
  OAI22_X1 U9108 ( .A1(n8128), .A2(n4341), .B1(n8129), .B2(n6799), .ZN(n7331)
         );
  XNOR2_X1 U9109 ( .A(n7331), .B(n8061), .ZN(n7399) );
  OR2_X1 U9110 ( .A1(n8128), .A2(n8050), .ZN(n7333) );
  NAND2_X1 U9111 ( .A1(n10011), .A2(n4318), .ZN(n7332) );
  NAND2_X1 U9112 ( .A1(n7333), .A2(n7332), .ZN(n7340) );
  NAND2_X1 U9113 ( .A1(n7399), .A2(n7340), .ZN(n7334) );
  AND2_X1 U9114 ( .A1(n7395), .A2(n7334), .ZN(n7335) );
  NAND2_X1 U9115 ( .A1(n7336), .A2(n7335), .ZN(n7343) );
  OAI22_X1 U9116 ( .A1(n8126), .A2(n4341), .B1(n10021), .B2(n6799), .ZN(n7337)
         );
  XNOR2_X1 U9117 ( .A(n7337), .B(n8048), .ZN(n7344) );
  OR2_X1 U9118 ( .A1(n8126), .A2(n8050), .ZN(n7339) );
  NAND2_X1 U9119 ( .A1(n9967), .A2(n4318), .ZN(n7338) );
  AND2_X1 U9120 ( .A1(n7339), .A2(n7338), .ZN(n7345) );
  NAND2_X1 U9121 ( .A1(n7344), .A2(n7345), .ZN(n7672) );
  INV_X1 U9122 ( .A(n7399), .ZN(n7397) );
  INV_X1 U9123 ( .A(n7340), .ZN(n7670) );
  NAND2_X1 U9124 ( .A1(n7397), .A2(n7670), .ZN(n7341) );
  AND2_X1 U9125 ( .A1(n7672), .A2(n7341), .ZN(n7342) );
  INV_X1 U9126 ( .A(n7344), .ZN(n7347) );
  INV_X1 U9127 ( .A(n7345), .ZN(n7346) );
  NAND2_X1 U9128 ( .A1(n7347), .A2(n7346), .ZN(n7664) );
  NAND2_X1 U9129 ( .A1(n7667), .A2(n7664), .ZN(n7766) );
  NAND2_X1 U9130 ( .A1(n10029), .A2(n7976), .ZN(n7350) );
  OAI21_X1 U9131 ( .B1(n7753), .B2(n4341), .A(n7350), .ZN(n7351) );
  XNOR2_X1 U9132 ( .A(n7351), .B(n8061), .ZN(n7772) );
  OR2_X1 U9133 ( .A1(n7753), .A2(n8050), .ZN(n7353) );
  NAND2_X1 U9134 ( .A1(n10029), .A2(n4318), .ZN(n7352) );
  NAND2_X1 U9135 ( .A1(n7353), .A2(n7352), .ZN(n7771) );
  XNOR2_X1 U9136 ( .A(n7772), .B(n7771), .ZN(n7354) );
  XNOR2_X1 U9137 ( .A(n7348), .B(n7354), .ZN(n7362) );
  OR2_X1 U9138 ( .A1(n8126), .A2(n9710), .ZN(n7356) );
  NAND2_X1 U9139 ( .A1(n9399), .A2(n9675), .ZN(n7355) );
  AND2_X1 U9140 ( .A1(n7356), .A2(n7355), .ZN(n7479) );
  INV_X1 U9141 ( .A(n7479), .ZN(n7357) );
  AOI22_X1 U9142 ( .A1(n7357), .A2(n9269), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7360) );
  INV_X1 U9143 ( .A(n7481), .ZN(n7358) );
  OR2_X1 U9144 ( .A1(n9349), .A2(n7358), .ZN(n7359) );
  OAI211_X1 U9145 ( .C1(n7483), .C2(n9366), .A(n7360), .B(n7359), .ZN(n7361)
         );
  AOI21_X1 U9146 ( .B1(n7362), .B2(n9312), .A(n7361), .ZN(n7363) );
  INV_X1 U9147 ( .A(n7363), .ZN(P1_U3213) );
  NAND2_X1 U9148 ( .A1(n7150), .A2(n7364), .ZN(n7378) );
  NAND2_X1 U9149 ( .A1(n7378), .A2(n7365), .ZN(n7366) );
  XNOR2_X1 U9150 ( .A(n7366), .B(n7367), .ZN(n9071) );
  XOR2_X1 U9151 ( .A(n7368), .B(n7367), .Z(n7369) );
  OAI222_X1 U9152 ( .A1(n8969), .A2(n7700), .B1(n8971), .B2(n7370), .C1(n8967), 
        .C2(n7369), .ZN(n9067) );
  INV_X1 U9153 ( .A(n9067), .ZN(n7371) );
  MUX2_X1 U9154 ( .A(n7372), .B(n7371), .S(n9008), .Z(n7375) );
  INV_X1 U9155 ( .A(n7373), .ZN(n8561) );
  AOI22_X1 U9156 ( .A1(n8977), .A2(n9068), .B1(n9003), .B2(n8561), .ZN(n7374)
         );
  OAI211_X1 U9157 ( .C1(n9071), .C2(n8980), .A(n7375), .B(n7374), .ZN(P2_U3227) );
  INV_X1 U9158 ( .A(n7376), .ZN(n7377) );
  NAND2_X1 U9159 ( .A1(n7378), .A2(n7377), .ZN(n7382) );
  INV_X1 U9160 ( .A(n7379), .ZN(n7380) );
  NOR2_X1 U9161 ( .A1(n7385), .A2(n7380), .ZN(n7381) );
  NAND2_X1 U9162 ( .A1(n7382), .A2(n7381), .ZN(n7384) );
  NAND2_X1 U9163 ( .A1(n7384), .A2(n7383), .ZN(n7391) );
  AOI22_X1 U9164 ( .A1(n8952), .A2(n8605), .B1(n8954), .B2(n8603), .ZN(n7389)
         );
  XNOR2_X1 U9165 ( .A(n7386), .B(n7385), .ZN(n7387) );
  NAND2_X1 U9166 ( .A1(n7387), .A2(n8949), .ZN(n7388) );
  OAI211_X1 U9167 ( .C1(n7391), .C2(n7687), .A(n7389), .B(n7388), .ZN(n7409)
         );
  MUX2_X1 U9168 ( .A(n7409), .B(P2_REG2_REG_7__SCAN_IN), .S(n8993), .Z(n7390)
         );
  INV_X1 U9169 ( .A(n7390), .ZN(n7394) );
  INV_X1 U9170 ( .A(n7391), .ZN(n7411) );
  INV_X1 U9171 ( .A(n7631), .ZN(n7408) );
  OAI22_X1 U9172 ( .A1(n8991), .A2(n7408), .B1(n7629), .B2(n8989), .ZN(n7392)
         );
  AOI21_X1 U9173 ( .B1(n7411), .B2(n8997), .A(n7392), .ZN(n7393) );
  NAND2_X1 U9174 ( .A1(n7394), .A2(n7393), .ZN(P2_U3226) );
  AND2_X1 U9175 ( .A1(n7396), .A2(n7395), .ZN(n7398) );
  NAND2_X1 U9176 ( .A1(n7398), .A2(n7397), .ZN(n7665) );
  INV_X1 U9177 ( .A(n7398), .ZN(n7400) );
  NAND2_X1 U9178 ( .A1(n7400), .A2(n7399), .ZN(n7669) );
  NAND2_X1 U9179 ( .A1(n7665), .A2(n7669), .ZN(n7401) );
  XNOR2_X1 U9180 ( .A(n7401), .B(n7670), .ZN(n7406) );
  OAI22_X1 U9181 ( .A1(n9366), .A2(n8129), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7402), .ZN(n7404) );
  OAI22_X1 U9182 ( .A1(n7491), .A2(n9359), .B1(n9375), .B2(n8126), .ZN(n7403)
         );
  AOI211_X1 U9183 ( .C1(n7496), .C2(n9372), .A(n7404), .B(n7403), .ZN(n7405)
         );
  OAI21_X1 U9184 ( .B1(n7406), .B2(n9380), .A(n7405), .ZN(P1_U3227) );
  NOR2_X1 U9185 ( .A1(n7408), .A2(n7407), .ZN(n7410) );
  AOI211_X1 U9186 ( .C1(n7411), .C2(n7689), .A(n7410), .B(n7409), .ZN(n10130)
         );
  NAND2_X1 U9187 ( .A1(n9073), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7412) );
  OAI21_X1 U9188 ( .B1(n10130), .B2(n9073), .A(n7412), .ZN(P2_U3466) );
  INV_X1 U9189 ( .A(n7413), .ZN(n7437) );
  OAI222_X1 U9190 ( .A1(n7852), .A2(n7437), .B1(n8387), .B2(n5399), .C1(
        P2_U3151), .C2(n7414), .ZN(P2_U3275) );
  INV_X1 U9191 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9899) );
  NAND2_X1 U9192 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9334) );
  OAI21_X1 U9193 ( .B1(n9960), .B2(n9899), .A(n9334), .ZN(n7420) );
  XNOR2_X1 U9194 ( .A(n7517), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7418) );
  AOI211_X1 U9195 ( .C1(n4413), .C2(n7418), .A(n9944), .B(n7518), .ZN(n7419)
         );
  AOI211_X1 U9196 ( .C1(n9947), .C2(n7517), .A(n7420), .B(n7419), .ZN(n7427)
         );
  INV_X1 U9197 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7423) );
  XOR2_X1 U9198 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7517), .Z(n7424) );
  OAI211_X1 U9199 ( .C1(n7425), .C2(n7424), .A(n7512), .B(n9951), .ZN(n7426)
         );
  NAND2_X1 U9200 ( .A1(n7427), .A2(n7426), .ZN(P1_U3254) );
  INV_X1 U9201 ( .A(n7428), .ZN(n7436) );
  INV_X1 U9202 ( .A(n9736), .ZN(n9972) );
  OAI22_X1 U9203 ( .A1(n9989), .A2(n6999), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9987), .ZN(n7429) );
  AOI21_X1 U9204 ( .B1(n9966), .B2(n7430), .A(n7429), .ZN(n7431) );
  OAI21_X1 U9205 ( .B1(n9982), .B2(n7432), .A(n7431), .ZN(n7433) );
  AOI21_X1 U9206 ( .B1(n7434), .B2(n9972), .A(n7433), .ZN(n7435) );
  OAI21_X1 U9207 ( .B1(n7436), .B2(n10001), .A(n7435), .ZN(P1_U3290) );
  OAI222_X1 U9208 ( .A1(n9866), .A2(n7438), .B1(n9864), .B2(n7437), .C1(n8358), 
        .C2(P1_U3086), .ZN(P1_U3335) );
  XOR2_X1 U9209 ( .A(n7440), .B(n7439), .Z(n7454) );
  XNOR2_X1 U9210 ( .A(n7442), .B(n7441), .ZN(n7452) );
  NAND2_X1 U9211 ( .A1(n10118), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7443) );
  NAND2_X1 U9212 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8435) );
  OAI211_X1 U9213 ( .C1(n10111), .C2(n7444), .A(n7443), .B(n8435), .ZN(n7451)
         );
  NAND3_X1 U9214 ( .A1(n7446), .A2(n7448), .A3(n7447), .ZN(n7449) );
  AOI21_X1 U9215 ( .B1(n4568), .B2(n7449), .A(n8668), .ZN(n7450) );
  AOI211_X1 U9216 ( .C1(n6751), .C2(n7452), .A(n7451), .B(n7450), .ZN(n7453)
         );
  OAI21_X1 U9217 ( .B1(n7454), .B2(n10106), .A(n7453), .ZN(P2_U3192) );
  NAND2_X1 U9218 ( .A1(n7383), .A2(n7455), .ZN(n7456) );
  XOR2_X1 U9219 ( .A(n7457), .B(n7456), .Z(n7510) );
  XNOR2_X1 U9220 ( .A(n7458), .B(n7457), .ZN(n7459) );
  AOI222_X1 U9221 ( .A1(n8949), .A2(n7459), .B1(n8602), .B2(n8954), .C1(n8604), 
        .C2(n8952), .ZN(n7505) );
  INV_X1 U9222 ( .A(n7505), .ZN(n7460) );
  NAND2_X1 U9223 ( .A1(n7460), .A2(n5734), .ZN(n7462) );
  AOI22_X1 U9224 ( .A1(n9167), .A2(n7701), .B1(P2_REG0_REG_8__SCAN_IN), .B2(
        n10292), .ZN(n7461) );
  OAI211_X1 U9225 ( .C1(n7510), .C2(n9173), .A(n7462), .B(n7461), .ZN(P2_U3414) );
  XNOR2_X1 U9226 ( .A(n7463), .B(n7728), .ZN(n7473) );
  OAI21_X1 U9227 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n4422), .A(n7446), .ZN(
        n7471) );
  NAND2_X1 U9228 ( .A1(n10118), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7464) );
  NAND2_X1 U9229 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8492) );
  OAI211_X1 U9230 ( .C1(n10111), .C2(n7465), .A(n7464), .B(n8492), .ZN(n7470)
         );
  XOR2_X1 U9231 ( .A(n7467), .B(n7466), .Z(n7468) );
  INV_X1 U9232 ( .A(n6751), .ZN(n10099) );
  NOR2_X1 U9233 ( .A1(n7468), .A2(n10099), .ZN(n7469) );
  AOI211_X1 U9234 ( .C1(n10114), .C2(n7471), .A(n7470), .B(n7469), .ZN(n7472)
         );
  OAI21_X1 U9235 ( .B1(n7473), .B2(n10106), .A(n7472), .ZN(P2_U3191) );
  XOR2_X1 U9236 ( .A(n7474), .B(n8135), .Z(n10032) );
  NOR2_X1 U9237 ( .A1(n4618), .A2(n6402), .ZN(n7478) );
  INV_X1 U9238 ( .A(n7475), .ZN(n7476) );
  NAND2_X1 U9239 ( .A1(n7476), .A2(n8145), .ZN(n7477) );
  AOI21_X1 U9240 ( .B1(n7477), .B2(n8124), .A(n8135), .ZN(n7549) );
  AOI21_X1 U9241 ( .B1(n7478), .B2(n7477), .A(n7549), .ZN(n7480) );
  OAI21_X1 U9242 ( .B1(n7480), .B2(n9708), .A(n7479), .ZN(n10033) );
  NAND2_X1 U9243 ( .A1(n10033), .A2(n9989), .ZN(n7486) );
  AOI211_X1 U9244 ( .C1(n10029), .C2(n9970), .A(n9724), .B(n7552), .ZN(n10028)
         );
  AOI22_X1 U9245 ( .A1(n10001), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7481), .B2(
        n9965), .ZN(n7482) );
  OAI21_X1 U9246 ( .B1(n7483), .B2(n9994), .A(n7482), .ZN(n7484) );
  AOI21_X1 U9247 ( .B1(n10028), .B2(n9991), .A(n7484), .ZN(n7485) );
  OAI211_X1 U9248 ( .C1(n10032), .C2(n9736), .A(n7486), .B(n7485), .ZN(
        P1_U3286) );
  XOR2_X1 U9249 ( .A(n8253), .B(n7487), .Z(n10016) );
  INV_X1 U9250 ( .A(n8142), .ZN(n8293) );
  NOR2_X1 U9251 ( .A1(n7488), .A2(n8293), .ZN(n7489) );
  AOI211_X1 U9252 ( .C1(n8253), .C2(n7490), .A(n9708), .B(n7489), .ZN(n7493)
         );
  OAI22_X1 U9253 ( .A1(n7491), .A2(n9710), .B1(n8126), .B2(n9712), .ZN(n7492)
         );
  NOR2_X1 U9254 ( .A1(n7493), .A2(n7492), .ZN(n10015) );
  MUX2_X1 U9255 ( .A(n7000), .B(n10015), .S(n9989), .Z(n7500) );
  INV_X1 U9256 ( .A(n7494), .ZN(n7495) );
  AOI21_X1 U9257 ( .B1(n10011), .B2(n7495), .A(n4425), .ZN(n10013) );
  INV_X1 U9258 ( .A(n7496), .ZN(n7497) );
  OAI22_X1 U9259 ( .A1(n9994), .A2(n8129), .B1(n9987), .B2(n7497), .ZN(n7498)
         );
  AOI21_X1 U9260 ( .B1(n10013), .B2(n9688), .A(n7498), .ZN(n7499) );
  OAI211_X1 U9261 ( .C1(n10016), .C2(n9736), .A(n7500), .B(n7499), .ZN(
        P1_U3288) );
  INV_X1 U9262 ( .A(n7501), .ZN(n9072) );
  MUX2_X1 U9263 ( .A(n7502), .B(n7505), .S(n4313), .Z(n7504) );
  NAND2_X1 U9264 ( .A1(n9054), .A2(n7701), .ZN(n7503) );
  OAI211_X1 U9265 ( .C1(n7510), .C2(n9061), .A(n7504), .B(n7503), .ZN(P2_U3467) );
  MUX2_X1 U9266 ( .A(n7506), .B(n7505), .S(n9008), .Z(n7509) );
  INV_X1 U9267 ( .A(n7507), .ZN(n7705) );
  AOI22_X1 U9268 ( .A1(n8977), .A2(n7701), .B1(n9003), .B2(n7705), .ZN(n7508)
         );
  OAI211_X1 U9269 ( .C1(n7510), .C2(n8980), .A(n7509), .B(n7508), .ZN(P2_U3225) );
  INV_X1 U9270 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7511) );
  MUX2_X1 U9271 ( .A(n7511), .B(P1_REG2_REG_12__SCAN_IN), .S(n9489), .Z(n7516)
         );
  INV_X1 U9272 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7513) );
  OAI21_X1 U9273 ( .B1(n7514), .B2(n7513), .A(n7512), .ZN(n7515) );
  AOI21_X1 U9274 ( .B1(n7516), .B2(n7515), .A(n9481), .ZN(n7526) );
  XOR2_X1 U9275 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9489), .Z(n7520) );
  OAI21_X1 U9276 ( .B1(n7520), .B2(n7519), .A(n9488), .ZN(n7521) );
  NAND2_X1 U9277 ( .A1(n7521), .A2(n9545), .ZN(n7525) );
  INV_X1 U9278 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7522) );
  NAND2_X1 U9279 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9229) );
  OAI21_X1 U9280 ( .B1(n9960), .B2(n7522), .A(n9229), .ZN(n7523) );
  AOI21_X1 U9281 ( .B1(n9489), .B2(n9947), .A(n7523), .ZN(n7524) );
  OAI211_X1 U9282 ( .C1(n7526), .C2(n9934), .A(n7525), .B(n7524), .ZN(P1_U3255) );
  INV_X1 U9283 ( .A(n7527), .ZN(n7602) );
  OAI222_X1 U9284 ( .A1(n7852), .A2(n7602), .B1(P2_U3151), .B2(n7529), .C1(
        n7528), .C2(n8387), .ZN(P2_U3274) );
  INV_X1 U9285 ( .A(n7530), .ZN(n7531) );
  OAI21_X1 U9286 ( .B1(n7531), .B2(n8169), .A(n8261), .ZN(n7532) );
  NAND2_X1 U9287 ( .A1(n7532), .A2(n7831), .ZN(n7533) );
  AOI222_X1 U9288 ( .A1(n9962), .A2(n7533), .B1(n9393), .B2(n9675), .C1(n9395), 
        .C2(n9673), .ZN(n9823) );
  OAI21_X1 U9289 ( .B1(n4454), .B2(n8261), .A(n7534), .ZN(n9819) );
  INV_X1 U9290 ( .A(n9820), .ZN(n9320) );
  AOI21_X1 U9291 ( .B1(n9820), .B2(n7570), .A(n7536), .ZN(n9821) );
  NAND2_X1 U9292 ( .A1(n9821), .A2(n9688), .ZN(n7538) );
  AOI22_X1 U9293 ( .A1(n10001), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9314), .B2(
        n9965), .ZN(n7537) );
  OAI211_X1 U9294 ( .C1(n9320), .C2(n9994), .A(n7538), .B(n7537), .ZN(n7539)
         );
  AOI21_X1 U9295 ( .B1(n9819), .B2(n9972), .A(n7539), .ZN(n7540) );
  OAI21_X1 U9296 ( .B1(n9823), .B2(n10001), .A(n7540), .ZN(P1_U3280) );
  INV_X1 U9297 ( .A(n7542), .ZN(n7543) );
  OR2_X1 U9298 ( .A1(n7544), .A2(n7543), .ZN(n7547) );
  XNOR2_X1 U9299 ( .A(n7541), .B(n7547), .ZN(n10042) );
  INV_X1 U9300 ( .A(n7547), .ZN(n7545) );
  NAND2_X1 U9301 ( .A1(n7545), .A2(n7546), .ZN(n7548) );
  OAI21_X1 U9302 ( .B1(n7549), .B2(n4929), .A(n7547), .ZN(n7649) );
  OAI21_X1 U9303 ( .B1(n7549), .B2(n7548), .A(n7649), .ZN(n7550) );
  INV_X1 U9304 ( .A(n7753), .ZN(n9400) );
  AOI222_X1 U9305 ( .A1(n9962), .A2(n7550), .B1(n9398), .B2(n9675), .C1(n9400), 
        .C2(n9673), .ZN(n10041) );
  MUX2_X1 U9306 ( .A(n7551), .B(n10041), .S(n9989), .Z(n7557) );
  INV_X1 U9307 ( .A(n7552), .ZN(n7553) );
  AOI211_X1 U9308 ( .C1(n10039), .C2(n7553), .A(n9724), .B(n7653), .ZN(n10038)
         );
  INV_X1 U9309 ( .A(n7554), .ZN(n7752) );
  OAI22_X1 U9310 ( .A1(n7758), .A2(n9994), .B1(n9987), .B2(n7752), .ZN(n7555)
         );
  AOI21_X1 U9311 ( .B1(n10038), .B2(n9991), .A(n7555), .ZN(n7556) );
  OAI211_X1 U9312 ( .C1(n9736), .C2(n10042), .A(n7557), .B(n7556), .ZN(
        P1_U3285) );
  NOR2_X1 U9313 ( .A1(n7567), .A2(n7558), .ZN(n7565) );
  NAND2_X1 U9314 ( .A1(n7596), .A2(n7560), .ZN(n7609) );
  NAND2_X1 U9315 ( .A1(n7609), .A2(n8245), .ZN(n7611) );
  INV_X1 U9316 ( .A(n7561), .ZN(n7563) );
  AOI21_X1 U9317 ( .B1(n7596), .B2(n7563), .A(n7562), .ZN(n7564) );
  AOI21_X1 U9318 ( .B1(n7565), .B2(n7611), .A(n7564), .ZN(n9829) );
  XNOR2_X1 U9319 ( .A(n7567), .B(n7566), .ZN(n7568) );
  AOI222_X1 U9320 ( .A1(n9962), .A2(n7568), .B1(n9394), .B2(n9675), .C1(n9396), 
        .C2(n9673), .ZN(n9828) );
  MUX2_X1 U9321 ( .A(n7511), .B(n9828), .S(n9989), .Z(n7575) );
  INV_X1 U9322 ( .A(n7570), .ZN(n7571) );
  AOI211_X1 U9323 ( .C1(n9826), .C2(n7619), .A(n9724), .B(n7571), .ZN(n9825)
         );
  INV_X1 U9324 ( .A(n9228), .ZN(n7572) );
  OAI22_X1 U9325 ( .A1(n6057), .A2(n9994), .B1(n7572), .B2(n9987), .ZN(n7573)
         );
  AOI21_X1 U9326 ( .B1(n9825), .B2(n9991), .A(n7573), .ZN(n7574) );
  OAI211_X1 U9327 ( .C1(n9829), .C2(n9736), .A(n7575), .B(n7574), .ZN(P1_U3281) );
  NAND2_X1 U9328 ( .A1(n7576), .A2(n7581), .ZN(n7577) );
  NAND2_X1 U9329 ( .A1(n7578), .A2(n7577), .ZN(n7585) );
  INV_X1 U9330 ( .A(n7585), .ZN(n8998) );
  NAND2_X1 U9331 ( .A1(n7580), .A2(n7579), .ZN(n7712) );
  XNOR2_X1 U9332 ( .A(n7712), .B(n5189), .ZN(n7582) );
  NAND2_X1 U9333 ( .A1(n7582), .A2(n8949), .ZN(n7584) );
  AOI22_X1 U9334 ( .A1(n8601), .A2(n8954), .B1(n8952), .B2(n8603), .ZN(n7583)
         );
  OAI211_X1 U9335 ( .C1(n7585), .C2(n7687), .A(n7584), .B(n7583), .ZN(n8994)
         );
  AOI21_X1 U9336 ( .B1(n7689), .B2(n8998), .A(n8994), .ZN(n7727) );
  AOI22_X1 U9337 ( .A1(n9167), .A2(n8502), .B1(n10292), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n7586) );
  OAI21_X1 U9338 ( .B1(n7727), .B2(n10292), .A(n7586), .ZN(P2_U3417) );
  INV_X1 U9339 ( .A(n7587), .ZN(n8291) );
  INV_X1 U9340 ( .A(n8294), .ZN(n7589) );
  OAI21_X1 U9341 ( .B1(n8291), .B2(n7589), .A(n7588), .ZN(n7590) );
  NAND2_X1 U9342 ( .A1(n7590), .A2(n7607), .ZN(n7591) );
  AOI222_X1 U9343 ( .A1(n9962), .A2(n7591), .B1(n9396), .B2(n9675), .C1(n9398), 
        .C2(n9673), .ZN(n9833) );
  INV_X1 U9344 ( .A(n7618), .ZN(n7593) );
  AOI21_X1 U9345 ( .B1(n7653), .B2(n7656), .A(n7795), .ZN(n7592) );
  NOR3_X1 U9346 ( .A1(n7593), .A2(n7592), .A3(n9724), .ZN(n9830) );
  AOI22_X1 U9347 ( .A1(n10001), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7788), .B2(
        n9965), .ZN(n7594) );
  OAI21_X1 U9348 ( .B1(n7795), .B2(n9994), .A(n7594), .ZN(n7600) );
  INV_X1 U9349 ( .A(n7595), .ZN(n7598) );
  INV_X1 U9350 ( .A(n7596), .ZN(n7597) );
  AOI21_X1 U9351 ( .B1(n7598), .B2(n8256), .A(n7597), .ZN(n9834) );
  NOR2_X1 U9352 ( .A1(n9834), .A2(n9736), .ZN(n7599) );
  AOI211_X1 U9353 ( .C1(n9830), .C2(n9991), .A(n7600), .B(n7599), .ZN(n7601)
         );
  OAI21_X1 U9354 ( .B1(n10001), .B2(n9833), .A(n7601), .ZN(P1_U3283) );
  OAI222_X1 U9355 ( .A1(n9866), .A2(n7603), .B1(n9864), .B2(n7602), .C1(n8286), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U9356 ( .A(n7644), .ZN(n7606) );
  AOI21_X1 U9357 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9183), .A(n7604), .ZN(
        n7605) );
  OAI21_X1 U9358 ( .B1(n7606), .B2(n7852), .A(n7605), .ZN(P2_U3272) );
  NAND2_X1 U9359 ( .A1(n7607), .A2(n8166), .ZN(n7608) );
  XNOR2_X1 U9360 ( .A(n7608), .B(n8245), .ZN(n7615) );
  OR2_X1 U9361 ( .A1(n7609), .A2(n8245), .ZN(n7610) );
  NAND2_X1 U9362 ( .A1(n7611), .A2(n7610), .ZN(n7731) );
  NAND2_X1 U9363 ( .A1(n7731), .A2(n10036), .ZN(n7614) );
  OAI22_X1 U9364 ( .A1(n9289), .A2(n9710), .B1(n9336), .B2(n9712), .ZN(n7612)
         );
  INV_X1 U9365 ( .A(n7612), .ZN(n7613) );
  OAI211_X1 U9366 ( .C1(n9708), .C2(n7615), .A(n7614), .B(n7613), .ZN(n7736)
         );
  INV_X1 U9367 ( .A(n7736), .ZN(n7625) );
  INV_X1 U9368 ( .A(n7616), .ZN(n7617) );
  NAND2_X1 U9369 ( .A1(n9989), .A2(n7617), .ZN(n7843) );
  INV_X1 U9370 ( .A(n7843), .ZN(n9998) );
  AOI21_X1 U9371 ( .B1(n7618), .B2(n6597), .A(n9724), .ZN(n7620) );
  NAND2_X1 U9372 ( .A1(n7620), .A2(n7619), .ZN(n7732) );
  AOI22_X1 U9373 ( .A1(n10001), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9333), .B2(
        n9965), .ZN(n7622) );
  NAND2_X1 U9374 ( .A1(n6597), .A2(n9966), .ZN(n7621) );
  OAI211_X1 U9375 ( .C1(n7732), .C2(n9982), .A(n7622), .B(n7621), .ZN(n7623)
         );
  AOI21_X1 U9376 ( .B1(n7731), .B2(n9998), .A(n7623), .ZN(n7624) );
  OAI21_X1 U9377 ( .B1(n7625), .B2(n10001), .A(n7624), .ZN(P1_U3282) );
  INV_X1 U9378 ( .A(n7695), .ZN(n7626) );
  AOI21_X1 U9379 ( .B1(n7628), .B2(n7627), .A(n7626), .ZN(n7637) );
  AND2_X1 U9380 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10108) );
  AOI21_X1 U9381 ( .B1(n8587), .B2(n8603), .A(n10108), .ZN(n7635) );
  INV_X1 U9382 ( .A(n7629), .ZN(n7630) );
  NAND2_X1 U9383 ( .A1(n8593), .A2(n7630), .ZN(n7634) );
  NAND2_X1 U9384 ( .A1(n8572), .A2(n8605), .ZN(n7633) );
  NAND2_X1 U9385 ( .A1(n8578), .A2(n7631), .ZN(n7632) );
  AND4_X1 U9386 ( .A1(n7635), .A2(n7634), .A3(n7633), .A4(n7632), .ZN(n7636)
         );
  OAI21_X1 U9387 ( .B1(n7637), .B2(n8581), .A(n7636), .ZN(P2_U3153) );
  INV_X1 U9388 ( .A(n7638), .ZN(n7642) );
  OAI222_X1 U9389 ( .A1(n9866), .A2(n7640), .B1(n9864), .B2(n7642), .C1(
        P1_U3086), .C2(n7639), .ZN(P1_U3333) );
  OAI222_X1 U9390 ( .A1(n8387), .A2(n7643), .B1(n7852), .B2(n7642), .C1(n7641), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  NAND2_X1 U9391 ( .A1(n7644), .A2(n9859), .ZN(n7645) );
  OAI211_X1 U9392 ( .C1(n7646), .C2(n9866), .A(n7645), .B(n8378), .ZN(P1_U3332) );
  NAND2_X1 U9393 ( .A1(n8743), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7647) );
  OAI21_X1 U9394 ( .B1(n8753), .B2(n8743), .A(n7647), .ZN(P2_U3522) );
  XOR2_X1 U9395 ( .A(n7648), .B(n7650), .Z(n10050) );
  NAND2_X1 U9396 ( .A1(n7649), .A2(n8151), .ZN(n7651) );
  XNOR2_X1 U9397 ( .A(n7651), .B(n7650), .ZN(n7652) );
  AOI22_X1 U9398 ( .A1(n7652), .A2(n9962), .B1(n9673), .B2(n9399), .ZN(n10049)
         );
  MUX2_X1 U9399 ( .A(n6996), .B(n10049), .S(n9989), .Z(n7659) );
  XNOR2_X1 U9400 ( .A(n7653), .B(n7656), .ZN(n7654) );
  OAI22_X1 U9401 ( .A1(n7654), .A2(n9724), .B1(n9289), .B2(n9712), .ZN(n10045)
         );
  INV_X1 U9402 ( .A(n9286), .ZN(n7655) );
  OAI22_X1 U9403 ( .A1(n7656), .A2(n9994), .B1(n9987), .B2(n7655), .ZN(n7657)
         );
  AOI21_X1 U9404 ( .B1(n10045), .B2(n9991), .A(n7657), .ZN(n7658) );
  OAI211_X1 U9405 ( .C1(n9736), .C2(n10050), .A(n7659), .B(n7658), .ZN(
        P1_U3284) );
  OR2_X1 U9406 ( .A1(n8128), .A2(n9710), .ZN(n7661) );
  OR2_X1 U9407 ( .A1(n7753), .A2(n9712), .ZN(n7660) );
  NAND2_X1 U9408 ( .A1(n7661), .A2(n7660), .ZN(n9961) );
  NOR2_X1 U9409 ( .A1(n7662), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9445) );
  AOI21_X1 U9410 ( .B1(n9269), .B2(n9961), .A(n9445), .ZN(n7663) );
  OAI21_X1 U9411 ( .B1(n9366), .B2(n10021), .A(n7663), .ZN(n7675) );
  INV_X1 U9412 ( .A(n7348), .ZN(n7747) );
  INV_X1 U9413 ( .A(n7664), .ZN(n7666) );
  OAI21_X1 U9414 ( .B1(n7667), .B2(n7666), .A(n7665), .ZN(n7668) );
  AOI21_X1 U9415 ( .B1(n7670), .B2(n7669), .A(n7668), .ZN(n7671) );
  AOI21_X1 U9416 ( .B1(n7747), .B2(n7672), .A(n7671), .ZN(n7673) );
  NOR2_X1 U9417 ( .A1(n7673), .A2(n9380), .ZN(n7674) );
  AOI211_X1 U9418 ( .C1(n9964), .C2(n9372), .A(n7675), .B(n7674), .ZN(n7676)
         );
  INV_X1 U9419 ( .A(n7676), .ZN(P1_U3239) );
  INV_X1 U9420 ( .A(n7678), .ZN(n7682) );
  XNOR2_X1 U9421 ( .A(n7677), .B(n7682), .ZN(n7688) );
  INV_X1 U9422 ( .A(n7688), .ZN(n8987) );
  NAND2_X1 U9423 ( .A1(n7712), .A2(n7679), .ZN(n7681) );
  NAND2_X1 U9424 ( .A1(n7681), .A2(n7680), .ZN(n7683) );
  XNOR2_X1 U9425 ( .A(n7683), .B(n7682), .ZN(n7684) );
  NAND2_X1 U9426 ( .A1(n7684), .A2(n8949), .ZN(n7686) );
  AOI22_X1 U9427 ( .A1(n8600), .A2(n8954), .B1(n8952), .B2(n8602), .ZN(n7685)
         );
  OAI211_X1 U9428 ( .C1(n7688), .C2(n7687), .A(n7686), .B(n7685), .ZN(n8984)
         );
  AOI21_X1 U9429 ( .B1(n7689), .B2(n8987), .A(n8984), .ZN(n9062) );
  AOI22_X1 U9430 ( .A1(n9167), .A2(n7690), .B1(n10292), .B2(
        P2_REG0_REG_10__SCAN_IN), .ZN(n7691) );
  OAI21_X1 U9431 ( .B1(n9062), .B2(n10292), .A(n7691), .ZN(P2_U3420) );
  AND3_X1 U9432 ( .A1(n7695), .A2(n7694), .A3(n7693), .ZN(n7696) );
  OAI21_X1 U9433 ( .B1(n7697), .B2(n7696), .A(n8557), .ZN(n7707) );
  NAND2_X1 U9434 ( .A1(n8587), .A2(n8602), .ZN(n7699) );
  OAI211_X1 U9435 ( .C1(n7700), .C2(n8590), .A(n7699), .B(n7698), .ZN(n7704)
         );
  INV_X1 U9436 ( .A(n7701), .ZN(n7702) );
  NOR2_X1 U9437 ( .A1(n8596), .A2(n7702), .ZN(n7703) );
  AOI211_X1 U9438 ( .C1(n7705), .C2(n8593), .A(n7704), .B(n7703), .ZN(n7706)
         );
  NAND2_X1 U9439 ( .A1(n7707), .A2(n7706), .ZN(P2_U3161) );
  NAND2_X1 U9440 ( .A1(n7708), .A2(n7709), .ZN(n7710) );
  XNOR2_X1 U9441 ( .A(n7710), .B(n8462), .ZN(n7726) );
  NAND2_X1 U9442 ( .A1(n7712), .A2(n7711), .ZN(n7714) );
  NAND2_X1 U9443 ( .A1(n7714), .A2(n7713), .ZN(n7715) );
  XNOR2_X1 U9444 ( .A(n7715), .B(n5612), .ZN(n7716) );
  AOI222_X1 U9445 ( .A1(n8949), .A2(n7716), .B1(n8951), .B2(n8954), .C1(n8601), 
        .C2(n8952), .ZN(n7722) );
  MUX2_X1 U9446 ( .A(n7717), .B(n7722), .S(n5734), .Z(n7719) );
  NAND2_X1 U9447 ( .A1(n9167), .A2(n8538), .ZN(n7718) );
  OAI211_X1 U9448 ( .C1(n7726), .C2(n9173), .A(n7719), .B(n7718), .ZN(P2_U3423) );
  INV_X1 U9449 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8645) );
  MUX2_X1 U9450 ( .A(n8645), .B(n7722), .S(n4313), .Z(n7721) );
  NAND2_X1 U9451 ( .A1(n9054), .A2(n8538), .ZN(n7720) );
  OAI211_X1 U9452 ( .C1(n9061), .C2(n7726), .A(n7721), .B(n7720), .ZN(P2_U3470) );
  MUX2_X1 U9453 ( .A(n10261), .B(n7722), .S(n9008), .Z(n7725) );
  INV_X1 U9454 ( .A(n7723), .ZN(n8542) );
  AOI22_X1 U9455 ( .A1(n8977), .A2(n8538), .B1(n9003), .B2(n8542), .ZN(n7724)
         );
  OAI211_X1 U9456 ( .C1(n7726), .C2(n8980), .A(n7725), .B(n7724), .ZN(P2_U3222) );
  INV_X1 U9457 ( .A(n8502), .ZN(n8992) );
  MUX2_X1 U9458 ( .A(n7728), .B(n7727), .S(n4313), .Z(n7729) );
  OAI21_X1 U9459 ( .B1(n8992), .B2(n9065), .A(n7729), .ZN(P2_U3468) );
  INV_X1 U9460 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10275) );
  INV_X1 U9461 ( .A(n6597), .ZN(n7734) );
  INV_X1 U9462 ( .A(n10031), .ZN(n7730) );
  NAND2_X1 U9463 ( .A1(n7731), .A2(n7730), .ZN(n7733) );
  OAI211_X1 U9464 ( .C1(n7734), .C2(n10020), .A(n7733), .B(n7732), .ZN(n7735)
         );
  NOR2_X1 U9465 ( .A1(n7736), .A2(n7735), .ZN(n7738) );
  MUX2_X1 U9466 ( .A(n10275), .B(n7738), .S(n10064), .Z(n7737) );
  INV_X1 U9467 ( .A(n7737), .ZN(P1_U3533) );
  INV_X1 U9468 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7739) );
  MUX2_X1 U9469 ( .A(n7739), .B(n7738), .S(n10055), .Z(n7740) );
  INV_X1 U9470 ( .A(n7740), .ZN(P1_U3486) );
  AND2_X1 U9471 ( .A1(n9399), .A2(n8063), .ZN(n7741) );
  AOI21_X1 U9472 ( .B1(n10039), .B2(n8058), .A(n7741), .ZN(n7775) );
  NAND2_X1 U9473 ( .A1(n10039), .A2(n7976), .ZN(n7743) );
  NAND2_X1 U9474 ( .A1(n9399), .A2(n8058), .ZN(n7742) );
  NAND2_X1 U9475 ( .A1(n7743), .A2(n7742), .ZN(n7744) );
  XNOR2_X1 U9476 ( .A(n7744), .B(n8048), .ZN(n7776) );
  INV_X1 U9477 ( .A(n7776), .ZN(n7749) );
  INV_X1 U9478 ( .A(n7771), .ZN(n7746) );
  OAI21_X1 U9479 ( .B1(n7348), .B2(n7771), .A(n7772), .ZN(n7745) );
  OAI21_X1 U9480 ( .B1(n7747), .B2(n7746), .A(n7745), .ZN(n7748) );
  NOR2_X1 U9481 ( .A1(n7748), .A2(n7749), .ZN(n9290) );
  AOI21_X1 U9482 ( .B1(n7749), .B2(n7748), .A(n9290), .ZN(n7750) );
  NAND2_X1 U9483 ( .A1(n7750), .A2(n7775), .ZN(n9293) );
  OAI21_X1 U9484 ( .B1(n7775), .B2(n7750), .A(n9293), .ZN(n7751) );
  NAND2_X1 U9485 ( .A1(n7751), .A2(n9312), .ZN(n7757) );
  NAND2_X1 U9486 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9472) );
  INV_X1 U9487 ( .A(n9472), .ZN(n7755) );
  OAI22_X1 U9488 ( .A1(n9359), .A2(n7753), .B1(n9349), .B2(n7752), .ZN(n7754)
         );
  AOI211_X1 U9489 ( .C1(n9317), .C2(n9398), .A(n7755), .B(n7754), .ZN(n7756)
         );
  OAI211_X1 U9490 ( .C1(n7758), .C2(n9366), .A(n7757), .B(n7756), .ZN(P1_U3221) );
  INV_X1 U9491 ( .A(n7759), .ZN(n7827) );
  OAI222_X1 U9492 ( .A1(P1_U3086), .A2(n7761), .B1(n9864), .B2(n7827), .C1(
        n7760), .C2(n9866), .ZN(P1_U3331) );
  NOR2_X1 U9493 ( .A1(n9289), .A2(n8050), .ZN(n7762) );
  AOI21_X1 U9494 ( .B1(n9831), .B2(n4318), .A(n7762), .ZN(n7915) );
  NAND2_X1 U9495 ( .A1(n7776), .A2(n7775), .ZN(n7773) );
  NOR2_X1 U9496 ( .A1(n7772), .A2(n7771), .ZN(n7763) );
  NAND2_X1 U9497 ( .A1(n7766), .A2(n7765), .ZN(n7779) );
  NAND2_X1 U9498 ( .A1(n10046), .A2(n7976), .ZN(n7768) );
  OR2_X1 U9499 ( .A1(n7790), .A2(n4341), .ZN(n7767) );
  NAND2_X1 U9500 ( .A1(n7768), .A2(n7767), .ZN(n7769) );
  XNOR2_X1 U9501 ( .A(n7769), .B(n8048), .ZN(n7781) );
  NOR2_X1 U9502 ( .A1(n7790), .A2(n8050), .ZN(n7770) );
  AOI21_X1 U9503 ( .B1(n10046), .B2(n8058), .A(n7770), .ZN(n7780) );
  XNOR2_X1 U9504 ( .A(n7781), .B(n7780), .ZN(n9292) );
  NAND3_X1 U9505 ( .A1(n7773), .A2(n7772), .A3(n7771), .ZN(n7774) );
  OAI21_X1 U9506 ( .B1(n7776), .B2(n7775), .A(n7774), .ZN(n7777) );
  NOR2_X1 U9507 ( .A1(n9292), .A2(n7777), .ZN(n7778) );
  NAND2_X1 U9508 ( .A1(n7779), .A2(n7778), .ZN(n9294) );
  NAND2_X1 U9509 ( .A1(n7781), .A2(n7780), .ZN(n7782) );
  NAND2_X1 U9510 ( .A1(n9831), .A2(n7976), .ZN(n7784) );
  OR2_X1 U9511 ( .A1(n9289), .A2(n4341), .ZN(n7783) );
  NAND2_X1 U9512 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  XNOR2_X1 U9513 ( .A(n7785), .B(n8048), .ZN(n7906) );
  INV_X1 U9514 ( .A(n7906), .ZN(n7917) );
  NOR2_X1 U9515 ( .A1(n4344), .A2(n7917), .ZN(n9337) );
  AOI21_X1 U9516 ( .B1(n4344), .B2(n7917), .A(n9337), .ZN(n7786) );
  NAND2_X1 U9517 ( .A1(n7786), .A2(n7915), .ZN(n9340) );
  OAI21_X1 U9518 ( .B1(n7915), .B2(n7786), .A(n9340), .ZN(n7787) );
  NAND2_X1 U9519 ( .A1(n7787), .A2(n9312), .ZN(n7794) );
  INV_X1 U9520 ( .A(n7788), .ZN(n7789) );
  OAI22_X1 U9521 ( .A1(n9359), .A2(n7790), .B1(n9349), .B2(n7789), .ZN(n7791)
         );
  AOI211_X1 U9522 ( .C1(n9317), .C2(n9396), .A(n7792), .B(n7791), .ZN(n7793)
         );
  OAI211_X1 U9523 ( .C1(n7795), .C2(n9366), .A(n7794), .B(n7793), .ZN(P1_U3217) );
  XOR2_X1 U9524 ( .A(n7797), .B(n7796), .Z(n7812) );
  NAND2_X1 U9525 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8469) );
  OAI21_X1 U9526 ( .B1(n10111), .B2(n7798), .A(n8469), .ZN(n7803) );
  AOI211_X1 U9527 ( .C1(n7801), .C2(n7800), .A(n10099), .B(n7799), .ZN(n7802)
         );
  AOI211_X1 U9528 ( .C1(n10118), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7803), .B(
        n7802), .ZN(n7811) );
  INV_X1 U9529 ( .A(n7804), .ZN(n7809) );
  NOR3_X1 U9530 ( .A1(n7807), .A2(n7805), .A3(n7806), .ZN(n7808) );
  OAI21_X1 U9531 ( .B1(n7809), .B2(n7808), .A(n10114), .ZN(n7810) );
  OAI211_X1 U9532 ( .C1(n7812), .C2(n10106), .A(n7811), .B(n7810), .ZN(
        P2_U3194) );
  XNOR2_X1 U9533 ( .A(n7813), .B(n8244), .ZN(n9813) );
  INV_X1 U9534 ( .A(n4447), .ZN(n7815) );
  AOI21_X1 U9535 ( .B1(n7816), .B2(n8244), .A(n7815), .ZN(n7817) );
  OAI222_X1 U9536 ( .A1(n9712), .A2(n9376), .B1(n9710), .B2(n7818), .C1(n9708), 
        .C2(n7817), .ZN(n9809) );
  INV_X1 U9537 ( .A(n9811), .ZN(n7823) );
  INV_X1 U9538 ( .A(n7865), .ZN(n7820) );
  AOI211_X1 U9539 ( .C1(n9811), .C2(n7819), .A(n9724), .B(n7820), .ZN(n9810)
         );
  NAND2_X1 U9540 ( .A1(n9810), .A2(n9991), .ZN(n7822) );
  AOI22_X1 U9541 ( .A1(n10001), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9373), .B2(
        n9965), .ZN(n7821) );
  OAI211_X1 U9542 ( .C1(n7823), .C2(n9994), .A(n7822), .B(n7821), .ZN(n7824)
         );
  AOI21_X1 U9543 ( .B1(n9809), .B2(n9989), .A(n7824), .ZN(n7825) );
  OAI21_X1 U9544 ( .B1(n9736), .B2(n9813), .A(n7825), .ZN(P1_U3278) );
  OAI222_X1 U9545 ( .A1(n7852), .A2(n7827), .B1(P2_U3151), .B2(n5703), .C1(
        n7826), .C2(n8387), .ZN(P2_U3271) );
  INV_X1 U9546 ( .A(n7828), .ZN(n7851) );
  OAI222_X1 U9547 ( .A1(P1_U3086), .A2(n7830), .B1(n9864), .B2(n7851), .C1(
        n7829), .C2(n9866), .ZN(P1_U3330) );
  NAND2_X1 U9548 ( .A1(n7831), .A2(n8185), .ZN(n7833) );
  XNOR2_X1 U9549 ( .A(n7833), .B(n8264), .ZN(n7838) );
  OAI22_X1 U9550 ( .A1(n9258), .A2(n9712), .B1(n9231), .B2(n9710), .ZN(n7837)
         );
  XNOR2_X1 U9551 ( .A(n7834), .B(n8264), .ZN(n9818) );
  NOR2_X1 U9552 ( .A1(n9818), .A2(n7835), .ZN(n7836) );
  AOI211_X1 U9553 ( .C1(n7838), .C2(n9962), .A(n7837), .B(n7836), .ZN(n9817)
         );
  INV_X1 U9554 ( .A(n7536), .ZN(n7840) );
  INV_X1 U9555 ( .A(n7819), .ZN(n7839) );
  AOI211_X1 U9556 ( .C1(n9815), .C2(n7840), .A(n9724), .B(n7839), .ZN(n9814)
         );
  AOI22_X1 U9557 ( .A1(n10001), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9193), .B2(
        n9965), .ZN(n7841) );
  OAI21_X1 U9558 ( .B1(n7842), .B2(n9994), .A(n7841), .ZN(n7845) );
  NOR2_X1 U9559 ( .A1(n9818), .A2(n7843), .ZN(n7844) );
  AOI211_X1 U9560 ( .C1(n9814), .C2(n9991), .A(n7845), .B(n7844), .ZN(n7846)
         );
  OAI21_X1 U9561 ( .B1(n9817), .B2(n10001), .A(n7846), .ZN(P1_U3279) );
  INV_X1 U9562 ( .A(n7847), .ZN(n7854) );
  OAI222_X1 U9563 ( .A1(n7852), .A2(n7854), .B1(P2_U3151), .B2(n7849), .C1(
        n7848), .C2(n8387), .ZN(P2_U3269) );
  OAI222_X1 U9564 ( .A1(n7852), .A2(n7851), .B1(P2_U3151), .B2(n8112), .C1(
        n7850), .C2(n8387), .ZN(P2_U3270) );
  OAI222_X1 U9565 ( .A1(P1_U3086), .A2(n7855), .B1(n9864), .B2(n7854), .C1(
        n7853), .C2(n9866), .ZN(P1_U3329) );
  INV_X1 U9566 ( .A(n7856), .ZN(n9863) );
  AOI21_X1 U9567 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9183), .A(n7857), .ZN(
        n7858) );
  OAI21_X1 U9568 ( .B1(n9863), .B2(n7852), .A(n7858), .ZN(P2_U3268) );
  NAND2_X1 U9569 ( .A1(n4447), .A2(n8181), .ZN(n7859) );
  XNOR2_X1 U9570 ( .A(n7859), .B(n8265), .ZN(n7860) );
  AOI222_X1 U9571 ( .A1(n9962), .A2(n7860), .B1(n9392), .B2(n9673), .C1(n9390), 
        .C2(n9675), .ZN(n9808) );
  NAND2_X1 U9572 ( .A1(n4453), .A2(n8265), .ZN(n9802) );
  NAND3_X1 U9573 ( .A1(n7861), .A2(n9802), .A3(n9972), .ZN(n7869) );
  INV_X1 U9574 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9507) );
  INV_X1 U9575 ( .A(n7863), .ZN(n9257) );
  OAI22_X1 U9576 ( .A1(n9989), .A2(n9507), .B1(n9257), .B2(n9987), .ZN(n7864)
         );
  AOI21_X1 U9577 ( .B1(n9803), .B2(n9966), .A(n7864), .ZN(n7868) );
  AND2_X1 U9578 ( .A1(n7865), .A2(n9803), .ZN(n7866) );
  NOR2_X1 U9579 ( .A1(n9723), .A2(n7866), .ZN(n9804) );
  NAND2_X1 U9580 ( .A1(n9804), .A2(n9688), .ZN(n7867) );
  AND3_X1 U9581 ( .A1(n7869), .A2(n7868), .A3(n7867), .ZN(n7870) );
  OAI21_X1 U9582 ( .B1(n9808), .B2(n10001), .A(n7870), .ZN(P1_U3277) );
  OAI222_X1 U9583 ( .A1(n9866), .A2(n7872), .B1(n9864), .B2(n7873), .C1(
        P1_U3086), .C2(n7871), .ZN(P1_U3352) );
  OAI222_X1 U9584 ( .A1(n8387), .A2(n7874), .B1(n7852), .B2(n7873), .C1(
        P2_U3151), .C2(n4790), .ZN(P2_U3292) );
  XNOR2_X1 U9585 ( .A(n7875), .B(n7882), .ZN(n9751) );
  INV_X1 U9586 ( .A(n9577), .ZN(n7877) );
  AOI211_X1 U9587 ( .C1(n9748), .C2(n7876), .A(n9724), .B(n7877), .ZN(n9747)
         );
  INV_X1 U9588 ( .A(n9748), .ZN(n8109) );
  INV_X1 U9589 ( .A(n8106), .ZN(n7878) );
  AOI22_X1 U9590 ( .A1(n7878), .A2(n9965), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n10001), .ZN(n7879) );
  OAI21_X1 U9591 ( .B1(n8109), .B2(n9994), .A(n7879), .ZN(n7887) );
  OAI21_X1 U9592 ( .B1(n7882), .B2(n7881), .A(n7880), .ZN(n7883) );
  INV_X1 U9593 ( .A(n9593), .ZN(n7890) );
  INV_X1 U9594 ( .A(n7876), .ZN(n7889) );
  AOI211_X1 U9595 ( .C1(n9753), .C2(n7890), .A(n9724), .B(n7889), .ZN(n9752)
         );
  AOI22_X1 U9596 ( .A1(n9363), .A2(n9965), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n10001), .ZN(n7891) );
  OAI21_X1 U9597 ( .B1(n9367), .B2(n9994), .A(n7891), .ZN(n7896) );
  OAI21_X1 U9598 ( .B1(n8272), .B2(n7893), .A(n7892), .ZN(n7894) );
  AOI222_X1 U9599 ( .A1(n9962), .A2(n7894), .B1(n9586), .B2(n9675), .C1(n9385), 
        .C2(n9673), .ZN(n9755) );
  NOR2_X1 U9600 ( .A1(n9755), .A2(n10001), .ZN(n7895) );
  OAI21_X1 U9601 ( .B1(n9756), .B2(n9736), .A(n7897), .ZN(P1_U3267) );
  XOR2_X1 U9602 ( .A(n7898), .B(n7899), .Z(n7905) );
  AOI22_X1 U9603 ( .A1(n9378), .A2(n7901), .B1(n9269), .B2(n7900), .ZN(n7904)
         );
  NAND2_X1 U9604 ( .A1(n7902), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7903) );
  OAI211_X1 U9605 ( .C1(n7905), .C2(n9380), .A(n7904), .B(n7903), .ZN(P1_U3237) );
  NAND2_X1 U9606 ( .A1(n6597), .A2(n7976), .ZN(n7908) );
  OR2_X1 U9607 ( .A1(n7910), .A2(n4341), .ZN(n7907) );
  NAND2_X1 U9608 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  XNOR2_X1 U9609 ( .A(n7909), .B(n8048), .ZN(n7913) );
  NOR2_X1 U9610 ( .A1(n7910), .A2(n8050), .ZN(n7911) );
  AOI21_X1 U9611 ( .B1(n6597), .B2(n8058), .A(n7911), .ZN(n7912) );
  NAND2_X1 U9612 ( .A1(n7913), .A2(n7912), .ZN(n9233) );
  OR2_X1 U9613 ( .A1(n7913), .A2(n7912), .ZN(n7914) );
  NAND2_X1 U9614 ( .A1(n9233), .A2(n7914), .ZN(n9339) );
  INV_X1 U9615 ( .A(n7915), .ZN(n7916) );
  AND2_X1 U9616 ( .A1(n7917), .A2(n7916), .ZN(n7918) );
  NOR2_X1 U9617 ( .A1(n9339), .A2(n7918), .ZN(n7919) );
  NAND2_X1 U9618 ( .A1(n9826), .A2(n7976), .ZN(n7921) );
  OR2_X1 U9619 ( .A1(n9336), .A2(n4341), .ZN(n7920) );
  NAND2_X1 U9620 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  XNOR2_X1 U9621 ( .A(n7922), .B(n8048), .ZN(n7925) );
  NOR2_X1 U9622 ( .A1(n9336), .A2(n8050), .ZN(n7923) );
  AOI21_X1 U9623 ( .B1(n9826), .B2(n4318), .A(n7923), .ZN(n7924) );
  NAND2_X1 U9624 ( .A1(n7925), .A2(n7924), .ZN(n7927) );
  OR2_X1 U9625 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  NAND2_X1 U9626 ( .A1(n9235), .A2(n7927), .ZN(n9310) );
  NAND2_X1 U9627 ( .A1(n9820), .A2(n7976), .ZN(n7929) );
  OR2_X1 U9628 ( .A1(n9231), .A2(n4341), .ZN(n7928) );
  NAND2_X1 U9629 ( .A1(n7929), .A2(n7928), .ZN(n7930) );
  XNOR2_X1 U9630 ( .A(n7930), .B(n8061), .ZN(n7932) );
  NOR2_X1 U9631 ( .A1(n9231), .A2(n8050), .ZN(n7931) );
  AOI21_X1 U9632 ( .B1(n9820), .B2(n8058), .A(n7931), .ZN(n7933) );
  XNOR2_X1 U9633 ( .A(n7932), .B(n7933), .ZN(n9311) );
  NAND2_X1 U9634 ( .A1(n9310), .A2(n9311), .ZN(n9309) );
  INV_X1 U9635 ( .A(n7932), .ZN(n7934) );
  NAND2_X1 U9636 ( .A1(n7934), .A2(n7933), .ZN(n7935) );
  NAND2_X1 U9637 ( .A1(n9309), .A2(n7935), .ZN(n7942) );
  INV_X1 U9638 ( .A(n7942), .ZN(n7940) );
  NAND2_X1 U9639 ( .A1(n9815), .A2(n7976), .ZN(n7937) );
  NAND2_X1 U9640 ( .A1(n9393), .A2(n4318), .ZN(n7936) );
  NAND2_X1 U9641 ( .A1(n7937), .A2(n7936), .ZN(n7938) );
  XNOR2_X1 U9642 ( .A(n7938), .B(n8048), .ZN(n7941) );
  INV_X1 U9643 ( .A(n7941), .ZN(n7939) );
  NAND2_X1 U9644 ( .A1(n7942), .A2(n7941), .ZN(n7947) );
  NAND2_X1 U9645 ( .A1(n9815), .A2(n4318), .ZN(n7945) );
  NAND2_X1 U9646 ( .A1(n9393), .A2(n8063), .ZN(n7944) );
  NAND2_X1 U9647 ( .A1(n7945), .A2(n7944), .ZN(n9192) );
  INV_X1 U9648 ( .A(n9192), .ZN(n7946) );
  INV_X1 U9649 ( .A(n9248), .ZN(n7953) );
  NAND2_X1 U9650 ( .A1(n9811), .A2(n7976), .ZN(n7949) );
  NAND2_X1 U9651 ( .A1(n9392), .A2(n8058), .ZN(n7948) );
  NAND2_X1 U9652 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  XNOR2_X1 U9653 ( .A(n7950), .B(n8048), .ZN(n9250) );
  NAND2_X1 U9654 ( .A1(n9811), .A2(n4318), .ZN(n7952) );
  NAND2_X1 U9655 ( .A1(n9392), .A2(n8063), .ZN(n7951) );
  NAND2_X1 U9656 ( .A1(n7953), .A2(n4374), .ZN(n7962) );
  NAND2_X1 U9657 ( .A1(n9803), .A2(n7976), .ZN(n7955) );
  OR2_X1 U9658 ( .A1(n9376), .A2(n4341), .ZN(n7954) );
  NAND2_X1 U9659 ( .A1(n7955), .A2(n7954), .ZN(n7956) );
  XNOR2_X1 U9660 ( .A(n7956), .B(n8061), .ZN(n7963) );
  NOR2_X1 U9661 ( .A1(n9376), .A2(n8050), .ZN(n7957) );
  AOI21_X1 U9662 ( .B1(n9803), .B2(n4318), .A(n7957), .ZN(n7964) );
  XNOR2_X1 U9663 ( .A(n7963), .B(n7964), .ZN(n9253) );
  INV_X1 U9664 ( .A(n9250), .ZN(n7959) );
  NAND2_X1 U9665 ( .A1(n7959), .A2(n9370), .ZN(n7960) );
  AND2_X1 U9666 ( .A1(n9253), .A2(n7960), .ZN(n7961) );
  INV_X1 U9667 ( .A(n7963), .ZN(n7965) );
  NAND2_X1 U9668 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  NAND2_X1 U9669 ( .A1(n9798), .A2(n7976), .ZN(n7968) );
  NAND2_X1 U9670 ( .A1(n9390), .A2(n4318), .ZN(n7967) );
  NAND2_X1 U9671 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  XNOR2_X1 U9672 ( .A(n7969), .B(n8061), .ZN(n7972) );
  NAND2_X1 U9673 ( .A1(n9798), .A2(n4318), .ZN(n7971) );
  NAND2_X1 U9674 ( .A1(n9390), .A2(n8063), .ZN(n7970) );
  NAND2_X1 U9675 ( .A1(n7971), .A2(n7970), .ZN(n7973) );
  NAND2_X1 U9676 ( .A1(n7972), .A2(n7973), .ZN(n9264) );
  INV_X1 U9677 ( .A(n7972), .ZN(n7975) );
  INV_X1 U9678 ( .A(n7973), .ZN(n7974) );
  NAND2_X1 U9679 ( .A1(n7975), .A2(n7974), .ZN(n9263) );
  NAND2_X1 U9680 ( .A1(n9789), .A2(n7976), .ZN(n7978) );
  NAND2_X1 U9681 ( .A1(n9674), .A2(n4318), .ZN(n7977) );
  NAND2_X1 U9682 ( .A1(n7978), .A2(n7977), .ZN(n7979) );
  XNOR2_X1 U9683 ( .A(n7979), .B(n8061), .ZN(n9212) );
  NAND2_X1 U9684 ( .A1(n9789), .A2(n4318), .ZN(n7981) );
  NAND2_X1 U9685 ( .A1(n9674), .A2(n8063), .ZN(n7980) );
  NAND2_X1 U9686 ( .A1(n7981), .A2(n7980), .ZN(n9211) );
  NAND2_X1 U9687 ( .A1(n9794), .A2(n7976), .ZN(n7983) );
  NAND2_X1 U9688 ( .A1(n9389), .A2(n4318), .ZN(n7982) );
  NAND2_X1 U9689 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  XNOR2_X1 U9690 ( .A(n7984), .B(n8061), .ZN(n7989) );
  NAND2_X1 U9691 ( .A1(n9794), .A2(n8058), .ZN(n7986) );
  NAND2_X1 U9692 ( .A1(n9389), .A2(n8063), .ZN(n7985) );
  NAND2_X1 U9693 ( .A1(n7986), .A2(n7985), .ZN(n9346) );
  OAI22_X1 U9694 ( .A1(n9212), .A2(n9211), .B1(n7989), .B2(n9346), .ZN(n7993)
         );
  INV_X1 U9695 ( .A(n7989), .ZN(n9210) );
  INV_X1 U9696 ( .A(n9346), .ZN(n7988) );
  INV_X1 U9697 ( .A(n9211), .ZN(n7987) );
  OAI21_X1 U9698 ( .B1(n9210), .B2(n7988), .A(n7987), .ZN(n7991) );
  AND2_X1 U9699 ( .A1(n9211), .A2(n9346), .ZN(n7990) );
  AOI22_X1 U9700 ( .A1(n9212), .A2(n7991), .B1(n7990), .B2(n7989), .ZN(n7992)
         );
  OAI21_X2 U9701 ( .B1(n9209), .B2(n7993), .A(n7992), .ZN(n9304) );
  NAND2_X1 U9702 ( .A1(n9782), .A2(n7976), .ZN(n7995) );
  NAND2_X1 U9703 ( .A1(n9221), .A2(n4318), .ZN(n7994) );
  NAND2_X1 U9704 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  XNOR2_X1 U9705 ( .A(n7996), .B(n8061), .ZN(n9302) );
  INV_X1 U9706 ( .A(n9302), .ZN(n7999) );
  NAND2_X1 U9707 ( .A1(n9782), .A2(n4318), .ZN(n7998) );
  NAND2_X1 U9708 ( .A1(n9221), .A2(n8063), .ZN(n7997) );
  NAND2_X1 U9709 ( .A1(n7998), .A2(n7997), .ZN(n8000) );
  INV_X1 U9710 ( .A(n8000), .ZN(n9301) );
  NAND2_X1 U9711 ( .A1(n7999), .A2(n9301), .ZN(n8001) );
  NAND2_X1 U9712 ( .A1(n9778), .A2(n7976), .ZN(n8003) );
  NAND2_X1 U9713 ( .A1(n9676), .A2(n8058), .ZN(n8002) );
  NAND2_X1 U9714 ( .A1(n8003), .A2(n8002), .ZN(n8004) );
  XNOR2_X1 U9715 ( .A(n8004), .B(n8061), .ZN(n8006) );
  AND2_X1 U9716 ( .A1(n9676), .A2(n8063), .ZN(n8005) );
  AOI21_X1 U9717 ( .B1(n9778), .B2(n4318), .A(n8005), .ZN(n8007) );
  XNOR2_X1 U9718 ( .A(n8006), .B(n8007), .ZN(n9220) );
  INV_X1 U9719 ( .A(n8006), .ZN(n8008) );
  AND2_X1 U9720 ( .A1(n8008), .A2(n8007), .ZN(n8009) );
  NAND2_X1 U9721 ( .A1(n9773), .A2(n8058), .ZN(n8011) );
  NAND2_X1 U9722 ( .A1(n9388), .A2(n8063), .ZN(n8010) );
  NAND2_X1 U9723 ( .A1(n9773), .A2(n7976), .ZN(n8013) );
  NAND2_X1 U9724 ( .A1(n9388), .A2(n4318), .ZN(n8012) );
  NAND2_X1 U9725 ( .A1(n8013), .A2(n8012), .ZN(n8014) );
  XNOR2_X1 U9726 ( .A(n8014), .B(n8048), .ZN(n9198) );
  NAND2_X1 U9727 ( .A1(n9769), .A2(n7976), .ZN(n8016) );
  NAND2_X1 U9728 ( .A1(n9387), .A2(n8058), .ZN(n8015) );
  NAND2_X1 U9729 ( .A1(n8016), .A2(n8015), .ZN(n8017) );
  XNOR2_X1 U9730 ( .A(n8017), .B(n8061), .ZN(n8020) );
  NAND2_X1 U9731 ( .A1(n9769), .A2(n4318), .ZN(n8019) );
  NAND2_X1 U9732 ( .A1(n9387), .A2(n8063), .ZN(n8018) );
  NAND2_X1 U9733 ( .A1(n8019), .A2(n8018), .ZN(n8021) );
  NAND2_X1 U9734 ( .A1(n8020), .A2(n8021), .ZN(n9201) );
  OAI21_X1 U9735 ( .B1(n9322), .B2(n9198), .A(n9201), .ZN(n8025) );
  NAND3_X1 U9736 ( .A1(n9201), .A2(n9322), .A3(n9198), .ZN(n8024) );
  INV_X1 U9737 ( .A(n8020), .ZN(n8023) );
  INV_X1 U9738 ( .A(n8021), .ZN(n8022) );
  NAND2_X1 U9739 ( .A1(n8023), .A2(n8022), .ZN(n9275) );
  NAND2_X1 U9740 ( .A1(n9764), .A2(n7976), .ZN(n8027) );
  NAND2_X1 U9741 ( .A1(n9386), .A2(n8058), .ZN(n8026) );
  NAND2_X1 U9742 ( .A1(n8027), .A2(n8026), .ZN(n8028) );
  XNOR2_X1 U9743 ( .A(n8028), .B(n8061), .ZN(n8032) );
  NAND2_X1 U9744 ( .A1(n9764), .A2(n4318), .ZN(n8030) );
  NAND2_X1 U9745 ( .A1(n9386), .A2(n8063), .ZN(n8029) );
  NAND2_X1 U9746 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  NOR2_X1 U9747 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  AOI21_X1 U9748 ( .B1(n8032), .B2(n8031), .A(n8033), .ZN(n9276) );
  INV_X1 U9749 ( .A(n8033), .ZN(n8034) );
  NAND2_X1 U9750 ( .A1(n9279), .A2(n8034), .ZN(n9239) );
  NAND2_X1 U9751 ( .A1(n9759), .A2(n7976), .ZN(n8036) );
  NAND2_X1 U9752 ( .A1(n9385), .A2(n4318), .ZN(n8035) );
  NAND2_X1 U9753 ( .A1(n8036), .A2(n8035), .ZN(n8037) );
  XNOR2_X1 U9754 ( .A(n8037), .B(n8061), .ZN(n8042) );
  AOI22_X1 U9755 ( .A1(n9759), .A2(n4318), .B1(n8063), .B2(n9385), .ZN(n8043)
         );
  XNOR2_X1 U9756 ( .A(n8042), .B(n8043), .ZN(n9240) );
  NAND2_X1 U9757 ( .A1(n9753), .A2(n7976), .ZN(n8039) );
  NAND2_X1 U9758 ( .A1(n9384), .A2(n4318), .ZN(n8038) );
  NAND2_X1 U9759 ( .A1(n8039), .A2(n8038), .ZN(n8040) );
  XNOR2_X1 U9760 ( .A(n8040), .B(n8061), .ZN(n8056) );
  AND2_X1 U9761 ( .A1(n8063), .A2(n9384), .ZN(n8041) );
  AOI21_X1 U9762 ( .B1(n9753), .B2(n4318), .A(n8041), .ZN(n8054) );
  XNOR2_X1 U9763 ( .A(n8056), .B(n8054), .ZN(n9355) );
  INV_X1 U9764 ( .A(n8042), .ZN(n8044) );
  NAND2_X1 U9765 ( .A1(n8044), .A2(n8043), .ZN(n9356) );
  NAND2_X1 U9766 ( .A1(n9748), .A2(n7976), .ZN(n8047) );
  NAND2_X1 U9767 ( .A1(n9586), .A2(n8058), .ZN(n8046) );
  NAND2_X1 U9768 ( .A1(n8047), .A2(n8046), .ZN(n8049) );
  XNOR2_X1 U9769 ( .A(n8049), .B(n8048), .ZN(n8053) );
  NOR2_X1 U9770 ( .A1(n9360), .A2(n8050), .ZN(n8051) );
  AOI21_X1 U9771 ( .B1(n9748), .B2(n4318), .A(n8051), .ZN(n8052) );
  NAND2_X1 U9772 ( .A1(n8053), .A2(n8052), .ZN(n8070) );
  OAI21_X1 U9773 ( .B1(n8053), .B2(n8052), .A(n8070), .ZN(n8100) );
  INV_X1 U9774 ( .A(n8054), .ZN(n8055) );
  NAND2_X1 U9775 ( .A1(n9742), .A2(n7976), .ZN(n8060) );
  NAND2_X1 U9776 ( .A1(n9383), .A2(n8058), .ZN(n8059) );
  NAND2_X1 U9777 ( .A1(n8060), .A2(n8059), .ZN(n8062) );
  XNOR2_X1 U9778 ( .A(n8062), .B(n8061), .ZN(n8065) );
  AOI22_X1 U9779 ( .A1(n9742), .A2(n8058), .B1(n8063), .B2(n9383), .ZN(n8064)
         );
  XNOR2_X1 U9780 ( .A(n8065), .B(n8064), .ZN(n8066) );
  INV_X1 U9781 ( .A(n8066), .ZN(n8071) );
  NAND3_X1 U9782 ( .A1(n8071), .A2(n9312), .A3(n8070), .ZN(n8076) );
  NAND3_X1 U9783 ( .A1(n8104), .A2(n9312), .A3(n8066), .ZN(n8075) );
  AOI22_X1 U9784 ( .A1(n9585), .A2(n9317), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8069) );
  NAND2_X1 U9785 ( .A1(n9578), .A2(n9372), .ZN(n8068) );
  OAI211_X1 U9786 ( .C1(n9360), .C2(n9359), .A(n8069), .B(n8068), .ZN(n8073)
         );
  NOR3_X1 U9787 ( .A1(n8071), .A2(n8070), .A3(n9380), .ZN(n8072) );
  AOI211_X1 U9788 ( .C1(n9742), .C2(n9378), .A(n8073), .B(n8072), .ZN(n8074)
         );
  OAI211_X1 U9789 ( .C1(n8104), .C2(n8076), .A(n8075), .B(n8074), .ZN(P1_U3220) );
  INV_X1 U9790 ( .A(n9084), .ZN(n8096) );
  OR2_X1 U9791 ( .A1(n8078), .A2(n4986), .ZN(n8082) );
  OR2_X1 U9792 ( .A1(n4986), .A2(n8079), .ZN(n8080) );
  XNOR2_X1 U9793 ( .A(n9090), .B(n8399), .ZN(n8084) );
  XNOR2_X1 U9794 ( .A(n8084), .B(n8803), .ZN(n8566) );
  NAND2_X1 U9795 ( .A1(n8084), .A2(n8092), .ZN(n8085) );
  NAND2_X1 U9796 ( .A1(n8569), .A2(n8085), .ZN(n8086) );
  XNOR2_X1 U9797 ( .A(n9084), .B(n8461), .ZN(n8405) );
  XNOR2_X1 U9798 ( .A(n8405), .B(n8786), .ZN(n8087) );
  AOI21_X1 U9799 ( .B1(n8086), .B2(n8087), .A(n8581), .ZN(n8090) );
  INV_X1 U9800 ( .A(n8086), .ZN(n8089) );
  INV_X1 U9801 ( .A(n8087), .ZN(n8088) );
  NAND2_X1 U9802 ( .A1(n8090), .A2(n8413), .ZN(n8095) );
  AOI22_X1 U9803 ( .A1(n8778), .A2(n8593), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8091) );
  OAI21_X1 U9804 ( .B1(n8092), .B2(n8590), .A(n8091), .ZN(n8093) );
  AOI21_X1 U9805 ( .B1(n8587), .B2(n8774), .A(n8093), .ZN(n8094) );
  OAI211_X1 U9806 ( .C1(n8096), .C2(n8596), .A(n8095), .B(n8094), .ZN(P2_U3154) );
  OAI222_X1 U9807 ( .A1(n8098), .A2(P1_U3086), .B1(n9864), .B2(n8398), .C1(
        n8097), .C2(n9866), .ZN(P1_U3326) );
  INV_X1 U9808 ( .A(n8099), .ZN(n8102) );
  INV_X1 U9809 ( .A(n8100), .ZN(n8101) );
  AOI21_X1 U9810 ( .B1(n9354), .B2(n8102), .A(n8101), .ZN(n8103) );
  AOI22_X1 U9811 ( .A1(n9384), .A2(n9371), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8105) );
  OAI21_X1 U9812 ( .B1(n9349), .B2(n8106), .A(n8105), .ZN(n8107) );
  AOI21_X1 U9813 ( .B1(n9317), .B2(n9383), .A(n8107), .ZN(n8108) );
  INV_X1 U9814 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8113) );
  NOR3_X1 U9815 ( .A1(n8111), .A2(n8110), .A3(P2_U3151), .ZN(n8381) );
  AOI22_X1 U9816 ( .A1(n8383), .A2(n8113), .B1(n8381), .B2(n8112), .ZN(
        P2_U3377) );
  INV_X1 U9817 ( .A(n8345), .ZN(n8326) );
  INV_X1 U9818 ( .A(n8325), .ZN(n8117) );
  INV_X1 U9819 ( .A(n8225), .ZN(n8116) );
  AOI21_X1 U9820 ( .B1(n8326), .B2(n8117), .A(n8116), .ZN(n8118) );
  OAI21_X1 U9821 ( .B1(n8118), .B2(n8238), .A(n8329), .ZN(n8119) );
  OAI21_X1 U9822 ( .B1(n8238), .B2(n8329), .A(n8119), .ZN(n8121) );
  NAND4_X1 U9823 ( .A1(n8226), .A2(n8238), .A3(n8345), .A4(n8225), .ZN(n8120)
         );
  OAI211_X1 U9824 ( .C1(n8238), .C2(n8226), .A(n8121), .B(n8120), .ZN(n8231)
         );
  INV_X1 U9825 ( .A(n8195), .ZN(n8198) );
  NOR2_X1 U9826 ( .A1(n6400), .A2(n4312), .ZN(n8127) );
  INV_X1 U9827 ( .A(n8127), .ZN(n8125) );
  OAI22_X1 U9828 ( .A1(n8129), .A2(n8125), .B1(n9401), .B2(n4312), .ZN(n8136)
         );
  AOI21_X1 U9829 ( .B1(n8127), .B2(n8126), .A(n8129), .ZN(n8133) );
  AOI21_X1 U9830 ( .B1(n8130), .B2(n9401), .A(n10011), .ZN(n8132) );
  AOI22_X1 U9831 ( .A1(n8130), .A2(n8129), .B1(n4312), .B2(n9401), .ZN(n8131)
         );
  OAI22_X1 U9832 ( .A1(n8133), .A2(n8132), .B1(n8131), .B2(n9967), .ZN(n8134)
         );
  AND2_X1 U9833 ( .A1(n8137), .A2(n8238), .ZN(n8144) );
  INV_X1 U9834 ( .A(n8138), .ZN(n8140) );
  OAI211_X1 U9835 ( .C1(n8141), .C2(n8140), .A(n6381), .B(n8139), .ZN(n8143)
         );
  NAND4_X1 U9836 ( .A1(n8145), .A2(n8144), .A3(n8143), .A4(n8142), .ZN(n8146)
         );
  AND2_X1 U9837 ( .A1(n8148), .A2(n8147), .ZN(n8150) );
  MUX2_X1 U9838 ( .A(n8150), .B(n8149), .S(n4312), .Z(n8155) );
  NAND2_X1 U9839 ( .A1(n8156), .A2(n8151), .ZN(n8153) );
  NAND2_X1 U9840 ( .A1(n8158), .A2(n8157), .ZN(n8162) );
  INV_X1 U9841 ( .A(n8159), .ZN(n8160) );
  NOR2_X1 U9842 ( .A1(n8162), .A2(n8160), .ZN(n8295) );
  OAI21_X1 U9843 ( .B1(n8168), .B2(n4513), .A(n8295), .ZN(n8164) );
  AND2_X1 U9844 ( .A1(n8170), .A2(n8166), .ZN(n8161) );
  OR2_X1 U9845 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  AND2_X1 U9846 ( .A1(n8163), .A2(n8171), .ZN(n8298) );
  NAND2_X1 U9847 ( .A1(n8164), .A2(n8298), .ZN(n8175) );
  INV_X1 U9848 ( .A(n8165), .ZN(n8167) );
  AOI21_X1 U9849 ( .B1(n8171), .B2(n8170), .A(n8169), .ZN(n8172) );
  AOI21_X1 U9850 ( .B1(n8173), .B2(n8295), .A(n8172), .ZN(n8174) );
  NAND2_X1 U9851 ( .A1(n8188), .A2(n8183), .ZN(n8179) );
  INV_X1 U9852 ( .A(n8184), .ZN(n8177) );
  NAND2_X1 U9853 ( .A1(n8189), .A2(n8176), .ZN(n8305) );
  INV_X1 U9854 ( .A(n8189), .ZN(n8180) );
  AOI21_X1 U9855 ( .B1(n8304), .B2(n9392), .A(n4312), .ZN(n8190) );
  INV_X1 U9856 ( .A(n8190), .ZN(n8182) );
  NAND2_X1 U9857 ( .A1(n8191), .A2(n8182), .ZN(n8192) );
  NAND2_X1 U9858 ( .A1(n8184), .A2(n8183), .ZN(n8297) );
  OR2_X1 U9859 ( .A1(n8297), .A2(n8185), .ZN(n8187) );
  AND2_X1 U9860 ( .A1(n8187), .A2(n8186), .ZN(n8300) );
  NAND2_X1 U9861 ( .A1(n8201), .A2(n8194), .ZN(n8307) );
  NAND2_X1 U9862 ( .A1(n8195), .A2(n8200), .ZN(n8311) );
  AND2_X1 U9863 ( .A1(n8200), .A2(n8199), .ZN(n8308) );
  NAND3_X1 U9864 ( .A1(n8310), .A2(n8238), .A3(n8201), .ZN(n8202) );
  AOI21_X1 U9865 ( .B1(n8203), .B2(n8308), .A(n8202), .ZN(n8204) );
  INV_X1 U9866 ( .A(n8205), .ZN(n9656) );
  INV_X1 U9867 ( .A(n8208), .ZN(n9631) );
  INV_X1 U9868 ( .A(n8313), .ZN(n8209) );
  NAND2_X1 U9869 ( .A1(n8209), .A2(n4312), .ZN(n8210) );
  OAI21_X1 U9870 ( .B1(n8280), .B2(n4312), .A(n8210), .ZN(n8211) );
  INV_X1 U9871 ( .A(n8242), .ZN(n8213) );
  AOI21_X1 U9872 ( .B1(n8214), .B2(n8285), .A(n8213), .ZN(n8215) );
  AOI21_X1 U9873 ( .B1(n9636), .B2(n9773), .A(n8281), .ZN(n8315) );
  OAI21_X1 U9874 ( .B1(n8215), .B2(n9646), .A(n8315), .ZN(n8217) );
  NAND4_X1 U9875 ( .A1(n8217), .A2(n4312), .A3(n8280), .A4(n8216), .ZN(n8223)
         );
  INV_X1 U9876 ( .A(n8219), .ZN(n8317) );
  AOI21_X1 U9877 ( .B1(n8282), .B2(n8324), .A(n8317), .ZN(n8221) );
  INV_X1 U9878 ( .A(n8324), .ZN(n8218) );
  AOI21_X1 U9879 ( .B1(n8219), .B2(n8316), .A(n8218), .ZN(n8220) );
  MUX2_X1 U9880 ( .A(n8221), .B(n8220), .S(n8238), .Z(n8222) );
  NAND2_X1 U9881 ( .A1(n8226), .A2(n8225), .ZN(n8349) );
  NAND2_X1 U9882 ( .A1(n8329), .A2(n8325), .ZN(n8227) );
  INV_X1 U9883 ( .A(n9382), .ZN(n8240) );
  NOR3_X1 U9884 ( .A1(n8234), .A2(n8240), .A3(n9740), .ZN(n8229) );
  NOR2_X1 U9885 ( .A1(n9740), .A2(n8238), .ZN(n8228) );
  INV_X1 U9886 ( .A(n8232), .ZN(n8233) );
  INV_X1 U9887 ( .A(n8234), .ZN(n8237) );
  INV_X1 U9888 ( .A(n8348), .ZN(n8235) );
  NAND2_X1 U9889 ( .A1(n8333), .A2(n8237), .ZN(n8351) );
  AOI21_X1 U9890 ( .B1(n8351), .B2(n8239), .A(n8238), .ZN(n8334) );
  NOR2_X1 U9891 ( .A1(n8334), .A2(n8286), .ZN(n8279) );
  INV_X1 U9892 ( .A(n8239), .ZN(n8355) );
  NAND2_X1 U9893 ( .A1(n8241), .A2(n8240), .ZN(n8330) );
  INV_X1 U9894 ( .A(n9609), .ZN(n8271) );
  NAND2_X1 U9895 ( .A1(n8243), .A2(n8242), .ZN(n9668) );
  XNOR2_X1 U9896 ( .A(n9782), .B(n9221), .ZN(n9684) );
  NOR2_X1 U9897 ( .A1(n8246), .A2(n7051), .ZN(n8252) );
  NOR2_X1 U9898 ( .A1(n8248), .A2(n8247), .ZN(n8251) );
  NAND4_X1 U9899 ( .A1(n8252), .A2(n8251), .A3(n8250), .A4(n8249), .ZN(n8254)
         );
  NOR3_X1 U9900 ( .A1(n8254), .A2(n6402), .A3(n8253), .ZN(n8255) );
  AND4_X1 U9901 ( .A1(n8257), .A2(n6599), .A3(n8256), .A4(n8255), .ZN(n8259)
         );
  NAND3_X1 U9902 ( .A1(n8260), .A2(n8259), .A3(n8258), .ZN(n8262) );
  NOR2_X1 U9903 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  NAND4_X1 U9904 ( .A1(n8265), .A2(n8264), .A3(n6443), .A4(n8263), .ZN(n8266)
         );
  NOR2_X1 U9905 ( .A1(n8307), .A2(n8266), .ZN(n8267) );
  NAND4_X1 U9906 ( .A1(n9684), .A2(n8308), .A3(n4367), .A4(n8267), .ZN(n8268)
         );
  NOR2_X1 U9907 ( .A1(n8269), .A2(n9646), .ZN(n8270) );
  NAND4_X1 U9908 ( .A1(n8275), .A2(n9583), .A3(n8330), .A4(n8274), .ZN(n8276)
         );
  NOR2_X1 U9909 ( .A1(n8358), .A2(n9550), .ZN(n8362) );
  OAI21_X1 U9910 ( .B1(n4312), .B2(n8286), .A(n8362), .ZN(n8278) );
  AOI211_X1 U9911 ( .C1(n8341), .C2(n8279), .A(n8361), .B(n8278), .ZN(n8371)
         );
  OAI21_X1 U9912 ( .B1(n4392), .B2(n8281), .A(n8280), .ZN(n8284) );
  INV_X1 U9913 ( .A(n8282), .ZN(n8283) );
  AOI21_X1 U9914 ( .B1(n8313), .B2(n8284), .A(n8283), .ZN(n8320) );
  NAND2_X1 U9915 ( .A1(n8320), .A2(n8285), .ZN(n8344) );
  INV_X1 U9916 ( .A(n8344), .ZN(n8323) );
  INV_X1 U9917 ( .A(n8287), .ZN(n8288) );
  NAND4_X1 U9918 ( .A1(n8290), .A2(n8289), .A3(n4411), .A4(n8288), .ZN(n8292)
         );
  OAI21_X1 U9919 ( .B1(n8293), .B2(n8292), .A(n8291), .ZN(n8296) );
  NAND3_X1 U9920 ( .A1(n8296), .A2(n8295), .A3(n8294), .ZN(n8299) );
  AOI21_X1 U9921 ( .B1(n8299), .B2(n8298), .A(n8297), .ZN(n8303) );
  INV_X1 U9922 ( .A(n8300), .ZN(n8301) );
  NOR3_X1 U9923 ( .A1(n8303), .A2(n8302), .A3(n8301), .ZN(n8306) );
  OAI21_X1 U9924 ( .B1(n8306), .B2(n8305), .A(n8304), .ZN(n8309) );
  AOI21_X1 U9925 ( .B1(n8309), .B2(n8308), .A(n8307), .ZN(n8312) );
  OAI21_X1 U9926 ( .B1(n8312), .B2(n8311), .A(n8310), .ZN(n8322) );
  NAND3_X1 U9927 ( .A1(n8315), .A2(n8314), .A3(n8313), .ZN(n8319) );
  INV_X1 U9928 ( .A(n8316), .ZN(n8318) );
  INV_X1 U9929 ( .A(n8343), .ZN(n8321) );
  AOI21_X1 U9930 ( .B1(n8323), .B2(n8322), .A(n8321), .ZN(n8328) );
  AND2_X1 U9931 ( .A1(n8325), .A2(n8324), .ZN(n8346) );
  INV_X1 U9932 ( .A(n8346), .ZN(n8327) );
  OAI21_X1 U9933 ( .B1(n8328), .B2(n8327), .A(n8326), .ZN(n8332) );
  INV_X1 U9934 ( .A(n8349), .ZN(n8331) );
  INV_X1 U9935 ( .A(n8334), .ZN(n8340) );
  INV_X1 U9936 ( .A(n8335), .ZN(n8356) );
  NOR2_X1 U9937 ( .A1(n8375), .A2(n8336), .ZN(n8337) );
  OAI21_X1 U9938 ( .B1(n8356), .B2(n9550), .A(n8337), .ZN(n8338) );
  INV_X1 U9939 ( .A(n8338), .ZN(n8339) );
  INV_X1 U9940 ( .A(n8342), .ZN(n9657) );
  OAI21_X1 U9941 ( .B1(n9657), .B2(n8344), .A(n8343), .ZN(n8347) );
  AOI21_X1 U9942 ( .B1(n8347), .B2(n8346), .A(n8345), .ZN(n8350) );
  OAI22_X1 U9943 ( .A1(n8350), .A2(n8349), .B1(n9740), .B2(n8348), .ZN(n8353)
         );
  OAI21_X1 U9944 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(n8357) );
  AOI211_X1 U9945 ( .C1(n8357), .C2(n8356), .A(n8355), .B(n8354), .ZN(n8359)
         );
  NOR2_X1 U9946 ( .A1(n8363), .A2(n8362), .ZN(n8364) );
  NOR3_X1 U9947 ( .A1(n8374), .A2(n8373), .A3(n8372), .ZN(n8377) );
  OAI21_X1 U9948 ( .B1(n8378), .B2(n8375), .A(P1_B_REG_SCAN_IN), .ZN(n8376) );
  INV_X1 U9949 ( .A(n8379), .ZN(n8385) );
  OAI222_X1 U9950 ( .A1(n9866), .A2(n8380), .B1(n9864), .B2(n8385), .C1(n6139), 
        .C2(P1_U3086), .ZN(P1_U3325) );
  INV_X1 U9951 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n8382) );
  AOI22_X1 U9952 ( .A1(n8383), .A2(n8382), .B1(n8381), .B2(n5703), .ZN(
        P2_U3376) );
  OAI222_X1 U9953 ( .A1(n8387), .A2(n8386), .B1(n7852), .B2(n8385), .C1(
        P2_U3151), .C2(n8384), .ZN(P2_U3265) );
  INV_X1 U9954 ( .A(n8388), .ZN(n9185) );
  OAI222_X1 U9955 ( .A1(n9866), .A2(n8389), .B1(n9864), .B2(n9185), .C1(n4319), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  NOR2_X1 U9956 ( .A1(n8390), .A2(n8989), .ZN(n8754) );
  NOR2_X1 U9957 ( .A1(n5732), .A2(n8991), .ZN(n8392) );
  AOI211_X1 U9958 ( .C1(n8993), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8754), .B(
        n8392), .ZN(n8395) );
  NAND2_X1 U9959 ( .A1(n8393), .A2(n8764), .ZN(n8394) );
  OAI211_X1 U9960 ( .C1(n8396), .C2(n8993), .A(n8395), .B(n8394), .ZN(P2_U3204) );
  OAI222_X1 U9961 ( .A1(n7852), .A2(n8398), .B1(n4779), .B2(P2_U3151), .C1(
        n8397), .C2(n8387), .ZN(P2_U3266) );
  XNOR2_X1 U9962 ( .A(n8774), .B(n8399), .ZN(n8400) );
  XNOR2_X1 U9963 ( .A(n8410), .B(n8400), .ZN(n8406) );
  INV_X1 U9964 ( .A(n8406), .ZN(n8401) );
  NAND2_X1 U9965 ( .A1(n8401), .A2(n8557), .ZN(n8414) );
  NAND2_X1 U9966 ( .A1(n8405), .A2(n8786), .ZN(n8402) );
  NAND2_X1 U9967 ( .A1(n8599), .A2(n8587), .ZN(n8404) );
  AOI22_X1 U9968 ( .A1(n8760), .A2(n8593), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8403) );
  OAI211_X1 U9969 ( .C1(n8576), .C2(n8590), .A(n8404), .B(n8403), .ZN(n8409)
         );
  INV_X1 U9970 ( .A(n8405), .ZN(n8407) );
  NOR4_X1 U9971 ( .A1(n8407), .A2(n8406), .A3(n8576), .A4(n8581), .ZN(n8408)
         );
  AOI211_X1 U9972 ( .C1(n8410), .C2(n8578), .A(n8409), .B(n8408), .ZN(n8411)
         );
  OAI211_X1 U9973 ( .C1(n8414), .C2(n8413), .A(n8412), .B(n8411), .ZN(P2_U3160) );
  XOR2_X1 U9974 ( .A(n8416), .B(n8415), .Z(n8421) );
  AOI22_X1 U9975 ( .A1(n8587), .A2(n8939), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8418) );
  NAND2_X1 U9976 ( .A1(n8593), .A2(n8941), .ZN(n8417) );
  OAI211_X1 U9977 ( .C1(n8968), .C2(n8590), .A(n8418), .B(n8417), .ZN(n8419)
         );
  AOI21_X1 U9978 ( .B1(n9160), .B2(n8578), .A(n8419), .ZN(n8420) );
  OAI21_X1 U9979 ( .B1(n8421), .B2(n8581), .A(n8420), .ZN(P2_U3155) );
  NOR2_X1 U9980 ( .A1(n8424), .A2(n8423), .ZN(n8430) );
  AOI22_X1 U9981 ( .A1(n8861), .A2(n8572), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8426) );
  NAND2_X1 U9982 ( .A1(n8829), .A2(n8593), .ZN(n8425) );
  OAI211_X1 U9983 ( .C1(n8427), .C2(n8575), .A(n8426), .B(n8425), .ZN(n8428)
         );
  AOI21_X1 U9984 ( .B1(n9107), .B2(n8578), .A(n8428), .ZN(n8429) );
  OAI21_X1 U9985 ( .B1(n8430), .B2(n8581), .A(n8429), .ZN(P2_U3156) );
  XNOR2_X1 U9986 ( .A(n8459), .B(n8537), .ZN(n8432) );
  NAND2_X1 U9987 ( .A1(n8432), .A2(n8433), .ZN(n8535) );
  OAI21_X1 U9988 ( .B1(n8433), .B2(n8432), .A(n8535), .ZN(n8434) );
  NAND2_X1 U9989 ( .A1(n8434), .A2(n8557), .ZN(n8441) );
  INV_X1 U9990 ( .A(n8983), .ZN(n8439) );
  NAND2_X1 U9991 ( .A1(n8587), .A2(n8600), .ZN(n8436) );
  OAI211_X1 U9992 ( .C1(n8437), .C2(n8590), .A(n8436), .B(n8435), .ZN(n8438)
         );
  AOI21_X1 U9993 ( .B1(n8439), .B2(n8593), .A(n8438), .ZN(n8440) );
  OAI211_X1 U9994 ( .C1(n9066), .C2(n8596), .A(n8441), .B(n8440), .ZN(P2_U3157) );
  XOR2_X1 U9995 ( .A(n8443), .B(n4439), .Z(n8450) );
  NAND2_X1 U9996 ( .A1(n8879), .A2(n8587), .ZN(n8445) );
  OAI211_X1 U9997 ( .C1(n8446), .C2(n8590), .A(n8445), .B(n8444), .ZN(n8447)
         );
  AOI21_X1 U9998 ( .B1(n8882), .B2(n8593), .A(n8447), .ZN(n8449) );
  NAND2_X1 U9999 ( .A1(n9130), .A2(n8578), .ZN(n8448) );
  OAI211_X1 U10000 ( .C1(n8450), .C2(n8581), .A(n8449), .B(n8448), .ZN(
        P2_U3159) );
  XOR2_X1 U10001 ( .A(n8452), .B(n8451), .Z(n8458) );
  AOI22_X1 U10002 ( .A1(n8861), .A2(n8587), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8454) );
  NAND2_X1 U10003 ( .A1(n8593), .A2(n8864), .ZN(n8453) );
  OAI211_X1 U10004 ( .C1(n8455), .C2(n8590), .A(n8454), .B(n8453), .ZN(n8456)
         );
  AOI21_X1 U10005 ( .B1(n9118), .B2(n8578), .A(n8456), .ZN(n8457) );
  OAI21_X1 U10006 ( .B1(n8458), .B2(n8581), .A(n8457), .ZN(P2_U3163) );
  INV_X1 U10007 ( .A(n8459), .ZN(n8460) );
  NAND2_X1 U10008 ( .A1(n8460), .A2(n8537), .ZN(n8534) );
  XNOR2_X1 U10009 ( .A(n8462), .B(n8461), .ZN(n8533) );
  NAND3_X1 U10010 ( .A1(n8535), .A2(n8534), .A3(n8533), .ZN(n8532) );
  NAND2_X1 U10011 ( .A1(n8532), .A2(n8463), .ZN(n8468) );
  INV_X1 U10012 ( .A(n8464), .ZN(n8465) );
  NOR2_X1 U10013 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  XNOR2_X1 U10014 ( .A(n8468), .B(n8467), .ZN(n8475) );
  NAND2_X1 U10015 ( .A1(n8587), .A2(n8938), .ZN(n8470) );
  OAI211_X1 U10016 ( .C1(n8970), .C2(n8590), .A(n8470), .B(n8469), .ZN(n8473)
         );
  INV_X1 U10017 ( .A(n9058), .ZN(n8471) );
  NOR2_X1 U10018 ( .A1(n8471), .A2(n8596), .ZN(n8472) );
  AOI211_X1 U10019 ( .C1(n8976), .C2(n8593), .A(n8473), .B(n8472), .ZN(n8474)
         );
  OAI21_X1 U10020 ( .B1(n8475), .B2(n8581), .A(n8474), .ZN(P2_U3164) );
  INV_X1 U10021 ( .A(n9148), .ZN(n8483) );
  OAI211_X1 U10022 ( .C1(n8478), .C2(n8477), .A(n8476), .B(n8557), .ZN(n8482)
         );
  NAND2_X1 U10023 ( .A1(n8587), .A2(n8889), .ZN(n8479) );
  NAND2_X1 U10024 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8712) );
  OAI211_X1 U10025 ( .C1(n8912), .C2(n8590), .A(n8479), .B(n8712), .ZN(n8480)
         );
  AOI21_X1 U10026 ( .B1(n8917), .B2(n8593), .A(n8480), .ZN(n8481) );
  OAI211_X1 U10027 ( .C1(n8483), .C2(n8596), .A(n8482), .B(n8481), .ZN(
        P2_U3166) );
  AOI21_X1 U10028 ( .B1(n8485), .B2(n8484), .A(n4343), .ZN(n8491) );
  NAND2_X1 U10029 ( .A1(n8587), .A2(n8899), .ZN(n8486) );
  NAND2_X1 U10030 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8725) );
  OAI211_X1 U10031 ( .C1(n8590), .C2(n8487), .A(n8486), .B(n8725), .ZN(n8488)
         );
  AOI21_X1 U10032 ( .B1(n8903), .B2(n8593), .A(n8488), .ZN(n8490) );
  NAND2_X1 U10033 ( .A1(n9142), .A2(n8578), .ZN(n8489) );
  OAI211_X1 U10034 ( .C1(n8491), .C2(n8581), .A(n8490), .B(n8489), .ZN(
        P2_U3168) );
  INV_X1 U10035 ( .A(n8492), .ZN(n8493) );
  AOI21_X1 U10036 ( .B1(n8587), .B2(n8601), .A(n8493), .ZN(n8497) );
  INV_X1 U10037 ( .A(n8990), .ZN(n8494) );
  NAND2_X1 U10038 ( .A1(n8593), .A2(n8494), .ZN(n8496) );
  NAND2_X1 U10039 ( .A1(n8572), .A2(n8603), .ZN(n8495) );
  NAND3_X1 U10040 ( .A1(n8497), .A2(n8496), .A3(n8495), .ZN(n8501) );
  AOI211_X1 U10041 ( .C1(n8499), .C2(n8498), .A(n8581), .B(n4414), .ZN(n8500)
         );
  AOI211_X1 U10042 ( .C1(n8502), .C2(n8578), .A(n8501), .B(n8500), .ZN(n8503)
         );
  INV_X1 U10043 ( .A(n8503), .ZN(P2_U3171) );
  NAND2_X1 U10044 ( .A1(n8505), .A2(n8504), .ZN(n8506) );
  XOR2_X1 U10045 ( .A(n8507), .B(n8506), .Z(n8513) );
  AOI22_X1 U10046 ( .A1(n8870), .A2(n8587), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8509) );
  NAND2_X1 U10047 ( .A1(n8593), .A2(n8873), .ZN(n8508) );
  OAI211_X1 U10048 ( .C1(n8510), .C2(n8590), .A(n8509), .B(n8508), .ZN(n8511)
         );
  AOI21_X1 U10049 ( .B1(n9124), .B2(n8578), .A(n8511), .ZN(n8512) );
  OAI21_X1 U10050 ( .B1(n8513), .B2(n8581), .A(n8512), .ZN(P2_U3173) );
  XOR2_X1 U10051 ( .A(n8515), .B(n8514), .Z(n8521) );
  NAND2_X1 U10052 ( .A1(n8587), .A2(n8953), .ZN(n8516) );
  NAND2_X1 U10053 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8663) );
  OAI211_X1 U10054 ( .C1(n8517), .C2(n8590), .A(n8516), .B(n8663), .ZN(n8518)
         );
  AOI21_X1 U10055 ( .B1(n8957), .B2(n8593), .A(n8518), .ZN(n8520) );
  NAND2_X1 U10056 ( .A1(n9166), .A2(n8578), .ZN(n8519) );
  OAI211_X1 U10057 ( .C1(n8521), .C2(n8581), .A(n8520), .B(n8519), .ZN(
        P2_U3174) );
  NAND2_X1 U10058 ( .A1(n8524), .A2(n8523), .ZN(n8525) );
  XNOR2_X1 U10059 ( .A(n8522), .B(n8525), .ZN(n8531) );
  AOI22_X1 U10060 ( .A1(n8870), .A2(n8572), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8527) );
  NAND2_X1 U10061 ( .A1(n8849), .A2(n8593), .ZN(n8526) );
  OAI211_X1 U10062 ( .C1(n8528), .C2(n8575), .A(n8527), .B(n8526), .ZN(n8529)
         );
  AOI21_X1 U10063 ( .B1(n9113), .B2(n8578), .A(n8529), .ZN(n8530) );
  OAI21_X1 U10064 ( .B1(n8531), .B2(n8581), .A(n8530), .ZN(P2_U3175) );
  NAND2_X1 U10065 ( .A1(n8532), .A2(n8557), .ZN(n8545) );
  AOI21_X1 U10066 ( .B1(n8535), .B2(n8534), .A(n8533), .ZN(n8544) );
  NAND2_X1 U10067 ( .A1(n8587), .A2(n8951), .ZN(n8536) );
  NAND2_X1 U10068 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8647) );
  OAI211_X1 U10069 ( .C1(n8537), .C2(n8590), .A(n8536), .B(n8647), .ZN(n8541)
         );
  INV_X1 U10070 ( .A(n8538), .ZN(n8539) );
  NOR2_X1 U10071 ( .A1(n8596), .A2(n8539), .ZN(n8540) );
  AOI211_X1 U10072 ( .C1(n8542), .C2(n8593), .A(n8541), .B(n8540), .ZN(n8543)
         );
  OAI21_X1 U10073 ( .B1(n8545), .B2(n8544), .A(n8543), .ZN(P2_U3176) );
  INV_X1 U10074 ( .A(n9136), .ZN(n8556) );
  INV_X1 U10075 ( .A(n8546), .ZN(n8548) );
  NOR3_X1 U10076 ( .A1(n4343), .A2(n8548), .A3(n8547), .ZN(n8551) );
  OAI21_X1 U10077 ( .B1(n8551), .B2(n4384), .A(n8557), .ZN(n8555) );
  NAND2_X1 U10078 ( .A1(n8890), .A2(n8587), .ZN(n8552) );
  NAND2_X1 U10079 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8746) );
  OAI211_X1 U10080 ( .C1(n8913), .C2(n8590), .A(n8552), .B(n8746), .ZN(n8553)
         );
  AOI21_X1 U10081 ( .B1(n8892), .B2(n8593), .A(n8553), .ZN(n8554) );
  OAI211_X1 U10082 ( .C1(n8556), .C2(n8596), .A(n8555), .B(n8554), .ZN(
        P2_U3178) );
  OAI211_X1 U10083 ( .C1(n8560), .C2(n8559), .A(n8558), .B(n8557), .ZN(n8565)
         );
  AND2_X1 U10084 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10089) );
  AOI21_X1 U10085 ( .B1(n8587), .B2(n8604), .A(n10089), .ZN(n8564) );
  AOI22_X1 U10086 ( .A1(n8572), .A2(n8606), .B1(n8578), .B2(n9068), .ZN(n8563)
         );
  NAND2_X1 U10087 ( .A1(n8593), .A2(n8561), .ZN(n8562) );
  NAND4_X1 U10088 ( .A1(n8565), .A2(n8564), .A3(n8563), .A4(n8562), .ZN(
        P2_U3179) );
  INV_X1 U10089 ( .A(n8566), .ZN(n8568) );
  INV_X1 U10090 ( .A(n8569), .ZN(n8570) );
  AOI21_X1 U10091 ( .B1(n8571), .B2(n4976), .A(n8570), .ZN(n8580) );
  AOI22_X1 U10092 ( .A1(n8815), .A2(n8572), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8574) );
  NAND2_X1 U10093 ( .A1(n8789), .A2(n8593), .ZN(n8573) );
  OAI211_X1 U10094 ( .C1(n8576), .C2(n8575), .A(n8574), .B(n8573), .ZN(n8577)
         );
  AOI21_X1 U10095 ( .B1(n9090), .B2(n8578), .A(n8577), .ZN(n8579) );
  OAI21_X1 U10096 ( .B1(n8580), .B2(n8581), .A(n8579), .ZN(P2_U3180) );
  INV_X1 U10097 ( .A(n9154), .ZN(n8597) );
  AOI21_X1 U10098 ( .B1(n8583), .B2(n8582), .A(n8581), .ZN(n8586) );
  NAND2_X1 U10099 ( .A1(n8586), .A2(n8585), .ZN(n8595) );
  NAND2_X1 U10100 ( .A1(n8587), .A2(n8930), .ZN(n8589) );
  NAND2_X1 U10101 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8698) );
  OAI211_X1 U10102 ( .C1(n8591), .C2(n8590), .A(n8589), .B(n8698), .ZN(n8592)
         );
  AOI21_X1 U10103 ( .B1(n8934), .B2(n8593), .A(n8592), .ZN(n8594) );
  OAI211_X1 U10104 ( .C1(n8597), .C2(n8596), .A(n8595), .B(n8594), .ZN(
        P2_U3181) );
  MUX2_X1 U10105 ( .A(n8598), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8743), .Z(
        P2_U3521) );
  MUX2_X1 U10106 ( .A(n8599), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8743), .Z(
        P2_U3520) );
  MUX2_X1 U10107 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8774), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10108 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8786), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10109 ( .A(n8803), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8743), .Z(
        P2_U3517) );
  MUX2_X1 U10110 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8815), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10111 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8826), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10112 ( .A(n8846), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8743), .Z(
        P2_U3514) );
  MUX2_X1 U10113 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8861), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10114 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8870), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10115 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8879), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10116 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8899), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8889), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10118 ( .A(n8930), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8743), .Z(
        P2_U3507) );
  MUX2_X1 U10119 ( .A(n8939), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8743), .Z(
        P2_U3506) );
  MUX2_X1 U10120 ( .A(n8953), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8743), .Z(
        P2_U3505) );
  MUX2_X1 U10121 ( .A(n8938), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8743), .Z(
        P2_U3504) );
  MUX2_X1 U10122 ( .A(n8951), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8743), .Z(
        P2_U3503) );
  MUX2_X1 U10123 ( .A(n8600), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8743), .Z(
        P2_U3502) );
  MUX2_X1 U10124 ( .A(n8601), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8743), .Z(
        P2_U3501) );
  MUX2_X1 U10125 ( .A(n8602), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8743), .Z(
        P2_U3500) );
  MUX2_X1 U10126 ( .A(n8603), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8743), .Z(
        P2_U3499) );
  MUX2_X1 U10127 ( .A(n8604), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8743), .Z(
        P2_U3498) );
  MUX2_X1 U10128 ( .A(n8605), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8743), .Z(
        P2_U3497) );
  MUX2_X1 U10129 ( .A(n8606), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8743), .Z(
        P2_U3496) );
  MUX2_X1 U10130 ( .A(n8607), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8743), .Z(
        P2_U3494) );
  MUX2_X1 U10131 ( .A(n8608), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8743), .Z(
        P2_U3493) );
  MUX2_X1 U10132 ( .A(n8609), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8743), .Z(
        P2_U3492) );
  MUX2_X1 U10133 ( .A(n8610), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8743), .Z(
        P2_U3491) );
  OAI22_X1 U10134 ( .A1(n10111), .A2(n6641), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8611), .ZN(n8612) );
  AOI21_X1 U10135 ( .B1(n10118), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n8612), .ZN(
        n8626) );
  OAI21_X1 U10136 ( .B1(n8615), .B2(n8614), .A(n8613), .ZN(n8620) );
  OAI21_X1 U10137 ( .B1(n8618), .B2(n8617), .A(n8616), .ZN(n8619) );
  AOI22_X1 U10138 ( .A1(n10095), .A2(n8620), .B1(n10114), .B2(n8619), .ZN(
        n8625) );
  OAI211_X1 U10139 ( .C1(n8623), .C2(n8622), .A(n6751), .B(n8621), .ZN(n8624)
         );
  NAND3_X1 U10140 ( .A1(n8626), .A2(n8625), .A3(n8624), .ZN(P2_U3184) );
  NOR2_X1 U10141 ( .A1(n8748), .A2(n9878), .ZN(n8627) );
  AOI211_X1 U10142 ( .C1(n8630), .C2(n8629), .A(n8628), .B(n8627), .ZN(n8644)
         );
  OAI211_X1 U10143 ( .C1(n8633), .C2(n8632), .A(n8631), .B(n6751), .ZN(n8643)
         );
  OAI21_X1 U10144 ( .B1(n8636), .B2(n8635), .A(n8634), .ZN(n8641) );
  OAI21_X1 U10145 ( .B1(n8639), .B2(n8638), .A(n8637), .ZN(n8640) );
  AOI22_X1 U10146 ( .A1(n10095), .A2(n8641), .B1(n10114), .B2(n8640), .ZN(
        n8642) );
  NAND3_X1 U10147 ( .A1(n8644), .A2(n8643), .A3(n8642), .ZN(P2_U3186) );
  XNOR2_X1 U10148 ( .A(n8646), .B(n8645), .ZN(n8658) );
  OAI21_X1 U10149 ( .B1(n10111), .B2(n8648), .A(n8647), .ZN(n8652) );
  AOI21_X1 U10150 ( .B1(n10261), .B2(n8649), .A(n7805), .ZN(n8650) );
  NOR2_X1 U10151 ( .A1(n8650), .A2(n8668), .ZN(n8651) );
  AOI211_X1 U10152 ( .C1(n10118), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n8652), .B(
        n8651), .ZN(n8657) );
  XNOR2_X1 U10153 ( .A(n8654), .B(n8653), .ZN(n8655) );
  NAND2_X1 U10154 ( .A1(n8655), .A2(n6751), .ZN(n8656) );
  OAI211_X1 U10155 ( .C1(n8658), .C2(n10106), .A(n8657), .B(n8656), .ZN(
        P2_U3193) );
  XNOR2_X1 U10156 ( .A(n8659), .B(n10237), .ZN(n8674) );
  OAI21_X1 U10157 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8672) );
  NAND2_X1 U10158 ( .A1(n10118), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8664) );
  OAI211_X1 U10159 ( .C1(n10111), .C2(n8665), .A(n8664), .B(n8663), .ZN(n8671)
         );
  NAND2_X1 U10160 ( .A1(n8667), .A2(n8962), .ZN(n8669) );
  AOI21_X1 U10161 ( .B1(n8666), .B2(n8669), .A(n8668), .ZN(n8670) );
  AOI211_X1 U10162 ( .C1(n6751), .C2(n8672), .A(n8671), .B(n8670), .ZN(n8673)
         );
  OAI21_X1 U10163 ( .B1(n8674), .B2(n10106), .A(n8673), .ZN(P2_U3195) );
  XOR2_X1 U10164 ( .A(n8676), .B(n8675), .Z(n8691) );
  AND3_X1 U10165 ( .A1(n8666), .A2(n8678), .A3(n8677), .ZN(n8679) );
  OAI21_X1 U10166 ( .B1(n8680), .B2(n8679), .A(n10114), .ZN(n8690) );
  OAI21_X1 U10167 ( .B1(n8683), .B2(n8682), .A(n8681), .ZN(n8688) );
  NAND2_X1 U10168 ( .A1(n10118), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U10169 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n8684) );
  OAI211_X1 U10170 ( .C1(n10111), .C2(n8686), .A(n8685), .B(n8684), .ZN(n8687)
         );
  AOI21_X1 U10171 ( .B1(n8688), .B2(n6751), .A(n8687), .ZN(n8689) );
  OAI211_X1 U10172 ( .C1(n8691), .C2(n10106), .A(n8690), .B(n8689), .ZN(
        P2_U3196) );
  XNOR2_X1 U10173 ( .A(n8692), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n8704) );
  OAI21_X1 U10174 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8694), .A(n8693), .ZN(
        n8695) );
  NAND2_X1 U10175 ( .A1(n8695), .A2(n10114), .ZN(n8703) );
  XNOR2_X1 U10176 ( .A(n8697), .B(n8696), .ZN(n8701) );
  NAND2_X1 U10177 ( .A1(n10118), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8699) );
  OAI211_X1 U10178 ( .C1(n10111), .C2(n4894), .A(n8699), .B(n8698), .ZN(n8700)
         );
  AOI21_X1 U10179 ( .B1(n8701), .B2(n6751), .A(n8700), .ZN(n8702) );
  OAI211_X1 U10180 ( .C1(n8704), .C2(n10106), .A(n8703), .B(n8702), .ZN(
        P2_U3197) );
  XOR2_X1 U10181 ( .A(n8706), .B(n8705), .Z(n8719) );
  NOR2_X1 U10182 ( .A1(n8708), .A2(n8707), .ZN(n8709) );
  OAI21_X1 U10183 ( .B1(n4390), .B2(n8709), .A(n10114), .ZN(n8718) );
  XNOR2_X1 U10184 ( .A(n8711), .B(n8710), .ZN(n8716) );
  NAND2_X1 U10185 ( .A1(n10118), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8713) );
  OAI211_X1 U10186 ( .C1(n8714), .C2(n10111), .A(n8713), .B(n8712), .ZN(n8715)
         );
  AOI21_X1 U10187 ( .B1(n8716), .B2(n6751), .A(n8715), .ZN(n8717) );
  OAI211_X1 U10188 ( .C1(n8719), .C2(n10106), .A(n8718), .B(n8717), .ZN(
        P2_U3198) );
  XNOR2_X1 U10189 ( .A(n8720), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8732) );
  OAI21_X1 U10190 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8721), .A(n8737), .ZN(
        n8722) );
  NAND2_X1 U10191 ( .A1(n8722), .A2(n10114), .ZN(n8731) );
  XNOR2_X1 U10192 ( .A(n8724), .B(n8723), .ZN(n8729) );
  NAND2_X1 U10193 ( .A1(n10118), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8726) );
  OAI211_X1 U10194 ( .C1(n10111), .C2(n8727), .A(n8726), .B(n8725), .ZN(n8728)
         );
  AOI21_X1 U10195 ( .B1(n8729), .B2(n6751), .A(n8728), .ZN(n8730) );
  OAI211_X1 U10196 ( .C1(n8732), .C2(n10106), .A(n8731), .B(n8730), .ZN(
        P2_U3199) );
  AND3_X1 U10197 ( .A1(n8737), .A2(n8736), .A3(n8735), .ZN(n8738) );
  INV_X1 U10198 ( .A(n8740), .ZN(n8742) );
  NAND2_X1 U10199 ( .A1(n8742), .A2(n8741), .ZN(n8745) );
  OAI21_X1 U10200 ( .B1(n8745), .B2(n8743), .A(n10111), .ZN(n8749) );
  INV_X1 U10201 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U10202 ( .A1(n9075), .A2(n8977), .ZN(n8755) );
  INV_X1 U10203 ( .A(n8751), .ZN(n8752) );
  AOI21_X1 U10204 ( .B1(n9076), .B2(n9008), .A(n8754), .ZN(n8758) );
  OAI211_X1 U10205 ( .C1(n9008), .C2(n8756), .A(n8755), .B(n8758), .ZN(
        P2_U3202) );
  NAND2_X1 U10206 ( .A1(n8993), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8757) );
  OAI211_X1 U10207 ( .C1(n9081), .C2(n8991), .A(n8758), .B(n8757), .ZN(
        P2_U3203) );
  INV_X1 U10208 ( .A(n8759), .ZN(n8767) );
  AOI22_X1 U10209 ( .A1(n8760), .A2(n9003), .B1(n8993), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8761) );
  OAI21_X1 U10210 ( .B1(n8762), .B2(n8991), .A(n8761), .ZN(n8763) );
  AOI21_X1 U10211 ( .B1(n8765), .B2(n8764), .A(n8763), .ZN(n8766) );
  OAI21_X1 U10212 ( .B1(n8767), .B2(n8993), .A(n8766), .ZN(P2_U3205) );
  XNOR2_X1 U10213 ( .A(n8769), .B(n8768), .ZN(n9087) );
  NAND2_X1 U10214 ( .A1(n8771), .A2(n8770), .ZN(n8772) );
  NAND3_X1 U10215 ( .A1(n8773), .A2(n8949), .A3(n8772), .ZN(n8776) );
  AOI22_X1 U10216 ( .A1(n8774), .A2(n8954), .B1(n8952), .B2(n8803), .ZN(n8775)
         );
  MUX2_X1 U10217 ( .A(n9082), .B(n8777), .S(n8993), .Z(n8780) );
  AOI22_X1 U10218 ( .A1(n9084), .A2(n8977), .B1(n9003), .B2(n8778), .ZN(n8779)
         );
  OAI211_X1 U10219 ( .C1(n9087), .C2(n8980), .A(n8780), .B(n8779), .ZN(
        P2_U3206) );
  XOR2_X1 U10220 ( .A(n8784), .B(n8781), .Z(n9093) );
  AND2_X1 U10221 ( .A1(n8783), .A2(n8782), .ZN(n8785) );
  XNOR2_X1 U10222 ( .A(n8785), .B(n8784), .ZN(n8787) );
  AOI222_X1 U10223 ( .A1(n8949), .A2(n8787), .B1(n8786), .B2(n8954), .C1(n8815), .C2(n8952), .ZN(n9088) );
  MUX2_X1 U10224 ( .A(n8788), .B(n9088), .S(n9008), .Z(n8791) );
  AOI22_X1 U10225 ( .A1(n9090), .A2(n8977), .B1(n9003), .B2(n8789), .ZN(n8790)
         );
  OAI211_X1 U10226 ( .C1(n9093), .C2(n8980), .A(n8791), .B(n8790), .ZN(
        P2_U3207) );
  XOR2_X1 U10227 ( .A(n8792), .B(n8798), .Z(n9097) );
  OR2_X1 U10228 ( .A1(n8793), .A2(n8794), .ZN(n8797) );
  NAND2_X1 U10229 ( .A1(n8797), .A2(n8795), .ZN(n8801) );
  NAND2_X1 U10230 ( .A1(n8797), .A2(n8796), .ZN(n8799) );
  NAND2_X1 U10231 ( .A1(n8799), .A2(n8798), .ZN(n8800) );
  NAND2_X1 U10232 ( .A1(n8801), .A2(n8800), .ZN(n8802) );
  NAND2_X1 U10233 ( .A1(n8802), .A2(n8949), .ZN(n8805) );
  AOI22_X1 U10234 ( .A1(n8803), .A2(n8954), .B1(n8826), .B2(n8952), .ZN(n8804)
         );
  NAND2_X1 U10235 ( .A1(n8805), .A2(n8804), .ZN(n9094) );
  NOR2_X1 U10236 ( .A1(n9096), .A2(n8817), .ZN(n8806) );
  OAI21_X1 U10237 ( .B1(n9094), .B2(n8806), .A(n9008), .ZN(n8809) );
  AOI22_X1 U10238 ( .A1(n8807), .A2(n9003), .B1(n8993), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8808) );
  OAI211_X1 U10239 ( .C1(n9097), .C2(n8980), .A(n8809), .B(n8808), .ZN(
        P2_U3208) );
  AOI21_X1 U10240 ( .B1(n8823), .B2(n8812), .A(n8811), .ZN(n8813) );
  XOR2_X1 U10241 ( .A(n8814), .B(n8813), .Z(n9105) );
  XNOR2_X1 U10242 ( .A(n8793), .B(n8814), .ZN(n8816) );
  AOI222_X1 U10243 ( .A1(n8949), .A2(n8816), .B1(n8815), .B2(n8954), .C1(n8846), .C2(n8952), .ZN(n9100) );
  OAI21_X1 U10244 ( .B1(n8818), .B2(n8817), .A(n9100), .ZN(n8819) );
  NAND2_X1 U10245 ( .A1(n8819), .A2(n9008), .ZN(n8822) );
  AOI22_X1 U10246 ( .A1(n8820), .A2(n9003), .B1(n8993), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8821) );
  OAI211_X1 U10247 ( .C1(n9105), .C2(n8980), .A(n8822), .B(n8821), .ZN(
        P2_U3209) );
  XOR2_X1 U10248 ( .A(n8825), .B(n8823), .Z(n9110) );
  INV_X1 U10249 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8828) );
  XOR2_X1 U10250 ( .A(n8825), .B(n8824), .Z(n8827) );
  AOI222_X1 U10251 ( .A1(n8949), .A2(n8827), .B1(n8826), .B2(n8954), .C1(n8861), .C2(n8952), .ZN(n9106) );
  MUX2_X1 U10252 ( .A(n8828), .B(n9106), .S(n9008), .Z(n8831) );
  AOI22_X1 U10253 ( .A1(n9107), .A2(n8977), .B1(n9003), .B2(n8829), .ZN(n8830)
         );
  OAI211_X1 U10254 ( .C1(n9110), .C2(n8980), .A(n8831), .B(n8830), .ZN(
        P2_U3210) );
  OR2_X1 U10255 ( .A1(n8867), .A2(n8833), .ZN(n8853) );
  NAND2_X1 U10256 ( .A1(n8853), .A2(n8834), .ZN(n8837) );
  NAND3_X1 U10257 ( .A1(n8837), .A2(n8836), .A3(n8835), .ZN(n8838) );
  NAND2_X1 U10258 ( .A1(n8839), .A2(n8838), .ZN(n9116) );
  INV_X1 U10259 ( .A(n8869), .ZN(n8840) );
  OAI21_X1 U10260 ( .B1(n8840), .B2(n8856), .A(n8854), .ZN(n8860) );
  INV_X1 U10261 ( .A(n8841), .ZN(n8842) );
  NAND3_X1 U10262 ( .A1(n8860), .A2(n8843), .A3(n8842), .ZN(n8845) );
  NAND2_X1 U10263 ( .A1(n8845), .A2(n8844), .ZN(n8847) );
  AOI222_X1 U10264 ( .A1(n8949), .A2(n8847), .B1(n8846), .B2(n8954), .C1(n8870), .C2(n8952), .ZN(n9111) );
  MUX2_X1 U10265 ( .A(n8848), .B(n9111), .S(n9008), .Z(n8851) );
  AOI22_X1 U10266 ( .A1(n9113), .A2(n8977), .B1(n9003), .B2(n8849), .ZN(n8850)
         );
  OAI211_X1 U10267 ( .C1(n9116), .C2(n8980), .A(n8851), .B(n8850), .ZN(
        P2_U3211) );
  NAND2_X1 U10268 ( .A1(n8853), .A2(n8852), .ZN(n8855) );
  XNOR2_X1 U10269 ( .A(n8855), .B(n8854), .ZN(n9121) );
  INV_X1 U10270 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8863) );
  INV_X1 U10271 ( .A(n8856), .ZN(n8857) );
  NAND3_X1 U10272 ( .A1(n8869), .A2(n8858), .A3(n8857), .ZN(n8859) );
  NAND2_X1 U10273 ( .A1(n8860), .A2(n8859), .ZN(n8862) );
  AOI222_X1 U10274 ( .A1(n8949), .A2(n8862), .B1(n8861), .B2(n8954), .C1(n8879), .C2(n8952), .ZN(n9117) );
  MUX2_X1 U10275 ( .A(n8863), .B(n9117), .S(n9008), .Z(n8866) );
  AOI22_X1 U10276 ( .A1(n9118), .A2(n8977), .B1(n9003), .B2(n8864), .ZN(n8865)
         );
  OAI211_X1 U10277 ( .C1(n9121), .C2(n8980), .A(n8866), .B(n8865), .ZN(
        P2_U3212) );
  XNOR2_X1 U10278 ( .A(n8867), .B(n8868), .ZN(n9127) );
  OAI21_X1 U10279 ( .B1(n4370), .B2(n4875), .A(n8869), .ZN(n8871) );
  AOI222_X1 U10280 ( .A1(n8949), .A2(n8871), .B1(n8870), .B2(n8954), .C1(n8890), .C2(n8952), .ZN(n9122) );
  MUX2_X1 U10281 ( .A(n8872), .B(n9122), .S(n9008), .Z(n8875) );
  AOI22_X1 U10282 ( .A1(n9124), .A2(n8977), .B1(n9003), .B2(n8873), .ZN(n8874)
         );
  OAI211_X1 U10283 ( .C1(n9127), .C2(n8980), .A(n8875), .B(n8874), .ZN(
        P2_U3213) );
  XNOR2_X1 U10284 ( .A(n8876), .B(n8878), .ZN(n9133) );
  INV_X1 U10285 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8881) );
  XNOR2_X1 U10286 ( .A(n8877), .B(n8878), .ZN(n8880) );
  AOI222_X1 U10287 ( .A1(n8949), .A2(n8880), .B1(n8879), .B2(n8954), .C1(n8899), .C2(n8952), .ZN(n9128) );
  MUX2_X1 U10288 ( .A(n8881), .B(n9128), .S(n9008), .Z(n8884) );
  AOI22_X1 U10289 ( .A1(n9130), .A2(n8977), .B1(n9003), .B2(n8882), .ZN(n8883)
         );
  OAI211_X1 U10290 ( .C1(n9133), .C2(n8980), .A(n8884), .B(n8883), .ZN(
        P2_U3214) );
  XNOR2_X1 U10291 ( .A(n8886), .B(n8885), .ZN(n9139) );
  XNOR2_X1 U10292 ( .A(n8888), .B(n8887), .ZN(n8891) );
  AOI222_X1 U10293 ( .A1(n8949), .A2(n8891), .B1(n8890), .B2(n8954), .C1(n8889), .C2(n8952), .ZN(n9134) );
  MUX2_X1 U10294 ( .A(n10246), .B(n9134), .S(n9008), .Z(n8894) );
  AOI22_X1 U10295 ( .A1(n9136), .A2(n8977), .B1(n9003), .B2(n8892), .ZN(n8893)
         );
  OAI211_X1 U10296 ( .C1(n9139), .C2(n8980), .A(n8894), .B(n8893), .ZN(
        P2_U3215) );
  XNOR2_X1 U10297 ( .A(n8895), .B(n8897), .ZN(n9145) );
  INV_X1 U10298 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8902) );
  OAI211_X1 U10299 ( .C1(n8898), .C2(n8897), .A(n8896), .B(n8949), .ZN(n8901)
         );
  AOI22_X1 U10300 ( .A1(n8899), .A2(n8954), .B1(n8952), .B2(n8930), .ZN(n8900)
         );
  MUX2_X1 U10301 ( .A(n8902), .B(n9140), .S(n9008), .Z(n8905) );
  AOI22_X1 U10302 ( .A1(n9142), .A2(n8977), .B1(n9003), .B2(n8903), .ZN(n8904)
         );
  OAI211_X1 U10303 ( .C1(n9145), .C2(n8980), .A(n8905), .B(n8904), .ZN(
        P2_U3216) );
  XNOR2_X1 U10304 ( .A(n8907), .B(n8906), .ZN(n9151) );
  NOR2_X1 U10305 ( .A1(n8908), .A2(n8926), .ZN(n8929) );
  NOR2_X1 U10306 ( .A1(n8929), .A2(n8909), .ZN(n8911) );
  XNOR2_X1 U10307 ( .A(n8911), .B(n8910), .ZN(n8915) );
  OAI22_X1 U10308 ( .A1(n8913), .A2(n8969), .B1(n8912), .B2(n8971), .ZN(n8914)
         );
  AOI21_X1 U10309 ( .B1(n8915), .B2(n8949), .A(n8914), .ZN(n9146) );
  MUX2_X1 U10310 ( .A(n8916), .B(n9146), .S(n9008), .Z(n8919) );
  AOI22_X1 U10311 ( .A1(n9148), .A2(n8977), .B1(n9003), .B2(n8917), .ZN(n8918)
         );
  OAI211_X1 U10312 ( .C1(n9151), .C2(n8980), .A(n8919), .B(n8918), .ZN(
        P2_U3217) );
  OR2_X1 U10313 ( .A1(n8920), .A2(n8921), .ZN(n8923) );
  NAND2_X1 U10314 ( .A1(n8923), .A2(n8922), .ZN(n8925) );
  INV_X1 U10315 ( .A(n8926), .ZN(n8924) );
  XNOR2_X1 U10316 ( .A(n8925), .B(n8924), .ZN(n9157) );
  INV_X1 U10317 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8933) );
  NAND2_X1 U10318 ( .A1(n8908), .A2(n8926), .ZN(n8927) );
  NAND2_X1 U10319 ( .A1(n8927), .A2(n8949), .ZN(n8928) );
  OR2_X1 U10320 ( .A1(n8929), .A2(n8928), .ZN(n8932) );
  AOI22_X1 U10321 ( .A1(n8930), .A2(n8954), .B1(n8952), .B2(n8953), .ZN(n8931)
         );
  MUX2_X1 U10322 ( .A(n8933), .B(n9152), .S(n9008), .Z(n8936) );
  AOI22_X1 U10323 ( .A1(n9154), .A2(n8977), .B1(n9003), .B2(n8934), .ZN(n8935)
         );
  OAI211_X1 U10324 ( .C1(n9157), .C2(n8980), .A(n8936), .B(n8935), .ZN(
        P2_U3218) );
  XNOR2_X1 U10325 ( .A(n8937), .B(n8943), .ZN(n8940) );
  AOI222_X1 U10326 ( .A1(n8949), .A2(n8940), .B1(n8939), .B2(n8954), .C1(n8938), .C2(n8952), .ZN(n9158) );
  AOI22_X1 U10327 ( .A1(n9160), .A2(n9002), .B1(n9003), .B2(n8941), .ZN(n8942)
         );
  AOI21_X1 U10328 ( .B1(n9158), .B2(n8942), .A(n8993), .ZN(n8946) );
  XOR2_X1 U10329 ( .A(n8920), .B(n8943), .Z(n9163) );
  OAI22_X1 U10330 ( .A1(n9163), .A2(n8980), .B1(n8944), .B2(n9008), .ZN(n8945)
         );
  OR2_X1 U10331 ( .A1(n8946), .A2(n8945), .ZN(P2_U3219) );
  INV_X1 U10332 ( .A(n8960), .ZN(n8947) );
  XNOR2_X1 U10333 ( .A(n8948), .B(n8947), .ZN(n8950) );
  NAND2_X1 U10334 ( .A1(n8950), .A2(n8949), .ZN(n8956) );
  AOI22_X1 U10335 ( .A1(n8954), .A2(n8953), .B1(n8952), .B2(n8951), .ZN(n8955)
         );
  AND2_X1 U10336 ( .A1(n8956), .A2(n8955), .ZN(n9164) );
  AOI22_X1 U10337 ( .A1(n9166), .A2(n9002), .B1(n9003), .B2(n8957), .ZN(n8958)
         );
  AOI21_X1 U10338 ( .B1(n9164), .B2(n8958), .A(n8993), .ZN(n8964) );
  CLKBUF_X1 U10339 ( .A(n8959), .Z(n8961) );
  XNOR2_X1 U10340 ( .A(n8961), .B(n8960), .ZN(n9170) );
  OAI22_X1 U10341 ( .A1(n9170), .A2(n8980), .B1(n8962), .B2(n9008), .ZN(n8963)
         );
  OR2_X1 U10342 ( .A1(n8964), .A2(n8963), .ZN(P2_U3220) );
  XOR2_X1 U10343 ( .A(n8972), .B(n8965), .Z(n8966) );
  OAI222_X1 U10344 ( .A1(n8971), .A2(n8970), .B1(n8969), .B2(n8968), .C1(n8967), .C2(n8966), .ZN(n9057) );
  OR2_X1 U10345 ( .A1(n8973), .A2(n8972), .ZN(n8974) );
  NAND2_X1 U10346 ( .A1(n8975), .A2(n8974), .ZN(n9174) );
  AOI22_X1 U10347 ( .A1(n8993), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n9003), .B2(
        n8976), .ZN(n8979) );
  NAND2_X1 U10348 ( .A1(n9058), .A2(n8977), .ZN(n8978) );
  OAI211_X1 U10349 ( .C1(n9174), .C2(n8980), .A(n8979), .B(n8978), .ZN(n8981)
         );
  AOI21_X1 U10350 ( .B1(n9057), .B2(n9008), .A(n8981), .ZN(n8982) );
  INV_X1 U10351 ( .A(n8982), .ZN(P2_U3221) );
  OAI22_X1 U10352 ( .A1(n8991), .A2(n9066), .B1(n8983), .B2(n8989), .ZN(n8986)
         );
  MUX2_X1 U10353 ( .A(n8984), .B(P2_REG2_REG_10__SCAN_IN), .S(n8993), .Z(n8985) );
  AOI211_X1 U10354 ( .C1(n8997), .C2(n8987), .A(n8986), .B(n8985), .ZN(n8988)
         );
  INV_X1 U10355 ( .A(n8988), .ZN(P2_U3223) );
  OAI22_X1 U10356 ( .A1(n8992), .A2(n8991), .B1(n8990), .B2(n8989), .ZN(n8996)
         );
  MUX2_X1 U10357 ( .A(n8994), .B(P2_REG2_REG_9__SCAN_IN), .S(n8993), .Z(n8995)
         );
  AOI211_X1 U10358 ( .C1(n8998), .C2(n8997), .A(n8996), .B(n8995), .ZN(n8999)
         );
  INV_X1 U10359 ( .A(n8999), .ZN(P2_U3224) );
  INV_X1 U10360 ( .A(n9000), .ZN(n9005) );
  AOI22_X1 U10361 ( .A1(n9003), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n9002), .B2(
        n9001), .ZN(n9004) );
  OAI211_X1 U10362 ( .C1(n9007), .C2(n9006), .A(n9005), .B(n9004), .ZN(n9009)
         );
  MUX2_X1 U10363 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9009), .S(n9008), .Z(
        P2_U3231) );
  INV_X1 U10364 ( .A(n9075), .ZN(n9011) );
  NAND2_X1 U10365 ( .A1(n9073), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9010) );
  NAND2_X1 U10366 ( .A1(n9076), .A2(n4313), .ZN(n9013) );
  OAI211_X1 U10367 ( .C1(n9011), .C2(n9065), .A(n9010), .B(n9013), .ZN(
        P2_U3490) );
  NAND2_X1 U10368 ( .A1(n9073), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9012) );
  OAI211_X1 U10369 ( .C1(n9081), .C2(n9065), .A(n9013), .B(n9012), .ZN(
        P2_U3489) );
  INV_X1 U10370 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9014) );
  MUX2_X1 U10371 ( .A(n9082), .B(n9014), .S(n9073), .Z(n9016) );
  NAND2_X1 U10372 ( .A1(n9084), .A2(n9054), .ZN(n9015) );
  OAI211_X1 U10373 ( .C1(n9087), .C2(n9061), .A(n9016), .B(n9015), .ZN(
        P2_U3486) );
  INV_X1 U10374 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9017) );
  MUX2_X1 U10375 ( .A(n9088), .B(n9017), .S(n9073), .Z(n9019) );
  NAND2_X1 U10376 ( .A1(n9090), .A2(n9054), .ZN(n9018) );
  OAI211_X1 U10377 ( .C1(n9093), .C2(n9061), .A(n9019), .B(n9018), .ZN(
        P2_U3485) );
  MUX2_X1 U10378 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9094), .S(n4313), .Z(n9021) );
  OAI22_X1 U10379 ( .A1(n9097), .A2(n9061), .B1(n9096), .B2(n9065), .ZN(n9020)
         );
  OR2_X1 U10380 ( .A1(n9021), .A2(n9020), .ZN(P2_U3484) );
  INV_X1 U10381 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9022) );
  MUX2_X1 U10382 ( .A(n9022), .B(n9100), .S(n4313), .Z(n9024) );
  NAND2_X1 U10383 ( .A1(n9102), .A2(n9054), .ZN(n9023) );
  OAI211_X1 U10384 ( .C1(n9061), .C2(n9105), .A(n9024), .B(n9023), .ZN(
        P2_U3483) );
  INV_X1 U10385 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9025) );
  MUX2_X1 U10386 ( .A(n9025), .B(n9106), .S(n4313), .Z(n9027) );
  NAND2_X1 U10387 ( .A1(n9107), .A2(n9054), .ZN(n9026) );
  OAI211_X1 U10388 ( .C1(n9110), .C2(n9061), .A(n9027), .B(n9026), .ZN(
        P2_U3482) );
  INV_X1 U10389 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9028) );
  MUX2_X1 U10390 ( .A(n9028), .B(n9111), .S(n4313), .Z(n9030) );
  NAND2_X1 U10391 ( .A1(n9113), .A2(n9054), .ZN(n9029) );
  OAI211_X1 U10392 ( .C1(n9061), .C2(n9116), .A(n9030), .B(n9029), .ZN(
        P2_U3481) );
  INV_X1 U10393 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9031) );
  MUX2_X1 U10394 ( .A(n9031), .B(n9117), .S(n4313), .Z(n9033) );
  NAND2_X1 U10395 ( .A1(n9118), .A2(n9054), .ZN(n9032) );
  OAI211_X1 U10396 ( .C1(n9061), .C2(n9121), .A(n9033), .B(n9032), .ZN(
        P2_U3480) );
  INV_X1 U10397 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9034) );
  MUX2_X1 U10398 ( .A(n9034), .B(n9122), .S(n4313), .Z(n9036) );
  NAND2_X1 U10399 ( .A1(n9124), .A2(n9054), .ZN(n9035) );
  OAI211_X1 U10400 ( .C1(n9127), .C2(n9061), .A(n9036), .B(n9035), .ZN(
        P2_U3479) );
  MUX2_X1 U10401 ( .A(n9037), .B(n9128), .S(n4313), .Z(n9039) );
  NAND2_X1 U10402 ( .A1(n9130), .A2(n9054), .ZN(n9038) );
  OAI211_X1 U10403 ( .C1(n9133), .C2(n9061), .A(n9039), .B(n9038), .ZN(
        P2_U3478) );
  INV_X1 U10404 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9040) );
  MUX2_X1 U10405 ( .A(n9040), .B(n9134), .S(n4313), .Z(n9042) );
  NAND2_X1 U10406 ( .A1(n9136), .A2(n9054), .ZN(n9041) );
  OAI211_X1 U10407 ( .C1(n9061), .C2(n9139), .A(n9042), .B(n9041), .ZN(
        P2_U3477) );
  MUX2_X1 U10408 ( .A(n9043), .B(n9140), .S(n4313), .Z(n9045) );
  NAND2_X1 U10409 ( .A1(n9142), .A2(n9054), .ZN(n9044) );
  OAI211_X1 U10410 ( .C1(n9145), .C2(n9061), .A(n9045), .B(n9044), .ZN(
        P2_U3476) );
  INV_X1 U10411 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9046) );
  MUX2_X1 U10412 ( .A(n9046), .B(n9146), .S(n4313), .Z(n9048) );
  NAND2_X1 U10413 ( .A1(n9148), .A2(n9054), .ZN(n9047) );
  OAI211_X1 U10414 ( .C1(n9151), .C2(n9061), .A(n9048), .B(n9047), .ZN(
        P2_U3475) );
  MUX2_X1 U10415 ( .A(n9049), .B(n9152), .S(n4313), .Z(n9051) );
  NAND2_X1 U10416 ( .A1(n9154), .A2(n9054), .ZN(n9050) );
  OAI211_X1 U10417 ( .C1(n9061), .C2(n9157), .A(n9051), .B(n9050), .ZN(
        P2_U3474) );
  MUX2_X1 U10418 ( .A(n10262), .B(n9158), .S(n4313), .Z(n9053) );
  NAND2_X1 U10419 ( .A1(n9160), .A2(n9054), .ZN(n9052) );
  OAI211_X1 U10420 ( .C1(n9163), .C2(n9061), .A(n9053), .B(n9052), .ZN(
        P2_U3473) );
  MUX2_X1 U10421 ( .A(n10237), .B(n9164), .S(n4313), .Z(n9056) );
  NAND2_X1 U10422 ( .A1(n9166), .A2(n9054), .ZN(n9055) );
  OAI211_X1 U10423 ( .C1(n9061), .C2(n9170), .A(n9056), .B(n9055), .ZN(
        P2_U3472) );
  AOI21_X1 U10424 ( .B1(n9069), .B2(n9058), .A(n9057), .ZN(n9171) );
  MUX2_X1 U10425 ( .A(n9059), .B(n9171), .S(n4313), .Z(n9060) );
  OAI21_X1 U10426 ( .B1(n9061), .B2(n9174), .A(n9060), .ZN(P2_U3471) );
  MUX2_X1 U10427 ( .A(n9063), .B(n9062), .S(n4313), .Z(n9064) );
  OAI21_X1 U10428 ( .B1(n9066), .B2(n9065), .A(n9064), .ZN(P2_U3469) );
  AOI21_X1 U10429 ( .B1(n9069), .B2(n9068), .A(n9067), .ZN(n9070) );
  OAI21_X1 U10430 ( .B1(n9072), .B2(n9071), .A(n9070), .ZN(n10291) );
  MUX2_X1 U10431 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10291), .S(n4313), .Z(
        P2_U3465) );
  MUX2_X1 U10432 ( .A(n9074), .B(P2_REG1_REG_0__SCAN_IN), .S(n9073), .Z(
        P2_U3459) );
  NAND2_X1 U10433 ( .A1(n9075), .A2(n9167), .ZN(n9077) );
  NAND2_X1 U10434 ( .A1(n9076), .A2(n5734), .ZN(n9080) );
  OAI211_X1 U10435 ( .C1(n9078), .C2(n5734), .A(n9077), .B(n9080), .ZN(
        P2_U3458) );
  NAND2_X1 U10436 ( .A1(n10292), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9079) );
  OAI211_X1 U10437 ( .C1(n9081), .C2(n9095), .A(n9080), .B(n9079), .ZN(
        P2_U3457) );
  INV_X1 U10438 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9083) );
  MUX2_X1 U10439 ( .A(n9083), .B(n9082), .S(n5734), .Z(n9086) );
  NAND2_X1 U10440 ( .A1(n9084), .A2(n9167), .ZN(n9085) );
  OAI211_X1 U10441 ( .C1(n9087), .C2(n9173), .A(n9086), .B(n9085), .ZN(
        P2_U3454) );
  INV_X1 U10442 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9089) );
  MUX2_X1 U10443 ( .A(n9089), .B(n9088), .S(n5734), .Z(n9092) );
  NAND2_X1 U10444 ( .A1(n9090), .A2(n9167), .ZN(n9091) );
  OAI211_X1 U10445 ( .C1(n9093), .C2(n9173), .A(n9092), .B(n9091), .ZN(
        P2_U3453) );
  MUX2_X1 U10446 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9094), .S(n5734), .Z(n9099) );
  OAI22_X1 U10447 ( .A1(n9097), .A2(n9173), .B1(n9096), .B2(n9095), .ZN(n9098)
         );
  OR2_X1 U10448 ( .A1(n9099), .A2(n9098), .ZN(P2_U3452) );
  INV_X1 U10449 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9101) );
  MUX2_X1 U10450 ( .A(n9101), .B(n9100), .S(n5734), .Z(n9104) );
  NAND2_X1 U10451 ( .A1(n9102), .A2(n9167), .ZN(n9103) );
  OAI211_X1 U10452 ( .C1(n9105), .C2(n9173), .A(n9104), .B(n9103), .ZN(
        P2_U3451) );
  MUX2_X1 U10453 ( .A(n10206), .B(n9106), .S(n5734), .Z(n9109) );
  NAND2_X1 U10454 ( .A1(n9107), .A2(n9167), .ZN(n9108) );
  OAI211_X1 U10455 ( .C1(n9110), .C2(n9173), .A(n9109), .B(n9108), .ZN(
        P2_U3450) );
  INV_X1 U10456 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9112) );
  MUX2_X1 U10457 ( .A(n9112), .B(n9111), .S(n5734), .Z(n9115) );
  NAND2_X1 U10458 ( .A1(n9113), .A2(n9167), .ZN(n9114) );
  OAI211_X1 U10459 ( .C1(n9116), .C2(n9173), .A(n9115), .B(n9114), .ZN(
        P2_U3449) );
  MUX2_X1 U10460 ( .A(n10218), .B(n9117), .S(n5734), .Z(n9120) );
  NAND2_X1 U10461 ( .A1(n9118), .A2(n9167), .ZN(n9119) );
  OAI211_X1 U10462 ( .C1(n9121), .C2(n9173), .A(n9120), .B(n9119), .ZN(
        P2_U3448) );
  INV_X1 U10463 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9123) );
  MUX2_X1 U10464 ( .A(n9123), .B(n9122), .S(n5734), .Z(n9126) );
  NAND2_X1 U10465 ( .A1(n9124), .A2(n9167), .ZN(n9125) );
  OAI211_X1 U10466 ( .C1(n9127), .C2(n9173), .A(n9126), .B(n9125), .ZN(
        P2_U3447) );
  INV_X1 U10467 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9129) );
  MUX2_X1 U10468 ( .A(n9129), .B(n9128), .S(n5734), .Z(n9132) );
  NAND2_X1 U10469 ( .A1(n9130), .A2(n9167), .ZN(n9131) );
  OAI211_X1 U10470 ( .C1(n9133), .C2(n9173), .A(n9132), .B(n9131), .ZN(
        P2_U3446) );
  INV_X1 U10471 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9135) );
  MUX2_X1 U10472 ( .A(n9135), .B(n9134), .S(n5734), .Z(n9138) );
  NAND2_X1 U10473 ( .A1(n9136), .A2(n9167), .ZN(n9137) );
  OAI211_X1 U10474 ( .C1(n9139), .C2(n9173), .A(n9138), .B(n9137), .ZN(
        P2_U3444) );
  INV_X1 U10475 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9141) );
  MUX2_X1 U10476 ( .A(n9141), .B(n9140), .S(n5734), .Z(n9144) );
  NAND2_X1 U10477 ( .A1(n9142), .A2(n9167), .ZN(n9143) );
  OAI211_X1 U10478 ( .C1(n9145), .C2(n9173), .A(n9144), .B(n9143), .ZN(
        P2_U3441) );
  INV_X1 U10479 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9147) );
  MUX2_X1 U10480 ( .A(n9147), .B(n9146), .S(n5734), .Z(n9150) );
  NAND2_X1 U10481 ( .A1(n9148), .A2(n9167), .ZN(n9149) );
  OAI211_X1 U10482 ( .C1(n9151), .C2(n9173), .A(n9150), .B(n9149), .ZN(
        P2_U3438) );
  INV_X1 U10483 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9153) );
  MUX2_X1 U10484 ( .A(n9153), .B(n9152), .S(n5734), .Z(n9156) );
  NAND2_X1 U10485 ( .A1(n9154), .A2(n9167), .ZN(n9155) );
  OAI211_X1 U10486 ( .C1(n9157), .C2(n9173), .A(n9156), .B(n9155), .ZN(
        P2_U3435) );
  MUX2_X1 U10487 ( .A(n9159), .B(n9158), .S(n5734), .Z(n9162) );
  NAND2_X1 U10488 ( .A1(n9160), .A2(n9167), .ZN(n9161) );
  OAI211_X1 U10489 ( .C1(n9163), .C2(n9173), .A(n9162), .B(n9161), .ZN(
        P2_U3432) );
  MUX2_X1 U10490 ( .A(n9165), .B(n9164), .S(n5734), .Z(n9169) );
  NAND2_X1 U10491 ( .A1(n9167), .A2(n9166), .ZN(n9168) );
  OAI211_X1 U10492 ( .C1(n9170), .C2(n9173), .A(n9169), .B(n9168), .ZN(
        P2_U3429) );
  MUX2_X1 U10493 ( .A(n10170), .B(n9171), .S(n5734), .Z(n9172) );
  OAI21_X1 U10494 ( .B1(n9174), .B2(n9173), .A(n9172), .ZN(P2_U3426) );
  NAND3_X1 U10495 ( .A1(n9176), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9178) );
  OAI22_X1 U10496 ( .A1(n9175), .A2(n9178), .B1(n9177), .B2(n8387), .ZN(n9179)
         );
  AOI21_X1 U10497 ( .B1(n9860), .B2(n9180), .A(n9179), .ZN(n9181) );
  INV_X1 U10498 ( .A(n9181), .ZN(P2_U3264) );
  AOI21_X1 U10499 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9183), .A(n9182), .ZN(
        n9184) );
  OAI21_X1 U10500 ( .B1(n9185), .B2(n7852), .A(n9184), .ZN(P2_U3267) );
  INV_X1 U10501 ( .A(n9186), .ZN(n9187) );
  MUX2_X1 U10502 ( .A(n9187), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10503 ( .A(n9189), .ZN(n9190) );
  AOI21_X1 U10504 ( .B1(n9192), .B2(n9191), .A(n9190), .ZN(n9197) );
  AOI22_X1 U10505 ( .A1(n9193), .A2(n9372), .B1(n9371), .B2(n9394), .ZN(n9194)
         );
  NAND2_X1 U10506 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9928) );
  OAI211_X1 U10507 ( .C1(n9258), .C2(n9375), .A(n9194), .B(n9928), .ZN(n9195)
         );
  AOI21_X1 U10508 ( .B1(n9815), .B2(n9378), .A(n9195), .ZN(n9196) );
  OAI21_X1 U10509 ( .B1(n9197), .B2(n9380), .A(n9196), .ZN(P1_U3215) );
  INV_X1 U10510 ( .A(n9198), .ZN(n9199) );
  NAND2_X1 U10511 ( .A1(n9200), .A2(n9199), .ZN(n9323) );
  NAND2_X1 U10512 ( .A1(n9323), .A2(n9322), .ZN(n9321) );
  OR2_X1 U10513 ( .A1(n9200), .A2(n9199), .ZN(n9325) );
  NAND2_X1 U10514 ( .A1(n9201), .A2(n9275), .ZN(n9202) );
  AND3_X1 U10515 ( .A1(n9321), .A2(n9325), .A3(n9202), .ZN(n9203) );
  OAI21_X1 U10516 ( .B1(n9278), .B2(n9203), .A(n9312), .ZN(n9208) );
  OAI22_X1 U10517 ( .A1(n9637), .A2(n9375), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9204), .ZN(n9206) );
  OAI22_X1 U10518 ( .A1(n9636), .A2(n9359), .B1(n9349), .B2(n9627), .ZN(n9205)
         );
  AOI211_X1 U10519 ( .C1(n9769), .C2(n9378), .A(n9206), .B(n9205), .ZN(n9207)
         );
  NAND2_X1 U10520 ( .A1(n9208), .A2(n9207), .ZN(P1_U3216) );
  XNOR2_X1 U10521 ( .A(n9209), .B(n9210), .ZN(n9347) );
  NOR2_X1 U10522 ( .A1(n9347), .A2(n9346), .ZN(n9345) );
  AOI21_X1 U10523 ( .B1(n9210), .B2(n9209), .A(n9345), .ZN(n9214) );
  XNOR2_X1 U10524 ( .A(n9212), .B(n9211), .ZN(n9213) );
  XNOR2_X1 U10525 ( .A(n9214), .B(n9213), .ZN(n9215) );
  NAND2_X1 U10526 ( .A1(n9215), .A2(n9312), .ZN(n9218) );
  AND2_X1 U10527 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9551) );
  OAI22_X1 U10528 ( .A1(n9359), .A2(n9700), .B1(n9349), .B2(n9695), .ZN(n9216)
         );
  AOI211_X1 U10529 ( .C1(n9317), .C2(n9221), .A(n9551), .B(n9216), .ZN(n9217)
         );
  OAI211_X1 U10530 ( .C1(n9694), .C2(n9366), .A(n9218), .B(n9217), .ZN(
        P1_U3219) );
  XOR2_X1 U10531 ( .A(n9220), .B(n9219), .Z(n9227) );
  NAND2_X1 U10532 ( .A1(n9388), .A2(n9675), .ZN(n9223) );
  NAND2_X1 U10533 ( .A1(n9221), .A2(n9673), .ZN(n9222) );
  NAND2_X1 U10534 ( .A1(n9223), .A2(n9222), .ZN(n9659) );
  AOI22_X1 U10535 ( .A1(n9659), .A2(n9269), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9224) );
  OAI21_X1 U10536 ( .B1(n9349), .B2(n9664), .A(n9224), .ZN(n9225) );
  AOI21_X1 U10537 ( .B1(n9778), .B2(n9378), .A(n9225), .ZN(n9226) );
  OAI21_X1 U10538 ( .B1(n9227), .B2(n9380), .A(n9226), .ZN(P1_U3223) );
  AOI22_X1 U10539 ( .A1(n9228), .A2(n9372), .B1(n9371), .B2(n9396), .ZN(n9230)
         );
  OAI211_X1 U10540 ( .C1(n9231), .C2(n9375), .A(n9230), .B(n9229), .ZN(n9237)
         );
  NAND3_X1 U10541 ( .A1(n9232), .A2(n9233), .A3(n4335), .ZN(n9234) );
  AOI21_X1 U10542 ( .B1(n9235), .B2(n9234), .A(n9380), .ZN(n9236) );
  AOI211_X1 U10543 ( .C1(n9826), .C2(n9378), .A(n9237), .B(n9236), .ZN(n9238)
         );
  INV_X1 U10544 ( .A(n9238), .ZN(P1_U3224) );
  OAI21_X1 U10545 ( .B1(n9240), .B2(n9239), .A(n9357), .ZN(n9241) );
  NAND2_X1 U10546 ( .A1(n9241), .A2(n9312), .ZN(n9247) );
  AND2_X1 U10547 ( .A1(n9386), .A2(n9673), .ZN(n9242) );
  AOI21_X1 U10548 ( .B1(n9384), .B2(n9675), .A(n9242), .ZN(n9602) );
  INV_X1 U10549 ( .A(n9602), .ZN(n9245) );
  OAI22_X1 U10550 ( .A1(n9595), .A2(n9349), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9243), .ZN(n9244) );
  AOI21_X1 U10551 ( .B1(n9245), .B2(n9269), .A(n9244), .ZN(n9246) );
  OAI211_X1 U10552 ( .C1(n4760), .C2(n9366), .A(n9247), .B(n9246), .ZN(
        P1_U3225) );
  INV_X1 U10553 ( .A(n9803), .ZN(n9262) );
  NAND2_X1 U10554 ( .A1(n9249), .A2(n9250), .ZN(n9251) );
  OAI21_X1 U10555 ( .B1(n9249), .B2(n9250), .A(n9251), .ZN(n9369) );
  NOR2_X1 U10556 ( .A1(n9369), .A2(n9370), .ZN(n9368) );
  INV_X1 U10557 ( .A(n9251), .ZN(n9252) );
  NOR3_X1 U10558 ( .A1(n9368), .A2(n9253), .A3(n9252), .ZN(n9256) );
  INV_X1 U10559 ( .A(n9254), .ZN(n9255) );
  OAI21_X1 U10560 ( .B1(n9256), .B2(n9255), .A(n9312), .ZN(n9261) );
  AND2_X1 U10561 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9512) );
  OAI22_X1 U10562 ( .A1(n9359), .A2(n9258), .B1(n9349), .B2(n9257), .ZN(n9259)
         );
  AOI211_X1 U10563 ( .C1(n9317), .C2(n9390), .A(n9512), .B(n9259), .ZN(n9260)
         );
  OAI211_X1 U10564 ( .C1(n9262), .C2(n9366), .A(n9261), .B(n9260), .ZN(
        P1_U3226) );
  NAND2_X1 U10565 ( .A1(n9264), .A2(n9263), .ZN(n9265) );
  XNOR2_X1 U10566 ( .A(n9266), .B(n9265), .ZN(n9274) );
  INV_X1 U10567 ( .A(n9726), .ZN(n9271) );
  NAND2_X1 U10568 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9527) );
  OR2_X1 U10569 ( .A1(n9376), .A2(n9710), .ZN(n9268) );
  NAND2_X1 U10570 ( .A1(n9389), .A2(n9675), .ZN(n9267) );
  NAND2_X1 U10571 ( .A1(n9268), .A2(n9267), .ZN(n9731) );
  NAND2_X1 U10572 ( .A1(n9269), .A2(n9731), .ZN(n9270) );
  OAI211_X1 U10573 ( .C1(n9349), .C2(n9271), .A(n9527), .B(n9270), .ZN(n9272)
         );
  AOI21_X1 U10574 ( .B1(n9798), .B2(n9378), .A(n9272), .ZN(n9273) );
  OAI21_X1 U10575 ( .B1(n9274), .B2(n9380), .A(n9273), .ZN(P1_U3228) );
  INV_X1 U10576 ( .A(n9275), .ZN(n9277) );
  NOR3_X1 U10577 ( .A1(n9278), .A2(n9277), .A3(n9276), .ZN(n9281) );
  INV_X1 U10578 ( .A(n9279), .ZN(n9280) );
  OAI21_X1 U10579 ( .B1(n9281), .B2(n9280), .A(n9312), .ZN(n9285) );
  AOI22_X1 U10580 ( .A1(n9385), .A2(n9317), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9284) );
  AOI22_X1 U10581 ( .A1(n9616), .A2(n9372), .B1(n9387), .B2(n9371), .ZN(n9283)
         );
  NAND2_X1 U10582 ( .A1(n9764), .A2(n9378), .ZN(n9282) );
  NAND4_X1 U10583 ( .A1(n9285), .A2(n9284), .A3(n9283), .A4(n9282), .ZN(
        P1_U3229) );
  AOI22_X1 U10584 ( .A1(n9286), .A2(n9372), .B1(n9371), .B2(n9399), .ZN(n9288)
         );
  OAI211_X1 U10585 ( .C1(n9289), .C2(n9375), .A(n9288), .B(n9287), .ZN(n9298)
         );
  INV_X1 U10586 ( .A(n9290), .ZN(n9291) );
  NAND3_X1 U10587 ( .A1(n9293), .A2(n9292), .A3(n9291), .ZN(n9296) );
  AOI21_X1 U10588 ( .B1(n9296), .B2(n9295), .A(n9380), .ZN(n9297) );
  AOI211_X1 U10589 ( .C1(n10046), .C2(n9378), .A(n9298), .B(n9297), .ZN(n9300)
         );
  INV_X1 U10590 ( .A(n9300), .ZN(P1_U3231) );
  XNOR2_X1 U10591 ( .A(n9302), .B(n9301), .ZN(n9303) );
  XNOR2_X1 U10592 ( .A(n9304), .B(n9303), .ZN(n9308) );
  OAI22_X1 U10593 ( .A1(n9375), .A2(n9648), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10160), .ZN(n9306) );
  OAI22_X1 U10594 ( .A1(n9359), .A2(n9711), .B1(n9349), .B2(n9680), .ZN(n9305)
         );
  AOI211_X1 U10595 ( .C1(n9782), .C2(n9378), .A(n9306), .B(n9305), .ZN(n9307)
         );
  OAI21_X1 U10596 ( .B1(n9308), .B2(n9380), .A(n9307), .ZN(P1_U3233) );
  OAI21_X1 U10597 ( .B1(n9311), .B2(n9310), .A(n9309), .ZN(n9313) );
  NAND2_X1 U10598 ( .A1(n9313), .A2(n9312), .ZN(n9319) );
  AND2_X1 U10599 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9486) );
  INV_X1 U10600 ( .A(n9314), .ZN(n9315) );
  OAI22_X1 U10601 ( .A1(n9359), .A2(n9336), .B1(n9349), .B2(n9315), .ZN(n9316)
         );
  AOI211_X1 U10602 ( .C1(n9317), .C2(n9393), .A(n9486), .B(n9316), .ZN(n9318)
         );
  OAI211_X1 U10603 ( .C1(n9320), .C2(n9366), .A(n9319), .B(n9318), .ZN(
        P1_U3234) );
  INV_X1 U10604 ( .A(n9321), .ZN(n9326) );
  AOI21_X1 U10605 ( .B1(n9325), .B2(n9323), .A(n9322), .ZN(n9324) );
  AOI21_X1 U10606 ( .B1(n9326), .B2(n9325), .A(n9324), .ZN(n9332) );
  OAI22_X1 U10607 ( .A1(n9649), .A2(n9375), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9327), .ZN(n9330) );
  INV_X1 U10608 ( .A(n9643), .ZN(n9328) );
  OAI22_X1 U10609 ( .A1(n9359), .A2(n9648), .B1(n9349), .B2(n9328), .ZN(n9329)
         );
  AOI211_X1 U10610 ( .C1(n9773), .C2(n9378), .A(n9330), .B(n9329), .ZN(n9331)
         );
  OAI21_X1 U10611 ( .B1(n9332), .B2(n9380), .A(n9331), .ZN(P1_U3235) );
  AOI22_X1 U10612 ( .A1(n9333), .A2(n9372), .B1(n9371), .B2(n9397), .ZN(n9335)
         );
  OAI211_X1 U10613 ( .C1(n9336), .C2(n9375), .A(n9335), .B(n9334), .ZN(n9343)
         );
  INV_X1 U10614 ( .A(n9337), .ZN(n9338) );
  NAND3_X1 U10615 ( .A1(n9340), .A2(n9339), .A3(n9338), .ZN(n9341) );
  AOI21_X1 U10616 ( .B1(n9341), .B2(n9232), .A(n9380), .ZN(n9342) );
  AOI211_X1 U10617 ( .C1(n6597), .C2(n9378), .A(n9343), .B(n9342), .ZN(n9344)
         );
  INV_X1 U10618 ( .A(n9344), .ZN(P1_U3236) );
  AOI21_X1 U10619 ( .B1(n9347), .B2(n9346), .A(n9345), .ZN(n9353) );
  OAI22_X1 U10620 ( .A1(n9375), .A2(n9711), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9348), .ZN(n9351) );
  OAI22_X1 U10621 ( .A1(n9359), .A2(n9709), .B1(n9349), .B2(n9715), .ZN(n9350)
         );
  AOI211_X1 U10622 ( .C1(n9794), .C2(n9378), .A(n9351), .B(n9350), .ZN(n9352)
         );
  OAI21_X1 U10623 ( .B1(n9353), .B2(n9380), .A(n9352), .ZN(P1_U3238) );
  OAI22_X1 U10624 ( .A1(n9612), .A2(n9359), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9358), .ZN(n9362) );
  NOR2_X1 U10625 ( .A1(n9360), .A2(n9375), .ZN(n9361) );
  AOI211_X1 U10626 ( .C1(n9363), .C2(n9372), .A(n9362), .B(n9361), .ZN(n9364)
         );
  OAI211_X1 U10627 ( .C1(n9367), .C2(n9366), .A(n9365), .B(n9364), .ZN(
        P1_U3240) );
  AOI21_X1 U10628 ( .B1(n9370), .B2(n9369), .A(n9368), .ZN(n9381) );
  AOI22_X1 U10629 ( .A1(n9373), .A2(n9372), .B1(n9371), .B2(n9393), .ZN(n9374)
         );
  NAND2_X1 U10630 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9941) );
  OAI211_X1 U10631 ( .C1(n9376), .C2(n9375), .A(n9374), .B(n9941), .ZN(n9377)
         );
  AOI21_X1 U10632 ( .B1(n9811), .B2(n9378), .A(n9377), .ZN(n9379) );
  OAI21_X1 U10633 ( .B1(n9381), .B2(n9380), .A(n9379), .ZN(P1_U3241) );
  MUX2_X1 U10634 ( .A(n9382), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9403), .Z(
        P1_U3584) );
  MUX2_X1 U10635 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9585), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10636 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9383), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10637 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9586), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10638 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9384), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10639 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9385), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10640 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9386), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10641 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9387), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10642 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9388), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10643 ( .A(n9676), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9403), .Z(
        P1_U3575) );
  MUX2_X1 U10644 ( .A(n9674), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9403), .Z(
        P1_U3573) );
  MUX2_X1 U10645 ( .A(n9389), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9403), .Z(
        P1_U3572) );
  MUX2_X1 U10646 ( .A(n9390), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9403), .Z(
        P1_U3571) );
  MUX2_X1 U10647 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9391), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10648 ( .A(n9392), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9403), .Z(
        P1_U3569) );
  MUX2_X1 U10649 ( .A(n9393), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9403), .Z(
        P1_U3568) );
  MUX2_X1 U10650 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9394), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10651 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9395), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10652 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9396), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10653 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9397), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10654 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9398), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10655 ( .A(n9399), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9403), .Z(
        P1_U3562) );
  MUX2_X1 U10656 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9400), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10657 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9401), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10658 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n6400), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10659 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9402), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10660 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n6380), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10661 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n7130), .S(P1_U3973), .Z(
        P1_U3556) );
  NAND2_X1 U10662 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9406) );
  AOI211_X1 U10663 ( .C1(n9406), .C2(n9405), .A(n9404), .B(n9944), .ZN(n9407)
         );
  INV_X1 U10664 ( .A(n9407), .ZN(n9416) );
  INV_X1 U10665 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9408) );
  OAI22_X1 U10666 ( .A1(n9960), .A2(n9408), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9988), .ZN(n9409) );
  AOI21_X1 U10667 ( .B1(n9410), .B2(n9947), .A(n9409), .ZN(n9415) );
  OAI211_X1 U10668 ( .C1(n9413), .C2(n9412), .A(n9951), .B(n9411), .ZN(n9414)
         );
  NAND3_X1 U10669 ( .A1(n9416), .A2(n9415), .A3(n9414), .ZN(P1_U3244) );
  AOI211_X1 U10670 ( .C1(n9419), .C2(n9418), .A(n9417), .B(n9944), .ZN(n9420)
         );
  INV_X1 U10671 ( .A(n9420), .ZN(n9429) );
  INV_X1 U10672 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9870) );
  OAI21_X1 U10673 ( .B1(n9960), .B2(n9870), .A(n9421), .ZN(n9422) );
  AOI21_X1 U10674 ( .B1(n9423), .B2(n9947), .A(n9422), .ZN(n9428) );
  OAI211_X1 U10675 ( .C1(n9426), .C2(n9425), .A(n9951), .B(n9424), .ZN(n9427)
         );
  NAND3_X1 U10676 ( .A1(n9429), .A2(n9428), .A3(n9427), .ZN(P1_U3246) );
  AOI211_X1 U10677 ( .C1(n9432), .C2(n9431), .A(n9944), .B(n9430), .ZN(n9433)
         );
  INV_X1 U10678 ( .A(n9433), .ZN(n9441) );
  INV_X1 U10679 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U10680 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9434) );
  OAI21_X1 U10681 ( .B1(n9960), .B2(n9881), .A(n9434), .ZN(n9435) );
  AOI21_X1 U10682 ( .B1(n6014), .B2(n9947), .A(n9435), .ZN(n9440) );
  OAI211_X1 U10683 ( .C1(n9438), .C2(n9437), .A(n9951), .B(n9436), .ZN(n9439)
         );
  NAND3_X1 U10684 ( .A1(n9441), .A2(n9440), .A3(n9439), .ZN(P1_U3248) );
  AOI211_X1 U10685 ( .C1(n9443), .C2(n9442), .A(n9944), .B(n4427), .ZN(n9444)
         );
  INV_X1 U10686 ( .A(n9444), .ZN(n9454) );
  INV_X1 U10687 ( .A(n9445), .ZN(n9446) );
  OAI21_X1 U10688 ( .B1(n9960), .B2(n9884), .A(n9446), .ZN(n9447) );
  AOI21_X1 U10689 ( .B1(n9448), .B2(n9947), .A(n9447), .ZN(n9453) );
  OAI211_X1 U10690 ( .C1(n9451), .C2(n9450), .A(n9951), .B(n9449), .ZN(n9452)
         );
  NAND3_X1 U10691 ( .A1(n9454), .A2(n9453), .A3(n9452), .ZN(P1_U3249) );
  AOI211_X1 U10692 ( .C1(n9457), .C2(n9456), .A(n9944), .B(n9455), .ZN(n9458)
         );
  INV_X1 U10693 ( .A(n9458), .ZN(n9467) );
  INV_X1 U10694 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U10695 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9459) );
  OAI21_X1 U10696 ( .B1(n9960), .B2(n9887), .A(n9459), .ZN(n9460) );
  AOI21_X1 U10697 ( .B1(n9461), .B2(n9947), .A(n9460), .ZN(n9466) );
  OAI211_X1 U10698 ( .C1(n9464), .C2(n9463), .A(n9951), .B(n9462), .ZN(n9465)
         );
  NAND3_X1 U10699 ( .A1(n9467), .A2(n9466), .A3(n9465), .ZN(P1_U3250) );
  AOI211_X1 U10700 ( .C1(n9470), .C2(n9469), .A(n9944), .B(n9468), .ZN(n9471)
         );
  INV_X1 U10701 ( .A(n9471), .ZN(n9480) );
  INV_X1 U10702 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9890) );
  OAI21_X1 U10703 ( .B1(n9960), .B2(n9890), .A(n9472), .ZN(n9473) );
  AOI21_X1 U10704 ( .B1(n9474), .B2(n9947), .A(n9473), .ZN(n9479) );
  OAI211_X1 U10705 ( .C1(n9477), .C2(n9476), .A(n9951), .B(n9475), .ZN(n9478)
         );
  NAND3_X1 U10706 ( .A1(n9480), .A2(n9479), .A3(n9478), .ZN(P1_U3251) );
  INV_X1 U10707 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9483) );
  MUX2_X1 U10708 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n9483), .S(n9501), .Z(n9484) );
  OAI21_X1 U10709 ( .B1(n9485), .B2(n9484), .A(n9951), .ZN(n9495) );
  INV_X1 U10710 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9904) );
  INV_X1 U10711 ( .A(n9486), .ZN(n9487) );
  OAI21_X1 U10712 ( .B1(n9960), .B2(n9904), .A(n9487), .ZN(n9493) );
  XNOR2_X1 U10713 ( .A(n9501), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9491) );
  OAI21_X1 U10714 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9489), .A(n9488), .ZN(
        n9490) );
  AOI211_X1 U10715 ( .C1(n9491), .C2(n9490), .A(n9944), .B(n9497), .ZN(n9492)
         );
  AOI211_X1 U10716 ( .C1(n9947), .C2(n9501), .A(n9493), .B(n9492), .ZN(n9494)
         );
  OAI21_X1 U10717 ( .B1(n9500), .B2(n9495), .A(n9494), .ZN(P1_U3256) );
  INV_X1 U10718 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9496) );
  XNOR2_X1 U10719 ( .A(n9522), .B(n9496), .ZN(n9517) );
  INV_X1 U10720 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9932) );
  AOI21_X1 U10721 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n9501), .A(n9497), .ZN(
        n9924) );
  XNOR2_X1 U10722 ( .A(n9927), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9923) );
  AND2_X1 U10723 ( .A1(n9927), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9498) );
  XOR2_X1 U10724 ( .A(n9517), .B(n9518), .Z(n9515) );
  INV_X1 U10725 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9502) );
  MUX2_X1 U10726 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n9502), .S(n9927), .Z(n9503) );
  INV_X1 U10727 ( .A(n9503), .ZN(n9920) );
  NOR2_X1 U10728 ( .A1(n9921), .A2(n9920), .ZN(n9919) );
  AOI21_X1 U10729 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9927), .A(n9919), .ZN(
        n9504) );
  NOR2_X1 U10730 ( .A1(n9504), .A2(n9505), .ZN(n9506) );
  INV_X1 U10731 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9936) );
  XNOR2_X1 U10732 ( .A(n9505), .B(n9504), .ZN(n9937) );
  MUX2_X1 U10733 ( .A(n9507), .B(P1_REG2_REG_16__SCAN_IN), .S(n9522), .Z(n9509) );
  INV_X1 U10734 ( .A(n9524), .ZN(n9508) );
  AOI211_X1 U10735 ( .C1(n9510), .C2(n9509), .A(n9508), .B(n9934), .ZN(n9511)
         );
  AOI211_X1 U10736 ( .C1(n9552), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9512), .B(
        n9511), .ZN(n9514) );
  NAND2_X1 U10737 ( .A1(n9947), .A2(n9522), .ZN(n9513) );
  OAI211_X1 U10738 ( .C1(n9515), .C2(n9944), .A(n9514), .B(n9513), .ZN(
        P1_U3259) );
  INV_X1 U10739 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9516) );
  XNOR2_X1 U10740 ( .A(n9540), .B(n9516), .ZN(n9538) );
  OR2_X1 U10741 ( .A1(n9522), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9519) );
  NAND2_X1 U10742 ( .A1(n9520), .A2(n9519), .ZN(n9539) );
  XOR2_X1 U10743 ( .A(n9538), .B(n9539), .Z(n9533) );
  INV_X1 U10744 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9521) );
  XNOR2_X1 U10745 ( .A(n9540), .B(n9521), .ZN(n9526) );
  NAND2_X1 U10746 ( .A1(n9522), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9523) );
  NAND2_X1 U10747 ( .A1(n9525), .A2(n9526), .ZN(n9535) );
  OAI21_X1 U10748 ( .B1(n9526), .B2(n9525), .A(n9535), .ZN(n9531) );
  INV_X1 U10749 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U10750 ( .A1(n9947), .A2(n9540), .ZN(n9528) );
  OAI211_X1 U10751 ( .C1(n9960), .C2(n9529), .A(n9528), .B(n9527), .ZN(n9530)
         );
  AOI21_X1 U10752 ( .B1(n9531), .B2(n9951), .A(n9530), .ZN(n9532) );
  OAI21_X1 U10753 ( .B1(n9533), .B2(n9944), .A(n9532), .ZN(P1_U3260) );
  OR2_X1 U10754 ( .A1(n9540), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9534) );
  AND2_X1 U10755 ( .A1(n9535), .A2(n9534), .ZN(n9954) );
  OR2_X1 U10756 ( .A1(n9948), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U10757 ( .A1(n9948), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9537) );
  AND2_X1 U10758 ( .A1(n9536), .A2(n9537), .ZN(n9953) );
  OR2_X1 U10759 ( .A1(n9540), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U10760 ( .A1(n9948), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9543) );
  OR2_X1 U10761 ( .A1(n9948), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U10762 ( .A1(n9543), .A2(n9542), .ZN(n9945) );
  XNOR2_X1 U10763 ( .A(n9544), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9548) );
  NOR2_X1 U10764 ( .A1(n10001), .A2(n9738), .ZN(n9559) );
  NOR2_X1 U10765 ( .A1(n8234), .A2(n9994), .ZN(n9553) );
  AOI211_X1 U10766 ( .C1(n10001), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9559), .B(
        n9553), .ZN(n9554) );
  OAI21_X1 U10767 ( .B1(n9555), .B2(n9982), .A(n9554), .ZN(P1_U3263) );
  OAI211_X1 U10768 ( .C1(n9740), .C2(n9557), .A(n10012), .B(n9556), .ZN(n9739)
         );
  NOR2_X1 U10769 ( .A1(n9740), .A2(n9994), .ZN(n9558) );
  AOI211_X1 U10770 ( .C1(n10001), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9559), .B(
        n9558), .ZN(n9560) );
  OAI21_X1 U10771 ( .B1(n9982), .B2(n9739), .A(n9560), .ZN(P1_U3264) );
  NAND2_X1 U10772 ( .A1(n9562), .A2(n9561), .ZN(n9563) );
  XNOR2_X1 U10773 ( .A(n9564), .B(n9563), .ZN(n9574) );
  NOR2_X1 U10774 ( .A1(n9565), .A2(n9982), .ZN(n9571) );
  NAND3_X1 U10775 ( .A1(n9566), .A2(P1_REG3_REG_28__SCAN_IN), .A3(n9965), .ZN(
        n9568) );
  NAND2_X1 U10776 ( .A1(n10001), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9567) );
  OAI211_X1 U10777 ( .C1(n9569), .C2(n9994), .A(n9568), .B(n9567), .ZN(n9570)
         );
  AOI211_X1 U10778 ( .C1(n9572), .C2(n9989), .A(n9571), .B(n9570), .ZN(n9573)
         );
  OAI21_X1 U10779 ( .B1(n9574), .B2(n9736), .A(n9573), .ZN(P1_U3356) );
  XNOR2_X1 U10780 ( .A(n9575), .B(n4918), .ZN(n9746) );
  AOI211_X1 U10781 ( .C1(n9742), .C2(n9577), .A(n9724), .B(n9576), .ZN(n9741)
         );
  INV_X1 U10782 ( .A(n9742), .ZN(n9580) );
  AOI22_X1 U10783 ( .A1(n9578), .A2(n9965), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n10001), .ZN(n9579) );
  OAI21_X1 U10784 ( .B1(n9580), .B2(n9994), .A(n9579), .ZN(n9590) );
  OAI21_X1 U10785 ( .B1(n9583), .B2(n9582), .A(n9581), .ZN(n9584) );
  AND2_X2 U10786 ( .A1(n9588), .A2(n9587), .ZN(n9744) );
  NOR2_X1 U10787 ( .A1(n9744), .A2(n10001), .ZN(n9589) );
  OAI21_X1 U10788 ( .B1(n9746), .B2(n9736), .A(n9591), .ZN(P1_U3265) );
  XNOR2_X1 U10789 ( .A(n9592), .B(n6522), .ZN(n9761) );
  AOI211_X1 U10790 ( .C1(n9759), .C2(n9614), .A(n9724), .B(n9593), .ZN(n9758)
         );
  NOR2_X1 U10791 ( .A1(n4760), .A2(n9994), .ZN(n9597) );
  OAI22_X1 U10792 ( .A1(n9595), .A2(n9987), .B1(n9594), .B2(n9989), .ZN(n9596)
         );
  AOI211_X1 U10793 ( .C1(n9758), .C2(n9991), .A(n9597), .B(n9596), .ZN(n9605)
         );
  INV_X1 U10794 ( .A(n9598), .ZN(n9599) );
  AOI21_X1 U10795 ( .B1(n9601), .B2(n9600), .A(n9599), .ZN(n9603) );
  OAI21_X1 U10796 ( .B1(n9603), .B2(n9708), .A(n9602), .ZN(n9757) );
  NAND2_X1 U10797 ( .A1(n9757), .A2(n9989), .ZN(n9604) );
  OAI211_X1 U10798 ( .C1(n9761), .C2(n9736), .A(n9605), .B(n9604), .ZN(
        P1_U3268) );
  XNOR2_X1 U10799 ( .A(n9606), .B(n9609), .ZN(n9766) );
  NAND2_X1 U10800 ( .A1(n9607), .A2(n9608), .ZN(n9610) );
  XNOR2_X1 U10801 ( .A(n9610), .B(n9609), .ZN(n9611) );
  OAI222_X1 U10802 ( .A1(n9712), .A2(n9612), .B1(n9710), .B2(n9649), .C1(n9611), .C2(n9708), .ZN(n9762) );
  INV_X1 U10803 ( .A(n9764), .ZN(n9619) );
  INV_X1 U10804 ( .A(n9614), .ZN(n9615) );
  AOI211_X1 U10805 ( .C1(n9764), .C2(n9613), .A(n9724), .B(n9615), .ZN(n9763)
         );
  NAND2_X1 U10806 ( .A1(n9763), .A2(n9991), .ZN(n9618) );
  AOI22_X1 U10807 ( .A1(n9616), .A2(n9965), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n10001), .ZN(n9617) );
  OAI211_X1 U10808 ( .C1(n9619), .C2(n9994), .A(n9618), .B(n9617), .ZN(n9620)
         );
  AOI21_X1 U10809 ( .B1(n9762), .B2(n9989), .A(n9620), .ZN(n9621) );
  OAI21_X1 U10810 ( .B1(n9766), .B2(n9736), .A(n9621), .ZN(P1_U3269) );
  XOR2_X1 U10811 ( .A(n9622), .B(n9634), .Z(n9771) );
  INV_X1 U10812 ( .A(n9641), .ZN(n9624) );
  INV_X1 U10813 ( .A(n9613), .ZN(n9623) );
  AOI211_X1 U10814 ( .C1(n9769), .C2(n9624), .A(n9724), .B(n9623), .ZN(n9768)
         );
  NOR2_X1 U10815 ( .A1(n9625), .A2(n9994), .ZN(n9629) );
  OAI22_X1 U10816 ( .A1(n9627), .A2(n9987), .B1(n9626), .B2(n9989), .ZN(n9628)
         );
  AOI211_X1 U10817 ( .C1(n9768), .C2(n9991), .A(n9629), .B(n9628), .ZN(n9639)
         );
  NAND2_X1 U10818 ( .A1(n9651), .A2(n9631), .ZN(n9633) );
  INV_X1 U10819 ( .A(n9607), .ZN(n9632) );
  AOI21_X1 U10820 ( .B1(n9634), .B2(n9633), .A(n9632), .ZN(n9635) );
  OAI222_X1 U10821 ( .A1(n9712), .A2(n9637), .B1(n9710), .B2(n9636), .C1(n9708), .C2(n9635), .ZN(n9767) );
  NAND2_X1 U10822 ( .A1(n9767), .A2(n9989), .ZN(n9638) );
  OAI211_X1 U10823 ( .C1(n9771), .C2(n9736), .A(n9639), .B(n9638), .ZN(
        P1_U3270) );
  XNOR2_X1 U10824 ( .A(n9640), .B(n9646), .ZN(n9776) );
  INV_X1 U10825 ( .A(n9663), .ZN(n9642) );
  AOI211_X1 U10826 ( .C1(n9773), .C2(n9642), .A(n9724), .B(n9641), .ZN(n9772)
         );
  AOI22_X1 U10827 ( .A1(n9643), .A2(n9965), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n10001), .ZN(n9644) );
  OAI21_X1 U10828 ( .B1(n9645), .B2(n9994), .A(n9644), .ZN(n9654) );
  AOI21_X1 U10829 ( .B1(n9647), .B2(n9646), .A(n9708), .ZN(n9652) );
  OAI22_X1 U10830 ( .A1(n9649), .A2(n9712), .B1(n9648), .B2(n9710), .ZN(n9650)
         );
  AOI21_X1 U10831 ( .B1(n9652), .B2(n9651), .A(n9650), .ZN(n9775) );
  NOR2_X1 U10832 ( .A1(n9775), .A2(n10001), .ZN(n9653) );
  AOI211_X1 U10833 ( .C1(n9772), .C2(n9991), .A(n9654), .B(n9653), .ZN(n9655)
         );
  OAI21_X1 U10834 ( .B1(n9776), .B2(n9736), .A(n9655), .ZN(P1_U3271) );
  AOI21_X1 U10835 ( .B1(n9657), .B2(n9684), .A(n9656), .ZN(n9658) );
  XOR2_X1 U10836 ( .A(n9668), .B(n9658), .Z(n9660) );
  AOI21_X1 U10837 ( .B1(n9660), .B2(n9962), .A(n9659), .ZN(n9780) );
  NAND2_X1 U10838 ( .A1(n9778), .A2(n4342), .ZN(n9661) );
  NAND2_X1 U10839 ( .A1(n9661), .A2(n10012), .ZN(n9662) );
  NOR2_X1 U10840 ( .A1(n9663), .A2(n9662), .ZN(n9777) );
  INV_X1 U10841 ( .A(n9778), .ZN(n9667) );
  INV_X1 U10842 ( .A(n9664), .ZN(n9665) );
  AOI22_X1 U10843 ( .A1(n9665), .A2(n9965), .B1(n10001), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9666) );
  OAI21_X1 U10844 ( .B1(n9667), .B2(n9994), .A(n9666), .ZN(n9671) );
  XOR2_X1 U10845 ( .A(n9669), .B(n9668), .Z(n9781) );
  NOR2_X1 U10846 ( .A1(n9781), .A2(n9736), .ZN(n9670) );
  AOI211_X1 U10847 ( .C1(n9777), .C2(n9991), .A(n9671), .B(n9670), .ZN(n9672)
         );
  OAI21_X1 U10848 ( .B1(n10001), .B2(n9780), .A(n9672), .ZN(P1_U3272) );
  XNOR2_X1 U10849 ( .A(n8342), .B(n9684), .ZN(n9677) );
  AOI222_X1 U10850 ( .A1(n9962), .A2(n9677), .B1(n9676), .B2(n9675), .C1(n9674), .C2(n9673), .ZN(n9785) );
  NAND2_X1 U10851 ( .A1(n9678), .A2(n9782), .ZN(n9679) );
  AND2_X1 U10852 ( .A1(n4342), .A2(n9679), .ZN(n9783) );
  INV_X1 U10853 ( .A(n9782), .ZN(n9683) );
  INV_X1 U10854 ( .A(n9680), .ZN(n9681) );
  AOI22_X1 U10855 ( .A1(n10001), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9681), 
        .B2(n9965), .ZN(n9682) );
  OAI21_X1 U10856 ( .B1(n9683), .B2(n9994), .A(n9682), .ZN(n9687) );
  XOR2_X1 U10857 ( .A(n9685), .B(n9684), .Z(n9786) );
  NOR2_X1 U10858 ( .A1(n9786), .A2(n9736), .ZN(n9686) );
  AOI211_X1 U10859 ( .C1(n9783), .C2(n9688), .A(n9687), .B(n9686), .ZN(n9689)
         );
  OAI21_X1 U10860 ( .B1(n10001), .B2(n9785), .A(n9689), .ZN(P1_U3273) );
  XNOR2_X1 U10861 ( .A(n9690), .B(n4367), .ZN(n9791) );
  INV_X1 U10862 ( .A(n9691), .ZN(n9693) );
  INV_X1 U10863 ( .A(n9678), .ZN(n9692) );
  AOI211_X1 U10864 ( .C1(n9789), .C2(n9693), .A(n9724), .B(n9692), .ZN(n9788)
         );
  NOR2_X1 U10865 ( .A1(n9694), .A2(n9994), .ZN(n9697) );
  OAI22_X1 U10866 ( .A1(n9989), .A2(n4510), .B1(n9695), .B2(n9987), .ZN(n9696)
         );
  AOI211_X1 U10867 ( .C1(n9788), .C2(n9991), .A(n9697), .B(n9696), .ZN(n9703)
         );
  XNOR2_X1 U10868 ( .A(n9698), .B(n4367), .ZN(n9699) );
  OAI222_X1 U10869 ( .A1(n9712), .A2(n9701), .B1(n9710), .B2(n9700), .C1(n9708), .C2(n9699), .ZN(n9787) );
  NAND2_X1 U10870 ( .A1(n9787), .A2(n9989), .ZN(n9702) );
  OAI211_X1 U10871 ( .C1(n9791), .C2(n9736), .A(n9703), .B(n9702), .ZN(
        P1_U3274) );
  XOR2_X1 U10872 ( .A(n9704), .B(n9706), .Z(n9796) );
  XNOR2_X1 U10873 ( .A(n9705), .B(n9706), .ZN(n9707) );
  OAI222_X1 U10874 ( .A1(n9712), .A2(n9711), .B1(n9710), .B2(n9709), .C1(n9708), .C2(n9707), .ZN(n9792) );
  INV_X1 U10875 ( .A(n9713), .ZN(n9714) );
  AOI211_X1 U10876 ( .C1(n9794), .C2(n9714), .A(n9724), .B(n9691), .ZN(n9793)
         );
  NAND2_X1 U10877 ( .A1(n9793), .A2(n9991), .ZN(n9718) );
  INV_X1 U10878 ( .A(n9715), .ZN(n9716) );
  AOI22_X1 U10879 ( .A1(n10001), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9716), 
        .B2(n9965), .ZN(n9717) );
  OAI211_X1 U10880 ( .C1(n9719), .C2(n9994), .A(n9718), .B(n9717), .ZN(n9720)
         );
  AOI21_X1 U10881 ( .B1(n9792), .B2(n9989), .A(n9720), .ZN(n9721) );
  OAI21_X1 U10882 ( .B1(n9796), .B2(n9736), .A(n9721), .ZN(P1_U3275) );
  XNOR2_X1 U10883 ( .A(n9722), .B(n9730), .ZN(n9801) );
  INV_X1 U10884 ( .A(n9723), .ZN(n9725) );
  AOI211_X1 U10885 ( .C1(n9798), .C2(n9725), .A(n9724), .B(n9713), .ZN(n9797)
         );
  AOI22_X1 U10886 ( .A1(n10001), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9726), 
        .B2(n9965), .ZN(n9727) );
  OAI21_X1 U10887 ( .B1(n9728), .B2(n9994), .A(n9727), .ZN(n9734) );
  XNOR2_X1 U10888 ( .A(n9729), .B(n9730), .ZN(n9732) );
  AOI21_X1 U10889 ( .B1(n9732), .B2(n9962), .A(n9731), .ZN(n9800) );
  NOR2_X1 U10890 ( .A1(n9800), .A2(n10001), .ZN(n9733) );
  AOI211_X1 U10891 ( .C1(n9797), .C2(n9991), .A(n9734), .B(n9733), .ZN(n9735)
         );
  OAI21_X1 U10892 ( .B1(n9736), .B2(n9801), .A(n9735), .ZN(P1_U3276) );
  MUX2_X1 U10893 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9737), .S(n10064), .Z(
        P1_U3553) );
  OAI211_X1 U10894 ( .C1(n9740), .C2(n10020), .A(n9739), .B(n9738), .ZN(n9836)
         );
  MUX2_X1 U10895 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9836), .S(n10064), .Z(
        P1_U3552) );
  AOI21_X1 U10896 ( .B1(n10047), .B2(n9742), .A(n9741), .ZN(n9743) );
  OAI21_X1 U10897 ( .B1(n9746), .B2(n10051), .A(n9745), .ZN(n9837) );
  MUX2_X1 U10898 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9837), .S(n10064), .Z(
        P1_U3550) );
  AOI21_X1 U10899 ( .B1(n10047), .B2(n9748), .A(n9747), .ZN(n9749) );
  OAI211_X1 U10900 ( .C1(n9751), .C2(n10051), .A(n9750), .B(n9749), .ZN(n9838)
         );
  MUX2_X1 U10901 ( .A(n9838), .B(P1_REG1_REG_27__SCAN_IN), .S(n10062), .Z(
        P1_U3549) );
  AOI21_X1 U10902 ( .B1(n10047), .B2(n9753), .A(n9752), .ZN(n9754) );
  OAI211_X1 U10903 ( .C1(n9756), .C2(n10051), .A(n9755), .B(n9754), .ZN(n9839)
         );
  MUX2_X1 U10904 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9839), .S(n10064), .Z(
        P1_U3548) );
  AOI211_X1 U10905 ( .C1(n10047), .C2(n9759), .A(n9758), .B(n9757), .ZN(n9760)
         );
  OAI21_X1 U10906 ( .B1(n9761), .B2(n10051), .A(n9760), .ZN(n9840) );
  MUX2_X1 U10907 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9840), .S(n10064), .Z(
        P1_U3547) );
  AOI211_X1 U10908 ( .C1(n10047), .C2(n9764), .A(n9763), .B(n9762), .ZN(n9765)
         );
  OAI21_X1 U10909 ( .B1(n9766), .B2(n10051), .A(n9765), .ZN(n9841) );
  MUX2_X1 U10910 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9841), .S(n10064), .Z(
        P1_U3546) );
  AOI211_X1 U10911 ( .C1(n10047), .C2(n9769), .A(n9768), .B(n9767), .ZN(n9770)
         );
  OAI21_X1 U10912 ( .B1(n10051), .B2(n9771), .A(n9770), .ZN(n9842) );
  MUX2_X1 U10913 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9842), .S(n10064), .Z(
        P1_U3545) );
  AOI21_X1 U10914 ( .B1(n10047), .B2(n9773), .A(n9772), .ZN(n9774) );
  OAI211_X1 U10915 ( .C1(n9776), .C2(n10051), .A(n9775), .B(n9774), .ZN(n9843)
         );
  MUX2_X1 U10916 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9843), .S(n10064), .Z(
        P1_U3544) );
  AOI21_X1 U10917 ( .B1(n10047), .B2(n9778), .A(n9777), .ZN(n9779) );
  OAI211_X1 U10918 ( .C1(n9781), .C2(n10051), .A(n9780), .B(n9779), .ZN(n9844)
         );
  MUX2_X1 U10919 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9844), .S(n10064), .Z(
        P1_U3543) );
  AOI22_X1 U10920 ( .A1(n9783), .A2(n10012), .B1(n10047), .B2(n9782), .ZN(
        n9784) );
  OAI211_X1 U10921 ( .C1(n9786), .C2(n10051), .A(n9785), .B(n9784), .ZN(n9845)
         );
  MUX2_X1 U10922 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9845), .S(n10064), .Z(
        P1_U3542) );
  AOI211_X1 U10923 ( .C1(n10047), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9790)
         );
  OAI21_X1 U10924 ( .B1(n10051), .B2(n9791), .A(n9790), .ZN(n9846) );
  MUX2_X1 U10925 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9846), .S(n10064), .Z(
        P1_U3541) );
  AOI211_X1 U10926 ( .C1(n10047), .C2(n9794), .A(n9793), .B(n9792), .ZN(n9795)
         );
  OAI21_X1 U10927 ( .B1(n10051), .B2(n9796), .A(n9795), .ZN(n9847) );
  MUX2_X1 U10928 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9847), .S(n10064), .Z(
        P1_U3540) );
  AOI21_X1 U10929 ( .B1(n10047), .B2(n9798), .A(n9797), .ZN(n9799) );
  OAI211_X1 U10930 ( .C1(n9801), .C2(n10051), .A(n9800), .B(n9799), .ZN(n9848)
         );
  MUX2_X1 U10931 ( .A(n9848), .B(P1_REG1_REG_17__SCAN_IN), .S(n10062), .Z(
        P1_U3539) );
  NAND3_X1 U10932 ( .A1(n7861), .A2(n10026), .A3(n9802), .ZN(n9807) );
  NAND2_X1 U10933 ( .A1(n9803), .A2(n10047), .ZN(n9806) );
  NAND2_X1 U10934 ( .A1(n9804), .A2(n10012), .ZN(n9805) );
  NAND4_X1 U10935 ( .A1(n9808), .A2(n9807), .A3(n9806), .A4(n9805), .ZN(n9849)
         );
  MUX2_X1 U10936 ( .A(n9849), .B(P1_REG1_REG_16__SCAN_IN), .S(n10062), .Z(
        P1_U3538) );
  AOI211_X1 U10937 ( .C1(n10047), .C2(n9811), .A(n9810), .B(n9809), .ZN(n9812)
         );
  OAI21_X1 U10938 ( .B1(n10051), .B2(n9813), .A(n9812), .ZN(n9850) );
  MUX2_X1 U10939 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9850), .S(n10064), .Z(
        P1_U3537) );
  AOI21_X1 U10940 ( .B1(n10047), .B2(n9815), .A(n9814), .ZN(n9816) );
  OAI211_X1 U10941 ( .C1(n9818), .C2(n10031), .A(n9817), .B(n9816), .ZN(n9851)
         );
  MUX2_X1 U10942 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9851), .S(n10064), .Z(
        P1_U3536) );
  INV_X1 U10943 ( .A(n9819), .ZN(n9824) );
  AOI22_X1 U10944 ( .A1(n9821), .A2(n10012), .B1(n10047), .B2(n9820), .ZN(
        n9822) );
  OAI211_X1 U10945 ( .C1(n10051), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9852)
         );
  MUX2_X1 U10946 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9852), .S(n10064), .Z(
        P1_U3535) );
  AOI21_X1 U10947 ( .B1(n10047), .B2(n9826), .A(n9825), .ZN(n9827) );
  OAI211_X1 U10948 ( .C1(n10051), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9853)
         );
  MUX2_X1 U10949 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9853), .S(n10064), .Z(
        P1_U3534) );
  AOI21_X1 U10950 ( .B1(n10047), .B2(n9831), .A(n9830), .ZN(n9832) );
  OAI211_X1 U10951 ( .C1(n10051), .C2(n9834), .A(n9833), .B(n9832), .ZN(n9854)
         );
  MUX2_X1 U10952 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9854), .S(n10064), .Z(
        P1_U3532) );
  MUX2_X1 U10953 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9835), .S(n10064), .Z(
        P1_U3523) );
  MUX2_X1 U10954 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9836), .S(n10055), .Z(
        P1_U3520) );
  MUX2_X1 U10955 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9837), .S(n10055), .Z(
        P1_U3518) );
  MUX2_X1 U10956 ( .A(n9838), .B(P1_REG0_REG_27__SCAN_IN), .S(n10053), .Z(
        P1_U3517) );
  MUX2_X1 U10957 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9839), .S(n10055), .Z(
        P1_U3516) );
  MUX2_X1 U10958 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9840), .S(n10055), .Z(
        P1_U3515) );
  MUX2_X1 U10959 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9841), .S(n10055), .Z(
        P1_U3514) );
  MUX2_X1 U10960 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9842), .S(n10055), .Z(
        P1_U3513) );
  MUX2_X1 U10961 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9843), .S(n10055), .Z(
        P1_U3512) );
  MUX2_X1 U10962 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9844), .S(n10055), .Z(
        P1_U3511) );
  MUX2_X1 U10963 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9845), .S(n10055), .Z(
        P1_U3510) );
  MUX2_X1 U10964 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9846), .S(n10055), .Z(
        P1_U3509) );
  MUX2_X1 U10965 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9847), .S(n10055), .Z(
        P1_U3507) );
  MUX2_X1 U10966 ( .A(n9848), .B(P1_REG0_REG_17__SCAN_IN), .S(n10053), .Z(
        P1_U3504) );
  MUX2_X1 U10967 ( .A(n9849), .B(P1_REG0_REG_16__SCAN_IN), .S(n10053), .Z(
        P1_U3501) );
  MUX2_X1 U10968 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9850), .S(n10055), .Z(
        P1_U3498) );
  MUX2_X1 U10969 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9851), .S(n10055), .Z(
        P1_U3495) );
  MUX2_X1 U10970 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9852), .S(n10055), .Z(
        P1_U3492) );
  MUX2_X1 U10971 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9853), .S(n10055), .Z(
        P1_U3489) );
  MUX2_X1 U10972 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n9854), .S(n10055), .Z(
        P1_U3483) );
  MUX2_X1 U10973 ( .A(n9855), .B(P1_D_REG_0__SCAN_IN), .S(n10003), .Z(P1_U3439) );
  NAND3_X1 U10974 ( .A1(n10193), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9857) );
  OAI22_X1 U10975 ( .A1(n6136), .A2(n9857), .B1(n9856), .B2(n9866), .ZN(n9858)
         );
  AOI21_X1 U10976 ( .B1(n9860), .B2(n9859), .A(n9858), .ZN(n9861) );
  INV_X1 U10977 ( .A(n9861), .ZN(P1_U3324) );
  OAI222_X1 U10978 ( .A1(n9866), .A2(n9865), .B1(n9864), .B2(n9863), .C1(n9862), .C2(P1_U3086), .ZN(P1_U3328) );
  MUX2_X1 U10979 ( .A(n9867), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U10980 ( .A1(n9868), .A2(n9869), .ZN(n9918) );
  NOR2_X1 U10981 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9914) );
  NOR2_X1 U10982 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9912) );
  NOR2_X1 U10983 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9910) );
  NOR2_X1 U10984 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9908) );
  NOR2_X1 U10985 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9906) );
  NOR2_X1 U10986 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9903) );
  NOR2_X1 U10987 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9901) );
  NOR2_X1 U10988 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9898) );
  NOR2_X1 U10989 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9895) );
  NOR2_X1 U10990 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9892) );
  NOR2_X1 U10991 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9889) );
  NOR2_X1 U10992 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9886) );
  NOR2_X1 U10993 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n9883) );
  NOR2_X1 U10994 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9880) );
  NAND2_X1 U10995 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9877) );
  XNOR2_X1 U10996 ( .A(n9870), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10308) );
  NAND2_X1 U10997 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9875) );
  AOI21_X1 U10998 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U10999 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9871) );
  NOR2_X1 U11000 ( .A1(n9408), .A2(n9871), .ZN(n10132) );
  NOR2_X1 U11001 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10132), .ZN(n9872) );
  NOR2_X1 U11002 ( .A1(n10133), .A2(n9872), .ZN(n10306) );
  INV_X1 U11003 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9873) );
  INV_X1 U11004 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U11005 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .B1(n9873), .B2(n10216), .ZN(n10305) );
  NAND2_X1 U11006 ( .A1(n10306), .A2(n10305), .ZN(n9874) );
  NAND2_X1 U11007 ( .A1(n9875), .A2(n9874), .ZN(n10307) );
  NAND2_X1 U11008 ( .A1(n10308), .A2(n10307), .ZN(n9876) );
  NAND2_X1 U11009 ( .A1(n9877), .A2(n9876), .ZN(n10310) );
  XOR2_X1 U11010 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n9878), .Z(n10309) );
  NOR2_X1 U11011 ( .A1(n10310), .A2(n10309), .ZN(n9879) );
  NOR2_X1 U11012 ( .A1(n9880), .A2(n9879), .ZN(n10298) );
  XOR2_X1 U11013 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n9881), .Z(n10297) );
  NOR2_X1 U11014 ( .A1(n10298), .A2(n10297), .ZN(n9882) );
  NOR2_X1 U11015 ( .A1(n9883), .A2(n9882), .ZN(n10296) );
  XOR2_X1 U11016 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n9884), .Z(n10295) );
  NOR2_X1 U11017 ( .A1(n10296), .A2(n10295), .ZN(n9885) );
  NOR2_X1 U11018 ( .A1(n9886), .A2(n9885), .ZN(n10302) );
  XOR2_X1 U11019 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n9887), .Z(n10301) );
  NOR2_X1 U11020 ( .A1(n10302), .A2(n10301), .ZN(n9888) );
  XOR2_X1 U11021 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9890), .Z(n10303) );
  NOR2_X1 U11022 ( .A1(n10304), .A2(n10303), .ZN(n9891) );
  XOR2_X1 U11023 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9893), .Z(n10299) );
  NOR2_X1 U11024 ( .A1(n10300), .A2(n10299), .ZN(n9894) );
  INV_X1 U11025 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U11026 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9896), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10192), .ZN(n10152) );
  XOR2_X1 U11027 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n9899), .Z(n10150) );
  INV_X1 U11028 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U11029 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7522), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10233), .ZN(n10148) );
  XOR2_X1 U11030 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n9904), .Z(n10146) );
  INV_X1 U11031 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9930) );
  XOR2_X1 U11032 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n9930), .Z(n10144) );
  INV_X1 U11033 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9943) );
  INV_X1 U11034 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U11035 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9943), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10203), .ZN(n10142) );
  NOR2_X1 U11036 ( .A1(n10143), .A2(n10142), .ZN(n9909) );
  NOR2_X1 U11037 ( .A1(n9910), .A2(n9909), .ZN(n10141) );
  XNOR2_X1 U11038 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10140) );
  NOR2_X1 U11039 ( .A1(n10141), .A2(n10140), .ZN(n9911) );
  NOR2_X1 U11040 ( .A1(n9912), .A2(n9911), .ZN(n10139) );
  XNOR2_X1 U11041 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10138) );
  NOR2_X1 U11042 ( .A1(n10139), .A2(n10138), .ZN(n9913) );
  NOR2_X1 U11043 ( .A1(n9914), .A2(n9913), .ZN(n9915) );
  NOR2_X1 U11044 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9915), .ZN(n10136) );
  AND2_X1 U11045 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9915), .ZN(n10135) );
  NOR2_X1 U11046 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10135), .ZN(n9916) );
  NOR2_X1 U11047 ( .A1(n10136), .A2(n9916), .ZN(n9917) );
  XOR2_X1 U11048 ( .A(n9918), .B(n9917), .Z(ADD_1068_U4) );
  INV_X1 U11049 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10205) );
  XOR2_X1 U11050 ( .A(n10205), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  AOI211_X1 U11051 ( .C1(n9921), .C2(n9920), .A(n9934), .B(n9919), .ZN(n9926)
         );
  AOI211_X1 U11052 ( .C1(n9924), .C2(n9923), .A(n9944), .B(n9922), .ZN(n9925)
         );
  AOI211_X1 U11053 ( .C1(n9947), .C2(n9927), .A(n9926), .B(n9925), .ZN(n9929)
         );
  OAI211_X1 U11054 ( .C1(n9960), .C2(n9930), .A(n9929), .B(n9928), .ZN(
        P1_U3257) );
  AOI211_X1 U11055 ( .C1(n9933), .C2(n9932), .A(n9931), .B(n9944), .ZN(n9939)
         );
  AOI211_X1 U11056 ( .C1(n9937), .C2(n9936), .A(n9935), .B(n9934), .ZN(n9938)
         );
  AOI211_X1 U11057 ( .C1(n9947), .C2(n9940), .A(n9939), .B(n9938), .ZN(n9942)
         );
  OAI211_X1 U11058 ( .C1(n9960), .C2(n9943), .A(n9942), .B(n9941), .ZN(
        P1_U3258) );
  INV_X1 U11059 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9959) );
  AOI21_X1 U11060 ( .B1(n9946), .B2(n9945), .A(n9944), .ZN(n9950) );
  AOI22_X1 U11061 ( .A1(n9950), .A2(n9949), .B1(n9948), .B2(n9947), .ZN(n9956)
         );
  OAI211_X1 U11062 ( .C1(n9954), .C2(n9953), .A(n9952), .B(n9951), .ZN(n9955)
         );
  AND2_X1 U11063 ( .A1(n9956), .A2(n9955), .ZN(n9958) );
  NAND2_X1 U11064 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9957) );
  OAI211_X1 U11065 ( .C1(n9960), .C2(n9959), .A(n9958), .B(n9957), .ZN(
        P1_U3261) );
  XNOR2_X1 U11066 ( .A(n9969), .B(n7475), .ZN(n9963) );
  AOI21_X1 U11067 ( .B1(n9963), .B2(n9962), .A(n9961), .ZN(n10022) );
  AOI222_X1 U11068 ( .A1(n9967), .A2(n9966), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n10001), .C1(n9965), .C2(n9964), .ZN(n9974) );
  XNOR2_X1 U11069 ( .A(n9969), .B(n9968), .ZN(n10025) );
  OAI211_X1 U11070 ( .C1(n4425), .C2(n10021), .A(n10012), .B(n9970), .ZN(
        n10019) );
  INV_X1 U11071 ( .A(n10019), .ZN(n9971) );
  AOI22_X1 U11072 ( .A1(n10025), .A2(n9972), .B1(n9991), .B2(n9971), .ZN(n9973) );
  OAI211_X1 U11073 ( .C1(n10001), .C2(n10022), .A(n9974), .B(n9973), .ZN(
        P1_U3287) );
  INV_X1 U11074 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9977) );
  INV_X1 U11075 ( .A(n9975), .ZN(n9976) );
  OAI22_X1 U11076 ( .A1(n9987), .A2(n9977), .B1(n6374), .B2(n9976), .ZN(n9979)
         );
  AOI211_X1 U11077 ( .C1(n9981), .C2(n9980), .A(n9979), .B(n9978), .ZN(n9984)
         );
  OAI22_X1 U11078 ( .A1(n9984), .A2(n10001), .B1(n9983), .B2(n9982), .ZN(n9985) );
  INV_X1 U11079 ( .A(n9985), .ZN(n9986) );
  OAI21_X1 U11080 ( .B1(n6998), .B2(n9989), .A(n9986), .ZN(P1_U3291) );
  OAI22_X1 U11081 ( .A1(n9989), .A2(n6997), .B1(n9988), .B2(n9987), .ZN(n9990)
         );
  AOI21_X1 U11082 ( .B1(n9992), .B2(n9991), .A(n9990), .ZN(n9993) );
  OAI21_X1 U11083 ( .B1(n9995), .B2(n9994), .A(n9993), .ZN(n9996) );
  AOI21_X1 U11084 ( .B1(n9998), .B2(n9997), .A(n9996), .ZN(n9999) );
  OAI21_X1 U11085 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(P1_U3292) );
  AND2_X1 U11086 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10003), .ZN(P1_U3294) );
  AND2_X1 U11087 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10003), .ZN(P1_U3295) );
  AND2_X1 U11088 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10003), .ZN(P1_U3296) );
  AND2_X1 U11089 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10003), .ZN(P1_U3297) );
  AND2_X1 U11090 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10003), .ZN(P1_U3298) );
  AND2_X1 U11091 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10003), .ZN(P1_U3299) );
  AND2_X1 U11092 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10003), .ZN(P1_U3300) );
  AND2_X1 U11093 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10003), .ZN(P1_U3301) );
  INV_X1 U11094 ( .A(n10003), .ZN(n10002) );
  INV_X1 U11095 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10271) );
  NOR2_X1 U11096 ( .A1(n10002), .A2(n10271), .ZN(P1_U3302) );
  AND2_X1 U11097 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10003), .ZN(P1_U3303) );
  AND2_X1 U11098 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10003), .ZN(P1_U3304) );
  AND2_X1 U11099 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10003), .ZN(P1_U3305) );
  AND2_X1 U11100 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10003), .ZN(P1_U3306) );
  INV_X1 U11101 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10258) );
  NOR2_X1 U11102 ( .A1(n10002), .A2(n10258), .ZN(P1_U3307) );
  AND2_X1 U11103 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10003), .ZN(P1_U3308) );
  AND2_X1 U11104 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10003), .ZN(P1_U3309) );
  AND2_X1 U11105 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10003), .ZN(P1_U3310) );
  AND2_X1 U11106 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10003), .ZN(P1_U3311) );
  AND2_X1 U11107 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10003), .ZN(P1_U3312) );
  AND2_X1 U11108 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10003), .ZN(P1_U3313) );
  AND2_X1 U11109 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10003), .ZN(P1_U3314) );
  INV_X1 U11110 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10274) );
  NOR2_X1 U11111 ( .A1(n10002), .A2(n10274), .ZN(P1_U3315) );
  AND2_X1 U11112 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10003), .ZN(P1_U3316) );
  AND2_X1 U11113 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10003), .ZN(P1_U3317) );
  AND2_X1 U11114 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10003), .ZN(P1_U3318) );
  AND2_X1 U11115 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10003), .ZN(P1_U3319) );
  AND2_X1 U11116 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10003), .ZN(P1_U3320) );
  AND2_X1 U11117 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10003), .ZN(P1_U3321) );
  AND2_X1 U11118 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10003), .ZN(P1_U3322) );
  AND2_X1 U11119 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10003), .ZN(P1_U3323) );
  AOI22_X1 U11120 ( .A1(n10005), .A2(n10012), .B1(n10047), .B2(n10004), .ZN(
        n10006) );
  OAI211_X1 U11121 ( .C1(n10051), .C2(n10008), .A(n10007), .B(n10006), .ZN(
        n10009) );
  INV_X1 U11122 ( .A(n10009), .ZN(n10056) );
  INV_X1 U11123 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10010) );
  AOI22_X1 U11124 ( .A1(n10055), .A2(n10056), .B1(n10010), .B2(n10053), .ZN(
        P1_U3465) );
  AOI22_X1 U11125 ( .A1(n10013), .A2(n10012), .B1(n10047), .B2(n10011), .ZN(
        n10014) );
  OAI211_X1 U11126 ( .C1(n10051), .C2(n10016), .A(n10015), .B(n10014), .ZN(
        n10017) );
  INV_X1 U11127 ( .A(n10017), .ZN(n10057) );
  INV_X1 U11128 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10018) );
  AOI22_X1 U11129 ( .A1(n10055), .A2(n10057), .B1(n10018), .B2(n10053), .ZN(
        P1_U3468) );
  OAI21_X1 U11130 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10024) );
  INV_X1 U11131 ( .A(n10022), .ZN(n10023) );
  AOI211_X1 U11132 ( .C1(n10026), .C2(n10025), .A(n10024), .B(n10023), .ZN(
        n10058) );
  INV_X1 U11133 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10027) );
  AOI22_X1 U11134 ( .A1(n10055), .A2(n10058), .B1(n10027), .B2(n10053), .ZN(
        P1_U3471) );
  INV_X1 U11135 ( .A(n10032), .ZN(n10035) );
  AOI21_X1 U11136 ( .B1(n10047), .B2(n10029), .A(n10028), .ZN(n10030) );
  OAI21_X1 U11137 ( .B1(n10032), .B2(n10031), .A(n10030), .ZN(n10034) );
  AOI211_X1 U11138 ( .C1(n10036), .C2(n10035), .A(n10034), .B(n10033), .ZN(
        n10060) );
  INV_X1 U11139 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10037) );
  AOI22_X1 U11140 ( .A1(n10055), .A2(n10060), .B1(n10037), .B2(n10053), .ZN(
        P1_U3474) );
  AOI21_X1 U11141 ( .B1(n10047), .B2(n10039), .A(n10038), .ZN(n10040) );
  OAI211_X1 U11142 ( .C1(n10051), .C2(n10042), .A(n10041), .B(n10040), .ZN(
        n10043) );
  INV_X1 U11143 ( .A(n10043), .ZN(n10061) );
  INV_X1 U11144 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U11145 ( .A1(n10055), .A2(n10061), .B1(n10044), .B2(n10053), .ZN(
        P1_U3477) );
  AOI21_X1 U11146 ( .B1(n10047), .B2(n10046), .A(n10045), .ZN(n10048) );
  OAI211_X1 U11147 ( .C1(n10051), .C2(n10050), .A(n10049), .B(n10048), .ZN(
        n10052) );
  INV_X1 U11148 ( .A(n10052), .ZN(n10063) );
  INV_X1 U11149 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U11150 ( .A1(n10055), .A2(n10063), .B1(n10054), .B2(n10053), .ZN(
        P1_U3480) );
  AOI22_X1 U11151 ( .A1(n10064), .A2(n10056), .B1(n7014), .B2(n10062), .ZN(
        P1_U3526) );
  AOI22_X1 U11152 ( .A1(n10064), .A2(n10057), .B1(n7016), .B2(n10062), .ZN(
        P1_U3527) );
  AOI22_X1 U11153 ( .A1(n10064), .A2(n10058), .B1(n7018), .B2(n10062), .ZN(
        P1_U3528) );
  INV_X1 U11154 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10059) );
  AOI22_X1 U11155 ( .A1(n10064), .A2(n10060), .B1(n10059), .B2(n10062), .ZN(
        P1_U3529) );
  AOI22_X1 U11156 ( .A1(n10064), .A2(n10061), .B1(n7019), .B2(n10062), .ZN(
        P1_U3530) );
  AOI22_X1 U11157 ( .A1(n10064), .A2(n10063), .B1(n7021), .B2(n10062), .ZN(
        P1_U3531) );
  XNOR2_X1 U11158 ( .A(n10066), .B(n10065), .ZN(n10071) );
  OAI21_X1 U11159 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n10068), .A(n10067), .ZN(
        n10069) );
  NAND2_X1 U11160 ( .A1(n10114), .A2(n10069), .ZN(n10070) );
  OAI21_X1 U11161 ( .B1(n10071), .B2(n10106), .A(n10070), .ZN(n10074) );
  OAI21_X1 U11162 ( .B1(n10111), .B2(n4790), .A(n10072), .ZN(n10073) );
  NOR2_X1 U11163 ( .A1(n10074), .A2(n10073), .ZN(n10081) );
  AOI21_X1 U11164 ( .B1(n10077), .B2(n10076), .A(n10075), .ZN(n10078) );
  NOR2_X1 U11165 ( .A1(n10078), .A2(n10099), .ZN(n10079) );
  AOI21_X1 U11166 ( .B1(n10118), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n10079), .ZN(
        n10080) );
  NAND2_X1 U11167 ( .A1(n10081), .A2(n10080), .ZN(P2_U3185) );
  OAI21_X1 U11168 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(n10094) );
  AND3_X1 U11169 ( .A1(n6922), .A2(n10086), .A3(n10085), .ZN(n10087) );
  OAI21_X1 U11170 ( .B1(n10088), .B2(n10087), .A(n10114), .ZN(n10091) );
  INV_X1 U11171 ( .A(n10089), .ZN(n10090) );
  OAI211_X1 U11172 ( .C1(n10111), .C2(n10092), .A(n10091), .B(n10090), .ZN(
        n10093) );
  AOI21_X1 U11173 ( .B1(n10095), .B2(n10094), .A(n10093), .ZN(n10103) );
  AOI21_X1 U11174 ( .B1(n10098), .B2(n10097), .A(n10096), .ZN(n10100) );
  NOR2_X1 U11175 ( .A1(n10100), .A2(n10099), .ZN(n10101) );
  AOI21_X1 U11176 ( .B1(n10118), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n10101), .ZN(
        n10102) );
  NAND2_X1 U11177 ( .A1(n10103), .A2(n10102), .ZN(P2_U3188) );
  OAI21_X1 U11178 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n10104), .A(n7181), .ZN(
        n10115) );
  XOR2_X1 U11179 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10105), .Z(n10107) );
  NOR2_X1 U11180 ( .A1(n10107), .A2(n10106), .ZN(n10113) );
  INV_X1 U11181 ( .A(n10108), .ZN(n10109) );
  OAI21_X1 U11182 ( .B1(n10111), .B2(n10110), .A(n10109), .ZN(n10112) );
  AOI211_X1 U11183 ( .C1(n10115), .C2(n10114), .A(n10113), .B(n10112), .ZN(
        n10121) );
  XNOR2_X1 U11184 ( .A(n10117), .B(n10116), .ZN(n10119) );
  AOI22_X1 U11185 ( .A1(n10119), .A2(n6751), .B1(n10118), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U11186 ( .A1(n10121), .A2(n10120), .ZN(P2_U3189) );
  AOI22_X1 U11187 ( .A1(n10292), .A2(n5014), .B1(n10122), .B2(n5734), .ZN(
        P2_U3393) );
  INV_X1 U11188 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U11189 ( .A1(n10292), .A2(n10124), .B1(n10123), .B2(n5734), .ZN(
        P2_U3396) );
  AOI22_X1 U11190 ( .A1(n10292), .A2(n5059), .B1(n10125), .B2(n5734), .ZN(
        P2_U3399) );
  INV_X1 U11191 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U11192 ( .A1(n10292), .A2(n10127), .B1(n10126), .B2(n5734), .ZN(
        P2_U3402) );
  INV_X1 U11193 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U11194 ( .A1(n10292), .A2(n10129), .B1(n10128), .B2(n5734), .ZN(
        P2_U3405) );
  INV_X1 U11195 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U11196 ( .A1(n10292), .A2(n10131), .B1(n10130), .B2(n5734), .ZN(
        P2_U3411) );
  NOR2_X1 U11197 ( .A1(n10133), .A2(n10132), .ZN(n10134) );
  XOR2_X1 U11198 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10134), .Z(ADD_1068_U5) );
  XOR2_X1 U11199 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11200 ( .A1(n10136), .A2(n10135), .ZN(n10137) );
  XOR2_X1 U11201 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10137), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11202 ( .A(n10139), .B(n10138), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11203 ( .A(n10141), .B(n10140), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11204 ( .A(n10143), .B(n10142), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11205 ( .A(n10145), .B(n10144), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11206 ( .A(n10147), .B(n10146), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11207 ( .A(n10149), .B(n10148), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11208 ( .A(n10151), .B(n10150), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11209 ( .A(n10153), .B(n10152), .ZN(ADD_1068_U63) );
  INV_X1 U11210 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10208) );
  NAND4_X1 U11211 ( .A1(P2_WR_REG_SCAN_IN), .A2(n10206), .A3(n10208), .A4(
        n7019), .ZN(n10159) );
  NAND4_X1 U11212 ( .A1(P2_D_REG_1__SCAN_IN), .A2(P1_REG2_REG_22__SCAN_IN), 
        .A3(n10218), .A4(n10203), .ZN(n10158) );
  NAND4_X1 U11213 ( .A1(SI_16_), .A2(P1_IR_REG_16__SCAN_IN), .A3(
        P1_REG0_REG_31__SCAN_IN), .A4(n10154), .ZN(n10155) );
  NOR2_X1 U11214 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(n10155), .ZN(n10156) );
  NAND4_X1 U11215 ( .A1(n10156), .A2(P2_REG0_REG_3__SCAN_IN), .A3(n10221), 
        .A4(P1_REG0_REG_30__SCAN_IN), .ZN(n10157) );
  NOR3_X1 U11216 ( .A1(n10159), .A2(n10158), .A3(n10157), .ZN(n10290) );
  NAND4_X1 U11217 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), 
        .A3(P1_D_REG_10__SCAN_IN), .A4(P1_REG1_REG_11__SCAN_IN), .ZN(n10180)
         );
  NAND4_X1 U11218 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .A3(
        P1_B_REG_SCAN_IN), .A4(n10160), .ZN(n10179) );
  NOR3_X1 U11219 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(P2_REG2_REG_11__SCAN_IN), 
        .A3(n10262), .ZN(n10162) );
  NOR3_X1 U11220 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        n10259), .ZN(n10161) );
  NAND4_X1 U11221 ( .A1(P2_B_REG_SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .A3(
        n10162), .A4(n10161), .ZN(n10178) );
  NOR4_X1 U11222 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG0_REG_1__SCAN_IN), 
        .A3(P1_REG2_REG_0__SCAN_IN), .A4(P2_ADDR_REG_2__SCAN_IN), .ZN(n10176)
         );
  NOR4_X1 U11223 ( .A1(SI_10_), .A2(P2_IR_REG_15__SCAN_IN), .A3(
        P1_DATAO_REG_0__SCAN_IN), .A4(n5098), .ZN(n10175) );
  NAND4_X1 U11224 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(SI_4_), .A3(
        P1_REG3_REG_8__SCAN_IN), .A4(n5336), .ZN(n10165) );
  NAND3_X1 U11225 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .A3(n10163), .ZN(n10164) );
  NOR3_X1 U11226 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(n10165), .A3(n10164), .ZN(
        n10174) );
  NAND4_X1 U11227 ( .A1(n10166), .A2(n10247), .A3(P1_REG3_REG_0__SCAN_IN), 
        .A4(P1_REG1_REG_4__SCAN_IN), .ZN(n10172) );
  NAND4_X1 U11228 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(P1_REG3_REG_13__SCAN_IN), 
        .A3(P1_REG2_REG_29__SCAN_IN), .A4(n10237), .ZN(n10169) );
  NAND4_X1 U11229 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), 
        .A3(n10167), .A4(n10233), .ZN(n10168) );
  OR4_X1 U11230 ( .A1(n10246), .A2(P1_IR_REG_9__SCAN_IN), .A3(n10169), .A4(
        n10168), .ZN(n10171) );
  NOR4_X1 U11231 ( .A1(n10172), .A2(n10171), .A3(P2_IR_REG_1__SCAN_IN), .A4(
        n10170), .ZN(n10173) );
  NAND4_X1 U11232 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  NOR4_X1 U11233 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10289) );
  AOI22_X1 U11234 ( .A1(n10182), .A2(keyinput16), .B1(n5014), .B2(keyinput63), 
        .ZN(n10181) );
  OAI221_X1 U11235 ( .B1(n10182), .B2(keyinput16), .C1(n5014), .C2(keyinput63), 
        .A(n10181), .ZN(n10190) );
  XNOR2_X1 U11236 ( .A(keyinput49), .B(n5336), .ZN(n10189) );
  XNOR2_X1 U11237 ( .A(keyinput55), .B(n5098), .ZN(n10188) );
  XNOR2_X1 U11238 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput25), .ZN(n10186)
         );
  XNOR2_X1 U11239 ( .A(SI_4_), .B(keyinput35), .ZN(n10185) );
  XNOR2_X1 U11240 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput14), .ZN(n10184) );
  XNOR2_X1 U11241 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput61), .ZN(n10183) );
  NAND4_X1 U11242 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10187) );
  NOR4_X1 U11243 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10231) );
  AOI22_X1 U11244 ( .A1(n5036), .A2(keyinput39), .B1(keyinput40), .B2(n10192), 
        .ZN(n10191) );
  OAI221_X1 U11245 ( .B1(n5036), .B2(keyinput39), .C1(n10192), .C2(keyinput40), 
        .A(n10191), .ZN(n10201) );
  XOR2_X1 U11246 ( .A(P1_REG0_REG_31__SCAN_IN), .B(keyinput10), .Z(n10200) );
  XNOR2_X1 U11247 ( .A(n10193), .B(keyinput21), .ZN(n10199) );
  XNOR2_X1 U11248 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput36), .ZN(n10197) );
  XNOR2_X1 U11249 ( .A(SI_10_), .B(keyinput30), .ZN(n10196) );
  XNOR2_X1 U11250 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput28), .ZN(n10195) );
  XNOR2_X1 U11251 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput38), .ZN(n10194) );
  NAND4_X1 U11252 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10198) );
  NOR4_X1 U11253 ( .A1(n10201), .A2(n10200), .A3(n10199), .A4(n10198), .ZN(
        n10230) );
  AOI22_X1 U11254 ( .A1(n7019), .A2(keyinput60), .B1(keyinput5), .B2(n10203), 
        .ZN(n10202) );
  OAI221_X1 U11255 ( .B1(n7019), .B2(keyinput60), .C1(n10203), .C2(keyinput5), 
        .A(n10202), .ZN(n10214) );
  AOI22_X1 U11256 ( .A1(n10206), .A2(keyinput2), .B1(keyinput13), .B2(n10205), 
        .ZN(n10204) );
  OAI221_X1 U11257 ( .B1(n10206), .B2(keyinput2), .C1(n10205), .C2(keyinput13), 
        .A(n10204), .ZN(n10213) );
  AOI22_X1 U11258 ( .A1(n5313), .A2(keyinput11), .B1(keyinput52), .B2(n10208), 
        .ZN(n10207) );
  OAI221_X1 U11259 ( .B1(n5313), .B2(keyinput11), .C1(n10208), .C2(keyinput52), 
        .A(n10207), .ZN(n10212) );
  XNOR2_X1 U11260 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput59), .ZN(n10210) );
  XNOR2_X1 U11261 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput45), .ZN(n10209)
         );
  NAND2_X1 U11262 ( .A1(n10210), .A2(n10209), .ZN(n10211) );
  NOR4_X1 U11263 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10229) );
  AOI22_X1 U11264 ( .A1(n6491), .A2(keyinput53), .B1(keyinput20), .B2(n10216), 
        .ZN(n10215) );
  OAI221_X1 U11265 ( .B1(n6491), .B2(keyinput53), .C1(n10216), .C2(keyinput20), 
        .A(n10215), .ZN(n10227) );
  AOI22_X1 U11266 ( .A1(n10218), .A2(keyinput27), .B1(n8113), .B2(keyinput3), 
        .ZN(n10217) );
  OAI221_X1 U11267 ( .B1(n10218), .B2(keyinput27), .C1(n8113), .C2(keyinput3), 
        .A(n10217), .ZN(n10226) );
  AOI22_X1 U11268 ( .A1(n10221), .A2(keyinput51), .B1(keyinput15), .B2(n10220), 
        .ZN(n10219) );
  OAI221_X1 U11269 ( .B1(n10221), .B2(keyinput51), .C1(n10220), .C2(keyinput15), .A(n10219), .ZN(n10225) );
  XOR2_X1 U11270 ( .A(n5059), .B(keyinput44), .Z(n10223) );
  XNOR2_X1 U11271 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput7), .ZN(n10222) );
  NAND2_X1 U11272 ( .A1(n10223), .A2(n10222), .ZN(n10224) );
  NOR4_X1 U11273 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n10228) );
  NAND4_X1 U11274 ( .A1(n10231), .A2(n10230), .A3(n10229), .A4(n10228), .ZN(
        n10288) );
  AOI22_X1 U11275 ( .A1(P1_U3086), .A2(keyinput41), .B1(keyinput43), .B2(
        n10233), .ZN(n10232) );
  OAI221_X1 U11276 ( .B1(P1_U3086), .B2(keyinput41), .C1(n10233), .C2(
        keyinput43), .A(n10232), .ZN(n10244) );
  AOI22_X1 U11277 ( .A1(n5142), .A2(keyinput24), .B1(keyinput23), .B2(n10235), 
        .ZN(n10234) );
  OAI221_X1 U11278 ( .B1(n5142), .B2(keyinput24), .C1(n10235), .C2(keyinput23), 
        .A(n10234), .ZN(n10243) );
  AOI22_X1 U11279 ( .A1(n10238), .A2(keyinput56), .B1(n10237), .B2(keyinput48), 
        .ZN(n10236) );
  OAI221_X1 U11280 ( .B1(n10238), .B2(keyinput56), .C1(n10237), .C2(keyinput48), .A(n10236), .ZN(n10242) );
  XNOR2_X1 U11281 ( .A(P2_REG0_REG_25__SCAN_IN), .B(keyinput1), .ZN(n10240) );
  XNOR2_X1 U11282 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput42), .ZN(n10239) );
  NAND2_X1 U11283 ( .A1(n10240), .A2(n10239), .ZN(n10241) );
  NOR4_X1 U11284 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10286) );
  AOI22_X1 U11285 ( .A1(n7014), .A2(keyinput50), .B1(n10246), .B2(keyinput12), 
        .ZN(n10245) );
  OAI221_X1 U11286 ( .B1(n7014), .B2(keyinput50), .C1(n10246), .C2(keyinput12), 
        .A(n10245), .ZN(n10256) );
  XNOR2_X1 U11287 ( .A(n10247), .B(keyinput46), .ZN(n10255) );
  XNOR2_X1 U11288 ( .A(keyinput8), .B(n10248), .ZN(n10254) );
  XNOR2_X1 U11289 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput9), .ZN(n10252) );
  XNOR2_X1 U11290 ( .A(SI_19_), .B(keyinput26), .ZN(n10251) );
  XNOR2_X1 U11291 ( .A(P2_REG0_REG_12__SCAN_IN), .B(keyinput29), .ZN(n10250)
         );
  XNOR2_X1 U11292 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput0), .ZN(n10249) );
  NAND4_X1 U11293 ( .A1(n10252), .A2(n10251), .A3(n10250), .A4(n10249), .ZN(
        n10253) );
  NOR4_X1 U11294 ( .A1(n10256), .A2(n10255), .A3(n10254), .A4(n10253), .ZN(
        n10285) );
  AOI22_X1 U11295 ( .A1(n10259), .A2(keyinput6), .B1(keyinput18), .B2(n10258), 
        .ZN(n10257) );
  OAI221_X1 U11296 ( .B1(n10259), .B2(keyinput6), .C1(n10258), .C2(keyinput18), 
        .A(n10257), .ZN(n10269) );
  AOI22_X1 U11297 ( .A1(n10262), .A2(keyinput47), .B1(keyinput17), .B2(n10261), 
        .ZN(n10260) );
  OAI221_X1 U11298 ( .B1(n10262), .B2(keyinput47), .C1(n10261), .C2(keyinput17), .A(n10260), .ZN(n10268) );
  XOR2_X1 U11299 ( .A(n5558), .B(keyinput22), .Z(n10266) );
  XNOR2_X1 U11300 ( .A(P2_B_REG_SCAN_IN), .B(keyinput19), .ZN(n10265) );
  XNOR2_X1 U11301 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput4), .ZN(n10264) );
  XNOR2_X1 U11302 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput58), .ZN(n10263) );
  NAND4_X1 U11303 ( .A1(n10266), .A2(n10265), .A3(n10264), .A4(n10263), .ZN(
        n10267) );
  NOR3_X1 U11304 ( .A1(n10269), .A2(n10268), .A3(n10267), .ZN(n10284) );
  AOI22_X1 U11305 ( .A1(n10272), .A2(keyinput57), .B1(keyinput33), .B2(n10271), 
        .ZN(n10270) );
  OAI221_X1 U11306 ( .B1(n10272), .B2(keyinput57), .C1(n10271), .C2(keyinput33), .A(n10270), .ZN(n10282) );
  AOI22_X1 U11307 ( .A1(n10275), .A2(keyinput37), .B1(n10274), .B2(keyinput31), 
        .ZN(n10273) );
  OAI221_X1 U11308 ( .B1(n10275), .B2(keyinput37), .C1(n10274), .C2(keyinput31), .A(n10273), .ZN(n10281) );
  XNOR2_X1 U11309 ( .A(P1_REG3_REG_20__SCAN_IN), .B(keyinput34), .ZN(n10279)
         );
  XNOR2_X1 U11310 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput32), .ZN(n10278) );
  XNOR2_X1 U11311 ( .A(P1_B_REG_SCAN_IN), .B(keyinput54), .ZN(n10277) );
  XNOR2_X1 U11312 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput62), .ZN(n10276)
         );
  NAND4_X1 U11313 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10280) );
  NOR3_X1 U11314 ( .A1(n10282), .A2(n10281), .A3(n10280), .ZN(n10283) );
  NAND4_X1 U11315 ( .A1(n10286), .A2(n10285), .A3(n10284), .A4(n10283), .ZN(
        n10287) );
  AOI211_X1 U11316 ( .C1(n10290), .C2(n10289), .A(n10288), .B(n10287), .ZN(
        n10294) );
  AOI22_X1 U11317 ( .A1(n10292), .A2(P2_REG0_REG_6__SCAN_IN), .B1(n10291), 
        .B2(n5734), .ZN(n10293) );
  XNOR2_X1 U11318 ( .A(n10294), .B(n10293), .ZN(P2_U3408) );
  XNOR2_X1 U11319 ( .A(n10296), .B(n10295), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11320 ( .A(n10298), .B(n10297), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11321 ( .A(n10300), .B(n10299), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11322 ( .A(n10302), .B(n10301), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11323 ( .A(n10304), .B(n10303), .ZN(ADD_1068_U48) );
  XOR2_X1 U11324 ( .A(n10306), .B(n10305), .Z(ADD_1068_U54) );
  XOR2_X1 U11325 ( .A(n10308), .B(n10307), .Z(ADD_1068_U53) );
  XNOR2_X1 U11326 ( .A(n10310), .B(n10309), .ZN(ADD_1068_U52) );
  NAND4_X1 U4862 ( .A1(n6367), .A2(n6366), .A3(n6365), .A4(n6364), .ZN(n7131)
         );
  NAND2_X1 U6351 ( .A1(n6009), .A2(n4379), .ZN(n10004) );
  CLKBUF_X1 U4825 ( .A(n8277), .Z(n4312) );
  CLKBUF_X1 U4847 ( .A(n5212), .Z(n5758) );
  CLKBUF_X1 U4848 ( .A(n5079), .Z(n5581) );
  CLKBUF_X3 U4863 ( .A(n6071), .Z(n6080) );
  CLKBUF_X1 U4972 ( .A(n5054), .Z(n5759) );
  XNOR2_X1 U5063 ( .A(n5013), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5015) );
  CLKBUF_X1 U6297 ( .A(n5600), .Z(n8609) );
endmodule

