

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9689, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349;

  INV_X1 U11133 ( .A(n18538), .ZN(n18216) );
  NAND2_X1 U11134 ( .A1(n10307), .A2(n9997), .ZN(n16172) );
  INV_X2 U11135 ( .A(n16808), .ZN(n13116) );
  NAND2_X1 U11136 ( .A1(n13695), .A2(n13255), .ZN(n13637) );
  INV_X1 U11137 ( .A(n15162), .ZN(n15287) );
  AND2_X2 U11138 ( .A1(n11140), .A2(n20101), .ZN(n11170) );
  CLKBUF_X2 U11140 ( .A(n12177), .Z(n17859) );
  CLKBUF_X2 U11141 ( .A(n10479), .Z(n14271) );
  CLKBUF_X2 U11142 ( .A(n12175), .Z(n17752) );
  AND2_X1 U11143 ( .A1(n10585), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10643) );
  CLKBUF_X2 U11144 ( .A(n12086), .Z(n17844) );
  CLKBUF_X2 U11145 ( .A(n14948), .Z(n15081) );
  INV_X2 U11146 ( .A(n11699), .ZN(n11753) );
  OR2_X1 U11147 ( .A1(n10573), .A2(n13387), .ZN(n11699) );
  CLKBUF_X2 U11148 ( .A(n12086), .Z(n9696) );
  INV_X1 U11149 ( .A(n11703), .ZN(n11748) );
  INV_X1 U11150 ( .A(n10670), .ZN(n11700) );
  CLKBUF_X2 U11151 ( .A(n14908), .Z(n15086) );
  NAND2_X1 U11152 ( .A1(n12765), .A2(n12978), .ZN(n13103) );
  INV_X1 U11153 ( .A(n9754), .ZN(n17879) );
  CLKBUF_X2 U11154 ( .A(n12095), .Z(n9698) );
  NOR2_X2 U11155 ( .A1(n12045), .A2(n19355), .ZN(n12105) );
  BUF_X1 U11156 ( .A(n15015), .Z(n15072) );
  BUF_X2 U11157 ( .A(n15074), .Z(n9694) );
  INV_X2 U11158 ( .A(n10483), .ZN(n10466) );
  INV_X1 U11159 ( .A(n12590), .ZN(n12780) );
  AND2_X1 U11161 ( .A1(n12440), .A2(n12869), .ZN(n14947) );
  AND2_X4 U11162 ( .A1(n12869), .A2(n14740), .ZN(n12560) );
  AND2_X2 U11163 ( .A1(n12442), .A2(n12868), .ZN(n15053) );
  INV_X2 U11164 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12777) );
  CLKBUF_X1 U11165 ( .A(n19084), .Z(n9689) );
  NOR2_X1 U11166 ( .A1(n19367), .A2(n19025), .ZN(n19084) );
  AND2_X1 U11168 ( .A1(n11768), .A2(n10578), .ZN(n11722) );
  INV_X1 U11169 ( .A(n15147), .ZN(n12765) );
  AND2_X1 U11170 ( .A1(n12440), .A2(n12869), .ZN(n9703) );
  NAND2_X1 U11171 ( .A1(n9943), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15214) );
  INV_X1 U11172 ( .A(n19656), .ZN(n16007) );
  AND2_X1 U11173 ( .A1(n9868), .A2(n9865), .ZN(n10489) );
  NOR2_X1 U11174 ( .A1(n18423), .A2(n18463), .ZN(n18440) );
  NAND2_X1 U11175 ( .A1(n19522), .A2(n19515), .ZN(n17603) );
  NAND2_X1 U11176 ( .A1(n12764), .A2(n13832), .ZN(n16636) );
  NOR2_X1 U11177 ( .A1(n16998), .A2(n17090), .ZN(n16997) );
  NOR2_X1 U11178 ( .A1(n18929), .A2(n18909), .ZN(n12300) );
  NOR2_X2 U11179 ( .A1(n17116), .A2(n12122), .ZN(n18463) );
  NAND2_X2 U11180 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19355) );
  INV_X1 U11181 ( .A(n13587), .ZN(n12764) );
  OAI21_X1 U11182 ( .B1(n16282), .B2(n16281), .A(n16236), .ZN(n16275) );
  NOR2_X1 U11183 ( .A1(n18334), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18333) );
  INV_X1 U11184 ( .A(n20604), .ZN(n20583) );
  AOI211_X1 U11186 ( .C1(n16441), .C2(n16440), .A(n16439), .B(n16438), .ZN(
        n16442) );
  INV_X2 U11187 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10346) );
  NOR2_X1 U11188 ( .A1(n18201), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16658) );
  NAND2_X2 U11189 ( .A1(n10000), .A2(n12880), .ZN(n13085) );
  INV_X4 U11190 ( .A(n9699), .ZN(n14265) );
  NAND2_X4 U11193 ( .A1(n10282), .A2(n10280), .ZN(n10474) );
  AND2_X2 U11194 ( .A1(n11595), .A2(n10541), .ZN(n9747) );
  AND2_X2 U11195 ( .A1(n10791), .A2(n10109), .ZN(n10845) );
  INV_X1 U11196 ( .A(n15162), .ZN(n9691) );
  AND2_X2 U11197 ( .A1(n13832), .A2(n13587), .ZN(n15162) );
  INV_X4 U11198 ( .A(n9746), .ZN(n16556) );
  BUF_X2 U11199 ( .A(n19699), .Z(n9706) );
  AND2_X2 U11200 ( .A1(n10578), .A2(n10346), .ZN(n9692) );
  XNOR2_X2 U11201 ( .A(n13809), .B(n13852), .ZN(n13808) );
  NAND2_X2 U11202 ( .A1(n13453), .A2(n13452), .ZN(n13809) );
  OR2_X2 U11205 ( .A1(n12041), .A2(n19355), .ZN(n9754) );
  NOR2_X4 U11206 ( .A1(n19355), .A2(n12044), .ZN(n12216) );
  XNOR2_X2 U11207 ( .A(n10839), .B(n11408), .ZN(n14037) );
  NAND2_X2 U11208 ( .A1(n9842), .A2(n14286), .ZN(n10839) );
  INV_X1 U11209 ( .A(n17877), .ZN(n9695) );
  INV_X1 U11210 ( .A(n19905), .ZN(n10400) );
  NAND2_X4 U11211 ( .A1(n10257), .A2(n10256), .ZN(n19905) );
  NOR2_X1 U11212 ( .A1(n12043), .A2(n12044), .ZN(n12086) );
  CLKBUF_X3 U11213 ( .A(n12095), .Z(n9697) );
  OR2_X1 U11214 ( .A1(n10266), .A2(n10268), .ZN(n10260) );
  XNOR2_X1 U11215 ( .A(n15249), .B(n15248), .ZN(n15534) );
  NOR2_X1 U11216 ( .A1(n15214), .A2(n10015), .ZN(n15216) );
  OR2_X1 U11217 ( .A1(n15214), .A2(n10020), .ZN(n15215) );
  NAND2_X1 U11218 ( .A1(n14436), .A2(n14435), .ZN(n9850) );
  NAND2_X1 U11219 ( .A1(n10085), .A2(n12162), .ZN(n18218) );
  OAI21_X2 U11220 ( .B1(n9876), .B2(n13484), .A(n10044), .ZN(n13670) );
  NAND2_X1 U11221 ( .A1(n11469), .A2(n10789), .ZN(n11457) );
  NAND2_X1 U11222 ( .A1(n9872), .A2(n13663), .ZN(n13662) );
  NAND3_X1 U11223 ( .A1(n9844), .A2(n10661), .A3(n9993), .ZN(n11454) );
  OR2_X1 U11224 ( .A1(n14400), .A2(n10318), .ZN(n14533) );
  NAND2_X1 U11225 ( .A1(n13254), .A2(n9934), .ZN(n13539) );
  INV_X1 U11226 ( .A(n10557), .ZN(n10555) );
  OR2_X2 U11227 ( .A1(n10565), .A2(n10564), .ZN(n10773) );
  OR2_X2 U11228 ( .A1(n10561), .A2(n10562), .ZN(n10767) );
  OAI21_X2 U11229 ( .B1(n12991), .B2(n12992), .A(n11592), .ZN(n13216) );
  NAND2_X1 U11230 ( .A1(n10009), .A2(n10007), .ZN(n13163) );
  BUF_X1 U11231 ( .A(n10545), .Z(n19869) );
  INV_X2 U11232 ( .A(n18601), .ZN(n19320) );
  NOR2_X1 U11233 ( .A1(n18488), .A2(n18808), .ZN(n18487) );
  AND3_X1 U11234 ( .A1(n10488), .A2(n10489), .A3(n10487), .ZN(n10246) );
  NOR2_X1 U11235 ( .A1(n11983), .A2(n16188), .ZN(n11982) );
  NAND2_X1 U11236 ( .A1(n9848), .A2(n9845), .ZN(n10522) );
  NAND2_X2 U11237 ( .A1(n11026), .A2(n10470), .ZN(n10483) );
  INV_X2 U11238 ( .A(n10474), .ZN(n10993) );
  INV_X1 U11239 ( .A(n11376), .ZN(n10218) );
  NOR2_X4 U11240 ( .A1(n19905), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11143) );
  AND2_X1 U11241 ( .A1(n9699), .A2(n13429), .ZN(n12019) );
  INV_X2 U11242 ( .A(n19896), .ZN(n12967) );
  CLKBUF_X2 U11243 ( .A(n12554), .Z(n15107) );
  BUF_X2 U11244 ( .A(n12092), .Z(n17855) );
  CLKBUF_X2 U11245 ( .A(n14947), .Z(n12885) );
  BUF_X1 U11246 ( .A(n12573), .Z(n9707) );
  CLKBUF_X2 U11247 ( .A(n12092), .Z(n17874) );
  BUF_X2 U11248 ( .A(n12573), .Z(n15082) );
  CLKBUF_X2 U11249 ( .A(n15084), .Z(n14991) );
  BUF_X2 U11250 ( .A(n13700), .Z(n14990) );
  NOR2_X2 U11251 ( .A1(n12042), .A2(n17603), .ZN(n12091) );
  AND2_X1 U11252 ( .A1(n12441), .A2(n12435), .ZN(n12573) );
  AND2_X2 U11253 ( .A1(n10052), .A2(n10346), .ZN(n10585) );
  NOR2_X4 U11254 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12869) );
  AND2_X1 U11256 ( .A1(n11549), .A2(n11548), .ZN(n10097) );
  OAI21_X1 U11257 ( .B1(n15385), .B2(n15373), .A(n15372), .ZN(n15681) );
  NAND2_X1 U11258 ( .A1(n12396), .A2(n10249), .ZN(n10248) );
  AND2_X1 U11259 ( .A1(n9982), .A2(n9980), .ZN(n12396) );
  NAND2_X1 U11260 ( .A1(n15397), .A2(n15399), .ZN(n15569) );
  OAI21_X1 U11261 ( .B1(n15103), .B2(n15104), .A(n15249), .ZN(n15624) );
  OR2_X2 U11262 ( .A1(n15414), .A2(n15398), .ZN(n15397) );
  AOI21_X1 U11263 ( .B1(n15300), .B2(n15299), .A(n15103), .ZN(n15635) );
  INV_X1 U11264 ( .A(n9897), .ZN(n15683) );
  NOR2_X1 U11265 ( .A1(n16275), .A2(n16237), .ZN(n16250) );
  AOI21_X1 U11266 ( .B1(n17132), .B2(n18464), .A(n10081), .ZN(n17136) );
  XNOR2_X1 U11267 ( .A(n9859), .B(n9858), .ZN(n16038) );
  XNOR2_X1 U11268 ( .A(n10082), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17132) );
  NAND2_X1 U11269 ( .A1(n16227), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16224) );
  OR2_X1 U11270 ( .A1(n16466), .A2(n17055), .ZN(n16998) );
  NOR2_X1 U11271 ( .A1(n11547), .A2(n11546), .ZN(n11548) );
  OAI22_X1 U11272 ( .A1(n16229), .A2(n10056), .B1(n10058), .B2(n16231), .ZN(
        n16291) );
  NOR2_X1 U11273 ( .A1(n15698), .A2(n15211), .ZN(n15691) );
  OAI22_X1 U11274 ( .A1(n16483), .A2(n10077), .B1(n16994), .B2(n10075), .ZN(
        n16989) );
  XNOR2_X1 U11275 ( .A(n12387), .B(n11135), .ZN(n15265) );
  NAND2_X1 U11276 ( .A1(n16047), .A2(n16046), .ZN(n16045) );
  NAND2_X1 U11277 ( .A1(n11476), .A2(n11475), .ZN(n14431) );
  CLKBUF_X1 U11278 ( .A(n14594), .Z(n14450) );
  NAND2_X1 U11279 ( .A1(n9944), .A2(n18205), .ZN(n18201) );
  NAND2_X1 U11280 ( .A1(n9945), .A2(n18218), .ZN(n9944) );
  AND3_X1 U11281 ( .A1(n15202), .A2(n15201), .A3(n15195), .ZN(n10006) );
  AND2_X1 U11282 ( .A1(n12161), .A2(n10086), .ZN(n10085) );
  AND2_X1 U11283 ( .A1(n18230), .A2(n10088), .ZN(n9945) );
  NOR2_X2 U11284 ( .A1(n15994), .A2(n15978), .ZN(n15979) );
  AOI21_X1 U11285 ( .B1(n10275), .B2(n10005), .A(n15209), .ZN(n10004) );
  XNOR2_X1 U11286 ( .A(n10165), .B(n10164), .ZN(n15484) );
  OAI21_X1 U11287 ( .B1(n10273), .B2(n14405), .A(n16761), .ZN(n10272) );
  XNOR2_X1 U11288 ( .A(n11477), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14433) );
  NAND2_X1 U11289 ( .A1(n11458), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11459) );
  AND2_X1 U11290 ( .A1(n15892), .A2(n15199), .ZN(n15756) );
  NAND2_X1 U11291 ( .A1(n10710), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13348) );
  NOR2_X1 U11292 ( .A1(n16103), .A2(n16102), .ZN(n15939) );
  NAND2_X1 U11293 ( .A1(n9979), .A2(n14505), .ZN(n10710) );
  NAND2_X1 U11294 ( .A1(n13476), .A2(n13468), .ZN(n13504) );
  INV_X1 U11295 ( .A(n15193), .ZN(n15209) );
  AOI21_X1 U11296 ( .B1(n14420), .B2(n14780), .A(n14109), .ZN(n14110) );
  NAND2_X1 U11297 ( .A1(n13709), .A2(n14101), .ZN(n13959) );
  XNOR2_X1 U11298 ( .A(n14533), .B(n14106), .ZN(n14420) );
  OR2_X1 U11299 ( .A1(n15997), .A2(n15981), .ZN(n15983) );
  NAND2_X2 U11300 ( .A1(n14533), .A2(n14532), .ZN(n9714) );
  AOI21_X1 U11301 ( .B1(n13812), .B2(n14780), .A(n13622), .ZN(n13624) );
  OR2_X1 U11302 ( .A1(n17130), .A2(n17131), .ZN(n10081) );
  NAND2_X1 U11303 ( .A1(n13289), .A2(n13295), .ZN(n13294) );
  AND2_X1 U11304 ( .A1(n10835), .A2(n10834), .ZN(n11470) );
  NAND2_X1 U11305 ( .A1(n9906), .A2(n9905), .ZN(n14400) );
  INV_X1 U11306 ( .A(n13254), .ZN(n9906) );
  NAND2_X1 U11307 ( .A1(n13167), .A2(n13166), .ZN(n13451) );
  NAND2_X1 U11308 ( .A1(n13172), .A2(n13146), .ZN(n13540) );
  AOI21_X1 U11309 ( .B1(n18296), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n19265), .ZN(n18388) );
  AND2_X1 U11310 ( .A1(n13320), .A2(n13319), .ZN(n13322) );
  NOR2_X1 U11311 ( .A1(n13640), .A2(n13694), .ZN(n9905) );
  INV_X1 U11312 ( .A(n13640), .ZN(n13253) );
  NAND2_X1 U11313 ( .A1(n10555), .A2(n10563), .ZN(n20205) );
  AND2_X1 U11314 ( .A1(n13252), .A2(n13251), .ZN(n13640) );
  CLKBUF_X1 U11315 ( .A(n10774), .Z(n13341) );
  NAND2_X1 U11316 ( .A1(n18462), .A2(n18463), .ZN(n18461) );
  OAI22_X1 U11317 ( .A1(n20257), .A2(n11803), .B1(n10779), .B2(n11217), .ZN(
        n10613) );
  NAND2_X1 U11318 ( .A1(n10555), .A2(n10546), .ZN(n20162) );
  NAND2_X1 U11319 ( .A1(n10014), .A2(n12910), .ZN(n13721) );
  INV_X1 U11320 ( .A(n13488), .ZN(n11057) );
  NAND2_X1 U11321 ( .A1(n9747), .A2(n10546), .ZN(n10779) );
  NAND2_X1 U11322 ( .A1(n9747), .A2(n10550), .ZN(n20257) );
  INV_X1 U11323 ( .A(n18547), .ZN(n18560) );
  INV_X1 U11324 ( .A(n18554), .ZN(n18526) );
  AND2_X1 U11325 ( .A1(n14304), .A2(n10221), .ZN(n16472) );
  OAI21_X2 U11326 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19534), .A(n17260), 
        .ZN(n18554) );
  OAI22_X1 U11327 ( .A1(n17390), .A2(n10175), .B1(n17547), .B2(n17381), .ZN(
        n17379) );
  NAND2_X1 U11328 ( .A1(n11191), .A2(n11190), .ZN(n14304) );
  INV_X1 U11329 ( .A(n10564), .ZN(n10546) );
  AND2_X1 U11330 ( .A1(n10202), .A2(n13174), .ZN(n10201) );
  NOR2_X1 U11331 ( .A1(n19359), .A2(n18060), .ZN(n18068) );
  AND2_X1 U11332 ( .A1(n10205), .A2(n12791), .ZN(n10200) );
  NOR3_X2 U11333 ( .A1(n10891), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n10116), .ZN(
        n10884) );
  AND2_X1 U11334 ( .A1(n11056), .A2(n11061), .ZN(n10130) );
  NOR2_X2 U11335 ( .A1(n14335), .A2(n20074), .ZN(n14253) );
  NAND2_X1 U11336 ( .A1(n19539), .A2(n18783), .ZN(n18601) );
  NOR2_X2 U11337 ( .A1(n19780), .A2(n20074), .ZN(n13231) );
  OAI21_X1 U11338 ( .B1(n12793), .B2(n12434), .A(n12798), .ZN(n13174) );
  OAI21_X2 U11339 ( .B1(n15264), .B2(n11574), .A(n11573), .ZN(n16533) );
  NAND2_X1 U11340 ( .A1(n10525), .A2(n9851), .ZN(n9882) );
  NOR2_X1 U11341 ( .A1(n13758), .A2(n13757), .ZN(n16854) );
  XNOR2_X1 U11342 ( .A(n11048), .B(n11049), .ZN(n11047) );
  INV_X2 U11343 ( .A(n19345), .ZN(n19358) );
  NOR2_X1 U11344 ( .A1(n12267), .A2(n18494), .ZN(n12269) );
  OR2_X1 U11345 ( .A1(n10511), .A2(n10513), .ZN(n10514) );
  AND2_X1 U11346 ( .A1(n10532), .A2(n10531), .ZN(n11049) );
  NAND2_X1 U11347 ( .A1(n10523), .A2(n10524), .ZN(n9881) );
  NOR2_X1 U11348 ( .A1(n18496), .A2(n18495), .ZN(n18494) );
  NAND2_X1 U11349 ( .A1(n10518), .A2(n10517), .ZN(n11582) );
  INV_X2 U11350 ( .A(n17921), .ZN(n17916) );
  AND2_X1 U11351 ( .A1(n9763), .A2(n10473), .ZN(n10538) );
  OAI21_X1 U11352 ( .B1(n10516), .B2(n10494), .A(n10493), .ZN(n10539) );
  CLKBUF_X3 U11353 ( .A(n11110), .Z(n11535) );
  AND2_X1 U11354 ( .A1(n12774), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12790) );
  AOI21_X1 U11355 ( .B1(n12965), .B2(n11166), .A(n11167), .ZN(n11174) );
  OR2_X1 U11356 ( .A1(n10854), .A2(n11966), .ZN(n10945) );
  AND3_X1 U11357 ( .A1(n10510), .A2(n10509), .A3(n10508), .ZN(n10512) );
  NOR2_X1 U11358 ( .A1(n12265), .A2(n18507), .ZN(n18496) );
  CLKBUF_X3 U11359 ( .A(n10522), .Z(n11110) );
  AND2_X1 U11360 ( .A1(n10536), .A2(n10500), .ZN(n10501) );
  NAND2_X1 U11361 ( .A1(n11020), .A2(n10486), .ZN(n11100) );
  NOR2_X1 U11362 ( .A1(n18044), .A2(n12123), .ZN(n12144) );
  NOR2_X1 U11363 ( .A1(n13403), .A2(n10483), .ZN(n13384) );
  INV_X2 U11364 ( .A(n18178), .ZN(n18171) );
  OAI211_X1 U11365 ( .C1(n16636), .C2(n13079), .A(n13103), .B(n12858), .ZN(
        n12782) );
  XNOR2_X1 U11366 ( .A(n12124), .B(n18047), .ZN(n12126) );
  AND2_X1 U11367 ( .A1(n15218), .A2(n12818), .ZN(n12857) );
  INV_X1 U11368 ( .A(n12818), .ZN(n10003) );
  AND2_X1 U11369 ( .A1(n10080), .A2(n12252), .ZN(n12124) );
  AND2_X1 U11370 ( .A1(n10467), .A2(n10466), .ZN(n10469) );
  OAI21_X1 U11371 ( .B1(n12853), .B2(n13097), .A(n9895), .ZN(n12599) );
  OR2_X1 U11372 ( .A1(n12758), .A2(n12760), .ZN(n12815) );
  INV_X1 U11373 ( .A(n16636), .ZN(n14536) );
  INV_X1 U11374 ( .A(n12853), .ZN(n12978) );
  NAND2_X1 U11375 ( .A1(n13079), .A2(n12554), .ZN(n12853) );
  INV_X1 U11376 ( .A(n13558), .ZN(n13097) );
  AND3_X1 U11377 ( .A1(n13547), .A2(n13832), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n13971) );
  INV_X1 U11378 ( .A(n12591), .ZN(n13079) );
  INV_X1 U11379 ( .A(n13832), .ZN(n12975) );
  CLKBUF_X1 U11380 ( .A(n12591), .Z(n13547) );
  OAI21_X1 U11381 ( .B1(n13564), .B2(n12591), .A(n13577), .ZN(n12597) );
  NAND3_X1 U11382 ( .A1(n12247), .A2(n12246), .A3(n12245), .ZN(n17562) );
  INV_X1 U11383 ( .A(n12713), .ZN(n10988) );
  INV_X1 U11384 ( .A(n12249), .ZN(n18056) );
  NAND3_X1 U11385 ( .A1(n12186), .A2(n12185), .A3(n12184), .ZN(n12326) );
  AND3_X1 U11386 ( .A1(n10335), .A2(n10659), .A3(n9760), .ZN(n11445) );
  NAND2_X1 U11388 ( .A1(n10338), .A2(n10319), .ZN(n18066) );
  OR2_X2 U11389 ( .A1(n12589), .A2(n12588), .ZN(n13571) );
  NAND2_X1 U11390 ( .A1(n9711), .A2(n13429), .ZN(n10694) );
  NAND2_X1 U11391 ( .A1(n9930), .A2(n9759), .ZN(n12591) );
  NAND2_X1 U11392 ( .A1(n10456), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10280) );
  INV_X4 U11393 ( .A(n10485), .ZN(n9699) );
  AND4_X1 U11394 ( .A1(n12453), .A2(n12452), .A3(n12451), .A4(n12450), .ZN(
        n12464) );
  AND4_X1 U11395 ( .A1(n12577), .A2(n12576), .A3(n12575), .A4(n12574), .ZN(
        n12578) );
  OR2_X1 U11396 ( .A1(n12496), .A2(n12495), .ZN(n12554) );
  NAND3_X1 U11397 ( .A1(n10420), .A2(n10419), .A3(n13387), .ZN(n10421) );
  AND4_X1 U11398 ( .A1(n12473), .A2(n12472), .A3(n12471), .A4(n12470), .ZN(
        n12484) );
  AND4_X1 U11399 ( .A1(n12457), .A2(n12456), .A3(n12455), .A4(n12454), .ZN(
        n12463) );
  AND4_X1 U11400 ( .A1(n12477), .A2(n12476), .A3(n12475), .A4(n12474), .ZN(
        n12483) );
  INV_X2 U11401 ( .A(U214), .ZN(n17212) );
  AND4_X1 U11402 ( .A1(n10418), .A2(n10417), .A3(n10416), .A4(n10415), .ZN(
        n10419) );
  NAND2_X1 U11403 ( .A1(n10191), .A2(n10190), .ZN(n18349) );
  AND2_X2 U11404 ( .A1(n11936), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11740) );
  AND2_X1 U11405 ( .A1(n10354), .A2(n10353), .ZN(n10359) );
  CLKBUF_X2 U11406 ( .A(n12573), .Z(n15040) );
  AND4_X1 U11407 ( .A1(n12469), .A2(n12468), .A3(n12467), .A4(n12466), .ZN(
        n12485) );
  AND2_X2 U11408 ( .A1(n11932), .A2(n13387), .ZN(n11747) );
  AND4_X1 U11409 ( .A1(n12481), .A2(n12480), .A3(n12479), .A4(n12478), .ZN(
        n12482) );
  INV_X2 U11410 ( .A(n18102), .ZN(n18119) );
  INV_X2 U11411 ( .A(n17245), .ZN(U215) );
  CLKBUF_X2 U11412 ( .A(n12573), .Z(n9708) );
  AND2_X1 U11413 ( .A1(n10348), .A2(n10347), .ZN(n10349) );
  AND2_X2 U11414 ( .A1(n12974), .A2(n15926), .ZN(n16764) );
  NAND2_X2 U11415 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20423), .ZN(n20445) );
  CLKBUF_X1 U11416 ( .A(n12694), .Z(n13223) );
  NAND2_X2 U11417 ( .A1(n20423), .A2(n20395), .ZN(n20444) );
  BUF_X2 U11418 ( .A(n12216), .Z(n17860) );
  NAND2_X2 U11419 ( .A1(n19552), .A2(n17110), .ZN(n18833) );
  NAND2_X2 U11420 ( .A1(n19484), .A2(n19421), .ZN(n19471) );
  INV_X2 U11421 ( .A(n10723), .ZN(n11760) );
  CLKBUF_X3 U11422 ( .A(n10591), .Z(n11932) );
  INV_X1 U11423 ( .A(n17877), .ZN(n12130) );
  INV_X2 U11424 ( .A(n17247), .ZN(n17249) );
  BUF_X2 U11425 ( .A(n15053), .Z(n15073) );
  AND2_X2 U11426 ( .A1(n12440), .A2(n12870), .ZN(n9710) );
  BUF_X2 U11427 ( .A(n12583), .Z(n14929) );
  NOR2_X1 U11428 ( .A1(n10159), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12435) );
  AND2_X2 U11429 ( .A1(n12440), .A2(n12439), .ZN(n12892) );
  AND2_X2 U11430 ( .A1(n12439), .A2(n14740), .ZN(n12555) );
  NOR2_X2 U11431 ( .A1(n9918), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12441) );
  CLKBUF_X1 U11432 ( .A(n20866), .Z(n15926) );
  NAND3_X1 U11433 ( .A1(n19522), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n16586), .ZN(n17877) );
  NAND2_X1 U11434 ( .A1(n12306), .A2(n19499), .ZN(n12042) );
  NAND2_X1 U11435 ( .A1(n19522), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12043) );
  AND2_X1 U11436 ( .A1(n13533), .A2(n12870), .ZN(n12583) );
  AND2_X1 U11437 ( .A1(n13262), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12439) );
  NOR2_X1 U11438 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12442) );
  CLKBUF_X1 U11439 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n19350) );
  INV_X1 U11440 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19499) );
  AND2_X1 U11441 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16586) );
  INV_X1 U11442 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19515) );
  NOR2_X2 U11443 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13533) );
  AND2_X1 U11444 ( .A1(n12870), .A2(n14740), .ZN(n9701) );
  AND2_X1 U11445 ( .A1(n12870), .A2(n14740), .ZN(n9702) );
  AND2_X2 U11446 ( .A1(n11022), .A2(n10504), .ZN(n11403) );
  OR2_X1 U11447 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  BUF_X4 U11448 ( .A(n15147), .Z(n15129) );
  NAND2_X2 U11449 ( .A1(n12967), .A2(n9704), .ZN(n11149) );
  NAND2_X1 U11450 ( .A1(n11466), .A2(n11189), .ZN(n9842) );
  MUX2_X1 U11451 ( .A(n10362), .B(n10361), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n9704) );
  XNOR2_X2 U11452 ( .A(n14396), .B(n13853), .ZN(n14395) );
  AND2_X2 U11453 ( .A1(n10052), .A2(n10346), .ZN(n9705) );
  OAI211_X2 U11454 ( .C1(n11467), .C2(n11465), .A(n11464), .B(n11463), .ZN(
        n14035) );
  AOI21_X2 U11455 ( .B1(n15386), .B2(n15397), .A(n15385), .ZN(n15688) );
  NAND2_X2 U11456 ( .A1(n12543), .A2(n12542), .ZN(n16614) );
  XNOR2_X1 U11457 ( .A(n10543), .B(n10542), .ZN(n19699) );
  OAI21_X2 U11458 ( .B1(n12792), .B2(n9712), .A(n12771), .ZN(n12775) );
  AND2_X1 U11459 ( .A1(n12440), .A2(n12870), .ZN(n9709) );
  MUX2_X1 U11460 ( .A(n10433), .B(n10432), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n9711) );
  NAND2_X1 U11461 ( .A1(n14533), .A2(n14532), .ZN(n9713) );
  NAND2_X1 U11462 ( .A1(n14533), .A2(n14532), .ZN(n15193) );
  AND2_X1 U11463 ( .A1(n11895), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11754) );
  AND2_X1 U11464 ( .A1(n11895), .A2(n13387), .ZN(n11755) );
  INV_X1 U11465 ( .A(n9857), .ZN(n9856) );
  NAND2_X1 U11466 ( .A1(n9854), .A2(n9857), .ZN(n9853) );
  NAND2_X1 U11467 ( .A1(n9974), .A2(n10988), .ZN(n9868) );
  NAND2_X1 U11468 ( .A1(n9866), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9865) );
  NOR2_X1 U11469 ( .A1(n14659), .A2(n14658), .ZN(n16581) );
  OAI211_X1 U11470 ( .C1(n16582), .C2(n19349), .A(n19324), .B(n19540), .ZN(
        n16679) );
  NOR2_X1 U11471 ( .A1(n12853), .A2(n13832), .ZN(n12600) );
  INV_X1 U11472 ( .A(n9983), .ZN(n9980) );
  BUF_X1 U11473 ( .A(n15015), .Z(n14985) );
  INV_X1 U11474 ( .A(n14400), .ZN(n13709) );
  NOR2_X1 U11475 ( .A1(n12857), .A2(n9926), .ZN(n9925) );
  NOR2_X1 U11476 ( .A1(n12782), .A2(n9766), .ZN(n9924) );
  NOR2_X1 U11477 ( .A1(n13085), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10277) );
  AND3_X1 U11478 ( .A1(n9699), .A2(n10468), .A3(n19905), .ZN(n11140) );
  NAND2_X1 U11479 ( .A1(n10484), .A2(n10470), .ZN(n10423) );
  AOI21_X1 U11480 ( .B1(n10039), .B2(n10038), .A(n10037), .ZN(n12312) );
  AND2_X1 U11481 ( .A1(n19366), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10037) );
  INV_X1 U11482 ( .A(n12313), .ZN(n10038) );
  NAND2_X2 U11483 ( .A1(n13571), .A2(n13097), .ZN(n12818) );
  AND2_X1 U11484 ( .A1(n9804), .A2(n15311), .ZN(n10216) );
  INV_X1 U11485 ( .A(n15591), .ZN(n14817) );
  INV_X1 U11486 ( .A(n15146), .ZN(n15159) );
  AND2_X1 U11487 ( .A1(n16762), .A2(n16768), .ZN(n10270) );
  OR2_X1 U11488 ( .A1(n13170), .A2(n14401), .ZN(n10328) );
  NOR2_X1 U11489 ( .A1(n10013), .A2(n14401), .ZN(n10012) );
  INV_X1 U11490 ( .A(n12910), .ZN(n10013) );
  NOR2_X1 U11491 ( .A1(n12905), .A2(n9922), .ZN(n14531) );
  NAND2_X1 U11492 ( .A1(n13908), .A2(n9922), .ZN(n13252) );
  INV_X1 U11493 ( .A(n13971), .ZN(n14103) );
  AND3_X1 U11494 ( .A1(n10733), .A2(n10732), .A3(n10731), .ZN(n11456) );
  AND4_X1 U11495 ( .A1(n10717), .A2(n10716), .A3(n10715), .A4(n10714), .ZN(
        n10733) );
  AND4_X1 U11496 ( .A1(n10730), .A2(n10729), .A3(n10728), .A4(n10727), .ZN(
        n10731) );
  INV_X1 U11497 ( .A(n13503), .ZN(n10125) );
  NAND2_X1 U11498 ( .A1(n16178), .A2(n10321), .ZN(n11500) );
  INV_X1 U11499 ( .A(n10305), .ZN(n10304) );
  OAI21_X1 U11500 ( .B1(n14433), .B2(n10306), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U11501 ( .A1(n9849), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9848) );
  AND2_X1 U11502 ( .A1(n12620), .A2(n12967), .ZN(n11836) );
  NAND3_X1 U11503 ( .A1(n10482), .A2(n10496), .A3(n10471), .ZN(n10477) );
  INV_X1 U11504 ( .A(n18308), .ZN(n10176) );
  BUF_X1 U11505 ( .A(n12177), .Z(n17878) );
  OR2_X1 U11506 ( .A1(n12044), .A2(n17603), .ZN(n10339) );
  NAND2_X1 U11507 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12306), .ZN(
        n12044) );
  OR2_X1 U11508 ( .A1(n18333), .A2(n18463), .ZN(n9961) );
  NAND2_X1 U11509 ( .A1(n12764), .A2(n12975), .ZN(n15286) );
  AND2_X1 U11510 ( .A1(n13078), .A2(n13077), .ZN(n13117) );
  INV_X1 U11511 ( .A(n11889), .ZN(n9858) );
  OR2_X1 U11512 ( .A1(n16924), .A2(n11189), .ZN(n11503) );
  NOR2_X1 U11513 ( .A1(n10327), .A2(n10076), .ZN(n10075) );
  OR2_X1 U11514 ( .A1(n16994), .A2(n9723), .ZN(n10077) );
  NAND2_X1 U11515 ( .A1(n9850), .A2(n9990), .ZN(n9989) );
  NOR2_X1 U11516 ( .A1(n9723), .A2(n9991), .ZN(n9990) );
  INV_X1 U11517 ( .A(n10258), .ZN(n9991) );
  NAND2_X1 U11518 ( .A1(n19749), .A2(n20487), .ZN(n20041) );
  OR2_X1 U11519 ( .A1(n19749), .A2(n20487), .ZN(n20130) );
  OAI21_X1 U11520 ( .B1(n16681), .B2(n16680), .A(n16679), .ZN(n16682) );
  INV_X1 U11521 ( .A(n10042), .ZN(n16680) );
  NAND2_X1 U11522 ( .A1(n18463), .A2(n18588), .ZN(n12160) );
  OR2_X1 U11523 ( .A1(n18231), .A2(n18463), .ZN(n12161) );
  NAND2_X1 U11524 ( .A1(n10095), .A2(n11527), .ZN(n10094) );
  NAND2_X1 U11525 ( .A1(n10248), .A2(n10096), .ZN(n10095) );
  OR2_X1 U11526 ( .A1(n17454), .A2(n9784), .ZN(n17808) );
  OAI22_X1 U11527 ( .A1(n10547), .A2(n10767), .B1(n10779), .B2(n11271), .ZN(
        n10548) );
  AOI21_X1 U11528 ( .B1(n12516), .B2(n12433), .A(n12432), .ZN(n12529) );
  INV_X1 U11529 ( .A(n12554), .ZN(n12772) );
  NAND2_X1 U11530 ( .A1(n13172), .A2(n13171), .ZN(n13193) );
  OR2_X1 U11531 ( .A1(n13170), .A2(n13169), .ZN(n13171) );
  OR2_X1 U11532 ( .A1(n13096), .A2(n13095), .ZN(n13195) );
  INV_X1 U11533 ( .A(n16957), .ZN(n10291) );
  AND4_X1 U11534 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        n10758) );
  OR2_X1 U11535 ( .A1(n16020), .A2(n11189), .ZN(n10915) );
  INV_X1 U11536 ( .A(n10788), .ZN(n10053) );
  INV_X1 U11537 ( .A(n10479), .ZN(n10468) );
  NAND2_X1 U11538 ( .A1(n10505), .A2(n11022), .ZN(n9849) );
  INV_X1 U11539 ( .A(n10470), .ZN(n11416) );
  OAI21_X1 U11540 ( .B1(n13393), .B2(n11679), .A(n10302), .ZN(n10301) );
  NAND2_X1 U11541 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10302) );
  NAND2_X1 U11542 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n9917) );
  INV_X1 U11543 ( .A(n18041), .ZN(n12145) );
  NAND2_X1 U11544 ( .A1(n18056), .A2(n18066), .ZN(n12140) );
  NAND2_X1 U11545 ( .A1(n12595), .A2(n13097), .ZN(n9895) );
  NOR2_X1 U11546 ( .A1(n15505), .A2(n15455), .ZN(n10209) );
  NOR2_X1 U11547 ( .A1(n12761), .A2(n9922), .ZN(n15067) );
  NAND2_X1 U11548 ( .A1(n10214), .A2(n14640), .ZN(n10213) );
  INV_X1 U11549 ( .A(n15466), .ZN(n10214) );
  NAND2_X1 U11550 ( .A1(n13959), .A2(n14780), .ZN(n10206) );
  INV_X1 U11551 ( .A(n15101), .ZN(n14983) );
  INV_X1 U11552 ( .A(n14797), .ZN(n14780) );
  AND2_X1 U11553 ( .A1(n9821), .A2(n10174), .ZN(n10173) );
  INV_X1 U11554 ( .A(n15343), .ZN(n10174) );
  INV_X1 U11555 ( .A(n15430), .ZN(n10171) );
  AND2_X1 U11556 ( .A1(n15207), .A2(n9834), .ZN(n9935) );
  NAND2_X1 U11557 ( .A1(n10006), .A2(n15778), .ZN(n9936) );
  AND2_X1 U11558 ( .A1(n14412), .A2(n14411), .ZN(n14413) );
  NAND2_X1 U11559 ( .A1(n9898), .A2(n14403), .ZN(n14404) );
  NAND2_X1 U11560 ( .A1(n13959), .A2(n9899), .ZN(n9898) );
  NAND2_X1 U11561 ( .A1(n12765), .A2(n15162), .ZN(n15165) );
  NOR2_X1 U11562 ( .A1(n10001), .A2(n12818), .ZN(n12814) );
  NOR2_X1 U11563 ( .A1(n12777), .A2(n9922), .ZN(n9921) );
  OR2_X1 U11564 ( .A1(n12911), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U11565 ( .A1(n12555), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15059), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12576) );
  NOR2_X1 U11566 ( .A1(n9932), .A2(n9931), .ZN(n9930) );
  AND2_X1 U11567 ( .A1(n9762), .A2(n9886), .ZN(n9929) );
  OAI21_X1 U11568 ( .B1(n21033), .B2(n21290), .A(n21010), .ZN(n13546) );
  AOI21_X1 U11569 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20463), .A(
        n10713), .ZN(n10984) );
  NOR2_X1 U11570 ( .A1(n10965), .A2(n10955), .ZN(n10100) );
  NAND2_X1 U11571 ( .A1(n9748), .A2(n10945), .ZN(n10948) );
  INV_X1 U11572 ( .A(n10948), .ZN(n11525) );
  AND2_X1 U11573 ( .A1(n10925), .A2(n10112), .ZN(n10942) );
  NOR2_X1 U11574 ( .A1(n10113), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10112) );
  INV_X1 U11575 ( .A(n10114), .ZN(n10113) );
  NAND2_X1 U11576 ( .A1(n10942), .A2(n10941), .ZN(n10947) );
  OR2_X1 U11577 ( .A1(n10889), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10927) );
  INV_X1 U11578 ( .A(n10893), .ZN(n10118) );
  INV_X1 U11579 ( .A(n10875), .ZN(n10117) );
  NOR2_X1 U11580 ( .A1(n10902), .A2(n10108), .ZN(n10107) );
  NAND2_X1 U11581 ( .A1(n10900), .A2(n10867), .ZN(n10108) );
  AND2_X1 U11582 ( .A1(n13302), .A2(n10104), .ZN(n10103) );
  AND3_X1 U11583 ( .A1(n10599), .A2(n10598), .A3(n10597), .ZN(n11178) );
  AND4_X1 U11584 ( .A1(n10596), .A2(n10595), .A3(n10594), .A4(n10593), .ZN(
        n10597) );
  AND4_X1 U11585 ( .A1(n10590), .A2(n10589), .A3(n10588), .A4(n10587), .ZN(
        n10598) );
  NOR2_X1 U11586 ( .A1(n10640), .A2(n10639), .ZN(n11446) );
  INV_X1 U11587 ( .A(n11755), .ZN(n11726) );
  INV_X1 U11588 ( .A(n11754), .ZN(n11697) );
  NAND2_X1 U11589 ( .A1(n10244), .A2(n10243), .ZN(n10242) );
  INV_X1 U11590 ( .A(n11508), .ZN(n10243) );
  INV_X1 U11591 ( .A(n16090), .ZN(n10244) );
  NAND2_X1 U11592 ( .A1(n16109), .A2(n10234), .ZN(n10233) );
  INV_X1 U11593 ( .A(n15967), .ZN(n10234) );
  INV_X1 U11594 ( .A(n16152), .ZN(n10237) );
  NAND2_X1 U11595 ( .A1(n10297), .A2(n14082), .ZN(n10296) );
  INV_X1 U11596 ( .A(n14175), .ZN(n10297) );
  INV_X1 U11597 ( .A(n13352), .ZN(n10229) );
  NAND2_X1 U11598 ( .A1(n12840), .A2(n12839), .ZN(n11161) );
  NOR2_X1 U11599 ( .A1(n16992), .A2(n10158), .ZN(n10157) );
  INV_X1 U11600 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10158) );
  NOR2_X1 U11601 ( .A1(n14295), .A2(n10155), .ZN(n10154) );
  AND4_X1 U11602 ( .A1(n10652), .A2(n10651), .A3(n10650), .A4(n10649), .ZN(
        n10659) );
  OAI22_X1 U11603 ( .A1(n10959), .A2(n9985), .B1(n10958), .B2(n9984), .ZN(
        n9983) );
  NAND2_X1 U11604 ( .A1(n11499), .A2(n10952), .ZN(n9985) );
  NAND2_X1 U11605 ( .A1(n11499), .A2(n12405), .ZN(n9984) );
  NAND2_X1 U11606 ( .A1(n11500), .A2(n9986), .ZN(n9982) );
  NOR2_X1 U11607 ( .A1(n10959), .A2(n9987), .ZN(n9986) );
  INV_X1 U11608 ( .A(n11499), .ZN(n9987) );
  OR2_X1 U11609 ( .A1(n16929), .A2(n11189), .ZN(n10960) );
  NOR2_X1 U11610 ( .A1(n10922), .A2(n10921), .ZN(n10923) );
  INV_X1 U11611 ( .A(n14171), .ZN(n10123) );
  INV_X1 U11612 ( .A(n16300), .ZN(n10059) );
  AND2_X1 U11613 ( .A1(n14434), .A2(n10852), .ZN(n10258) );
  INV_X1 U11614 ( .A(n10794), .ZN(n9977) );
  AND2_X1 U11615 ( .A1(n10833), .A2(n10832), .ZN(n11185) );
  NOR2_X1 U11616 ( .A1(n10485), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10219) );
  INV_X1 U11617 ( .A(n13304), .ZN(n11061) );
  NAND2_X1 U11618 ( .A1(n10527), .A2(n10526), .ZN(n11048) );
  NOR2_X1 U11619 ( .A1(n10628), .A2(n10627), .ZN(n11447) );
  INV_X1 U11620 ( .A(n11574), .ZN(n11596) );
  NOR2_X1 U11621 ( .A1(n10470), .A2(n19880), .ZN(n10480) );
  OR2_X1 U11622 ( .A1(n12042), .A2(n19355), .ZN(n9746) );
  OR2_X1 U11623 ( .A1(n12046), .A2(n12042), .ZN(n12215) );
  NOR2_X1 U11624 ( .A1(n12046), .A2(n12044), .ZN(n12092) );
  NAND2_X1 U11625 ( .A1(n9972), .A2(n9971), .ZN(n16558) );
  INV_X1 U11626 ( .A(n12041), .ZN(n9972) );
  INV_X1 U11627 ( .A(n12043), .ZN(n9971) );
  NOR2_X1 U11628 ( .A1(n12271), .A2(n18487), .ZN(n12274) );
  INV_X1 U11629 ( .A(n12154), .ZN(n9964) );
  AND2_X1 U11630 ( .A1(n10090), .A2(n10324), .ZN(n10089) );
  NAND2_X1 U11631 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18472), .ZN(
        n12277) );
  NAND2_X1 U11632 ( .A1(n12124), .A2(n12125), .ZN(n12123) );
  INV_X1 U11633 ( .A(n10039), .ZN(n12320) );
  AOI21_X1 U11634 ( .B1(n12312), .B2(n12311), .A(n12310), .ZN(n12322) );
  NAND2_X1 U11635 ( .A1(n13328), .A2(n13326), .ZN(n13268) );
  INV_X1 U11636 ( .A(n15286), .ZN(n12779) );
  AND2_X1 U11637 ( .A1(n14046), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15245) );
  INV_X1 U11638 ( .A(n13616), .ZN(n15246) );
  INV_X1 U11639 ( .A(n15300), .ZN(n10215) );
  INV_X1 U11640 ( .A(n15207), .ZN(n10005) );
  AND2_X1 U11641 ( .A1(n15515), .A2(n9820), .ZN(n10210) );
  NAND2_X1 U11642 ( .A1(n13974), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13973) );
  NAND2_X1 U11643 ( .A1(n13618), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13688) );
  NAND2_X1 U11644 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13256) );
  AND2_X1 U11645 ( .A1(n15456), .A2(n9829), .ZN(n15402) );
  INV_X1 U11646 ( .A(n15400), .ZN(n10169) );
  NAND2_X1 U11647 ( .A1(n15456), .A2(n9815), .ZN(n15432) );
  NAND2_X1 U11648 ( .A1(n15456), .A2(n9816), .ZN(n15418) );
  NAND2_X1 U11649 ( .A1(n9936), .A2(n15207), .ZN(n15724) );
  NAND2_X1 U11650 ( .A1(n9714), .A2(n14538), .ZN(n14585) );
  AOI21_X1 U11651 ( .B1(n10012), .B2(n13138), .A(n12976), .ZN(n10010) );
  INV_X1 U11652 ( .A(n10012), .ZN(n10011) );
  NAND2_X1 U11653 ( .A1(n13085), .A2(n9999), .ZN(n12911) );
  OR2_X1 U11654 ( .A1(n10000), .A2(n12880), .ZN(n9999) );
  INV_X1 U11655 ( .A(n13539), .ZN(n13639) );
  NAND2_X1 U11656 ( .A1(n12790), .A2(n12789), .ZN(n12791) );
  INV_X1 U11657 ( .A(n12854), .ZN(n13519) );
  INV_X1 U11658 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20737) );
  INV_X1 U11659 ( .A(n13761), .ZN(n20694) );
  NOR2_X1 U11660 ( .A1(n13637), .A2(n13639), .ZN(n13865) );
  INV_X1 U11661 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20779) );
  NAND2_X1 U11662 ( .A1(n9922), .A2(n13546), .ZN(n14128) );
  AND4_X1 U11663 ( .A1(n12449), .A2(n12448), .A3(n12447), .A4(n12446), .ZN(
        n12465) );
  AOI21_X1 U11664 ( .B1(n9703), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A(n12461), .ZN(n12462) );
  NOR2_X1 U11665 ( .A1(n14547), .A2(n20694), .ZN(n14043) );
  NAND2_X1 U11666 ( .A1(n12540), .A2(n12539), .ZN(n12543) );
  NOR2_X1 U11667 ( .A1(n16898), .A2(n16899), .ZN(n16897) );
  NAND2_X1 U11668 ( .A1(n10884), .A2(n10885), .ZN(n10889) );
  NAND2_X1 U11669 ( .A1(n10927), .A2(n10945), .ZN(n10925) );
  AND2_X1 U11670 ( .A1(n9726), .A2(n10110), .ZN(n10109) );
  NAND2_X1 U11671 ( .A1(n11605), .A2(n10300), .ZN(n10299) );
  INV_X1 U11672 ( .A(n13478), .ZN(n10300) );
  NOR2_X1 U11673 ( .A1(n9852), .A2(n11889), .ZN(n16027) );
  INV_X1 U11674 ( .A(n11838), .ZN(n11839) );
  AND2_X1 U11675 ( .A1(n9795), .A2(n10222), .ZN(n10221) );
  INV_X1 U11676 ( .A(n16494), .ZN(n10222) );
  NAND2_X1 U11677 ( .A1(n10225), .A2(n10228), .ZN(n13490) );
  NAND2_X1 U11678 ( .A1(n13429), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12713) );
  OR2_X1 U11679 ( .A1(n13434), .A2(n12017), .ZN(n12629) );
  NOR2_X1 U11680 ( .A1(n10151), .A2(n10148), .ZN(n10146) );
  INV_X1 U11681 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10151) );
  NAND2_X1 U11682 ( .A1(n11996), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12005) );
  NAND2_X1 U11683 ( .A1(n11998), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12004) );
  NAND2_X1 U11684 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12001) );
  OR2_X1 U11685 ( .A1(n10310), .A2(n12406), .ZN(n10309) );
  OR2_X1 U11686 ( .A1(n16912), .A2(n11189), .ZN(n11505) );
  INV_X1 U11687 ( .A(n11503), .ZN(n11501) );
  AND2_X1 U11688 ( .A1(n16405), .A2(n11430), .ZN(n16374) );
  AOI21_X1 U11689 ( .B1(n16291), .B2(n16290), .A(n16234), .ZN(n16282) );
  AND3_X1 U11690 ( .A1(n11089), .A2(n11088), .A3(n11087), .ZN(n14083) );
  OR3_X1 U11691 ( .A1(n14328), .A2(n11189), .A3(n16459), .ZN(n16300) );
  NOR2_X1 U11692 ( .A1(n16228), .A2(n10064), .ZN(n10063) );
  AND2_X1 U11693 ( .A1(n10856), .A2(n16492), .ZN(n16484) );
  OR2_X1 U11694 ( .A1(n11478), .A2(n11189), .ZN(n11477) );
  AND3_X1 U11695 ( .A1(n11064), .A2(n11063), .A3(n11062), .ZN(n13128) );
  NAND2_X1 U11696 ( .A1(n13485), .A2(n13675), .ZN(n10044) );
  AND2_X1 U11697 ( .A1(n11454), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9877) );
  OR2_X1 U11698 ( .A1(n11536), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10493) );
  AND2_X1 U11699 ( .A1(n11041), .A2(n13124), .ZN(n11482) );
  XNOR2_X1 U11700 ( .A(n16533), .B(n11575), .ZN(n12962) );
  AND2_X1 U11701 ( .A1(n20466), .A2(n20478), .ZN(n20454) );
  NAND2_X1 U11702 ( .A1(n10372), .A2(n13387), .ZN(n10373) );
  NAND2_X1 U11703 ( .A1(n17095), .A2(n13220), .ZN(n20320) );
  NAND2_X1 U11704 ( .A1(n10457), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10257) );
  NAND2_X1 U11705 ( .A1(n10460), .A2(n13387), .ZN(n10256) );
  INV_X1 U11706 ( .A(n20320), .ZN(n20074) );
  NOR2_X1 U11707 ( .A1(n18904), .A2(n12282), .ZN(n12333) );
  NAND2_X1 U11708 ( .A1(n10186), .A2(n10182), .ZN(n10181) );
  INV_X1 U11709 ( .A(n17139), .ZN(n10182) );
  OR2_X1 U11710 ( .A1(n17301), .A2(n10183), .ZN(n10180) );
  OR2_X1 U11711 ( .A1(n18194), .A2(n17139), .ZN(n10183) );
  INV_X1 U11712 ( .A(n18257), .ZN(n10187) );
  NAND2_X1 U11713 ( .A1(n10176), .A2(n18297), .ZN(n10175) );
  NAND2_X1 U11714 ( .A1(n10177), .A2(n10176), .ZN(n10178) );
  INV_X1 U11715 ( .A(n17390), .ZN(n10177) );
  NOR2_X1 U11716 ( .A1(n18469), .A2(n18457), .ZN(n17504) );
  AOI211_X1 U11717 ( .C1(n12175), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n12244), .B(n12243), .ZN(n12245) );
  OR2_X1 U11718 ( .A1(n16581), .A2(n10043), .ZN(n10042) );
  AND2_X1 U11719 ( .A1(n14661), .A2(n14660), .ZN(n10043) );
  AND2_X1 U11720 ( .A1(n9698), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12096) );
  NOR2_X1 U11721 ( .A1(n9968), .A2(n9966), .ZN(n9965) );
  INV_X1 U11722 ( .A(n12131), .ZN(n9968) );
  NAND2_X1 U11723 ( .A1(n12093), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n9967) );
  INV_X1 U11724 ( .A(n18236), .ZN(n12361) );
  NOR2_X1 U11725 ( .A1(n18389), .A2(n21325), .ZN(n10190) );
  INV_X1 U11726 ( .A(n18387), .ZN(n10191) );
  NAND2_X1 U11728 ( .A1(n9959), .A2(n18463), .ZN(n17119) );
  NOR2_X1 U11729 ( .A1(n10087), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10086) );
  INV_X1 U11730 ( .A(n12160), .ZN(n10087) );
  OR2_X1 U11731 ( .A1(n18344), .A2(n18246), .ZN(n12159) );
  NOR2_X1 U11732 ( .A1(n12296), .A2(n12326), .ZN(n19336) );
  NAND2_X1 U11733 ( .A1(n18511), .A2(n12143), .ZN(n18498) );
  NAND2_X1 U11734 ( .A1(n18512), .A2(n18513), .ZN(n18511) );
  NOR2_X1 U11735 ( .A1(n18917), .A2(n12326), .ZN(n12329) );
  INV_X1 U11736 ( .A(n16683), .ZN(n18553) );
  NOR2_X2 U11737 ( .A1(n12174), .A2(n12173), .ZN(n19539) );
  INV_X1 U11738 ( .A(n17562), .ZN(n18893) );
  NAND2_X1 U11739 ( .A1(n12831), .A2(n12668), .ZN(n21026) );
  AND2_X1 U11740 ( .A1(n15180), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20593) );
  INV_X1 U11741 ( .A(n20592), .ZN(n20602) );
  XNOR2_X1 U11742 ( .A(n13829), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15252) );
  NAND2_X1 U11743 ( .A1(n10264), .A2(n10263), .ZN(n10259) );
  INV_X1 U11744 ( .A(n16774), .ZN(n16759) );
  OR2_X1 U11745 ( .A1(n16628), .A2(n20508), .ZN(n20516) );
  NAND2_X1 U11746 ( .A1(n10268), .A2(n10262), .ZN(n10261) );
  AND2_X1 U11747 ( .A1(n10267), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10262) );
  INV_X1 U11748 ( .A(n15220), .ZN(n10164) );
  INV_X1 U11749 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16622) );
  NOR2_X1 U11750 ( .A1(n9753), .A2(n12013), .ZN(n16890) );
  OR2_X1 U11751 ( .A1(n12034), .A2(n10317), .ZN(n12037) );
  NOR2_X1 U11752 ( .A1(n9693), .A2(n19687), .ZN(n12036) );
  NAND2_X1 U11753 ( .A1(n11533), .A2(n11532), .ZN(n11541) );
  NAND2_X1 U11754 ( .A1(n19712), .A2(n10284), .ZN(n10287) );
  INV_X1 U11755 ( .A(n19713), .ZN(n16970) );
  INV_X1 U11756 ( .A(n20487), .ZN(n19776) );
  INV_X1 U11757 ( .A(n16322), .ZN(n10049) );
  NAND2_X1 U11758 ( .A1(n17074), .A2(n19828), .ZN(n9885) );
  NAND2_X1 U11759 ( .A1(n17072), .A2(n19848), .ZN(n9884) );
  INV_X1 U11760 ( .A(n17038), .ZN(n19840) );
  INV_X1 U11761 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17047) );
  NAND2_X1 U11762 ( .A1(n19848), .A2(n10284), .ZN(n10290) );
  AND2_X1 U11763 ( .A1(n17046), .A2(n15261), .ZN(n17038) );
  AND2_X1 U11764 ( .A1(n17046), .A2(n20472), .ZN(n19848) );
  NAND2_X1 U11765 ( .A1(n10094), .A2(n10093), .ZN(n11550) );
  XNOR2_X1 U11766 ( .A(n11528), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11488) );
  NAND2_X1 U11767 ( .A1(n10051), .A2(n16172), .ZN(n16333) );
  NAND2_X1 U11768 ( .A1(n9769), .A2(n16327), .ZN(n10051) );
  XNOR2_X1 U11769 ( .A(n10073), .B(n16251), .ZN(n16393) );
  NAND2_X1 U11770 ( .A1(n10074), .A2(n16249), .ZN(n10073) );
  INV_X1 U11771 ( .A(n16250), .ZN(n10074) );
  XNOR2_X1 U11772 ( .A(n16997), .B(n17068), .ZN(n17073) );
  INV_X1 U11773 ( .A(n19854), .ZN(n17070) );
  INV_X1 U11774 ( .A(n19870), .ZN(n17086) );
  AND2_X1 U11775 ( .A1(n16436), .A2(n16431), .ZN(n16432) );
  INV_X1 U11776 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20492) );
  XNOR2_X1 U11777 ( .A(n13215), .B(n13218), .ZN(n19749) );
  INV_X1 U11778 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n17100) );
  NAND2_X1 U11779 ( .A1(n17674), .A2(n9831), .ZN(n17665) );
  NAND2_X1 U11780 ( .A1(n17684), .A2(n9837), .ZN(n17672) );
  NAND2_X1 U11781 ( .A1(n17672), .A2(n17916), .ZN(n17674) );
  NOR2_X1 U11782 ( .A1(n17627), .A2(n17679), .ZN(n17684) );
  NOR2_X1 U11783 ( .A1(n17969), .A2(n10029), .ZN(n10028) );
  INV_X1 U11784 ( .A(n10030), .ZN(n10029) );
  NOR2_X1 U11785 ( .A1(n17393), .A2(n17739), .ZN(n17716) );
  NOR3_X1 U11786 ( .A1(n17808), .A2(n17812), .A3(n17431), .ZN(n17796) );
  INV_X1 U11787 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n10023) );
  AND2_X1 U11788 ( .A1(n17924), .A2(n10040), .ZN(n17899) );
  INV_X1 U11789 ( .A(n17903), .ZN(n10040) );
  INV_X1 U11790 ( .A(n17924), .ZN(n17911) );
  INV_X1 U11791 ( .A(n17940), .ZN(n17936) );
  NAND2_X1 U11792 ( .A1(n18043), .A2(P3_EAX_REG_7__SCAN_IN), .ZN(n18037) );
  INV_X1 U11793 ( .A(n12250), .ZN(n18044) );
  CLKBUF_X1 U11794 ( .A(n12362), .Z(n17547) );
  AND2_X1 U11795 ( .A1(n18396), .A2(n17160), .ZN(n9948) );
  INV_X1 U11796 ( .A(n18467), .ZN(n18396) );
  INV_X1 U11797 ( .A(n18399), .ZN(n18464) );
  NAND2_X1 U11798 ( .A1(n9955), .A2(n9949), .ZN(n17159) );
  NAND2_X1 U11799 ( .A1(n17119), .A2(n9956), .ZN(n9955) );
  NAND2_X1 U11800 ( .A1(n9950), .A2(n17122), .ZN(n9949) );
  INV_X1 U11801 ( .A(n9957), .ZN(n9956) );
  OR2_X1 U11802 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11006), .ZN(
        n10670) );
  OAI21_X1 U11803 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n12306), .A(
        n12307), .ZN(n12308) );
  OR2_X1 U11804 ( .A1(n12311), .A2(n12312), .ZN(n12307) );
  AND2_X1 U11805 ( .A1(n12529), .A2(n12528), .ZN(n12531) );
  AOI21_X1 U11806 ( .B1(n12499), .B2(n12504), .A(n12431), .ZN(n12516) );
  OR2_X1 U11807 ( .A1(n13706), .A2(n13705), .ZN(n14408) );
  NOR2_X1 U11808 ( .A1(n13184), .A2(n13183), .ZN(n13197) );
  INV_X1 U11809 ( .A(n12754), .ZN(n12755) );
  INV_X1 U11810 ( .A(n12767), .ZN(n12756) );
  NAND2_X1 U11811 ( .A1(n9906), .A2(n13253), .ZN(n13695) );
  BUF_X4 U11812 ( .A(n12892), .Z(n15071) );
  NAND2_X1 U11813 ( .A1(n12555), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n9886) );
  NAND2_X1 U11814 ( .A1(n12438), .A2(n12444), .ZN(n9932) );
  NAND2_X1 U11815 ( .A1(n12436), .A2(n12443), .ZN(n9931) );
  AOI21_X1 U11816 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20737), .A(
        n12531), .ZN(n12526) );
  AND2_X1 U11817 ( .A1(n12486), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13972) );
  AND2_X1 U11818 ( .A1(n11149), .A2(n10993), .ZN(n11023) );
  INV_X1 U11819 ( .A(n16045), .ZN(n9854) );
  NAND2_X1 U11820 ( .A1(n9861), .A2(n16041), .ZN(n9860) );
  NOR2_X1 U11821 ( .A1(n9823), .A2(n9861), .ZN(n9857) );
  AND2_X1 U11822 ( .A1(n11503), .A2(n16312), .ZN(n10952) );
  NAND2_X1 U11823 ( .A1(n10055), .A2(n10054), .ZN(n10788) );
  OR2_X1 U11824 ( .A1(n11182), .A2(n14265), .ZN(n10054) );
  NAND2_X1 U11825 ( .A1(n9771), .A2(n11024), .ZN(n9867) );
  INV_X1 U11826 ( .A(n9881), .ZN(n9851) );
  INV_X1 U11827 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11668) );
  INV_X1 U11828 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11662) );
  INV_X1 U11829 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11661) );
  OAI21_X1 U11830 ( .B1(n13393), .B2(n11686), .A(n10279), .ZN(n10381) );
  NAND2_X1 U11831 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10279) );
  AND2_X1 U11832 ( .A1(n10688), .A2(n10689), .ZN(n10713) );
  AND2_X1 U11833 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10356) );
  NAND2_X1 U11834 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10353) );
  NAND2_X1 U11835 ( .A1(n19350), .A2(n19499), .ZN(n12041) );
  INV_X1 U11836 ( .A(n12140), .ZN(n10080) );
  INV_X1 U11837 ( .A(n15325), .ZN(n10217) );
  OR2_X1 U11838 ( .A1(n15009), .A2(n15370), .ZN(n15354) );
  AND2_X1 U11839 ( .A1(n15723), .A2(n9835), .ZN(n10275) );
  AND2_X1 U11840 ( .A1(n10006), .A2(n10275), .ZN(n9894) );
  INV_X1 U11841 ( .A(n15067), .ZN(n15099) );
  INV_X1 U11842 ( .A(n10213), .ZN(n10211) );
  NAND2_X1 U11843 ( .A1(n10021), .A2(n15232), .ZN(n10020) );
  INV_X1 U11844 ( .A(n15826), .ZN(n10021) );
  INV_X1 U11845 ( .A(n15416), .ZN(n10170) );
  OR2_X1 U11846 ( .A1(n15527), .A2(n10167), .ZN(n10166) );
  NAND2_X1 U11847 ( .A1(n10168), .A2(n15517), .ZN(n10167) );
  INV_X1 U11848 ( .A(n15468), .ZN(n10168) );
  OR2_X1 U11849 ( .A1(n12902), .A2(n12901), .ZN(n14535) );
  AND2_X1 U11850 ( .A1(n15162), .A2(n15147), .ZN(n15146) );
  AND2_X1 U11851 ( .A1(n15107), .A2(n13587), .ZN(n14530) );
  OR2_X1 U11852 ( .A1(n13250), .A2(n13249), .ZN(n13813) );
  NAND2_X1 U11853 ( .A1(n13085), .A2(n9922), .ZN(n10278) );
  NAND2_X1 U11854 ( .A1(n9756), .A2(n13519), .ZN(n12864) );
  OR2_X1 U11855 ( .A1(n12823), .A2(n12822), .ZN(n16616) );
  OR2_X1 U11856 ( .A1(n13515), .A2(n13983), .ZN(n20869) );
  NAND2_X1 U11857 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12458) );
  INV_X1 U11858 ( .A(n14530), .ZN(n14401) );
  AND2_X1 U11859 ( .A1(n10853), .A2(n10101), .ZN(n10866) );
  AND2_X1 U11860 ( .A1(n10103), .A2(n10102), .ZN(n10101) );
  INV_X1 U11861 ( .A(n10836), .ZN(n10111) );
  NOR2_X1 U11862 ( .A1(n10735), .A2(n10734), .ZN(n10791) );
  INV_X1 U11863 ( .A(n10695), .ZN(n10696) );
  NAND2_X1 U11864 ( .A1(n10703), .A2(n10696), .ZN(n10735) );
  NAND2_X1 U11865 ( .A1(n11966), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10682) );
  INV_X1 U11866 ( .A(n11014), .ZN(n10683) );
  NAND2_X1 U11867 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10575), .ZN(
        n11703) );
  CLKBUF_X1 U11868 ( .A(n11841), .Z(n11911) );
  NAND2_X1 U11869 ( .A1(n11936), .A2(n13387), .ZN(n11735) );
  INV_X1 U11870 ( .A(n13491), .ZN(n10227) );
  NOR2_X1 U11871 ( .A1(n16173), .A2(n10150), .ZN(n10149) );
  INV_X1 U11872 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10150) );
  NOR2_X1 U11873 ( .A1(n10145), .A2(n10142), .ZN(n10141) );
  INV_X1 U11874 ( .A(n10143), .ZN(n10142) );
  NOR2_X1 U11875 ( .A1(n12008), .A2(n10144), .ZN(n10143) );
  INV_X1 U11876 ( .A(n11990), .ZN(n11490) );
  NAND2_X1 U11877 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10310) );
  AND2_X1 U11878 ( .A1(n9833), .A2(n16323), .ZN(n9997) );
  AND2_X1 U11879 ( .A1(n15965), .A2(n16063), .ZN(n10133) );
  NAND2_X1 U11880 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10308) );
  NOR3_X1 U11881 ( .A1(n15983), .A2(n10236), .A3(n15967), .ZN(n16120) );
  NOR2_X1 U11882 ( .A1(n15983), .A2(n15967), .ZN(n16118) );
  AND2_X1 U11883 ( .A1(n9722), .A2(n9832), .ZN(n9994) );
  AND2_X1 U11884 ( .A1(n15987), .A2(n10880), .ZN(n10919) );
  NOR2_X1 U11885 ( .A1(n16427), .A2(n16441), .ZN(n10312) );
  AND2_X1 U11886 ( .A1(n9749), .A2(n10883), .ZN(n10914) );
  NOR2_X1 U11887 ( .A1(n14331), .A2(n10239), .ZN(n10238) );
  INV_X1 U11888 ( .A(n14179), .ZN(n10239) );
  AND2_X1 U11889 ( .A1(n10304), .A2(n11481), .ZN(n9722) );
  INV_X1 U11890 ( .A(n13504), .ZN(n10124) );
  INV_X1 U11891 ( .A(n16980), .ZN(n10064) );
  NOR2_X1 U11892 ( .A1(n14442), .A2(n10224), .ZN(n10223) );
  INV_X1 U11893 ( .A(n14303), .ZN(n10224) );
  AND4_X1 U11894 ( .A1(n10665), .A2(n10664), .A3(n10663), .A4(n10662), .ZN(
        n10679) );
  AND4_X1 U11895 ( .A1(n10669), .A2(n10668), .A3(n10667), .A4(n10666), .ZN(
        n10678) );
  NAND2_X1 U11896 ( .A1(n11471), .A2(n11470), .ZN(n11478) );
  INV_X1 U11897 ( .A(n11469), .ZN(n11471) );
  XNOR2_X1 U11898 ( .A(n11478), .B(n11189), .ZN(n11473) );
  INV_X1 U11899 ( .A(n13670), .ZN(n11462) );
  AND2_X1 U11900 ( .A1(n9798), .A2(n10742), .ZN(n9993) );
  NAND2_X1 U11901 ( .A1(n11455), .A2(n11456), .ZN(n9878) );
  OR2_X1 U11902 ( .A1(n19834), .A2(n11451), .ZN(n11452) );
  NAND2_X1 U11903 ( .A1(n10046), .A2(n10047), .ZN(n10045) );
  NAND4_X1 U11904 ( .A1(n10400), .A2(n10474), .A3(n10468), .A4(n19896), .ZN(
        n10484) );
  AOI21_X1 U11905 ( .B1(n10699), .B2(n19693), .A(n9757), .ZN(n10704) );
  NAND2_X1 U11906 ( .A1(n10491), .A2(n10486), .ZN(n9863) );
  INV_X1 U11907 ( .A(n10694), .ZN(n11423) );
  AOI21_X1 U11908 ( .B1(n9851), .B2(n11582), .A(n11581), .ZN(n11583) );
  OR2_X1 U11909 ( .A1(n10544), .A2(n15264), .ZN(n10562) );
  NOR2_X1 U11910 ( .A1(n10391), .A2(n10281), .ZN(n10456) );
  NAND2_X1 U11911 ( .A1(n20471), .A2(n20320), .ZN(n13224) );
  AOI22_X1 U11912 ( .A1(n10591), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n10584), .ZN(n10394) );
  AND2_X1 U11913 ( .A1(n20492), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10973) );
  AND2_X1 U11914 ( .A1(n21291), .A2(n10984), .ZN(n10999) );
  NOR2_X1 U11915 ( .A1(n18125), .A2(n18893), .ZN(n12283) );
  NOR2_X1 U11916 ( .A1(n12192), .A2(n9916), .ZN(n9915) );
  NAND2_X1 U11917 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19515), .ZN(
        n12046) );
  INV_X1 U11918 ( .A(n16586), .ZN(n12045) );
  NAND2_X1 U11919 ( .A1(n19539), .A2(n18893), .ZN(n16681) );
  AND2_X1 U11921 ( .A1(n9818), .A2(n10091), .ZN(n10090) );
  INV_X1 U11922 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U11923 ( .A1(n18475), .A2(n12150), .ZN(n12151) );
  AND2_X1 U11924 ( .A1(n19336), .A2(n12280), .ZN(n14661) );
  NOR2_X1 U11925 ( .A1(n19539), .A2(n18124), .ZN(n16582) );
  NOR2_X1 U11926 ( .A1(n17259), .A2(n19542), .ZN(n16579) );
  INV_X1 U11927 ( .A(n19343), .ZN(n19346) );
  AND2_X1 U11928 ( .A1(n15389), .A2(n9828), .ZN(n15326) );
  INV_X1 U11929 ( .A(n15327), .ZN(n10172) );
  AND2_X1 U11930 ( .A1(n15389), .A2(n15375), .ZN(n15377) );
  AND2_X1 U11931 ( .A1(n15402), .A2(n15387), .ZN(n15389) );
  AND2_X1 U11932 ( .A1(n16646), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13077) );
  NAND2_X1 U11933 ( .A1(n12603), .A2(n12602), .ZN(n20619) );
  OR2_X1 U11934 ( .A1(n15050), .A2(n15633), .ZN(n15070) );
  NAND2_X1 U11935 ( .A1(n15029), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15050) );
  OR2_X1 U11936 ( .A1(n14902), .A2(n15344), .ZN(n15012) );
  NAND2_X1 U11937 ( .A1(n14969), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14973) );
  AND2_X1 U11938 ( .A1(n13828), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14969) );
  INV_X1 U11939 ( .A(n15006), .ZN(n13828) );
  NOR2_X1 U11940 ( .A1(n14855), .A2(n14854), .ZN(n14883) );
  NAND2_X1 U11941 ( .A1(n14883), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14888) );
  INV_X1 U11942 ( .A(n10329), .ZN(n10207) );
  NAND2_X1 U11943 ( .A1(n14835), .A2(n9789), .ZN(n15427) );
  NAND2_X1 U11944 ( .A1(n14836), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14855) );
  NOR2_X1 U11945 ( .A1(n14783), .A2(n16704), .ZN(n14801) );
  NAND2_X1 U11946 ( .A1(n14801), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14829) );
  AND2_X1 U11947 ( .A1(n14750), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14768) );
  NOR2_X1 U11948 ( .A1(n14626), .A2(n14645), .ZN(n14750) );
  INV_X1 U11949 ( .A(n14641), .ZN(n10212) );
  NOR2_X1 U11950 ( .A1(n14367), .A2(n15785), .ZN(n14595) );
  AND2_X1 U11951 ( .A1(n10198), .A2(n14611), .ZN(n10197) );
  OR2_X1 U11952 ( .A1(n14593), .A2(n10199), .ZN(n10198) );
  NAND2_X1 U11953 ( .A1(n10196), .A2(n14598), .ZN(n10195) );
  NAND2_X1 U11954 ( .A1(n14594), .A2(n14593), .ZN(n10196) );
  NAND2_X1 U11955 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n14351), .ZN(
        n14367) );
  NOR2_X1 U11956 ( .A1(n21296), .A2(n14223), .ZN(n14351) );
  INV_X1 U11957 ( .A(n13973), .ZN(n14107) );
  NAND2_X1 U11958 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n14107), .ZN(
        n14223) );
  OAI211_X1 U11959 ( .C1(n13616), .C2(n13977), .A(n13976), .B(n13975), .ZN(
        n13979) );
  NOR2_X1 U11960 ( .A1(n20559), .A2(n13688), .ZN(n13974) );
  NAND2_X1 U11961 ( .A1(n13713), .A2(n13712), .ZN(n13714) );
  NAND2_X1 U11962 ( .A1(n10206), .A2(n13710), .ZN(n13713) );
  INV_X1 U11963 ( .A(n13624), .ZN(n13625) );
  CLKBUF_X1 U11964 ( .A(n13623), .Z(n13266) );
  NOR2_X1 U11965 ( .A1(n13257), .A2(n13256), .ZN(n13618) );
  NAND2_X1 U11966 ( .A1(n13150), .A2(n13149), .ZN(n13156) );
  NAND2_X1 U11967 ( .A1(n13615), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13148) );
  NAND2_X1 U11968 ( .A1(n10016), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10015) );
  INV_X1 U11969 ( .A(n10017), .ZN(n10016) );
  NOR2_X1 U11970 ( .A1(n15629), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10267) );
  NAND2_X1 U11971 ( .A1(n10019), .A2(n10018), .ZN(n10017) );
  INV_X1 U11972 ( .A(n10020), .ZN(n10018) );
  INV_X1 U11973 ( .A(n15628), .ZN(n10019) );
  AND2_X1 U11974 ( .A1(n15326), .A2(n15312), .ZN(n15314) );
  NAND2_X1 U11975 ( .A1(n15314), .A2(n15296), .ZN(n15298) );
  NAND2_X1 U11976 ( .A1(n15389), .A2(n10173), .ZN(n15341) );
  NAND2_X1 U11977 ( .A1(n15389), .A2(n9821), .ZN(n15361) );
  OAI21_X1 U11978 ( .B1(n15212), .B2(n9941), .A(n9939), .ZN(n15658) );
  NAND2_X1 U11979 ( .A1(n9714), .A2(n9942), .ZN(n9940) );
  NAND2_X1 U11980 ( .A1(n9943), .A2(n9938), .ZN(n9897) );
  OR2_X1 U11981 ( .A1(n15212), .A2(n15213), .ZN(n9938) );
  NAND2_X1 U11982 ( .A1(n15209), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9896) );
  AND2_X1 U11983 ( .A1(n15508), .A2(n15132), .ZN(n15456) );
  NOR2_X1 U11984 ( .A1(n9717), .A2(n15507), .ZN(n15508) );
  NOR3_X1 U11985 ( .A1(n15469), .A2(n15527), .A3(n15468), .ZN(n15525) );
  NOR2_X1 U11986 ( .A1(n15469), .A2(n15468), .ZN(n15524) );
  OR2_X1 U11987 ( .A1(n14649), .A2(n14648), .ZN(n15469) );
  NAND2_X1 U11988 ( .A1(n14620), .A2(n14619), .ZN(n14649) );
  AOI21_X1 U11989 ( .B1(n9724), .B2(n14587), .A(n9768), .ZN(n9892) );
  NOR2_X1 U11990 ( .A1(n16835), .A2(n14376), .ZN(n14620) );
  INV_X1 U11991 ( .A(n14242), .ZN(n10162) );
  INV_X1 U11992 ( .A(n14241), .ZN(n10163) );
  AND2_X1 U11993 ( .A1(n14375), .A2(n14374), .ZN(n16832) );
  NAND2_X1 U11994 ( .A1(n10161), .A2(n10160), .ZN(n16835) );
  INV_X1 U11995 ( .A(n16832), .ZN(n10160) );
  INV_X1 U11996 ( .A(n10272), .ZN(n10271) );
  NAND2_X1 U11997 ( .A1(n16856), .A2(n14119), .ZN(n14241) );
  AND2_X1 U11998 ( .A1(n16854), .A2(n16853), .ZN(n16856) );
  AND2_X1 U11999 ( .A1(n13756), .A2(n13755), .ZN(n13757) );
  NAND2_X1 U12000 ( .A1(n13631), .A2(n13630), .ZN(n13758) );
  NAND2_X1 U12001 ( .A1(n9756), .A2(n9727), .ZN(n13107) );
  NAND2_X1 U12002 ( .A1(n10003), .A2(n12597), .ZN(n10002) );
  AND2_X1 U12003 ( .A1(n13270), .A2(n13269), .ZN(n13278) );
  NAND2_X1 U12004 ( .A1(n13117), .A2(n15278), .ZN(n15863) );
  OR2_X1 U12005 ( .A1(n20657), .A2(n20656), .ZN(n15224) );
  OR2_X1 U12006 ( .A1(n20657), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13210) );
  INV_X1 U12007 ( .A(n15863), .ZN(n15914) );
  NAND2_X1 U12008 ( .A1(n12769), .A2(n12768), .ZN(n13082) );
  NAND2_X1 U12009 ( .A1(n12766), .A2(n12764), .ZN(n12769) );
  AOI21_X1 U12010 ( .B1(n10010), .B2(n10011), .A(n10008), .ZN(n10007) );
  NAND2_X1 U12011 ( .A1(n12909), .A2(n12908), .ZN(n10014) );
  AOI21_X1 U12012 ( .B1(n13141), .B2(n13140), .A(n14531), .ZN(n13143) );
  OR2_X1 U12013 ( .A1(n13718), .A2(n13085), .ZN(n13086) );
  NAND2_X1 U12014 ( .A1(n13085), .A2(n12791), .ZN(n10202) );
  XNOR2_X1 U12015 ( .A(n13173), .B(n13544), .ZN(n13908) );
  NAND2_X1 U12016 ( .A1(n13577), .A2(n12591), .ZN(n12596) );
  CLKBUF_X1 U12017 ( .A(n13533), .Z(n14739) );
  NAND2_X1 U12018 ( .A1(n13637), .A2(n13539), .ZN(n20695) );
  AND2_X1 U12019 ( .A1(n13540), .A2(n15927), .ZN(n13764) );
  NAND2_X1 U12020 ( .A1(n10344), .A2(n12578), .ZN(n13558) );
  AND3_X1 U12021 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n9922), .A3(n13546), 
        .ZN(n13596) );
  NAND2_X1 U12022 ( .A1(n16764), .A2(n15109), .ZN(n13592) );
  AND2_X1 U12023 ( .A1(n21133), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16646) );
  AND2_X1 U12024 ( .A1(n14265), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12620) );
  NAND2_X1 U12025 ( .A1(n12019), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12622) );
  CLKBUF_X1 U12026 ( .A(n11010), .Z(n11011) );
  NOR2_X1 U12027 ( .A1(n11410), .A2(n11409), .ZN(n13427) );
  NOR2_X1 U12028 ( .A1(n10099), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10098) );
  INV_X1 U12029 ( .A(n10100), .ZN(n10099) );
  NOR2_X1 U12030 ( .A1(n16908), .A2(n19656), .ZN(n16898) );
  NOR2_X1 U12031 ( .A1(n19656), .A2(n16920), .ZN(n16909) );
  NOR2_X1 U12032 ( .A1(n16909), .A2(n16910), .ZN(n16908) );
  NAND2_X1 U12033 ( .A1(n10948), .A2(n10949), .ZN(n10956) );
  NAND2_X1 U12034 ( .A1(n11525), .A2(n10938), .ZN(n10939) );
  NOR2_X1 U12035 ( .A1(n19656), .A2(n16933), .ZN(n15935) );
  NOR2_X1 U12036 ( .A1(n10136), .A2(n10135), .ZN(n16934) );
  OAI21_X1 U12037 ( .B1(n10138), .B2(n16007), .A(n16007), .ZN(n10136) );
  NOR2_X1 U12038 ( .A1(n16944), .A2(n10138), .ZN(n10135) );
  OAI21_X1 U12039 ( .B1(n19656), .B2(n10140), .A(n10139), .ZN(n10138) );
  INV_X1 U12040 ( .A(n16945), .ZN(n10140) );
  INV_X1 U12041 ( .A(n16201), .ZN(n10139) );
  NOR2_X1 U12042 ( .A1(n10929), .A2(n10115), .ZN(n10114) );
  AND2_X1 U12043 ( .A1(n15949), .A2(n10931), .ZN(n10933) );
  NOR2_X1 U12044 ( .A1(n16944), .A2(n16945), .ZN(n16943) );
  AND2_X1 U12045 ( .A1(n14277), .A2(n12011), .ZN(n15973) );
  INV_X1 U12046 ( .A(n10914), .ZN(n19590) );
  AND2_X1 U12047 ( .A1(n9735), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10156) );
  NOR2_X1 U12048 ( .A1(n10902), .A2(n10106), .ZN(n10105) );
  INV_X1 U12049 ( .A(n10867), .ZN(n10106) );
  NAND2_X1 U12050 ( .A1(n10853), .A2(n10103), .ZN(n10859) );
  NAND2_X1 U12051 ( .A1(n10791), .A2(n10790), .ZN(n10837) );
  XNOR2_X1 U12052 ( .A(n11161), .B(n11160), .ZN(n12965) );
  NOR3_X1 U12053 ( .A1(n16033), .A2(n9817), .A3(n16032), .ZN(n11533) );
  INV_X1 U12054 ( .A(n12388), .ZN(n10127) );
  AND2_X1 U12055 ( .A1(n10128), .A2(n10126), .ZN(n12389) );
  INV_X1 U12056 ( .A(n11507), .ZN(n10126) );
  AND3_X1 U12057 ( .A1(n11080), .A2(n11079), .A3(n11078), .ZN(n13503) );
  NAND2_X1 U12058 ( .A1(n19666), .A2(n9803), .ZN(n13287) );
  NOR3_X1 U12059 ( .A1(n10242), .A2(n10241), .A3(n10245), .ZN(n10240) );
  INV_X1 U12060 ( .A(n15938), .ZN(n10241) );
  INV_X1 U12061 ( .A(n12402), .ZN(n10245) );
  NOR2_X1 U12062 ( .A1(n11401), .A2(n11402), .ZN(n11554) );
  AOI21_X1 U12063 ( .B1(n16027), .B2(n9741), .A(n9825), .ZN(n9870) );
  NOR2_X1 U12064 ( .A1(n15937), .A2(n10242), .ZN(n12401) );
  NAND2_X1 U12065 ( .A1(n10232), .A2(n10231), .ZN(n10230) );
  NOR2_X1 U12066 ( .A1(n10236), .A2(n15952), .ZN(n10231) );
  INV_X1 U12067 ( .A(n10233), .ZN(n10232) );
  NAND2_X1 U12068 ( .A1(n11794), .A2(n10293), .ZN(n10292) );
  AOI211_X1 U12069 ( .C1(n16955), .C2(n11813), .A(n19668), .B(n11816), .ZN(
        n16957) );
  NAND2_X1 U12070 ( .A1(n16054), .A2(n16053), .ZN(n16052) );
  CLKBUF_X1 U12071 ( .A(n16068), .Z(n16128) );
  AND2_X1 U12072 ( .A1(n11382), .A2(n11381), .ZN(n16152) );
  NOR2_X1 U12073 ( .A1(n9814), .A2(n10295), .ZN(n10294) );
  INV_X1 U12074 ( .A(n13662), .ZN(n9871) );
  INV_X1 U12075 ( .A(n16072), .ZN(n10295) );
  AND2_X1 U12076 ( .A1(n11308), .A2(n11307), .ZN(n17080) );
  NAND2_X1 U12077 ( .A1(n16472), .A2(n16473), .ZN(n17079) );
  AND2_X1 U12078 ( .A1(n11261), .A2(n11260), .ZN(n16494) );
  NAND2_X1 U12079 ( .A1(n14304), .A2(n14303), .ZN(n14441) );
  INV_X1 U12080 ( .A(n19561), .ZN(n13124) );
  NOR2_X1 U12081 ( .A1(n12989), .A2(n10226), .ZN(n13681) );
  NAND2_X1 U12082 ( .A1(n10228), .A2(n10227), .ZN(n10226) );
  INV_X1 U12083 ( .A(n11836), .ZN(n19668) );
  AND2_X1 U12084 ( .A1(n19744), .A2(n11956), .ZN(n12959) );
  NAND2_X1 U12085 ( .A1(n11152), .A2(n11151), .ZN(n12840) );
  NAND2_X1 U12086 ( .A1(n10220), .A2(n10218), .ZN(n11152) );
  INV_X1 U12087 ( .A(n11447), .ZN(n10220) );
  OAI21_X1 U12088 ( .B1(n11965), .B2(n11964), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12694) );
  NOR2_X1 U12089 ( .A1(n12629), .A2(n12035), .ZN(n19819) );
  XNOR2_X1 U12090 ( .A(n11544), .B(n11543), .ZN(n11977) );
  OR2_X1 U12091 ( .A1(n11985), .A2(n16211), .ZN(n11986) );
  OR2_X1 U12092 ( .A1(n11986), .A2(n16199), .ZN(n11983) );
  NAND2_X1 U12093 ( .A1(n15979), .A2(n10133), .ZN(n16062) );
  AND2_X1 U12094 ( .A1(n11490), .A2(n10141), .ZN(n11989) );
  NAND2_X1 U12095 ( .A1(n11490), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12009) );
  NOR2_X1 U12096 ( .A1(n16011), .A2(n16010), .ZN(n16074) );
  AND3_X1 U12097 ( .A1(n11086), .A2(n11085), .A3(n11084), .ZN(n14171) );
  NAND2_X1 U12098 ( .A1(n10124), .A2(n9790), .ZN(n14172) );
  NAND2_X1 U12099 ( .A1(n11996), .A2(n9735), .ZN(n12006) );
  AND2_X1 U12100 ( .A1(n13313), .A2(n13312), .ZN(n13474) );
  AND2_X1 U12101 ( .A1(n9721), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10153) );
  AND3_X1 U12102 ( .A1(n11072), .A2(n11071), .A3(n11070), .ZN(n13297) );
  NOR2_X1 U12103 ( .A1(n13296), .A2(n13297), .ZN(n13312) );
  INV_X1 U12104 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14295) );
  NAND2_X1 U12105 ( .A1(n11999), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12003) );
  AND3_X1 U12106 ( .A1(n11060), .A2(n11059), .A3(n11058), .ZN(n13304) );
  NAND2_X1 U12107 ( .A1(n10134), .A2(n9767), .ZN(n12002) );
  INV_X1 U12108 ( .A(n12001), .ZN(n10134) );
  XNOR2_X1 U12109 ( .A(n9881), .B(n11582), .ZN(n10533) );
  NOR2_X1 U12110 ( .A1(n9983), .A2(n10250), .ZN(n9981) );
  NAND2_X1 U12111 ( .A1(n12033), .A2(n10967), .ZN(n11518) );
  INV_X1 U12112 ( .A(n10128), .ZN(n16035) );
  AND2_X1 U12113 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n16348), .ZN(
        n16335) );
  AND2_X1 U12114 ( .A1(n10961), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16186) );
  NAND2_X1 U12115 ( .A1(n16198), .A2(n16195), .ZN(n9843) );
  NAND2_X1 U12116 ( .A1(n15979), .A2(n10131), .ZN(n16057) );
  AND2_X1 U12117 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  INV_X1 U12118 ( .A(n16055), .ZN(n10132) );
  NOR2_X1 U12119 ( .A1(n16057), .A2(n15950), .ZN(n16049) );
  NAND2_X1 U12120 ( .A1(n9989), .A2(n9988), .ZN(n10253) );
  AND2_X1 U12121 ( .A1(n9992), .A2(n10078), .ZN(n9988) );
  AND2_X1 U12122 ( .A1(n10923), .A2(n16993), .ZN(n9992) );
  AND2_X1 U12123 ( .A1(n15979), .A2(n15965), .ZN(n16064) );
  OR2_X1 U12124 ( .A1(n15986), .A2(n10909), .ZN(n16247) );
  AND3_X1 U12125 ( .A1(n11099), .A2(n11098), .A3(n11097), .ZN(n15992) );
  NAND2_X1 U12126 ( .A1(n10120), .A2(n10119), .ZN(n15994) );
  INV_X1 U12127 ( .A(n15992), .ZN(n10119) );
  INV_X1 U12128 ( .A(n15991), .ZN(n10120) );
  AND2_X1 U12129 ( .A1(n11429), .A2(n11481), .ZN(n16405) );
  AND2_X1 U12130 ( .A1(n10919), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16262) );
  OR3_X1 U12131 ( .A1(n19590), .A2(n11189), .A3(n16420), .ZN(n16260) );
  NAND2_X1 U12132 ( .A1(n14321), .A2(n10238), .ZN(n16153) );
  NAND2_X1 U12133 ( .A1(n9995), .A2(n9722), .ZN(n16295) );
  AND2_X1 U12134 ( .A1(n17049), .A2(n14320), .ZN(n14321) );
  NAND2_X1 U12135 ( .A1(n14321), .A2(n14179), .ZN(n14332) );
  NAND2_X1 U12136 ( .A1(n9791), .A2(n10122), .ZN(n10121) );
  INV_X1 U12137 ( .A(n14083), .ZN(n10122) );
  NAND2_X1 U12138 ( .A1(n10124), .A2(n9791), .ZN(n14174) );
  NAND2_X1 U12139 ( .A1(n10060), .A2(n16301), .ZN(n10056) );
  AOI21_X1 U12140 ( .B1(n10060), .B2(n10062), .A(n10059), .ZN(n10058) );
  CLKBUF_X1 U12141 ( .A(n16295), .Z(n16296) );
  NOR2_X1 U12142 ( .A1(n17051), .A2(n17050), .ZN(n17049) );
  NOR2_X1 U12143 ( .A1(n17079), .A2(n17080), .ZN(n17078) );
  NAND2_X1 U12144 ( .A1(n17078), .A2(n14491), .ZN(n17051) );
  AND2_X1 U12145 ( .A1(n14304), .A2(n10223), .ZN(n14469) );
  NAND2_X1 U12146 ( .A1(n14304), .A2(n9795), .ZN(n16495) );
  INV_X1 U12147 ( .A(n14443), .ZN(n14306) );
  NAND2_X1 U12148 ( .A1(n13322), .A2(n13285), .ZN(n13296) );
  NOR2_X1 U12149 ( .A1(n10069), .A2(n9977), .ZN(n9976) );
  NAND2_X1 U12150 ( .A1(n13679), .A2(n11186), .ZN(n14092) );
  AND2_X1 U12151 ( .A1(n11057), .A2(n9777), .ZN(n13320) );
  INV_X1 U12152 ( .A(n13128), .ZN(n10129) );
  NAND2_X1 U12153 ( .A1(n11057), .A2(n10130), .ZN(n13306) );
  AND3_X1 U12154 ( .A1(n11055), .A2(n11054), .A3(n11053), .ZN(n13487) );
  NAND2_X1 U12155 ( .A1(n11057), .A2(n11056), .ZN(n13303) );
  NAND2_X1 U12156 ( .A1(n9878), .A2(n11454), .ZN(n13485) );
  INV_X1 U12157 ( .A(n10710), .ZN(n10711) );
  NAND2_X1 U12158 ( .A1(n11042), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10487) );
  NAND2_X1 U12159 ( .A1(n11536), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10488) );
  CLKBUF_X1 U12160 ( .A(n11136), .Z(n13413) );
  NAND2_X1 U12161 ( .A1(n11568), .A2(n20101), .ZN(n11593) );
  OAI21_X1 U12162 ( .B1(n11977), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11978), 
        .ZN(n14277) );
  NAND2_X1 U12163 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U12164 ( .A1(n10990), .A2(n10989), .ZN(n13219) );
  AND2_X1 U12165 ( .A1(n19749), .A2(n19776), .ZN(n20067) );
  AND2_X1 U12166 ( .A1(n20466), .A2(n14255), .ZN(n20097) );
  INV_X1 U12167 ( .A(n20097), .ZN(n20132) );
  INV_X1 U12168 ( .A(n20454), .ZN(n20209) );
  INV_X1 U12169 ( .A(n20260), .ZN(n13646) );
  NOR2_X1 U12170 ( .A1(n10410), .A2(n13387), .ZN(n10411) );
  INV_X1 U12171 ( .A(n20316), .ZN(n20068) );
  INV_X1 U12172 ( .A(n20130), .ZN(n14254) );
  OR2_X1 U12173 ( .A1(n19749), .A2(n19776), .ZN(n20166) );
  NOR2_X2 U12174 ( .A1(n13225), .A2(n13224), .ZN(n19909) );
  NOR2_X2 U12175 ( .A1(n13223), .A2(n13224), .ZN(n19910) );
  OR2_X1 U12176 ( .A1(n20466), .A2(n14255), .ZN(n20316) );
  INV_X1 U12177 ( .A(n19909), .ZN(n19900) );
  INV_X1 U12178 ( .A(n19910), .ZN(n19902) );
  INV_X1 U12179 ( .A(n19890), .ZN(n19904) );
  NOR2_X1 U12180 ( .A1(n12283), .A2(n12291), .ZN(n19542) );
  AOI21_X1 U12181 ( .B1(n12322), .B2(n12317), .A(n12321), .ZN(n19324) );
  NOR3_X1 U12182 ( .A1(n16579), .A2(n16582), .A3(n19349), .ZN(n19323) );
  OAI21_X1 U12184 ( .B1(n17357), .B2(n10186), .A(n10185), .ZN(n17340) );
  NAND2_X1 U12185 ( .A1(n17547), .A2(n18257), .ZN(n10185) );
  NOR2_X1 U12188 ( .A1(n17703), .A2(n10031), .ZN(n10030) );
  INV_X1 U12189 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U12190 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .ZN(n10036) );
  NAND2_X1 U12191 ( .A1(n10025), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n10024) );
  NOR2_X1 U12192 ( .A1(n17481), .A2(n17854), .ZN(n10025) );
  NAND2_X1 U12193 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17899), .ZN(n17896) );
  NOR2_X1 U12194 ( .A1(n18080), .A2(n9908), .ZN(n9907) );
  INV_X1 U12195 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n9908) );
  AND2_X1 U12196 ( .A1(n18255), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18234) );
  INV_X1 U12198 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n21325) );
  NAND2_X1 U12199 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18389) );
  NAND2_X1 U12200 ( .A1(n17511), .A2(n10326), .ZN(n18387) );
  NAND2_X1 U12201 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18415) );
  NOR2_X1 U12202 ( .A1(n12279), .A2(n18459), .ZN(n18731) );
  NOR2_X1 U12203 ( .A1(n12273), .A2(n12277), .ZN(n12279) );
  XNOR2_X1 U12204 ( .A(n12149), .B(n9970), .ZN(n18476) );
  INV_X1 U12205 ( .A(n12148), .ZN(n9970) );
  NAND2_X1 U12206 ( .A1(n18476), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18475) );
  NAND2_X1 U12207 ( .A1(n9836), .A2(n9728), .ZN(n18481) );
  INV_X1 U12208 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17566) );
  INV_X1 U12209 ( .A(n19539), .ZN(n18125) );
  INV_X1 U12210 ( .A(n17161), .ZN(n9951) );
  NAND2_X1 U12211 ( .A1(n9954), .A2(n9953), .ZN(n9952) );
  NAND2_X1 U12212 ( .A1(n19505), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9953) );
  NOR2_X1 U12213 ( .A1(n18382), .A2(n18200), .ZN(n16595) );
  NAND2_X1 U12214 ( .A1(n10083), .A2(n18218), .ZN(n18200) );
  AND2_X1 U12215 ( .A1(n18230), .A2(n10084), .ZN(n10083) );
  NOR2_X1 U12216 ( .A1(n12164), .A2(n18205), .ZN(n10084) );
  NOR3_X1 U12217 ( .A1(n18322), .A2(n12156), .A3(n18321), .ZN(n18252) );
  INV_X1 U12218 ( .A(n9961), .ZN(n18302) );
  AND2_X1 U12219 ( .A1(n9961), .A2(n9960), .ZN(n18322) );
  INV_X1 U12220 ( .A(n18281), .ZN(n9960) );
  NAND2_X1 U12221 ( .A1(n9963), .A2(n9962), .ZN(n18334) );
  AND2_X1 U12222 ( .A1(n12153), .A2(n9806), .ZN(n9962) );
  NAND2_X1 U12223 ( .A1(n9964), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9963) );
  NOR2_X1 U12224 ( .A1(n12155), .A2(n12154), .ZN(n18344) );
  NOR2_X1 U12225 ( .A1(n18729), .A2(n18700), .ZN(n18374) );
  NOR2_X1 U12226 ( .A1(n18731), .A2(n18718), .ZN(n18368) );
  NAND2_X1 U12227 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18368), .ZN(
        n18367) );
  NAND2_X1 U12228 ( .A1(n18440), .A2(n9818), .ZN(n18403) );
  INV_X1 U12229 ( .A(n18036), .ZN(n17116) );
  AOI21_X1 U12230 ( .B1(n12278), .B2(n12277), .A(n12276), .ZN(n18460) );
  AOI21_X1 U12231 ( .B1(n9730), .B2(n9947), .A(n9946), .ZN(n18484) );
  NOR2_X1 U12232 ( .A1(n18499), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9946) );
  INV_X1 U12233 ( .A(n18498), .ZN(n9947) );
  NAND2_X1 U12234 ( .A1(n18484), .A2(n18483), .ZN(n18482) );
  AOI211_X1 U12235 ( .C1(n17839), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n12183), .B(n12182), .ZN(n12184) );
  AOI211_X1 U12236 ( .C1(n12324), .C2(n12323), .A(n12322), .B(n12321), .ZN(
        n19321) );
  INV_X1 U12237 ( .A(n19331), .ZN(n19360) );
  NOR2_X1 U12238 ( .A1(n9909), .A2(n16579), .ZN(n19343) );
  OR2_X1 U12239 ( .A1(n16582), .A2(n9910), .ZN(n9909) );
  AND2_X1 U12240 ( .A1(n12290), .A2(n14661), .ZN(n9910) );
  INV_X1 U12241 ( .A(n19334), .ZN(n19353) );
  NOR2_X1 U12242 ( .A1(n19550), .A2(n14658), .ZN(n19334) );
  NOR2_X1 U12243 ( .A1(n12372), .A2(n19346), .ZN(n19349) );
  NOR2_X1 U12244 ( .A1(n12204), .A2(n12203), .ZN(n18914) );
  INV_X1 U12245 ( .A(n17926), .ZN(n18922) );
  NOR2_X1 U12246 ( .A1(n12214), .A2(n12213), .ZN(n18917) );
  NAND2_X1 U12247 ( .A1(n17110), .A2(n18891), .ZN(n19001) );
  AOI22_X1 U12248 ( .A1(n19321), .A2(n19320), .B1(n19325), .B2(n17109), .ZN(
        n19329) );
  INV_X1 U12249 ( .A(n15476), .ZN(n20554) );
  INV_X1 U12250 ( .A(n20578), .ZN(n20596) );
  INV_X1 U12251 ( .A(n20595), .ZN(n20580) );
  AND2_X1 U12252 ( .A1(n13831), .A2(n15476), .ZN(n20585) );
  INV_X1 U12253 ( .A(n20618), .ZN(n21041) );
  AND2_X1 U12254 ( .A1(n20618), .A2(n15533), .ZN(n21040) );
  NAND2_X2 U12255 ( .A1(n13053), .A2(n13052), .ZN(n20618) );
  CLKBUF_X1 U12256 ( .A(n15529), .Z(n15513) );
  INV_X1 U12257 ( .A(n21040), .ZN(n16730) );
  INV_X1 U12258 ( .A(n15594), .ZN(n15587) );
  CLKBUF_X1 U12259 ( .A(n15110), .Z(n15600) );
  INV_X1 U12260 ( .A(n15608), .ZN(n15612) );
  OR2_X1 U12261 ( .A1(n15610), .A2(n12923), .ZN(n15608) );
  BUF_X1 U12262 ( .A(n20647), .Z(n21029) );
  NOR2_X1 U12263 ( .A1(n20619), .A2(n21029), .ZN(n20644) );
  BUF_X1 U12264 ( .A(n20644), .Z(n20646) );
  INV_X1 U12265 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15785) );
  NAND2_X1 U12266 ( .A1(n9891), .A2(n14587), .ZN(n15194) );
  OR2_X1 U12267 ( .A1(n9919), .A2(n9724), .ZN(n9891) );
  INV_X1 U12268 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21296) );
  INV_X1 U12269 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20559) );
  INV_X1 U12270 ( .A(n20516), .ZN(n16772) );
  XNOR2_X1 U12271 ( .A(n9901), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15835) );
  NAND2_X1 U12272 ( .A1(n9902), .A2(n9943), .ZN(n9901) );
  OAI21_X1 U12273 ( .B1(n15683), .B2(n9904), .A(n9903), .ZN(n9902) );
  NAND2_X1 U12274 ( .A1(n15676), .A2(n15858), .ZN(n9904) );
  NAND2_X1 U12275 ( .A1(n16767), .A2(n16768), .ZN(n10274) );
  NOR2_X1 U12276 ( .A1(n15224), .A2(n15914), .ZN(n15871) );
  INV_X1 U12277 ( .A(n15228), .ZN(n20658) );
  AND2_X1 U12278 ( .A1(n13117), .A2(n14742), .ZN(n20657) );
  AND2_X1 U12279 ( .A1(n13538), .A2(n14128), .ZN(n20663) );
  INV_X1 U12280 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13262) );
  NOR2_X1 U12281 ( .A1(n20695), .A2(n14546), .ZN(n20769) );
  OAI21_X1 U12282 ( .B1(n20785), .B2(n20784), .A(n20783), .ZN(n20803) );
  OAI211_X1 U12283 ( .C1(n12826), .C2(n14133), .A(n14129), .B(n20700), .ZN(
        n14162) );
  NOR2_X1 U12284 ( .A1(n14547), .A2(n13989), .ZN(n20925) );
  OAI211_X1 U12285 ( .C1(n14047), .C2(n14052), .A(n20818), .B(n20876), .ZN(
        n14074) );
  INV_X1 U12286 ( .A(n14007), .ZN(n20885) );
  INV_X1 U12287 ( .A(n13997), .ZN(n20891) );
  INV_X1 U12288 ( .A(n14016), .ZN(n20897) );
  INV_X1 U12289 ( .A(n13992), .ZN(n20909) );
  INV_X1 U12290 ( .A(n14027), .ZN(n20915) );
  INV_X1 U12291 ( .A(n14012), .ZN(n20921) );
  OAI211_X1 U12292 ( .C1(n15926), .C2(n14556), .A(n20744), .B(n14555), .ZN(
        n14578) );
  INV_X1 U12293 ( .A(n14021), .ZN(n20931) );
  NOR2_X1 U12295 ( .A1(n16943), .A2(n19656), .ZN(n15957) );
  NAND2_X1 U12296 ( .A1(n10925), .A2(n10114), .ZN(n15949) );
  NOR2_X1 U12297 ( .A1(n19656), .A2(n15962), .ZN(n16605) );
  NAND2_X1 U12298 ( .A1(n10878), .A2(n10877), .ZN(n15972) );
  OR2_X1 U12299 ( .A1(n10891), .A2(n10875), .ZN(n10894) );
  OR2_X1 U12300 ( .A1(n19557), .A2(n12023), .ZN(n19676) );
  NAND2_X1 U12301 ( .A1(n10853), .A2(n13302), .ZN(n10857) );
  INV_X1 U12302 ( .A(n19676), .ZN(n19697) );
  NOR2_X1 U12303 ( .A1(n12989), .A2(n11175), .ZN(n13353) );
  NAND2_X1 U12304 ( .A1(n10284), .A2(n19698), .ZN(n14508) );
  INV_X1 U12305 ( .A(n19698), .ZN(n19687) );
  AND2_X1 U12306 ( .A1(n19557), .A2(n12020), .ZN(n19671) );
  AND2_X1 U12307 ( .A1(n19819), .A2(n21150), .ZN(n19698) );
  AND3_X1 U12308 ( .A1(n11373), .A2(n11372), .A3(n11371), .ZN(n14175) );
  AND3_X1 U12309 ( .A1(n11283), .A2(n11282), .A3(n11281), .ZN(n13478) );
  INV_X1 U12310 ( .A(n13294), .ZN(n11606) );
  AND3_X1 U12311 ( .A1(n11212), .A2(n10336), .A3(n11211), .ZN(n13290) );
  CLKBUF_X1 U12312 ( .A(n13287), .Z(n13288) );
  AND2_X1 U12313 ( .A1(n19666), .A2(n11604), .ZN(n19665) );
  OAI21_X1 U12314 ( .B1(n16036), .B2(n16027), .A(n11906), .ZN(n16022) );
  XNOR2_X1 U12315 ( .A(n9862), .B(n11864), .ZN(n16042) );
  NAND2_X1 U12316 ( .A1(n11840), .A2(n16045), .ZN(n9862) );
  AND2_X1 U12317 ( .A1(n12959), .A2(n12694), .ZN(n19717) );
  INV_X1 U12318 ( .A(n19719), .ZN(n16156) );
  NAND2_X1 U12319 ( .A1(n19744), .A2(n11967), .ZN(n16155) );
  OR2_X1 U12320 ( .A1(n16973), .A2(n12959), .ZN(n19746) );
  AND2_X1 U12321 ( .A1(n19744), .A2(n10400), .ZN(n19772) );
  INV_X1 U12322 ( .A(n19821), .ZN(n12708) );
  NOR2_X1 U12323 ( .A1(n11521), .A2(n10250), .ZN(n10249) );
  NOR2_X1 U12324 ( .A1(n11527), .A2(n9758), .ZN(n10247) );
  NOR2_X1 U12325 ( .A1(n16483), .A2(n16484), .ZN(n16468) );
  INV_X1 U12326 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17036) );
  INV_X1 U12327 ( .A(n19848), .ZN(n16307) );
  XNOR2_X1 U12328 ( .A(n9841), .B(n11506), .ZN(n16163) );
  NAND2_X1 U12329 ( .A1(n10057), .A2(n10060), .ZN(n16303) );
  NAND2_X1 U12330 ( .A1(n16229), .A2(n10061), .ZN(n10057) );
  NAND2_X1 U12331 ( .A1(n16229), .A2(n16986), .ZN(n10065) );
  AND2_X1 U12332 ( .A1(n9989), .A2(n10078), .ZN(n16996) );
  NAND2_X1 U12333 ( .A1(n14431), .A2(n14433), .ZN(n10303) );
  CLKBUF_X1 U12334 ( .A(n14431), .Z(n14432) );
  INV_X1 U12335 ( .A(n10284), .ZN(n13359) );
  AND2_X1 U12336 ( .A1(n11482), .A2(n11405), .ZN(n19854) );
  INV_X1 U12337 ( .A(n16432), .ZN(n17054) );
  NAND2_X1 U12338 ( .A1(n12969), .A2(n12968), .ZN(n20487) );
  INV_X1 U12339 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20481) );
  INV_X1 U12340 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20463) );
  NAND2_X1 U12341 ( .A1(n12960), .A2(n12963), .ZN(n20478) );
  INV_X1 U12342 ( .A(n16552), .ZN(n16542) );
  XNOR2_X1 U12343 ( .A(n12991), .B(n12992), .ZN(n20466) );
  AOI21_X1 U12344 ( .B1(n10284), .B2(n13409), .A(n10285), .ZN(n16551) );
  NAND2_X1 U12345 ( .A1(n10286), .A2(n11273), .ZN(n10285) );
  INV_X1 U12346 ( .A(n13390), .ZN(n10286) );
  INV_X1 U12347 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21165) );
  INV_X1 U12348 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11842) );
  INV_X1 U12349 ( .A(n20370), .ZN(n19907) );
  OAI21_X1 U12350 ( .B1(n14260), .B2(n14263), .A(n14259), .ZN(n19911) );
  AND2_X1 U12351 ( .A1(n20067), .A2(n20454), .ZN(n20011) );
  NOR2_X2 U12352 ( .A1(n20316), .A2(n20041), .ZN(n20093) );
  OAI21_X1 U12353 ( .B1(n20124), .B2(n20103), .A(n20320), .ZN(n20126) );
  NOR2_X1 U12354 ( .A1(n20130), .A2(n20132), .ZN(n20167) );
  INV_X1 U12355 ( .A(n20330), .ZN(n20285) );
  INV_X1 U12356 ( .A(n20336), .ZN(n20288) );
  INV_X1 U12357 ( .A(n20342), .ZN(n20291) );
  INV_X1 U12358 ( .A(n20348), .ZN(n20294) );
  OAI21_X1 U12359 ( .B1(n13657), .B2(n13656), .A(n13655), .ZN(n20306) );
  INV_X1 U12360 ( .A(n20371), .ZN(n20304) );
  INV_X1 U12361 ( .A(n20176), .ZN(n20322) );
  INV_X1 U12362 ( .A(n20179), .ZN(n20327) );
  AND2_X1 U12363 ( .A1(n14265), .A2(n19904), .ZN(n20326) );
  INV_X1 U12364 ( .A(n20182), .ZN(n20333) );
  OAI22_X1 U12365 ( .A1(n19885), .A2(n19902), .B1(n21078), .B2(n19900), .ZN(
        n20339) );
  AND2_X1 U12366 ( .A1(n10479), .A2(n19904), .ZN(n20349) );
  INV_X1 U12367 ( .A(n20191), .ZN(n20351) );
  NOR2_X2 U12368 ( .A1(n20166), .A2(n20316), .ZN(n20366) );
  NOR3_X1 U12369 ( .A1(n13448), .A2(n13447), .A3(n13446), .ZN(n17101) );
  INV_X1 U12370 ( .A(n19555), .ZN(n19551) );
  NOR2_X1 U12371 ( .A1(n18122), .A2(n12333), .ZN(n17259) );
  AND2_X1 U12372 ( .A1(n10180), .A2(n9827), .ZN(n17286) );
  INV_X1 U12373 ( .A(n10188), .ZN(n17347) );
  AND2_X1 U12374 ( .A1(n10178), .A2(n17547), .ZN(n17380) );
  NOR2_X1 U12375 ( .A1(n17401), .A2(n10186), .ZN(n17390) );
  INV_X1 U12376 ( .A(n10178), .ZN(n17389) );
  INV_X1 U12377 ( .A(n17598), .ZN(n17605) );
  NOR2_X1 U12378 ( .A1(n19553), .A2(n19385), .ZN(n17600) );
  INV_X1 U12379 ( .A(n17620), .ZN(n17604) );
  INV_X1 U12380 ( .A(n17616), .ZN(n17615) );
  INV_X1 U12381 ( .A(n17388), .ZN(n17619) );
  AND2_X1 U12382 ( .A1(n17716), .A2(n10027), .ZN(n17685) );
  AND2_X1 U12383 ( .A1(n10028), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n10027) );
  NOR2_X1 U12384 ( .A1(n17808), .A2(n10033), .ZN(n17743) );
  NAND2_X1 U12385 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  INV_X1 U12386 ( .A(n10036), .ZN(n10035) );
  NOR2_X1 U12387 ( .A1(n17812), .A2(n17412), .ZN(n10034) );
  NOR2_X1 U12388 ( .A1(n17891), .A2(n10024), .ZN(n17838) );
  NOR3_X1 U12389 ( .A1(n17891), .A2(n10026), .A3(n17854), .ZN(n17852) );
  NOR2_X1 U12390 ( .A1(n17891), .A2(n17854), .ZN(n17853) );
  NOR3_X1 U12391 ( .A1(n17530), .A2(n17890), .A3(n17896), .ZN(n17895) );
  AND2_X1 U12392 ( .A1(n10042), .A2(n10041), .ZN(n17924) );
  NOR2_X1 U12393 ( .A1(n18893), .A2(n9799), .ZN(n10041) );
  NAND2_X1 U12394 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17936), .ZN(n17935) );
  NAND2_X1 U12395 ( .A1(n17954), .A2(n9743), .ZN(n17940) );
  NAND2_X1 U12396 ( .A1(n17954), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17950) );
  NOR2_X1 U12397 ( .A1(n21123), .A2(n17959), .ZN(n17954) );
  NOR2_X1 U12398 ( .A1(n17964), .A2(n17969), .ZN(n17960) );
  NAND2_X1 U12399 ( .A1(n17960), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17959) );
  NOR2_X1 U12400 ( .A1(n18002), .A2(n9914), .ZN(n17965) );
  NAND2_X1 U12401 ( .A1(n17965), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17964) );
  INV_X1 U12402 ( .A(n17985), .ZN(n17981) );
  OR3_X1 U12403 ( .A1(n17969), .A2(n18002), .A3(n18129), .ZN(n17995) );
  NAND2_X1 U12404 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18006), .ZN(n18002) );
  INV_X1 U12405 ( .A(n17994), .ZN(n18000) );
  INV_X1 U12406 ( .A(n17975), .ZN(n18001) );
  NOR2_X1 U12407 ( .A1(n18177), .A2(n18011), .ZN(n18006) );
  NOR2_X1 U12408 ( .A1(n18037), .A2(n9911), .ZN(n18012) );
  NAND2_X1 U12409 ( .A1(n18012), .A2(P3_EAX_REG_14__SCAN_IN), .ZN(n18011) );
  NOR2_X1 U12410 ( .A1(n12121), .A2(n12120), .ZN(n18041) );
  AND2_X1 U12411 ( .A1(n9913), .A2(n9912), .ZN(n18043) );
  NOR2_X1 U12412 ( .A1(n17925), .A2(n18040), .ZN(n9912) );
  NAND2_X1 U12413 ( .A1(n19359), .A2(n9913), .ZN(n18052) );
  NOR2_X1 U12414 ( .A1(n18058), .A2(n18929), .ZN(n18063) );
  AND3_X1 U12415 ( .A1(n12100), .A2(n12099), .A3(n12098), .ZN(n10319) );
  NOR2_X1 U12416 ( .A1(n12097), .A2(n12096), .ZN(n12099) );
  INV_X1 U12417 ( .A(n12135), .ZN(n9969) );
  INV_X1 U12418 ( .A(n18052), .ZN(n18067) );
  INV_X1 U12419 ( .A(n18180), .ZN(n18174) );
  NAND2_X1 U12421 ( .A1(n18255), .A2(n9734), .ZN(n18212) );
  OR2_X1 U12422 ( .A1(n18349), .A2(n10189), .ZN(n18336) );
  NAND2_X1 U12423 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10189) );
  NAND2_X1 U12424 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18374), .ZN(
        n18697) );
  INV_X1 U12425 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18457) );
  INV_X1 U12426 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18469) );
  INV_X1 U12427 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18492) );
  AND3_X1 U12428 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18493) );
  NAND2_X1 U12429 ( .A1(n17119), .A2(n9954), .ZN(n10082) );
  AND2_X1 U12430 ( .A1(n12162), .A2(n9778), .ZN(n18219) );
  INV_X1 U12431 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19393) );
  NOR2_X1 U12432 ( .A1(n18498), .A2(n18499), .ZN(n18497) );
  NOR2_X1 U12433 ( .A1(n19326), .A2(n18871), .ZN(n18868) );
  INV_X1 U12434 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19364) );
  INV_X1 U12435 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19366) );
  INV_X1 U12436 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19371) );
  INV_X1 U12437 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19419) );
  CLKBUF_X1 U12438 ( .A(n19480), .Z(n19474) );
  CLKBUF_X1 U12439 ( .A(n17239), .Z(n17245) );
  AOI21_X1 U12440 ( .B1(n15484), .B2(n20595), .A(n15293), .ZN(n15294) );
  AOI21_X1 U12441 ( .B1(n15534), .B2(n16764), .A(n15253), .ZN(n15254) );
  OAI21_X1 U12442 ( .B1(n15624), .B2(n16770), .A(n15623), .ZN(n15625) );
  NAND2_X1 U12443 ( .A1(n9927), .A2(n15244), .ZN(P1_U3000) );
  INV_X1 U12444 ( .A(n12014), .ZN(n12039) );
  NOR2_X1 U12445 ( .A1(n12037), .A2(n12036), .ZN(n12038) );
  AOI21_X1 U12446 ( .B1(n9753), .B2(n12013), .A(n19704), .ZN(n12014) );
  OAI21_X1 U12447 ( .B1(n19712), .B2(n10288), .A(n10287), .ZN(n13281) );
  INV_X1 U12448 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10288) );
  OR2_X1 U12449 ( .A1(n11488), .A2(n17039), .ZN(n11497) );
  NAND2_X1 U12450 ( .A1(n9720), .A2(n19828), .ZN(n12398) );
  NAND2_X1 U12451 ( .A1(n9840), .A2(n9838), .ZN(P2_U2986) );
  INV_X1 U12452 ( .A(n9839), .ZN(n9838) );
  NAND2_X1 U12453 ( .A1(n16163), .A2(n19828), .ZN(n9840) );
  OAI21_X1 U12454 ( .B1(n16170), .B2(n17039), .A(n16169), .ZN(n9839) );
  OAI211_X1 U12455 ( .C1(n17039), .C2(n16333), .A(n10050), .B(n10048), .ZN(
        P2_U2988) );
  AOI21_X1 U12456 ( .B1(n16330), .B2(n19848), .A(n16183), .ZN(n10050) );
  NAND2_X1 U12457 ( .A1(n10049), .A2(n19828), .ZN(n10048) );
  AOI21_X1 U12458 ( .B1(n17073), .B2(n11531), .A(n9883), .ZN(n16990) );
  NAND2_X1 U12459 ( .A1(n9885), .A2(n9884), .ZN(n9883) );
  NOR2_X1 U12460 ( .A1(n17043), .A2(n10289), .ZN(n17044) );
  NAND2_X1 U12461 ( .A1(n9794), .A2(n10290), .ZN(n10289) );
  INV_X1 U12462 ( .A(n11564), .ZN(n11565) );
  OR2_X1 U12463 ( .A1(n11488), .A2(n19859), .ZN(n11483) );
  NAND2_X1 U12464 ( .A1(n9720), .A2(n19866), .ZN(n12414) );
  OR2_X1 U12465 ( .A1(n16322), .A2(n16500), .ZN(n16332) );
  OAI21_X1 U12466 ( .B1(n16393), .B2(n16500), .A(n10071), .ZN(P2_U3026) );
  INV_X1 U12467 ( .A(n10072), .ZN(n10071) );
  OAI21_X1 U12468 ( .B1(n16403), .B2(n19859), .A(n16402), .ZN(n10072) );
  AOI21_X1 U12469 ( .B1(n17665), .B2(P3_EBX_REG_29__SCAN_IN), .A(n10022), .ZN(
        n17666) );
  AND2_X1 U12470 ( .A1(n17921), .A2(n17934), .ZN(n10022) );
  NAND2_X1 U12471 ( .A1(n17716), .A2(n10028), .ZN(n17701) );
  NAND2_X1 U12472 ( .A1(n17716), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n17702) );
  NOR2_X1 U12473 ( .A1(n17808), .A2(n17812), .ZN(n17784) );
  AOI21_X1 U12474 ( .B1(n17159), .B2(n18464), .A(n9948), .ZN(n17123) );
  NOR2_X1 U12475 ( .A1(n12041), .A2(n17603), .ZN(n12095) );
  INV_X2 U12476 ( .A(n14277), .ZN(n19656) );
  NAND2_X1 U12478 ( .A1(n11999), .A2(n9721), .ZN(n11997) );
  OR2_X1 U12479 ( .A1(n13662), .A2(n10296), .ZN(n9715) );
  OR2_X1 U12480 ( .A1(n10063), .A2(n16230), .ZN(n10060) );
  AND4_X1 U12481 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n9716)
         );
  INV_X1 U12482 ( .A(n15193), .ZN(n15782) );
  INV_X1 U12483 ( .A(n10573), .ZN(n10574) );
  INV_X1 U12484 ( .A(n11766), .ZN(n10573) );
  NAND2_X1 U12485 ( .A1(n9995), .A2(n10304), .ZN(n16466) );
  OR3_X1 U12486 ( .A1(n15469), .A2(n10166), .A3(n15883), .ZN(n9717) );
  NAND2_X1 U12487 ( .A1(n10868), .A2(n10105), .ZN(n9718) );
  AND2_X1 U12488 ( .A1(n9995), .A2(n9994), .ZN(n16254) );
  NOR2_X1 U12489 ( .A1(n10212), .A2(n10213), .ZN(n15465) );
  OR2_X1 U12490 ( .A1(n16172), .A2(n10310), .ZN(n9719) );
  AND2_X1 U12491 ( .A1(n15338), .A2(n9810), .ZN(n15103) );
  XNOR2_X1 U12492 ( .A(n12397), .B(n12396), .ZN(n9720) );
  AND2_X1 U12493 ( .A1(n10154), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9721) );
  OR2_X1 U12494 ( .A1(n9824), .A2(n16484), .ZN(n9723) );
  AND2_X1 U12495 ( .A1(n14585), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9724) );
  INV_X2 U12496 ( .A(n13429), .ZN(n11024) );
  NAND2_X1 U12497 ( .A1(n14594), .A2(n9796), .ZN(n14624) );
  OR3_X1 U12498 ( .A1(n15983), .A2(n10233), .A3(n10236), .ZN(n9725) );
  AND2_X1 U12499 ( .A1(n10111), .A2(n10790), .ZN(n9726) );
  INV_X1 U12500 ( .A(n10208), .ZN(n15441) );
  AND2_X1 U12501 ( .A1(n13519), .A2(n9937), .ZN(n9727) );
  AND2_X1 U12502 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9728) );
  INV_X1 U12503 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18350) );
  AND2_X1 U12504 ( .A1(n10228), .A2(n9802), .ZN(n9729) );
  NAND2_X1 U12505 ( .A1(n18499), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9730) );
  AND2_X1 U12506 ( .A1(n14641), .A2(n9820), .ZN(n9731) );
  AND2_X1 U12507 ( .A1(n10065), .A2(n16987), .ZN(n9732) );
  AND3_X2 U12508 ( .A1(n10679), .A2(n10678), .A3(n10677), .ZN(n11189) );
  NAND2_X1 U12509 ( .A1(n14236), .A2(n14235), .ZN(n9733) );
  NOR2_X1 U12511 ( .A1(n13662), .A2(n9814), .ZN(n14329) );
  NOR2_X1 U12512 ( .A1(n13294), .A2(n10299), .ZN(n13464) );
  INV_X1 U12513 ( .A(n11459), .ZN(n13671) );
  AND2_X1 U12514 ( .A1(n12361), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9734) );
  AND2_X1 U12515 ( .A1(n10157), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9735) );
  OR2_X1 U12516 ( .A1(n10299), .A2(n10298), .ZN(n9736) );
  AND2_X1 U12517 ( .A1(n9734), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9737) );
  AND2_X1 U12518 ( .A1(n10238), .A2(n10237), .ZN(n9738) );
  AND2_X1 U12519 ( .A1(n10141), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9739) );
  NAND2_X1 U12520 ( .A1(n10578), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13393) );
  AND2_X1 U12521 ( .A1(n11982), .A2(n10149), .ZN(n9740) );
  NOR2_X1 U12522 ( .A1(n16021), .A2(n16028), .ZN(n9741) );
  AND4_X1 U12523 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(P3_EAX_REG_8__SCAN_IN), .ZN(n9742) );
  AND2_X1 U12524 ( .A1(n9907), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9743) );
  AND2_X1 U12525 ( .A1(n10312), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9744) );
  AND2_X1 U12526 ( .A1(n9997), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9745) );
  INV_X1 U12527 ( .A(n11722), .ZN(n10829) );
  INV_X1 U12528 ( .A(n10585), .ZN(n11876) );
  NAND2_X1 U12529 ( .A1(n10307), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16205) );
  NAND2_X1 U12530 ( .A1(n15724), .A2(n15723), .ZN(n15699) );
  OR2_X1 U12531 ( .A1(n10947), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n9748) );
  AND2_X1 U12532 ( .A1(n10937), .A2(n9843), .ZN(n16178) );
  OR2_X1 U12533 ( .A1(n10891), .A2(n10116), .ZN(n9749) );
  XNOR2_X1 U12534 ( .A(n17126), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12362) );
  NAND2_X1 U12535 ( .A1(n10311), .A2(n10312), .ZN(n16276) );
  INV_X1 U12536 ( .A(n12395), .ZN(n10250) );
  NAND2_X1 U12537 ( .A1(n9890), .A2(n9892), .ZN(n15778) );
  NOR2_X1 U12538 ( .A1(n16224), .A2(n10308), .ZN(n16193) );
  NOR2_X1 U12539 ( .A1(n12002), .A2(n17036), .ZN(n11999) );
  AND3_X1 U12540 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12000) );
  AND2_X1 U12541 ( .A1(n11999), .A2(n10154), .ZN(n9750) );
  AND2_X1 U12542 ( .A1(n10307), .A2(n9745), .ZN(n9751) );
  INV_X1 U12543 ( .A(n9852), .ZN(n9859) );
  OAI211_X1 U12544 ( .C1(n11840), .C2(n9856), .A(n9855), .B(n9853), .ZN(n9852)
         );
  OR3_X1 U12545 ( .A1(n10891), .A2(n10893), .A3(n10875), .ZN(n9752) );
  INV_X1 U12546 ( .A(n11100), .ZN(n11042) );
  INV_X1 U12547 ( .A(n17121), .ZN(n9954) );
  NOR2_X1 U12548 ( .A1(n16897), .A2(n19656), .ZN(n9753) );
  NOR2_X2 U12549 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10586) );
  AND4_X1 U12550 ( .A1(n12547), .A2(n12546), .A3(n12545), .A4(n12544), .ZN(
        n9755) );
  AND3_X1 U12551 ( .A1(n12764), .A2(n12975), .A3(n12772), .ZN(n9756) );
  NOR2_X1 U12552 ( .A1(n11446), .A2(n11966), .ZN(n9757) );
  NAND2_X1 U12553 ( .A1(n15778), .A2(n15195), .ZN(n15731) );
  OR2_X1 U12554 ( .A1(n11520), .A2(n11519), .ZN(n9758) );
  NAND2_X1 U12555 ( .A1(n16052), .A2(n10292), .ZN(n16954) );
  INV_X1 U12556 ( .A(n18047), .ZN(n12125) );
  NOR2_X1 U12557 ( .A1(n12111), .A2(n12110), .ZN(n18047) );
  NAND2_X1 U12558 ( .A1(n10203), .A2(n10201), .ZN(n13173) );
  AND3_X1 U12559 ( .A1(n12437), .A2(n12445), .A3(n9929), .ZN(n9759) );
  NOR2_X1 U12560 ( .A1(n10384), .A2(n10283), .ZN(n10459) );
  AND4_X1 U12561 ( .A1(n10337), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(
        n9760) );
  OR2_X1 U12562 ( .A1(n16295), .A2(n16427), .ZN(n9761) );
  NAND2_X1 U12563 ( .A1(n10303), .A2(n11480), .ZN(n16502) );
  INV_X1 U12564 ( .A(n10327), .ZN(n10078) );
  AND3_X1 U12565 ( .A1(n9889), .A2(n9888), .A3(n9887), .ZN(n9762) );
  OR2_X1 U12566 ( .A1(n9706), .A2(n14520), .ZN(n10566) );
  NAND2_X1 U12567 ( .A1(n10988), .A2(n10485), .ZN(n10492) );
  INV_X1 U12568 ( .A(n10492), .ZN(n10486) );
  NAND2_X1 U12569 ( .A1(n14835), .A2(n10209), .ZN(n10208) );
  NAND2_X1 U12570 ( .A1(n10311), .A2(n9744), .ZN(n10314) );
  INV_X1 U12571 ( .A(n16295), .ZN(n10311) );
  OR2_X1 U12572 ( .A1(n11412), .A2(n17100), .ZN(n9763) );
  AND2_X1 U12573 ( .A1(n14400), .A2(n14399), .ZN(n9764) );
  INV_X1 U12574 ( .A(n11480), .ZN(n10306) );
  OAI211_X1 U12575 ( .C1(n11577), .C2(n11588), .A(n11587), .B(n11586), .ZN(
        n12992) );
  NAND2_X1 U12576 ( .A1(n10858), .A2(n10945), .ZN(n10868) );
  NAND2_X1 U12577 ( .A1(n14835), .A2(n14834), .ZN(n15454) );
  XOR2_X1 U12578 ( .A(n11530), .B(n11529), .Z(n9765) );
  INV_X1 U12579 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11865) );
  AND2_X1 U12580 ( .A1(n12815), .A2(n12761), .ZN(n9766) );
  AND2_X1 U12581 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n9767) );
  AND2_X1 U12582 ( .A1(n15209), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9768) );
  OR2_X1 U12583 ( .A1(n15213), .A2(n15209), .ZN(n9943) );
  OR2_X1 U12584 ( .A1(n16194), .A2(n16339), .ZN(n9769) );
  NAND2_X1 U12585 ( .A1(n10195), .A2(n14624), .ZN(n9770) );
  NAND2_X1 U12586 ( .A1(n11149), .A2(n9699), .ZN(n9771) );
  NAND2_X1 U12587 ( .A1(n10868), .A2(n10867), .ZN(n10872) );
  INV_X1 U12588 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18360) );
  NAND2_X1 U12589 ( .A1(n9850), .A2(n14434), .ZN(n16503) );
  OR2_X1 U12590 ( .A1(n15937), .A2(n16090), .ZN(n9772) );
  OR2_X1 U12591 ( .A1(n15214), .A2(n15826), .ZN(n9773) );
  AND2_X1 U12592 ( .A1(n12188), .A2(n12189), .ZN(n9774) );
  AND2_X1 U12593 ( .A1(n10783), .A2(n10785), .ZN(n9775) );
  AND2_X1 U12594 ( .A1(n10184), .A2(n17547), .ZN(n9776) );
  AND2_X1 U12595 ( .A1(n10130), .A2(n10129), .ZN(n9777) );
  INV_X1 U12596 ( .A(n11582), .ZN(n10525) );
  INV_X1 U12597 ( .A(n16762), .ZN(n10273) );
  AND2_X1 U12598 ( .A1(n12161), .A2(n12160), .ZN(n9778) );
  AND2_X1 U12599 ( .A1(n9994), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9779) );
  NAND2_X1 U12600 ( .A1(n9875), .A2(n11468), .ZN(n11472) );
  AND2_X1 U12601 ( .A1(n9897), .A2(n9896), .ZN(n9780) );
  AND2_X1 U12602 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U12603 ( .A1(n10334), .A2(n10255), .ZN(n9782) );
  CLKBUF_X1 U12604 ( .A(n13960), .Z(n15035) );
  CLKBUF_X3 U12605 ( .A(n13700), .Z(n14930) );
  NAND2_X1 U12606 ( .A1(n16682), .A2(n19535), .ZN(n18058) );
  INV_X1 U12607 ( .A(n18058), .ZN(n9913) );
  NOR2_X1 U12608 ( .A1(n10002), .A2(n10001), .ZN(n12810) );
  INV_X1 U12609 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12434) );
  INV_X1 U12610 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U12611 ( .A1(n14271), .A2(n10219), .ZN(n11376) );
  NOR2_X1 U12612 ( .A1(n11989), .A2(n11988), .ZN(n9783) );
  OR3_X1 U12613 ( .A1(n17891), .A2(n10024), .A3(n10023), .ZN(n9784) );
  NAND2_X1 U12614 ( .A1(n12960), .A2(n11576), .ZN(n12991) );
  NAND2_X1 U12615 ( .A1(n10791), .A2(n9726), .ZN(n10844) );
  NOR2_X1 U12616 ( .A1(n12007), .A2(n16285), .ZN(n11992) );
  NOR2_X1 U12617 ( .A1(n13662), .A2(n14175), .ZN(n14081) );
  NAND2_X1 U12618 ( .A1(n16074), .A2(n16073), .ZN(n15991) );
  NAND2_X1 U12619 ( .A1(n18440), .A2(n10090), .ZN(n9785) );
  NOR2_X1 U12620 ( .A1(n12004), .A2(n17006), .ZN(n11996) );
  AND2_X1 U12621 ( .A1(n11999), .A2(n10153), .ZN(n11998) );
  AND2_X1 U12622 ( .A1(n11996), .A2(n10157), .ZN(n11995) );
  NAND2_X1 U12623 ( .A1(n15456), .A2(n15444), .ZN(n15429) );
  AND2_X1 U12624 ( .A1(n17716), .A2(n10030), .ZN(n9786) );
  AND2_X1 U12625 ( .A1(n17954), .A2(n9907), .ZN(n9787) );
  AND2_X1 U12626 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9788) );
  AND2_X1 U12627 ( .A1(n10209), .A2(n15440), .ZN(n9789) );
  AND2_X1 U12628 ( .A1(n10125), .A2(n13664), .ZN(n9790) );
  AND2_X1 U12629 ( .A1(n9790), .A2(n10123), .ZN(n9791) );
  NAND2_X1 U12630 ( .A1(n12961), .A2(n12962), .ZN(n12960) );
  NAND2_X1 U12631 ( .A1(n9871), .A2(n10294), .ZN(n16071) );
  NOR2_X1 U12632 ( .A1(n13504), .A2(n13503), .ZN(n13505) );
  AND2_X1 U12633 ( .A1(n14321), .A2(n9738), .ZN(n9792) );
  INV_X1 U12634 ( .A(n13467), .ZN(n10298) );
  AND2_X1 U12635 ( .A1(n11457), .A2(n21051), .ZN(n13669) );
  AND2_X1 U12636 ( .A1(n11490), .A2(n10143), .ZN(n9793) );
  INV_X1 U12637 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20470) );
  NAND2_X1 U12638 ( .A1(n9978), .A2(n10794), .ZN(n14036) );
  OR3_X1 U12639 ( .A1(n17041), .A2(n17040), .A3(n17039), .ZN(n9794) );
  INV_X1 U12640 ( .A(n16215), .ZN(n10252) );
  AND2_X1 U12641 ( .A1(n10223), .A2(n14468), .ZN(n9795) );
  INV_X1 U12642 ( .A(n16994), .ZN(n10255) );
  XNOR2_X1 U12643 ( .A(n11472), .B(n11473), .ZN(n14291) );
  INV_X1 U12644 ( .A(n10843), .ZN(n10110) );
  NAND2_X1 U12645 ( .A1(n13361), .A2(n11453), .ZN(n13484) );
  NAND2_X1 U12646 ( .A1(n10274), .A2(n14405), .ZN(n16760) );
  AND2_X1 U12647 ( .A1(n14593), .A2(n10199), .ZN(n9796) );
  INV_X1 U12648 ( .A(n16993), .ZN(n10076) );
  AND2_X1 U12649 ( .A1(n10045), .A2(n11455), .ZN(n9797) );
  AND2_X1 U12650 ( .A1(n11996), .A2(n10156), .ZN(n11994) );
  AND2_X1 U12651 ( .A1(n10660), .A2(n10600), .ZN(n9798) );
  OR2_X1 U12652 ( .A1(n19539), .A2(n19391), .ZN(n9799) );
  OR2_X1 U12653 ( .A1(n15469), .A2(n10166), .ZN(n9800) );
  OR2_X1 U12654 ( .A1(n15972), .A2(n10918), .ZN(n9801) );
  NAND2_X1 U12655 ( .A1(n13564), .A2(n13577), .ZN(n15108) );
  INV_X1 U12656 ( .A(n15108), .ZN(n9937) );
  INV_X1 U12657 ( .A(n10062), .ZN(n10061) );
  NAND2_X1 U12658 ( .A1(n16979), .A2(n16986), .ZN(n10062) );
  NOR2_X1 U12659 ( .A1(n15983), .A2(n10230), .ZN(n10235) );
  AND2_X1 U12660 ( .A1(n10227), .A2(n13680), .ZN(n9802) );
  AND2_X1 U12661 ( .A1(n9788), .A2(n10332), .ZN(n9803) );
  INV_X1 U12662 ( .A(n11090), .ZN(n16011) );
  NOR2_X1 U12663 ( .A1(n13504), .A2(n10121), .ZN(n11090) );
  AND2_X1 U12664 ( .A1(n15011), .A2(n10217), .ZN(n9804) );
  AND2_X1 U12665 ( .A1(n18440), .A2(n18435), .ZN(n9805) );
  OR2_X1 U12666 ( .A1(n18382), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9806) );
  NOR2_X1 U12667 ( .A1(n12967), .A2(n21165), .ZN(n9807) );
  AND2_X1 U12668 ( .A1(n10188), .A2(n10187), .ZN(n9808) );
  AND2_X1 U12669 ( .A1(n9789), .A2(n10207), .ZN(n9809) );
  AOI21_X1 U12670 ( .B1(n16944), .B2(n16007), .A(n10138), .ZN(n10137) );
  AND2_X1 U12671 ( .A1(n10216), .A2(n10215), .ZN(n9810) );
  AND2_X1 U12672 ( .A1(n9737), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9811) );
  NOR2_X1 U12673 ( .A1(n11175), .A2(n10229), .ZN(n10228) );
  NAND2_X1 U12674 ( .A1(n19666), .A2(n9788), .ZN(n13127) );
  NAND2_X1 U12675 ( .A1(n21165), .A2(n11006), .ZN(n9812) );
  NOR2_X1 U12676 ( .A1(n16856), .A2(n16855), .ZN(n9813) );
  INV_X1 U12677 ( .A(n19866), .ZN(n16500) );
  AND2_X1 U12678 ( .A1(n11482), .A2(n20495), .ZN(n19866) );
  NAND2_X1 U12679 ( .A1(n11982), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11981) );
  NAND2_X1 U12680 ( .A1(n11606), .A2(n11605), .ZN(n13311) );
  NAND2_X1 U12681 ( .A1(n18255), .A2(n9737), .ZN(n10179) );
  OR2_X1 U12682 ( .A1(n13084), .A2(n13083), .ZN(n20653) );
  INV_X1 U12683 ( .A(n20653), .ZN(n16861) );
  OR2_X1 U12684 ( .A1(n10296), .A2(n14330), .ZN(n9814) );
  AND2_X1 U12685 ( .A1(n10171), .A2(n15444), .ZN(n9815) );
  AND2_X1 U12686 ( .A1(n9815), .A2(n10170), .ZN(n9816) );
  OR2_X1 U12687 ( .A1(n10127), .A2(n11507), .ZN(n9817) );
  INV_X1 U12688 ( .A(n18463), .ZN(n18382) );
  AND2_X1 U12689 ( .A1(n18435), .A2(n18413), .ZN(n9818) );
  OR3_X1 U12690 ( .A1(n11815), .A2(n16955), .A3(n11814), .ZN(n9819) );
  AND2_X1 U12691 ( .A1(n10211), .A2(n15521), .ZN(n9820) );
  AND2_X1 U12692 ( .A1(n15375), .A2(n15359), .ZN(n9821) );
  AND2_X1 U12693 ( .A1(n16957), .A2(n16053), .ZN(n9822) );
  INV_X1 U12694 ( .A(n10924), .ZN(n10115) );
  AND2_X1 U12695 ( .A1(n11864), .A2(n16041), .ZN(n9823) );
  NAND2_X1 U12696 ( .A1(n11884), .A2(n11862), .ZN(n11864) );
  AND2_X1 U12697 ( .A1(n10862), .A2(n16478), .ZN(n9824) );
  NAND2_X1 U12698 ( .A1(n11982), .A2(n10147), .ZN(n10152) );
  NAND2_X1 U12699 ( .A1(n10163), .A2(n10162), .ZN(n16833) );
  INV_X1 U12700 ( .A(n16833), .ZN(n10161) );
  INV_X1 U12701 ( .A(n12164), .ZN(n10088) );
  NOR2_X1 U12702 ( .A1(n18382), .A2(n12303), .ZN(n12164) );
  AND2_X1 U12703 ( .A1(n14833), .A2(n14832), .ZN(n15505) );
  INV_X1 U12704 ( .A(n13507), .ZN(n9872) );
  NOR2_X1 U12705 ( .A1(n11924), .A2(n11923), .ZN(n9825) );
  INV_X1 U12706 ( .A(n10032), .ZN(n17782) );
  NOR3_X1 U12707 ( .A1(n17808), .A2(n10036), .A3(n17812), .ZN(n10032) );
  NAND2_X1 U12708 ( .A1(n14481), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9826) );
  INV_X1 U12709 ( .A(n10148), .ZN(n10147) );
  NAND2_X1 U12710 ( .A1(n10149), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10148) );
  AND2_X1 U12711 ( .A1(n10181), .A2(n17547), .ZN(n9827) );
  AND2_X1 U12712 ( .A1(n10173), .A2(n10172), .ZN(n9828) );
  AND2_X1 U12713 ( .A1(n9816), .A2(n10169), .ZN(n9829) );
  AND2_X1 U12714 ( .A1(n9738), .A2(n15995), .ZN(n9830) );
  INV_X1 U12715 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10104) );
  INV_X1 U12716 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10008) );
  INV_X1 U12717 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10144) );
  NOR2_X2 U12718 ( .A1(n12227), .A2(n12226), .ZN(n18929) );
  AND2_X1 U12720 ( .A1(n11982), .A2(n10146), .ZN(n11542) );
  OR2_X1 U12721 ( .A1(n17918), .A2(n17660), .ZN(n9831) );
  INV_X1 U12722 ( .A(n14598), .ZN(n10199) );
  INV_X1 U12723 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n10026) );
  INV_X1 U12724 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10102) );
  AND2_X1 U12725 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n9744), .ZN(
        n9832) );
  INV_X1 U12726 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10145) );
  NOR2_X1 U12727 ( .A1(n10308), .A2(n16195), .ZN(n9833) );
  AND2_X1 U12728 ( .A1(n21206), .A2(n16786), .ZN(n9834) );
  AND2_X1 U12729 ( .A1(n15208), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9835) );
  INV_X1 U12731 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10155) );
  INV_X1 U12732 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10313) );
  INV_X1 U12733 ( .A(n16323), .ZN(n9998) );
  AND2_X1 U12734 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .ZN(n9837) );
  INV_X1 U12735 ( .A(n15639), .ZN(n9942) );
  INV_X1 U12736 ( .A(n17591), .ZN(n19399) );
  INV_X1 U12737 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19503) );
  AND2_X2 U12738 ( .A1(n9874), .A2(n11768), .ZN(n11742) );
  NOR2_X1 U12739 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11768) );
  AND2_X1 U12740 ( .A1(n10345), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9874) );
  NAND4_X1 U12741 ( .A1(n18833), .A2(n19551), .A3(n19399), .A4(n19389), .ZN(
        n17620) );
  OAI22_X2 U12742 ( .A1(n17189), .A2(n13592), .B1(n13556), .B2(n13593), .ZN(
        n20893) );
  OAI22_X2 U12743 ( .A1(n17182), .A2(n13592), .B1(n13563), .B2(n13593), .ZN(
        n20917) );
  OAI22_X2 U12744 ( .A1(n13576), .A2(n13593), .B1(n17180), .B2(n13592), .ZN(
        n20924) );
  OAI22_X2 U12745 ( .A1(n21227), .A2(n13592), .B1(n21176), .B2(n13593), .ZN(
        n20875) );
  OAI22_X2 U12746 ( .A1(n21269), .A2(n13592), .B1(n13543), .B2(n13593), .ZN(
        n20905) );
  OAI22_X2 U12747 ( .A1(n17187), .A2(n13592), .B1(n13569), .B2(n13593), .ZN(
        n20899) );
  OAI22_X2 U12748 ( .A1(n13594), .A2(n13593), .B1(n17184), .B2(n13592), .ZN(
        n20911) );
  NOR4_X2 U12749 ( .A1(n20527), .A2(n20526), .A3(n20525), .A4(n20524), .ZN(
        n21020) );
  AOI22_X2 U12750 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19407), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19419), .ZN(n19489) );
  OAI22_X2 U12751 ( .A1(n13585), .A2(n13593), .B1(n17191), .B2(n13592), .ZN(
        n20887) );
  NOR4_X2 U12752 ( .A1(n17269), .A2(n17268), .A3(n17267), .A4(n17266), .ZN(
        n19530) );
  NOR2_X2 U12753 ( .A1(n10474), .A2(n19890), .ZN(n20343) );
  OAI22_X2 U12754 ( .A1(n16171), .A2(n16312), .B1(n11504), .B2(n11503), .ZN(
        n9841) );
  XNOR2_X2 U12755 ( .A(n11469), .B(n11470), .ZN(n11466) );
  NAND2_X2 U12756 ( .A1(n11500), .A2(n11499), .ZN(n11502) );
  NAND4_X1 U12757 ( .A1(n10572), .A2(n10571), .A3(n10569), .A4(n10570), .ZN(
        n9844) );
  NAND3_X1 U12758 ( .A1(n9844), .A2(n10661), .A3(n9798), .ZN(n11455) );
  NAND2_X1 U12759 ( .A1(n9844), .A2(n10600), .ZN(n10046) );
  INV_X1 U12760 ( .A(n9846), .ZN(n9845) );
  OAI21_X1 U12761 ( .B1(n12622), .B2(n13445), .A(n9847), .ZN(n9846) );
  NAND4_X1 U12762 ( .A1(n11947), .A2(n10465), .A3(n10466), .A4(n10464), .ZN(
        n9847) );
  NAND2_X2 U12763 ( .A1(n10472), .A2(n11024), .ZN(n11022) );
  NAND2_X1 U12764 ( .A1(n10469), .A2(n11140), .ZN(n10505) );
  NAND2_X1 U12765 ( .A1(n9850), .A2(n10258), .ZN(n16483) );
  NAND3_X1 U12766 ( .A1(n16045), .A2(n11840), .A3(n9860), .ZN(n9855) );
  INV_X1 U12767 ( .A(n11864), .ZN(n9861) );
  NAND2_X2 U12768 ( .A1(n10542), .A2(n10540), .ZN(n15264) );
  NAND2_X2 U12769 ( .A1(n10503), .A2(n10502), .ZN(n10542) );
  NAND2_X2 U12770 ( .A1(n10489), .A2(n9863), .ZN(n10516) );
  NAND2_X1 U12771 ( .A1(n9864), .A2(n10423), .ZN(n10491) );
  NAND2_X1 U12772 ( .A1(n11414), .A2(n11416), .ZN(n9864) );
  NAND2_X1 U12773 ( .A1(n11413), .A2(n9867), .ZN(n9866) );
  AND2_X2 U12774 ( .A1(n10070), .A2(n13445), .ZN(n9974) );
  NAND2_X1 U12775 ( .A1(n9870), .A2(n9869), .ZN(n11946) );
  NAND2_X1 U12776 ( .A1(n16036), .A2(n9741), .ZN(n9869) );
  NOR2_X2 U12777 ( .A1(n13287), .A2(n13290), .ZN(n13289) );
  NAND2_X2 U12778 ( .A1(n11603), .A2(n11602), .ZN(n19666) );
  AOI21_X2 U12779 ( .B1(n16054), .B2(n9822), .A(n9873), .ZN(n11838) );
  OAI21_X2 U12780 ( .B1(n10292), .B2(n10291), .A(n9819), .ZN(n9873) );
  XNOR2_X2 U12781 ( .A(n11794), .B(n11815), .ZN(n16054) );
  XNOR2_X2 U12782 ( .A(n11838), .B(n10315), .ZN(n16047) );
  AND2_X2 U12783 ( .A1(n16060), .A2(n10316), .ZN(n11794) );
  NAND2_X2 U12784 ( .A1(n9874), .A2(n10346), .ZN(n10387) );
  AND2_X4 U12785 ( .A1(n9874), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10591) );
  NAND2_X1 U12786 ( .A1(n14291), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11476) );
  NAND2_X1 U12787 ( .A1(n14035), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9875) );
  AND2_X1 U12788 ( .A1(n9877), .A2(n9878), .ZN(n9876) );
  NAND2_X2 U12789 ( .A1(n9879), .A2(n9882), .ZN(n11046) );
  NAND2_X1 U12790 ( .A1(n9880), .A2(n11577), .ZN(n9879) );
  NAND2_X1 U12791 ( .A1(n11582), .A2(n9881), .ZN(n9880) );
  XNOR2_X2 U12792 ( .A(n11046), .B(n11047), .ZN(n11595) );
  OR2_X2 U12793 ( .A1(n19869), .A2(n11595), .ZN(n10565) );
  OR2_X2 U12794 ( .A1(n13192), .A2(n13193), .ZN(n13254) );
  XNOR2_X1 U12795 ( .A(n13191), .B(n13190), .ZN(n13192) );
  NAND3_X1 U12796 ( .A1(n12442), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A3(
        n12868), .ZN(n9888) );
  NAND3_X1 U12797 ( .A1(n12868), .A2(n12777), .A3(n9781), .ZN(n9887) );
  AND3_X2 U12798 ( .A1(n12868), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n12777), .ZN(n15074) );
  AND2_X2 U12799 ( .A1(n12435), .A2(n12869), .ZN(n15059) );
  NAND3_X1 U12800 ( .A1(n12435), .A2(n12869), .A3(
        P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U12801 ( .A1(n9919), .A2(n14587), .ZN(n9890) );
  NAND2_X1 U12802 ( .A1(n9894), .A2(n15778), .ZN(n9893) );
  NAND2_X1 U12803 ( .A1(n9893), .A2(n10004), .ZN(n15690) );
  NAND3_X1 U12804 ( .A1(n12598), .A2(n12600), .A3(n12599), .ZN(n12766) );
  NOR2_X1 U12805 ( .A1(n9764), .A2(n14401), .ZN(n9899) );
  NAND2_X1 U12806 ( .A1(n12567), .A2(n12568), .ZN(n10192) );
  NAND4_X2 U12807 ( .A1(n9900), .A2(n10003), .A3(n13832), .A4(n12597), .ZN(
        n12767) );
  INV_X1 U12808 ( .A(n10192), .ZN(n9900) );
  NAND2_X1 U12809 ( .A1(n9714), .A2(n15670), .ZN(n9903) );
  OR2_X1 U12810 ( .A1(n15213), .A2(n15639), .ZN(n9941) );
  NAND3_X1 U12811 ( .A1(n9742), .A2(P3_EAX_REG_10__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .ZN(n9911) );
  NAND3_X1 U12812 ( .A1(n9716), .A2(P3_EAX_REG_19__SCAN_IN), .A3(
        P3_EAX_REG_22__SCAN_IN), .ZN(n9914) );
  NAND4_X1 U12813 ( .A1(n9915), .A2(n12194), .A3(n12193), .A4(n9774), .ZN(
        n17926) );
  NAND3_X1 U12814 ( .A1(n12190), .A2(n12191), .A3(n9917), .ZN(n9916) );
  INV_X2 U12815 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12306) );
  INV_X1 U12816 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9918) );
  AND2_X2 U12817 ( .A1(n12441), .A2(n13533), .ZN(n15084) );
  XNOR2_X1 U12818 ( .A(n9919), .B(n14539), .ZN(n16847) );
  NAND2_X1 U12819 ( .A1(n14529), .A2(n14528), .ZN(n9919) );
  NAND2_X1 U12820 ( .A1(n9923), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U12821 ( .A1(n9920), .A2(n12776), .ZN(n10000) );
  NAND2_X1 U12822 ( .A1(n9923), .A2(n9921), .ZN(n9920) );
  INV_X1 U12823 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n9922) );
  NAND4_X1 U12824 ( .A1(n9925), .A2(n13082), .A3(n9924), .A4(n12762), .ZN(
        n9923) );
  INV_X1 U12825 ( .A(n12773), .ZN(n9926) );
  NAND3_X1 U12826 ( .A1(n10260), .A2(n9928), .A3(n10261), .ZN(n9927) );
  AND2_X1 U12827 ( .A1(n10259), .A2(n16861), .ZN(n9928) );
  NAND2_X1 U12828 ( .A1(n13254), .A2(n9933), .ZN(n13202) );
  AND2_X1 U12829 ( .A1(n9934), .A2(n14530), .ZN(n9933) );
  NAND2_X1 U12830 ( .A1(n13193), .A2(n13192), .ZN(n9934) );
  NAND2_X1 U12831 ( .A1(n9936), .A2(n9935), .ZN(n15698) );
  NAND2_X1 U12832 ( .A1(n15214), .A2(n15658), .ZN(n15647) );
  OR2_X1 U12833 ( .A1(n15213), .A2(n9940), .ZN(n9939) );
  OAI21_X1 U12834 ( .B1(n17120), .B2(n9952), .A(n9951), .ZN(n9950) );
  OAI21_X1 U12835 ( .B1(n17121), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n9958), .ZN(n9957) );
  INV_X1 U12836 ( .A(n17122), .ZN(n9958) );
  INV_X1 U12837 ( .A(n17120), .ZN(n9959) );
  NAND4_X1 U12838 ( .A1(n9969), .A2(n12133), .A3(n12137), .A4(n9965), .ZN(
        n16683) );
  NAND4_X1 U12839 ( .A1(n12134), .A2(n12132), .A3(n12136), .A4(n9967), .ZN(
        n9966) );
  NAND2_X2 U12840 ( .A1(n12151), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18729) );
  INV_X2 U12841 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19522) );
  AND2_X2 U12842 ( .A1(n9973), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10052) );
  INV_X1 U12843 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9973) );
  NOR2_X1 U12844 ( .A1(n13403), .A2(n9974), .ZN(n13423) );
  NAND2_X1 U12845 ( .A1(n10067), .A2(n9975), .ZN(n14436) );
  NAND2_X1 U12846 ( .A1(n9978), .A2(n9976), .ZN(n9975) );
  NAND2_X1 U12847 ( .A1(n13667), .A2(n13668), .ZN(n9978) );
  NAND3_X1 U12848 ( .A1(n10045), .A2(n11455), .A3(n11189), .ZN(n9979) );
  NAND2_X1 U12849 ( .A1(n9982), .A2(n9981), .ZN(n11522) );
  INV_X1 U12850 ( .A(n10565), .ZN(n10079) );
  INV_X1 U12851 ( .A(n14431), .ZN(n9996) );
  AND2_X2 U12852 ( .A1(n9995), .A2(n9779), .ZN(n16227) );
  NAND2_X2 U12853 ( .A1(n9996), .A2(n11480), .ZN(n9995) );
  NAND2_X1 U12854 ( .A1(n10307), .A2(n9833), .ZN(n16194) );
  CLKBUF_X1 U12855 ( .A(n10192), .Z(n10001) );
  OAI21_X1 U12856 ( .B1(n12909), .B2(n10011), .A(n10010), .ZN(n12977) );
  NAND2_X1 U12857 ( .A1(n12909), .A2(n10010), .ZN(n10009) );
  NOR2_X1 U12858 ( .A1(n15214), .A2(n10017), .ZN(n15616) );
  MUX2_X1 U12859 ( .A(n19366), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10039) );
  AND2_X4 U12860 ( .A1(n10052), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10584) );
  NAND3_X1 U12861 ( .A1(n10045), .A2(n11455), .A3(n13360), .ZN(n13361) );
  NAND2_X1 U12862 ( .A1(n10661), .A2(n10660), .ZN(n10047) );
  AND2_X1 U12863 ( .A1(n10052), .A2(n11768), .ZN(n11718) );
  NAND2_X2 U12864 ( .A1(n10787), .A2(n10053), .ZN(n11469) );
  NAND3_X1 U12865 ( .A1(n10784), .A2(n10786), .A3(n9775), .ZN(n10055) );
  NAND2_X1 U12866 ( .A1(n10066), .A2(n10840), .ZN(n14294) );
  NAND2_X1 U12867 ( .A1(n14036), .A2(n14037), .ZN(n10066) );
  INV_X1 U12868 ( .A(n10068), .ZN(n10067) );
  OAI21_X1 U12869 ( .B1(n14037), .B2(n10069), .A(n14292), .ZN(n10068) );
  NAND2_X1 U12870 ( .A1(n10840), .A2(n9826), .ZN(n10069) );
  NAND3_X1 U12871 ( .A1(n11010), .A2(n11026), .A3(n10485), .ZN(n10070) );
  NAND3_X1 U12872 ( .A1(n10482), .A2(n10480), .A3(n10481), .ZN(n11010) );
  NAND2_X2 U12873 ( .A1(n10079), .A2(n10551), .ZN(n19991) );
  NAND2_X1 U12874 ( .A1(n18482), .A2(n12147), .ZN(n12149) );
  INV_X1 U12875 ( .A(n12252), .ZN(n18051) );
  NAND3_X1 U12876 ( .A1(n12073), .A2(n12075), .A3(n12074), .ZN(n12252) );
  NAND2_X1 U12877 ( .A1(n18440), .A2(n10089), .ZN(n12152) );
  AND2_X4 U12878 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10578) );
  NAND2_X1 U12879 ( .A1(n10247), .A2(n10248), .ZN(n10093) );
  INV_X1 U12880 ( .A(n9758), .ZN(n10096) );
  NAND3_X1 U12881 ( .A1(n10247), .A2(n10248), .A3(n19828), .ZN(n10092) );
  OAI211_X1 U12882 ( .C1(n10094), .C2(n19845), .A(n10097), .B(n10092), .ZN(
        P2_U2983) );
  AND2_X1 U12883 ( .A1(n10953), .A2(n10098), .ZN(n11524) );
  NAND2_X1 U12884 ( .A1(n10953), .A2(n10954), .ZN(n10964) );
  NAND2_X1 U12885 ( .A1(n10953), .A2(n10100), .ZN(n11523) );
  NAND2_X1 U12886 ( .A1(n10868), .A2(n10107), .ZN(n10898) );
  NAND2_X1 U12887 ( .A1(n10925), .A2(n10924), .ZN(n10930) );
  NAND3_X1 U12888 ( .A1(n10118), .A2(n10117), .A3(n10881), .ZN(n10116) );
  INV_X2 U12889 ( .A(n10387), .ZN(n11765) );
  NOR2_X1 U12890 ( .A1(n16033), .A2(n16032), .ZN(n10128) );
  INV_X1 U12891 ( .A(n11533), .ZN(n12387) );
  NAND2_X1 U12892 ( .A1(n11490), .A2(n9739), .ZN(n11985) );
  INV_X1 U12893 ( .A(n10152), .ZN(n11980) );
  MUX2_X1 U12894 ( .A(n15219), .B(n15129), .S(n15298), .Z(n10165) );
  NAND2_X1 U12895 ( .A1(n18255), .A2(n9811), .ZN(n18191) );
  INV_X1 U12896 ( .A(n10179), .ZN(n18185) );
  NAND2_X1 U12897 ( .A1(n10180), .A2(n10181), .ZN(n17284) );
  INV_X1 U12899 ( .A(n10184), .ZN(n17300) );
  OR2_X1 U12900 ( .A1(n17357), .A2(n10186), .ZN(n10188) );
  OAI21_X1 U12901 ( .B1(n12856), .B2(n10192), .A(n13587), .ZN(n12861) );
  INV_X1 U12902 ( .A(n14237), .ZN(n14222) );
  NAND2_X2 U12903 ( .A1(n14237), .A2(n9733), .ZN(n14355) );
  AND2_X2 U12904 ( .A1(n10194), .A2(n10193), .ZN(n14237) );
  INV_X1 U12905 ( .A(n14110), .ZN(n10193) );
  INV_X1 U12906 ( .A(n14098), .ZN(n10194) );
  NOR2_X2 U12907 ( .A1(n12777), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12440) );
  OAI211_X1 U12908 ( .C1(n14594), .C2(n10199), .A(n14624), .B(n10197), .ZN(
        n14625) );
  NAND2_X1 U12909 ( .A1(n13086), .A2(n10200), .ZN(n10204) );
  NAND2_X1 U12910 ( .A1(n13718), .A2(n12791), .ZN(n10203) );
  OAI22_X2 U12911 ( .A1(n13515), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13197), 
        .B2(n13186), .ZN(n13191) );
  NAND2_X2 U12912 ( .A1(n10204), .A2(n13173), .ZN(n13515) );
  INV_X1 U12913 ( .A(n13174), .ZN(n10205) );
  AND2_X2 U12914 ( .A1(n14835), .A2(n9809), .ZN(n15413) );
  NAND2_X1 U12915 ( .A1(n14641), .A2(n10210), .ZN(n15514) );
  NAND2_X1 U12916 ( .A1(n14641), .A2(n14640), .ZN(n14767) );
  NAND2_X1 U12917 ( .A1(n15338), .A2(n10216), .ZN(n15299) );
  AND2_X1 U12918 ( .A1(n15338), .A2(n9804), .ZN(n15310) );
  NAND2_X1 U12919 ( .A1(n15338), .A2(n15011), .ZN(n15324) );
  INV_X1 U12920 ( .A(n12989), .ZN(n10225) );
  NAND2_X1 U12921 ( .A1(n10225), .A2(n9729), .ZN(n13679) );
  INV_X1 U12922 ( .A(n10235), .ZN(n16103) );
  INV_X1 U12923 ( .A(n16117), .ZN(n10236) );
  NAND2_X1 U12924 ( .A1(n14321), .A2(n9830), .ZN(n15997) );
  NAND2_X1 U12925 ( .A1(n15939), .A2(n10240), .ZN(n11401) );
  NAND2_X1 U12926 ( .A1(n15939), .A2(n15938), .ZN(n15937) );
  NAND3_X1 U12927 ( .A1(n10538), .A2(n10246), .A3(n10535), .ZN(n10503) );
  NAND4_X1 U12928 ( .A1(n10538), .A2(n10539), .A3(n10246), .A4(n10537), .ZN(
        n10540) );
  NAND2_X2 U12929 ( .A1(n10515), .A2(n10514), .ZN(n11577) );
  NAND2_X1 U12930 ( .A1(n10251), .A2(n16216), .ZN(n16209) );
  NAND3_X1 U12931 ( .A1(n10253), .A2(n10254), .A3(n10252), .ZN(n10251) );
  NAND2_X1 U12932 ( .A1(n10923), .A2(n9782), .ZN(n10254) );
  NAND2_X1 U12933 ( .A1(n10254), .A2(n10253), .ZN(n16218) );
  AOI21_X2 U12934 ( .B1(n16209), .B2(n16208), .A(n10934), .ZN(n16198) );
  NAND4_X1 U12935 ( .A1(n10394), .A2(n10392), .A3(n10393), .A4(n10395), .ZN(
        n10460) );
  NAND4_X1 U12936 ( .A1(n10398), .A2(n10399), .A3(n10396), .A4(n10397), .ZN(
        n10457) );
  NAND4_X1 U12937 ( .A1(n10616), .A2(n10614), .A3(n10617), .A4(n10615), .ZN(
        n10661) );
  NAND3_X1 U12938 ( .A1(n10260), .A2(n10259), .A3(n10261), .ZN(n15255) );
  NAND2_X1 U12939 ( .A1(n15216), .A2(n15217), .ZN(n10263) );
  OR2_X1 U12940 ( .A1(n15216), .A2(n10265), .ZN(n10264) );
  NOR2_X1 U12941 ( .A1(n10267), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10265) );
  OR2_X1 U12942 ( .A1(n15216), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10266) );
  INV_X1 U12943 ( .A(n15627), .ZN(n10268) );
  NAND2_X1 U12944 ( .A1(n16767), .A2(n10270), .ZN(n10269) );
  NAND2_X1 U12945 ( .A1(n10269), .A2(n10271), .ZN(n14525) );
  NAND2_X1 U12946 ( .A1(n12599), .A2(n12598), .ZN(n12778) );
  MUX2_X1 U12947 ( .A(n20698), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12499) );
  NAND2_X1 U12948 ( .A1(n13086), .A2(n13984), .ZN(n13840) );
  NAND2_X1 U12949 ( .A1(n13718), .A2(n13085), .ZN(n13984) );
  OAI211_X1 U12950 ( .C1(n13718), .C2(n10278), .A(n10333), .B(n10276), .ZN(
        n13170) );
  NAND2_X1 U12951 ( .A1(n13718), .A2(n10277), .ZN(n10276) );
  AND2_X4 U12952 ( .A1(n10586), .A2(n10346), .ZN(n11766) );
  AND2_X2 U12953 ( .A1(n10474), .A2(n19905), .ZN(n10482) );
  NAND3_X1 U12954 ( .A1(n10390), .A2(n10323), .A3(n10331), .ZN(n10281) );
  NAND2_X1 U12955 ( .A1(n10459), .A2(n13387), .ZN(n10282) );
  NAND2_X1 U12956 ( .A1(n10382), .A2(n10383), .ZN(n10283) );
  NAND2_X1 U12957 ( .A1(n11595), .A2(n11596), .ZN(n11600) );
  CLKBUF_X1 U12958 ( .A(n11595), .Z(n10284) );
  INV_X1 U12959 ( .A(n11794), .ZN(n16061) );
  INV_X1 U12960 ( .A(n11815), .ZN(n10293) );
  NOR2_X2 U12961 ( .A1(n13294), .A2(n9736), .ZN(n13465) );
  INV_X1 U12962 ( .A(n10301), .ZN(n10390) );
  INV_X2 U12963 ( .A(n16224), .ZN(n10307) );
  NOR2_X2 U12964 ( .A1(n16172), .A2(n10309), .ZN(n11528) );
  INV_X1 U12965 ( .A(n10314), .ZN(n16266) );
  INV_X1 U12966 ( .A(n11515), .ZN(n11516) );
  NAND2_X1 U12967 ( .A1(n13142), .A2(n13143), .ZN(n13172) );
  OAI21_X1 U12968 ( .B1(n16170), .B2(n19859), .A(n11514), .ZN(n11515) );
  AOI21_X1 U12969 ( .B1(n13215), .B2(n11601), .A(n9807), .ZN(n11602) );
  NAND2_X1 U12970 ( .A1(n11600), .A2(n11599), .ZN(n13215) );
  NAND2_X1 U12971 ( .A1(n10555), .A2(n10551), .ZN(n20100) );
  OR2_X2 U12972 ( .A1(n10561), .A2(n10564), .ZN(n10760) );
  OR2_X2 U12973 ( .A1(n10557), .A2(n10556), .ZN(n20136) );
  OAI22_X1 U12974 ( .A1(n11223), .A2(n10773), .B1(n10778), .B2(n11219), .ZN(
        n10606) );
  AOI21_X1 U12975 ( .B1(n10401), .B2(n10474), .A(n10400), .ZN(n10403) );
  NAND2_X1 U12976 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10348) );
  OR2_X2 U12977 ( .A1(n11595), .A2(n10541), .ZN(n10561) );
  MUX2_X2 U12978 ( .A(n10362), .B(n10361), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10479) );
  INV_X1 U12979 ( .A(n12105), .ZN(n12221) );
  AND3_X1 U12980 ( .A1(n11861), .A2(n11836), .A3(n11835), .ZN(n10315) );
  OR4_X1 U12981 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(
        n10316) );
  AND3_X1 U12982 ( .A1(n11349), .A2(n11348), .A3(n11347), .ZN(n13661) );
  AND2_X1 U12983 ( .A1(n12033), .A2(n19679), .ZN(n10317) );
  INV_X1 U12984 ( .A(n19859), .ZN(n11551) );
  NAND2_X1 U12985 ( .A1(n14101), .A2(n14100), .ZN(n10318) );
  NOR2_X1 U12986 ( .A1(n16012), .A2(n16074), .ZN(n10320) );
  AND2_X1 U12987 ( .A1(n16180), .A2(n16184), .ZN(n10321) );
  OR2_X1 U12988 ( .A1(n17426), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10322) );
  AND2_X1 U12989 ( .A1(n10386), .A2(n10385), .ZN(n10323) );
  AND3_X1 U12990 ( .A1(n18699), .A2(n18749), .A3(n18721), .ZN(n10324) );
  AND2_X1 U12991 ( .A1(n12362), .A2(n10322), .ZN(n10325) );
  AND3_X1 U12992 ( .A1(n17504), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n17473), .ZN(n10326) );
  OR2_X1 U12993 ( .A1(n16469), .A2(n16467), .ZN(n10327) );
  NAND2_X1 U12994 ( .A1(n14887), .A2(n14886), .ZN(n10329) );
  INV_X2 U12995 ( .A(n18085), .ZN(n18118) );
  AND2_X1 U12996 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10330) );
  AND2_X1 U12997 ( .A1(n10389), .A2(n10388), .ZN(n10331) );
  INV_X1 U12998 ( .A(n10566), .ZN(n10551) );
  AND2_X1 U12999 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10332) );
  NAND2_X1 U13000 ( .A1(n13185), .A2(n13195), .ZN(n10333) );
  NAND2_X1 U13001 ( .A1(n16049), .A2(n16048), .ZN(n15930) );
  BUF_X4 U13002 ( .A(n12128), .Z(n17826) );
  XNOR2_X1 U13003 ( .A(n13164), .B(n13163), .ZN(n13162) );
  AND3_X1 U13004 ( .A1(n16240), .A2(n16249), .A3(n10906), .ZN(n10334) );
  INV_X1 U13005 ( .A(n15427), .ZN(n15442) );
  AND4_X1 U13006 ( .A1(n10647), .A2(n10646), .A3(n10645), .A4(n10644), .ZN(
        n10335) );
  AND4_X1 U13007 ( .A1(n11206), .A2(n11205), .A3(n11204), .A4(n11203), .ZN(
        n10336) );
  AND3_X1 U13008 ( .A1(n11256), .A2(n11255), .A3(n11254), .ZN(n13310) );
  AND3_X1 U13009 ( .A1(n10655), .A2(n10654), .A3(n10653), .ZN(n10337) );
  AND4_X1 U13010 ( .A1(n12090), .A2(n12089), .A3(n12088), .A4(n12087), .ZN(
        n10338) );
  NOR2_X1 U13011 ( .A1(n18555), .A2(n18526), .ZN(n18296) );
  AND3_X1 U13012 ( .A1(n20737), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10340) );
  AND3_X1 U13013 ( .A1(n10673), .A2(n10672), .A3(n10671), .ZN(n10341) );
  OAI21_X1 U13014 ( .B1(n11457), .B2(n10880), .A(n14458), .ZN(n10793) );
  AND2_X1 U13015 ( .A1(n12159), .A2(n12158), .ZN(n10342) );
  NOR2_X1 U13016 ( .A1(n12383), .A2(n12382), .ZN(n10343) );
  OR2_X1 U13017 ( .A1(n19563), .A2(n14265), .ZN(n17039) );
  INV_X1 U13018 ( .A(n17039), .ZN(n11531) );
  INV_X1 U13019 ( .A(n19845), .ZN(n19828) );
  BUF_X1 U13020 ( .A(n10534), .Z(n10543) );
  XNOR2_X1 U13021 ( .A(n11577), .B(n10533), .ZN(n10545) );
  NAND2_X1 U13022 ( .A1(n11595), .A2(n19869), .ZN(n10557) );
  AND4_X1 U13023 ( .A1(n12572), .A2(n12571), .A3(n12570), .A4(n12569), .ZN(
        n10344) );
  INV_X1 U13024 ( .A(n13958), .ZN(n13616) );
  OAI22_X1 U13025 ( .A1(n11662), .A2(n20205), .B1(n20257), .B2(n11851), .ZN(
        n10554) );
  INV_X1 U13026 ( .A(n11028), .ZN(n10401) );
  OR2_X1 U13027 ( .A1(n13970), .A2(n13969), .ZN(n14416) );
  AND3_X1 U13028 ( .A1(n13137), .A2(n13136), .A3(n13135), .ZN(n13168) );
  AND2_X1 U13029 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10355) );
  AND4_X1 U13030 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10383) );
  AND2_X1 U13031 ( .A1(n12434), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12432) );
  NAND2_X1 U13032 ( .A1(n12553), .A2(n13079), .ZN(n12568) );
  INV_X1 U13033 ( .A(n16196), .ZN(n10936) );
  OAI22_X1 U13034 ( .A1(n11841), .A2(n10724), .B1(n11898), .B2(n11680), .ZN(
        n10391) );
  INV_X1 U13035 ( .A(n14888), .ZN(n13827) );
  INV_X1 U13036 ( .A(n14829), .ZN(n13826) );
  OR2_X1 U13037 ( .A1(n12891), .A2(n12890), .ZN(n13194) );
  AND4_X1 U13038 ( .A1(n12551), .A2(n12550), .A3(n12549), .A4(n12548), .ZN(
        n12552) );
  OAI21_X1 U13039 ( .B1(n16198), .B2(n16195), .A(n10936), .ZN(n10937) );
  AND4_X1 U13040 ( .A1(n10341), .A2(n10676), .A3(n10675), .A4(n10674), .ZN(
        n10677) );
  AND4_X1 U13041 ( .A1(n10497), .A2(n12967), .A3(n10993), .A4(n19905), .ZN(
        n10498) );
  OR2_X2 U13042 ( .A1(n10565), .A2(n10562), .ZN(n10759) );
  INV_X1 U13043 ( .A(n10562), .ZN(n10563) );
  AND2_X1 U13044 ( .A1(n20779), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12504) );
  NOR2_X1 U13045 ( .A1(n15012), .A2(n15652), .ZN(n15029) );
  AND2_X1 U13046 ( .A1(n13827), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15003) );
  AND2_X1 U13047 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n13826), .ZN(
        n14836) );
  INV_X1 U13048 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13257) );
  OR2_X1 U13049 ( .A1(n13514), .A2(n13513), .ZN(n13534) );
  INV_X1 U13050 ( .A(n13138), .ZN(n12908) );
  INV_X1 U13051 ( .A(n10956), .ZN(n10953) );
  OAI21_X1 U13052 ( .B1(n10683), .B2(n11966), .A(n10682), .ZN(n10705) );
  INV_X1 U13053 ( .A(n13310), .ZN(n11605) );
  OR2_X1 U13054 ( .A1(n11834), .A2(n11837), .ZN(n11861) );
  AND4_X1 U13055 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10757) );
  AND3_X1 U13056 ( .A1(n11093), .A2(n11092), .A3(n11091), .ZN(n16010) );
  INV_X1 U13057 ( .A(n12394), .ZN(n11519) );
  NAND2_X1 U13058 ( .A1(n9801), .A2(n10920), .ZN(n10921) );
  NAND2_X1 U13059 ( .A1(n10412), .A2(n10411), .ZN(n10422) );
  NAND2_X1 U13060 ( .A1(n9747), .A2(n10563), .ZN(n10772) );
  NOR2_X1 U13061 ( .A1(n18917), .A2(n18922), .ZN(n12285) );
  INV_X1 U13062 ( .A(n12091), .ZN(n17745) );
  AOI21_X1 U13063 ( .B1(n12339), .B2(n18730), .A(n16592), .ZN(n12340) );
  AND2_X1 U13064 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12266), .ZN(
        n12267) );
  AND2_X1 U13065 ( .A1(n12538), .A2(n12537), .ZN(n12539) );
  AND2_X1 U13066 ( .A1(n14114), .A2(n14113), .ZN(n16853) );
  AND2_X1 U13067 ( .A1(n15340), .A2(n15339), .ZN(n15011) );
  NAND2_X1 U13068 ( .A1(n15083), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12456) );
  NOR2_X1 U13069 ( .A1(n15070), .A2(n15187), .ZN(n13829) );
  OR2_X1 U13070 ( .A1(n14973), .A2(n15667), .ZN(n14902) );
  NAND2_X1 U13071 ( .A1(n15003), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15006) );
  NAND2_X1 U13072 ( .A1(n14768), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14783) );
  NOR2_X1 U13073 ( .A1(n13577), .A2(n14046), .ZN(n13958) );
  INV_X1 U13074 ( .A(n15744), .ZN(n15201) );
  INV_X1 U13075 ( .A(n13633), .ZN(n13631) );
  NAND2_X1 U13076 ( .A1(n12767), .A2(n13587), .ZN(n12768) );
  AND3_X1 U13077 ( .A1(n11103), .A2(n11102), .A3(n11101), .ZN(n15978) );
  INV_X1 U13078 ( .A(n13487), .ZN(n11056) );
  NAND2_X1 U13079 ( .A1(n11839), .A2(n10315), .ZN(n11840) );
  INV_X1 U13080 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11543) );
  OR2_X1 U13081 ( .A1(n16262), .A2(n16272), .ZN(n16237) );
  INV_X1 U13082 ( .A(n11532), .ZN(n11135) );
  AOI21_X1 U13083 ( .B1(n19699), .B2(n11596), .A(n11571), .ZN(n12961) );
  AND2_X1 U13084 ( .A1(n18917), .A2(n17926), .ZN(n12280) );
  INV_X1 U13085 ( .A(n12355), .ZN(n18255) );
  NAND2_X1 U13086 ( .A1(n12144), .A2(n12145), .ZN(n12122) );
  NOR2_X1 U13087 ( .A1(n18929), .A2(n16681), .ZN(n12290) );
  AND2_X1 U13088 ( .A1(n15281), .A2(n12614), .ZN(n15282) );
  INV_X1 U13089 ( .A(n20593), .ZN(n20581) );
  OR2_X1 U13090 ( .A1(n13846), .A2(n13845), .ZN(n20578) );
  AND2_X1 U13091 ( .A1(n14766), .A2(n14765), .ZN(n15466) );
  AND3_X1 U13092 ( .A1(n14354), .A2(n14353), .A3(n14352), .ZN(n14451) );
  INV_X1 U13093 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15217) );
  OR3_X1 U13094 ( .A1(n15852), .A2(n15826), .A3(n15239), .ZN(n15821) );
  OR2_X1 U13095 ( .A1(n16783), .A2(n16775), .ZN(n15852) );
  XNOR2_X1 U13096 ( .A(n13451), .B(n13211), .ZN(n13449) );
  AND2_X1 U13097 ( .A1(n13119), .A2(n13118), .ZN(n15228) );
  NAND2_X1 U13098 ( .A1(n12803), .A2(n12802), .ZN(n13544) );
  AND3_X1 U13099 ( .A1(n12867), .A2(n13102), .A3(n12866), .ZN(n14744) );
  INV_X1 U13100 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20698) );
  OR2_X1 U13101 ( .A1(n13539), .A2(n13253), .ZN(n13722) );
  NAND2_X1 U13102 ( .A1(n13865), .A2(n13906), .ZN(n20859) );
  AND2_X1 U13103 ( .A1(n13540), .A2(n13721), .ZN(n13761) );
  OR2_X1 U13104 ( .A1(n13540), .A2(n15927), .ZN(n13989) );
  AOI21_X1 U13105 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20779), .A(n14128), 
        .ZN(n20744) );
  INV_X1 U13106 ( .A(n13906), .ZN(n13988) );
  INV_X1 U13107 ( .A(n13764), .ZN(n14546) );
  INV_X1 U13108 ( .A(n11536), .ZN(n11134) );
  AND3_X1 U13109 ( .A1(n11116), .A2(n11115), .A3(n11114), .ZN(n15950) );
  INV_X1 U13110 ( .A(n11215), .ZN(n14442) );
  AND2_X1 U13111 ( .A1(n11148), .A2(n11147), .ZN(n13491) );
  AOI211_X1 U13112 ( .C1(n19718), .C2(n19854), .A(n11559), .B(n11558), .ZN(
        n11563) );
  NAND2_X1 U13113 ( .A1(n10711), .A2(n13355), .ZN(n13349) );
  INV_X1 U13114 ( .A(n19863), .ZN(n16436) );
  INV_X1 U13115 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20101) );
  INV_X1 U13116 ( .A(n20478), .ZN(n14255) );
  OR2_X1 U13117 ( .A1(n20466), .A2(n20478), .ZN(n20260) );
  INV_X1 U13119 ( .A(n17600), .ZN(n17609) );
  NAND2_X1 U13120 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17743), .ZN(n17739) );
  NOR2_X1 U13121 ( .A1(n12085), .A2(n12084), .ZN(n12249) );
  INV_X1 U13122 ( .A(n18234), .ZN(n18235) );
  INV_X1 U13123 ( .A(n18401), .ZN(n18393) );
  INV_X1 U13124 ( .A(n18415), .ZN(n17473) );
  NOR2_X1 U13125 ( .A1(n18302), .A2(n10342), .ZN(n18248) );
  NOR2_X1 U13126 ( .A1(n18344), .A2(n18662), .ZN(n18281) );
  NOR2_X1 U13127 ( .A1(n18367), .A2(n18699), .ZN(n18705) );
  AOI21_X1 U13128 ( .B1(n19336), .B2(n19343), .A(n19335), .ZN(n19345) );
  NOR2_X1 U13129 ( .A1(n18811), .A2(n18508), .ZN(n18507) );
  XNOR2_X1 U13130 ( .A(n18066), .B(n18056), .ZN(n12127) );
  INV_X2 U13131 ( .A(n12221), .ZN(n17763) );
  NOR2_X1 U13132 ( .A1(n12237), .A2(n12236), .ZN(n18909) );
  OR3_X1 U13133 ( .A1(n21026), .A2(n13116), .A3(n13825), .ZN(n15180) );
  AND2_X1 U13134 ( .A1(n15180), .A2(n13841), .ZN(n20604) );
  AND2_X1 U13135 ( .A1(n21026), .A2(n13837), .ZN(n20595) );
  OR2_X1 U13136 ( .A1(n13050), .A2(n20508), .ZN(n13053) );
  INV_X1 U13137 ( .A(n15606), .ZN(n15610) );
  INV_X1 U13138 ( .A(n12926), .ZN(n13030) );
  INV_X1 U13139 ( .A(n13001), .ZN(n13042) );
  NAND2_X1 U13140 ( .A1(n14595), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14626) );
  INV_X1 U13141 ( .A(n16769), .ZN(n16742) );
  NOR2_X1 U13142 ( .A1(n15222), .A2(n15846), .ZN(n15234) );
  AND2_X1 U13143 ( .A1(n13117), .A2(n13108), .ZN(n16857) );
  AND2_X1 U13144 ( .A1(n13117), .A2(n13104), .ZN(n20656) );
  NAND2_X1 U13145 ( .A1(n16614), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21010) );
  NOR2_X2 U13146 ( .A1(n20695), .A2(n13989), .ZN(n20689) );
  NOR2_X1 U13147 ( .A1(n13540), .A2(n13721), .ZN(n13906) );
  OAI21_X1 U13148 ( .B1(n20705), .B2(n20704), .A(n20703), .ZN(n20729) );
  NOR2_X2 U13149 ( .A1(n20695), .A2(n20694), .ZN(n20770) );
  OAI21_X1 U13150 ( .B1(n14189), .B2(n14192), .A(n20876), .ZN(n14214) );
  NOR2_X1 U13151 ( .A1(n13722), .A2(n13989), .ZN(n14218) );
  NOR2_X2 U13152 ( .A1(n13722), .A2(n13988), .ZN(n20801) );
  NOR2_X2 U13153 ( .A1(n13722), .A2(n20694), .ZN(n20802) );
  NOR2_X1 U13154 ( .A1(n13722), .A2(n14546), .ZN(n14166) );
  AND2_X1 U13155 ( .A1(n13865), .A2(n13864), .ZN(n14126) );
  OAI21_X1 U13156 ( .B1(n20823), .B2(n20822), .A(n20821), .ZN(n20862) );
  AND2_X1 U13157 ( .A1(n13865), .A2(n13761), .ZN(n20861) );
  AND2_X1 U13158 ( .A1(n13865), .A2(n13764), .ZN(n20926) );
  OAI21_X1 U13159 ( .B1(n20881), .B2(n20880), .A(n20879), .ZN(n20928) );
  NOR2_X2 U13160 ( .A1(n14547), .A2(n14546), .ZN(n20688) );
  INV_X1 U13161 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21133) );
  AND2_X1 U13162 ( .A1(n12032), .A2(n12031), .ZN(n19679) );
  INV_X1 U13163 ( .A(n19690), .ZN(n19672) );
  XNOR2_X1 U13164 ( .A(n13216), .B(n13217), .ZN(n13218) );
  INV_X1 U13165 ( .A(n16533), .ZN(n12969) );
  AND2_X1 U13166 ( .A1(n12959), .A2(n13225), .ZN(n19719) );
  INV_X1 U13167 ( .A(n19754), .ZN(n19773) );
  INV_X1 U13168 ( .A(n12694), .ZN(n13225) );
  INV_X1 U13169 ( .A(n17046), .ZN(n19837) );
  AND2_X1 U13170 ( .A1(n11482), .A2(n11426), .ZN(n19863) );
  NAND2_X1 U13171 ( .A1(n13219), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16552) );
  NOR2_X2 U13172 ( .A1(n20132), .A2(n20041), .ZN(n19937) );
  INV_X1 U13173 ( .A(n19989), .ZN(n19981) );
  INV_X1 U13174 ( .A(n19998), .ZN(n20016) );
  NOR2_X1 U13175 ( .A1(n20041), .A2(n20260), .ZN(n20022) );
  OR3_X1 U13176 ( .A1(n20046), .A2(n20074), .A3(n20045), .ZN(n20063) );
  INV_X1 U13177 ( .A(n20161), .ZN(n20153) );
  OAI21_X1 U13178 ( .B1(n20172), .B2(n20195), .A(n20320), .ZN(n20197) );
  NOR2_X2 U13179 ( .A1(n20166), .A2(n20209), .ZN(n20229) );
  INV_X1 U13180 ( .A(n20233), .ZN(n20250) );
  AND2_X1 U13181 ( .A1(n20261), .A2(n20258), .ZN(n20279) );
  INV_X1 U13182 ( .A(n20284), .ZN(n20305) );
  AND2_X1 U13183 ( .A1(n13429), .A2(n19904), .ZN(n20314) );
  INV_X1 U13184 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20312) );
  OR2_X1 U13185 ( .A1(n17290), .A2(n17289), .ZN(n17291) );
  INV_X1 U13186 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17906) );
  NOR2_X1 U13187 ( .A1(n18131), .A2(n17995), .ZN(n17990) );
  INV_X1 U13188 ( .A(n18063), .ZN(n18060) );
  NOR2_X1 U13189 ( .A1(n18123), .A2(n18072), .ZN(n18104) );
  NAND2_X1 U13190 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18236) );
  INV_X1 U13191 ( .A(n18356), .ZN(n18340) );
  INV_X1 U13192 ( .A(n18705), .ZN(n18623) );
  NOR2_X2 U13193 ( .A1(n19503), .A2(n18549), .ZN(n18401) );
  NOR2_X1 U13194 ( .A1(n17260), .A2(n19539), .ZN(n18502) );
  INV_X1 U13195 ( .A(n18792), .ZN(n18725) );
  NAND2_X1 U13196 ( .A1(n19353), .A2(n19360), .ZN(n18763) );
  INV_X1 U13197 ( .A(n18740), .ZN(n18788) );
  NOR2_X1 U13198 ( .A1(n18828), .A2(n18854), .ZN(n18873) );
  INV_X1 U13199 ( .A(U212), .ZN(n17207) );
  NAND2_X1 U13200 ( .A1(n16614), .A2(n12592), .ZN(n12831) );
  OR2_X1 U13201 ( .A1(n15412), .A2(n15178), .ZN(n15384) );
  NAND2_X1 U13202 ( .A1(n15180), .A2(n13830), .ZN(n15476) );
  OR2_X1 U13203 ( .A1(n13846), .A2(n13834), .ZN(n20592) );
  NAND2_X1 U13204 ( .A1(n12922), .A2(n12921), .ZN(n15606) );
  INV_X1 U13205 ( .A(n20619), .ZN(n20649) );
  NOR2_X1 U13206 ( .A1(n12831), .A2(n12830), .ZN(n12931) );
  OR2_X1 U13207 ( .A1(n13015), .A2(n13587), .ZN(n13001) );
  INV_X1 U13208 ( .A(n16689), .ZN(n15743) );
  NAND2_X1 U13209 ( .A1(n16774), .A2(n13158), .ZN(n16769) );
  NAND2_X1 U13210 ( .A1(n20516), .A2(n12982), .ZN(n16774) );
  INV_X1 U13211 ( .A(n16857), .ZN(n20652) );
  AOI22_X1 U13212 ( .A1(n20666), .A2(n20671), .B1(n20665), .B2(n20811), .ZN(
        n20693) );
  NAND2_X1 U13213 ( .A1(n20734), .A2(n13906), .ZN(n20727) );
  AOI22_X1 U13214 ( .A1(n20697), .A2(n20704), .B1(n20811), .B2(n20777), .ZN(
        n20732) );
  AOI22_X1 U13215 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20742), .B1(n20741), 
        .B2(n20745), .ZN(n20774) );
  INV_X1 U13216 ( .A(n20769), .ZN(n14221) );
  INV_X1 U13217 ( .A(n14218), .ZN(n13603) );
  AOI22_X1 U13218 ( .A1(n20778), .A2(n20784), .B1(n20871), .B2(n20777), .ZN(
        n20806) );
  INV_X1 U13219 ( .A(n14166), .ZN(n13752) );
  INV_X1 U13220 ( .A(n14126), .ZN(n14170) );
  INV_X1 U13221 ( .A(n13863), .ZN(n13905) );
  AOI22_X1 U13222 ( .A1(n20813), .A2(n20822), .B1(n20812), .B2(n20811), .ZN(
        n20865) );
  INV_X1 U13223 ( .A(n20861), .ZN(n13806) );
  INV_X1 U13224 ( .A(n14002), .ZN(n20903) );
  AOI22_X1 U13225 ( .A1(n20872), .A2(n20880), .B1(n20871), .B2(n20870), .ZN(
        n20932) );
  INV_X1 U13226 ( .A(n14043), .ZN(n14584) );
  NAND2_X1 U13227 ( .A1(n20312), .A2(n20101), .ZN(n20133) );
  AOI22_X1 U13228 ( .A1(n16890), .A2(n19636), .B1(n19671), .B2(n19718), .ZN(
        n16891) );
  INV_X1 U13229 ( .A(n19679), .ZN(n19692) );
  INV_X1 U13230 ( .A(n19671), .ZN(n19703) );
  OR2_X1 U13231 ( .A1(n13434), .A2(n12709), .ZN(n19688) );
  AND2_X1 U13232 ( .A1(n11975), .A2(n11974), .ZN(n11976) );
  NAND2_X1 U13233 ( .A1(n11162), .A2(n19744), .ZN(n19754) );
  AND2_X2 U13234 ( .A1(n11955), .A2(n13124), .ZN(n19744) );
  NOR2_X1 U13235 ( .A1(n19773), .A2(n19772), .ZN(n19758) );
  INV_X1 U13236 ( .A(n19746), .ZN(n19779) );
  NAND2_X1 U13237 ( .A1(n12712), .A2(n12711), .ZN(n19816) );
  INV_X1 U13238 ( .A(n19822), .ZN(n12707) );
  OR2_X1 U13239 ( .A1(n19563), .A2(n9699), .ZN(n19845) );
  INV_X1 U13240 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17022) );
  NAND2_X1 U13241 ( .A1(n19563), .A2(n11489), .ZN(n17046) );
  INV_X1 U13242 ( .A(n11443), .ZN(n11484) );
  NAND2_X1 U13243 ( .A1(n11482), .A2(n20496), .ZN(n19859) );
  INV_X1 U13244 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21126) );
  NAND2_X1 U13245 ( .A1(n20097), .A2(n20067), .ZN(n19968) );
  OR2_X1 U13246 ( .A1(n20041), .A2(n20209), .ZN(n19989) );
  INV_X1 U13247 ( .A(n20011), .ZN(n20019) );
  INV_X1 U13248 ( .A(n20022), .ZN(n20038) );
  NAND2_X1 U13249 ( .A1(n20067), .A2(n13646), .ZN(n20066) );
  NAND2_X1 U13250 ( .A1(n20068), .A2(n20067), .ZN(n20129) );
  NAND2_X1 U13251 ( .A1(n20098), .A2(n20097), .ZN(n20161) );
  INV_X1 U13252 ( .A(n20339), .ZN(n20185) );
  INV_X1 U13253 ( .A(n20167), .ZN(n20200) );
  NAND2_X1 U13254 ( .A1(n14254), .A2(n20454), .ZN(n20233) );
  AOI21_X1 U13255 ( .B1(n13340), .B2(n13339), .A(n13338), .ZN(n20254) );
  NAND2_X1 U13256 ( .A1(n14254), .A2(n13646), .ZN(n20284) );
  NAND2_X1 U13257 ( .A1(n14254), .A2(n20068), .ZN(n20370) );
  NOR2_X1 U13258 ( .A1(n19323), .A2(n18123), .ZN(n19555) );
  OR2_X1 U13259 ( .A1(n19329), .A2(n19391), .ZN(n17260) );
  NAND2_X1 U13260 ( .A1(n12384), .A2(n10343), .ZN(n12385) );
  INV_X1 U13261 ( .A(n17617), .ZN(n17608) );
  NOR2_X1 U13262 ( .A1(n17633), .A2(n17632), .ZN(n17658) );
  NAND2_X1 U13263 ( .A1(n18102), .A2(n18121), .ZN(n18085) );
  INV_X1 U13264 ( .A(n18104), .ZN(n18121) );
  INV_X1 U13265 ( .A(n18173), .ZN(n18176) );
  NAND2_X1 U13266 ( .A1(n18036), .A2(n18502), .ZN(n18399) );
  NOR2_X1 U13267 ( .A1(n18296), .A2(n18401), .ZN(n18538) );
  OR2_X1 U13268 ( .A1(n18615), .A2(n18199), .ZN(n12351) );
  INV_X1 U13269 ( .A(n18854), .ZN(n18871) );
  INV_X1 U13270 ( .A(n18462), .ZN(n18793) );
  INV_X1 U13271 ( .A(n18873), .ZN(n18841) );
  INV_X1 U13272 ( .A(n18864), .ZN(n18878) );
  INV_X1 U13273 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19375) );
  INV_X1 U13274 ( .A(n18940), .ZN(n19281) );
  INV_X1 U13275 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19492) );
  INV_X1 U13276 ( .A(n17214), .ZN(n17209) );
  OR2_X1 U13277 ( .A1(n12386), .A2(n12385), .ZN(P3_U2642) );
  INV_X1 U13278 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10581) );
  INV_X1 U13279 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13280 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10585), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U13281 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10351) );
  AND2_X4 U13282 ( .A1(n10578), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10449) );
  AND2_X4 U13283 ( .A1(n10578), .A2(n10346), .ZN(n10592) );
  AOI22_X1 U13284 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10350) );
  AND2_X4 U13285 ( .A1(n10586), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11895) );
  NAND2_X1 U13286 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10347) );
  NAND4_X1 U13287 ( .A1(n10352), .A2(n10351), .A3(n10350), .A4(n10349), .ZN(
        n10362) );
  AOI22_X1 U13288 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10360) );
  NAND2_X1 U13289 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10354) );
  NOR2_X1 U13290 ( .A1(n10356), .A2(n10355), .ZN(n10358) );
  AOI22_X1 U13291 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10357) );
  NAND4_X1 U13292 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10361) );
  AOI22_X1 U13293 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13294 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10365) );
  INV_X2 U13295 ( .A(n10387), .ZN(n11912) );
  AOI22_X1 U13296 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10585), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13297 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10363) );
  NAND4_X1 U13298 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n10367) );
  NAND2_X1 U13299 ( .A1(n10367), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10374) );
  AOI22_X1 U13300 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13301 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13302 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10585), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13303 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10368) );
  NAND4_X1 U13304 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        n10372) );
  NAND2_X2 U13305 ( .A1(n10374), .A2(n10373), .ZN(n19896) );
  XNOR2_X1 U13306 ( .A(n9704), .B(n19896), .ZN(n11028) );
  INV_X1 U13307 ( .A(n11895), .ZN(n11841) );
  INV_X1 U13308 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10376) );
  INV_X1 U13309 ( .A(n10592), .ZN(n11898) );
  INV_X1 U13310 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10375) );
  OAI22_X1 U13311 ( .A1(n11841), .A2(n10376), .B1(n11898), .B2(n10375), .ZN(
        n10384) );
  NAND2_X1 U13312 ( .A1(n10591), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10380) );
  NAND2_X1 U13313 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10379) );
  INV_X1 U13314 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11682) );
  OR2_X1 U13315 ( .A1(n10387), .A2(n11682), .ZN(n10378) );
  NAND2_X1 U13316 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10377) );
  INV_X1 U13317 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11686) );
  INV_X1 U13318 ( .A(n10381), .ZN(n10382) );
  NAND2_X1 U13319 ( .A1(n10591), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10386) );
  NAND2_X1 U13320 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10385) );
  INV_X1 U13321 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11873) );
  INV_X1 U13322 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11679) );
  NAND2_X1 U13323 ( .A1(n10585), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10389) );
  INV_X1 U13324 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11286) );
  OR2_X1 U13325 ( .A1(n10387), .A2(n11286), .ZN(n10388) );
  INV_X1 U13326 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10724) );
  INV_X1 U13327 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U13328 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U13329 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10585), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U13330 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U13331 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U13332 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U13333 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13334 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10396) );
  INV_X1 U13335 ( .A(n11023), .ZN(n10402) );
  NAND2_X1 U13336 ( .A1(n10403), .A2(n10402), .ZN(n11414) );
  INV_X1 U13337 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10552) );
  OAI22_X1 U13338 ( .A1(n10573), .A2(n10552), .B1(n13393), .B2(n11661), .ZN(
        n10405) );
  OAI22_X1 U13339 ( .A1(n11841), .A2(n21045), .B1(n11898), .B2(n11662), .ZN(
        n10404) );
  NOR2_X1 U13340 ( .A1(n10405), .A2(n10404), .ZN(n10412) );
  NAND2_X1 U13341 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10409) );
  NAND2_X1 U13342 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10408) );
  NAND2_X1 U13343 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10407) );
  NAND2_X1 U13344 ( .A1(n10591), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10406) );
  NAND4_X1 U13345 ( .A1(n10409), .A2(n10408), .A3(n10407), .A4(n10406), .ZN(
        n10410) );
  OAI22_X1 U13346 ( .A1(n10573), .A2(n11842), .B1(n13393), .B2(n11668), .ZN(
        n10414) );
  INV_X1 U13347 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10558) );
  INV_X1 U13348 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10547) );
  OAI22_X1 U13349 ( .A1(n11841), .A2(n10558), .B1(n11898), .B2(n10547), .ZN(
        n10413) );
  NOR2_X1 U13350 ( .A1(n10414), .A2(n10413), .ZN(n10420) );
  NAND2_X1 U13351 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10418) );
  NAND2_X1 U13352 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10417) );
  NAND2_X1 U13353 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10416) );
  NAND2_X1 U13354 ( .A1(n10591), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10415) );
  NAND2_X2 U13355 ( .A1(n10422), .A2(n10421), .ZN(n10470) );
  AOI22_X1 U13356 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11895), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13357 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10585), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13358 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13359 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10424) );
  NAND4_X1 U13360 ( .A1(n10427), .A2(n10426), .A3(n10425), .A4(n10424), .ZN(
        n10433) );
  AOI22_X1 U13361 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13362 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10585), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U13363 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11895), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13364 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10428) );
  NAND4_X1 U13365 ( .A1(n10431), .A2(n10430), .A3(n10429), .A4(n10428), .ZN(
        n10432) );
  MUX2_X2 U13366 ( .A(n10433), .B(n10432), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10485) );
  NAND2_X1 U13367 ( .A1(n10491), .A2(n9771), .ZN(n11412) );
  AOI22_X1 U13368 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10585), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U13369 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13370 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U13371 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10434) );
  NAND4_X1 U13372 ( .A1(n10437), .A2(n10436), .A3(n10435), .A4(n10434), .ZN(
        n10443) );
  AOI22_X1 U13373 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10585), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U13374 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13375 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13376 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10438) );
  NAND4_X1 U13377 ( .A1(n10441), .A2(n10440), .A3(n10439), .A4(n10438), .ZN(
        n10442) );
  MUX2_X2 U13378 ( .A(n10443), .B(n10442), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19880) );
  NOR2_X1 U13379 ( .A1(n10479), .A2(n19896), .ZN(n10444) );
  NAND3_X2 U13380 ( .A1(n10482), .A2(n10480), .A3(n10444), .ZN(n13445) );
  AOI22_X1 U13381 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13382 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13383 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13384 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10445) );
  NAND4_X1 U13385 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10455) );
  AOI22_X1 U13386 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10585), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U13387 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13388 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11895), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13389 ( .A1(n10584), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10450) );
  NAND4_X1 U13390 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10454) );
  MUX2_X2 U13391 ( .A(n10455), .B(n10454), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13429) );
  NAND2_X1 U13392 ( .A1(n10694), .A2(n10470), .ZN(n10495) );
  INV_X1 U13393 ( .A(n10495), .ZN(n10465) );
  NAND2_X1 U13394 ( .A1(n9699), .A2(n11024), .ZN(n11951) );
  NAND2_X2 U13395 ( .A1(n11951), .A2(n10694), .ZN(n11947) );
  INV_X1 U13397 ( .A(n10456), .ZN(n10458) );
  NAND4_X1 U13398 ( .A1(n10458), .A2(n10457), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10463) );
  INV_X1 U13399 ( .A(n10459), .ZN(n10461) );
  NAND4_X1 U13400 ( .A1(n10461), .A2(n10460), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n13387), .ZN(n10462) );
  AOI21_X1 U13401 ( .B1(n10463), .B2(n10462), .A(n10479), .ZN(n10464) );
  AND2_X1 U13402 ( .A1(n11024), .A2(n19896), .ZN(n10467) );
  AND2_X1 U13403 ( .A1(n10470), .A2(n10479), .ZN(n10496) );
  AND2_X1 U13404 ( .A1(n19896), .A2(n19880), .ZN(n10471) );
  INV_X1 U13405 ( .A(n10477), .ZN(n10472) );
  NAND2_X1 U13406 ( .A1(n10522), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10473) );
  OAI21_X1 U13407 ( .B1(n9704), .B2(n11416), .A(n11149), .ZN(n10476) );
  AOI21_X1 U13408 ( .B1(n10474), .B2(n12967), .A(n19880), .ZN(n10475) );
  NAND3_X1 U13409 ( .A1(n19905), .A2(n10476), .A3(n10475), .ZN(n10478) );
  NAND3_X1 U13410 ( .A1(n10478), .A2(n10477), .A3(n11024), .ZN(n11413) );
  AND2_X1 U13411 ( .A1(n19896), .A2(n10479), .ZN(n10481) );
  NOR2_X2 U13412 ( .A1(n10484), .A2(n10483), .ZN(n11953) );
  AND2_X4 U13413 ( .A1(n11953), .A2(n10486), .ZN(n11536) );
  INV_X2 U13414 ( .A(n13445), .ZN(n11020) );
  INV_X1 U13415 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U13416 ( .A1(n11007), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19558) );
  INV_X1 U13417 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14513) );
  NAND2_X1 U13418 ( .A1(n14513), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U13419 ( .A1(n19558), .A2(n10490), .ZN(n10535) );
  NOR2_X1 U13420 ( .A1(n10492), .A2(n10483), .ZN(n10494) );
  INV_X4 U13421 ( .A(n10479), .ZN(n11966) );
  NAND2_X1 U13422 ( .A1(n10495), .A2(n11966), .ZN(n10499) );
  INV_X1 U13423 ( .A(n10496), .ZN(n10497) );
  NAND3_X1 U13424 ( .A1(n11947), .A2(n10499), .A3(n10498), .ZN(n13403) );
  NAND2_X1 U13425 ( .A1(n13384), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10536) );
  NOR2_X1 U13426 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12616) );
  NAND2_X1 U13427 ( .A1(n12616), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10500) );
  NAND2_X1 U13428 ( .A1(n10539), .A2(n10501), .ZN(n10502) );
  NAND2_X1 U13429 ( .A1(n10516), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10507) );
  NAND2_X1 U13430 ( .A1(n11020), .A2(n13429), .ZN(n10504) );
  NAND2_X1 U13431 ( .A1(n11403), .A2(n10505), .ZN(n11136) );
  AOI22_X1 U13432 ( .A1(n11136), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12616), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U13433 ( .A1(n10507), .A2(n10506), .ZN(n10511) );
  AOI22_X1 U13434 ( .A1(n11042), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10510) );
  NAND2_X1 U13435 ( .A1(n10522), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10509) );
  NAND2_X1 U13436 ( .A1(n11536), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10508) );
  XNOR2_X1 U13437 ( .A(n10511), .B(n10512), .ZN(n10534) );
  NAND2_X1 U13438 ( .A1(n10542), .A2(n10534), .ZN(n10515) );
  INV_X1 U13439 ( .A(n10512), .ZN(n10513) );
  NAND2_X1 U13440 ( .A1(n10516), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10518) );
  AOI21_X1 U13441 ( .B1(n17100), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10517) );
  INV_X1 U13442 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19857) );
  NAND2_X1 U13443 ( .A1(n11536), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10520) );
  NAND2_X1 U13444 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10519) );
  OAI211_X1 U13445 ( .C1(n11100), .C2(n19857), .A(n10520), .B(n10519), .ZN(
        n10521) );
  INV_X1 U13446 ( .A(n10521), .ZN(n10524) );
  NAND2_X1 U13447 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10523) );
  NAND2_X1 U13448 ( .A1(n10516), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10527) );
  NAND2_X1 U13449 ( .A1(n12616), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10526) );
  INV_X1 U13450 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13356) );
  NAND2_X1 U13451 ( .A1(n11536), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10529) );
  NAND2_X1 U13452 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10528) );
  OAI211_X1 U13453 ( .C1(n11100), .C2(n13356), .A(n10529), .B(n10528), .ZN(
        n10530) );
  INV_X1 U13454 ( .A(n10530), .ZN(n10532) );
  NAND2_X1 U13455 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10531) );
  AND2_X1 U13456 ( .A1(n10536), .A2(n10535), .ZN(n10537) );
  OR2_X1 U13457 ( .A1(n10543), .A2(n15264), .ZN(n10556) );
  OR2_X2 U13458 ( .A1(n10565), .A2(n10556), .ZN(n10764) );
  INV_X1 U13459 ( .A(n10545), .ZN(n10541) );
  INV_X1 U13460 ( .A(n15264), .ZN(n14520) );
  OR2_X2 U13461 ( .A1(n10561), .A2(n10566), .ZN(n10765) );
  OAI22_X1 U13462 ( .A1(n10581), .A2(n10764), .B1(n10765), .B2(n11842), .ZN(
        n10549) );
  INV_X1 U13463 ( .A(n10543), .ZN(n10544) );
  NAND2_X1 U13464 ( .A1(n9706), .A2(n15264), .ZN(n10564) );
  INV_X1 U13465 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11271) );
  NOR2_X1 U13466 ( .A1(n10549), .A2(n10548), .ZN(n10572) );
  INV_X1 U13467 ( .A(n10556), .ZN(n10550) );
  INV_X1 U13468 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11851) );
  INV_X1 U13469 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11267) );
  OR2_X2 U13470 ( .A1(n10561), .A2(n10556), .ZN(n10778) );
  OAI22_X1 U13471 ( .A1(n11267), .A2(n10778), .B1(n20100), .B2(n10552), .ZN(
        n10553) );
  NOR2_X1 U13472 ( .A1(n10554), .A2(n10553), .ZN(n10571) );
  INV_X1 U13473 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11274) );
  OAI22_X1 U13474 ( .A1(n11668), .A2(n10759), .B1(n20162), .B2(n11274), .ZN(
        n10560) );
  INV_X1 U13475 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11272) );
  OAI22_X1 U13476 ( .A1(n10558), .A2(n19991), .B1(n20136), .B2(n11272), .ZN(
        n10559) );
  NOR2_X1 U13477 ( .A1(n10560), .A2(n10559), .ZN(n10570) );
  INV_X1 U13478 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11664) );
  OAI22_X1 U13479 ( .A1(n11664), .A2(n10760), .B1(n10772), .B2(n11661), .ZN(
        n10568) );
  INV_X1 U13480 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11844) );
  NAND2_X1 U13481 ( .A1(n9747), .A2(n10551), .ZN(n10774) );
  OAI22_X1 U13482 ( .A1(n10773), .A2(n11844), .B1(n10774), .B2(n21045), .ZN(
        n10567) );
  NOR2_X1 U13483 ( .A1(n10568), .A2(n10567), .ZN(n10569) );
  OAI22_X1 U13484 ( .A1(n11272), .A2(n11699), .B1(n11697), .B2(n11851), .ZN(
        n10583) );
  NAND3_X1 U13485 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11006) );
  INV_X1 U13486 ( .A(n11006), .ZN(n10575) );
  NAND2_X1 U13487 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n11700), .ZN(
        n10576) );
  OAI21_X1 U13488 ( .B1(n11703), .B2(n11842), .A(n10576), .ZN(n10577) );
  AOI21_X1 U13489 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n10577), .ZN(n10580) );
  NAND2_X1 U13490 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10579) );
  OAI211_X1 U13491 ( .C1(n11726), .C2(n10581), .A(n10580), .B(n10579), .ZN(
        n10582) );
  NOR2_X1 U13492 ( .A1(n10583), .A2(n10582), .ZN(n10599) );
  BUF_X4 U13493 ( .A(n10584), .Z(n11936) );
  NAND2_X1 U13494 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10590) );
  NAND2_X1 U13495 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10589) );
  NAND2_X1 U13496 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10588) );
  AND2_X1 U13497 ( .A1(n10586), .A2(n11768), .ZN(n11729) );
  AOI22_X1 U13498 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10587) );
  AND2_X2 U13499 ( .A1(n11912), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10648) );
  NAND2_X1 U13500 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10596) );
  NAND2_X1 U13501 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10595) );
  NAND2_X1 U13502 ( .A1(n9692), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10723) );
  NAND2_X1 U13503 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10594) );
  NAND2_X1 U13504 ( .A1(n10449), .A2(n13387), .ZN(n11273) );
  INV_X2 U13505 ( .A(n11273), .ZN(n13391) );
  NAND2_X1 U13506 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10593) );
  NAND2_X1 U13507 ( .A1(n9699), .A2(n11178), .ZN(n10600) );
  INV_X1 U13508 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11796) );
  INV_X1 U13509 ( .A(n10774), .ZN(n10601) );
  NAND2_X1 U13510 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10602) );
  OAI211_X1 U13511 ( .C1(n10764), .C2(n11796), .A(n10602), .B(n14265), .ZN(
        n10604) );
  INV_X1 U13512 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14268) );
  INV_X1 U13513 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11625) );
  OAI22_X1 U13514 ( .A1(n14268), .A2(n10765), .B1(n10772), .B2(n11625), .ZN(
        n10603) );
  NOR2_X1 U13515 ( .A1(n10604), .A2(n10603), .ZN(n10617) );
  INV_X1 U13516 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11223) );
  INV_X1 U13517 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11219) );
  INV_X1 U13518 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11632) );
  INV_X1 U13519 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11626) );
  OAI22_X1 U13520 ( .A1(n11632), .A2(n10759), .B1(n20205), .B2(n11626), .ZN(
        n10605) );
  NOR2_X1 U13521 ( .A1(n10606), .A2(n10605), .ZN(n10616) );
  INV_X1 U13522 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11628) );
  INV_X1 U13523 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11216) );
  OAI22_X1 U13524 ( .A1(n11628), .A2(n10760), .B1(n20162), .B2(n11216), .ZN(
        n10610) );
  INV_X1 U13525 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10608) );
  INV_X1 U13526 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10607) );
  OAI22_X1 U13527 ( .A1(n10608), .A2(n10767), .B1(n20136), .B2(n10607), .ZN(
        n10609) );
  NOR2_X1 U13528 ( .A1(n10610), .A2(n10609), .ZN(n10615) );
  INV_X1 U13529 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11803) );
  INV_X1 U13530 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11217) );
  INV_X1 U13531 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10611) );
  INV_X1 U13532 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10629) );
  OAI22_X1 U13533 ( .A1(n10611), .A2(n19991), .B1(n20100), .B2(n10629), .ZN(
        n10612) );
  NOR2_X1 U13534 ( .A1(n10613), .A2(n10612), .ZN(n10614) );
  AOI22_X1 U13535 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11748), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13536 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13537 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11755), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13538 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10618) );
  NAND4_X1 U13539 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10628) );
  AOI22_X1 U13540 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13541 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13542 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11747), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10624) );
  INV_X1 U13543 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13347) );
  INV_X1 U13544 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11607) );
  OAI22_X1 U13545 ( .A1(n10723), .A2(n13347), .B1(n10670), .B2(n11607), .ZN(
        n10622) );
  INV_X1 U13546 ( .A(n10622), .ZN(n10623) );
  NAND4_X1 U13547 ( .A1(n10626), .A2(n10625), .A3(n10624), .A4(n10623), .ZN(
        n10627) );
  OR2_X1 U13548 ( .A1(n11447), .A2(n14265), .ZN(n12844) );
  INV_X1 U13549 ( .A(n12844), .ZN(n10642) );
  AOI22_X1 U13550 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10648), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13551 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11754), .B1(
        n11760), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10633) );
  OAI22_X1 U13552 ( .A1(n11273), .A2(n10629), .B1(n14268), .B2(n11703), .ZN(
        n10630) );
  INV_X1 U13553 ( .A(n10630), .ZN(n10632) );
  AOI22_X1 U13554 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n11700), .ZN(n10631) );
  NAND4_X1 U13555 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10631), .ZN(
        n10640) );
  AOI22_X1 U13556 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11742), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13557 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11718), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13558 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11747), .B1(
        n10643), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10636) );
  INV_X2 U13559 ( .A(n11735), .ZN(n11741) );
  AOI22_X1 U13560 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11741), .B1(
        n11755), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10635) );
  NAND4_X1 U13561 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .ZN(
        n10639) );
  INV_X1 U13562 ( .A(n11446), .ZN(n10641) );
  NAND2_X1 U13563 ( .A1(n10642), .A2(n10641), .ZN(n11444) );
  NAND2_X1 U13564 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10647) );
  NAND2_X1 U13565 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10646) );
  NAND2_X1 U13566 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10645) );
  AOI22_X1 U13567 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10644) );
  NAND2_X1 U13568 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10652) );
  NAND2_X1 U13569 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10651) );
  NAND2_X1 U13570 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10650) );
  NAND2_X1 U13571 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10649) );
  NAND2_X1 U13572 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10655) );
  AOI22_X1 U13573 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n11700), .ZN(n10654) );
  NAND2_X1 U13574 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10653) );
  NAND2_X1 U13575 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10658) );
  NAND2_X1 U13576 ( .A1(n11755), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10657) );
  NAND2_X1 U13577 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10656) );
  NAND2_X1 U13578 ( .A1(n11444), .A2(n11445), .ZN(n10660) );
  NAND2_X1 U13579 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10665) );
  NAND2_X1 U13580 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10664) );
  NAND2_X1 U13581 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10663) );
  AOI22_X1 U13582 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10662) );
  NAND2_X1 U13583 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10669) );
  NAND2_X1 U13584 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10668) );
  NAND2_X1 U13585 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10667) );
  NAND2_X1 U13586 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10666) );
  NAND2_X1 U13587 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10673) );
  AOI22_X1 U13588 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n11700), .ZN(n10672) );
  NAND2_X1 U13589 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10671) );
  NAND2_X1 U13590 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10676) );
  NAND2_X1 U13591 ( .A1(n11755), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10675) );
  NAND2_X1 U13592 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10674) );
  INV_X1 U13593 ( .A(n11189), .ZN(n10880) );
  NOR2_X1 U13594 ( .A1(n14271), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10699) );
  INV_X1 U13595 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n19693) );
  XNOR2_X1 U13596 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U13597 ( .A1(n10976), .A2(n10973), .ZN(n10681) );
  NAND2_X1 U13598 ( .A1(n20481), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10680) );
  NAND2_X1 U13599 ( .A1(n10681), .A2(n10680), .ZN(n10685) );
  MUX2_X1 U13600 ( .A(n20470), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10684) );
  XNOR2_X1 U13601 ( .A(n10685), .B(n10684), .ZN(n10978) );
  MUX2_X1 U13602 ( .A(n10978), .B(n11445), .S(n11423), .Z(n11014) );
  NOR2_X2 U13603 ( .A1(n10704), .A2(n10705), .ZN(n10703) );
  NAND2_X1 U13604 ( .A1(n10685), .A2(n10684), .ZN(n10687) );
  NAND2_X1 U13605 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20470), .ZN(
        n10686) );
  NAND2_X1 U13606 ( .A1(n10687), .A2(n10686), .ZN(n10688) );
  XNOR2_X1 U13607 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10689) );
  INV_X1 U13608 ( .A(n10713), .ZN(n10693) );
  INV_X1 U13609 ( .A(n10688), .ZN(n10691) );
  INV_X1 U13610 ( .A(n10689), .ZN(n10690) );
  NAND2_X1 U13611 ( .A1(n10691), .A2(n10690), .ZN(n10692) );
  NAND2_X1 U13612 ( .A1(n10693), .A2(n10692), .ZN(n10995) );
  MUX2_X1 U13613 ( .A(n11178), .B(n10995), .S(n10694), .Z(n10971) );
  MUX2_X1 U13614 ( .A(n10971), .B(P2_EBX_REG_3__SCAN_IN), .S(n11966), .Z(
        n10695) );
  OAI21_X1 U13615 ( .B1(n10703), .B2(n10696), .A(n10735), .ZN(n14505) );
  INV_X1 U13616 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13411) );
  AND2_X1 U13617 ( .A1(n13411), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10697) );
  NOR2_X1 U13618 ( .A1(n10973), .A2(n10697), .ZN(n11003) );
  INV_X1 U13619 ( .A(n11003), .ZN(n10698) );
  MUX2_X1 U13620 ( .A(n10698), .B(n11447), .S(n11423), .Z(n10700) );
  AOI21_X1 U13621 ( .B1(n10700), .B2(n14271), .A(n10699), .ZN(n14515) );
  NAND2_X1 U13622 ( .A1(n14515), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12837) );
  NAND3_X1 U13623 ( .A1(n11966), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10701) );
  NAND2_X1 U13624 ( .A1(n10704), .A2(n10701), .ZN(n19691) );
  NOR2_X1 U13625 ( .A1(n12837), .A2(n19691), .ZN(n10702) );
  NAND2_X1 U13626 ( .A1(n12837), .A2(n19691), .ZN(n12730) );
  OAI21_X1 U13627 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10702), .A(
        n12730), .ZN(n19842) );
  INV_X1 U13628 ( .A(n10703), .ZN(n10707) );
  NAND2_X1 U13629 ( .A1(n10705), .A2(n10704), .ZN(n10706) );
  NAND2_X1 U13630 ( .A1(n10707), .A2(n10706), .ZN(n14382) );
  INV_X1 U13631 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19876) );
  XNOR2_X1 U13632 ( .A(n14382), .B(n19876), .ZN(n19841) );
  OR2_X1 U13633 ( .A1(n19842), .A2(n19841), .ZN(n19844) );
  INV_X1 U13634 ( .A(n14382), .ZN(n10708) );
  NAND2_X1 U13635 ( .A1(n10708), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10709) );
  AND2_X1 U13636 ( .A1(n19844), .A2(n10709), .ZN(n13350) );
  NAND2_X1 U13637 ( .A1(n13348), .A2(n13350), .ZN(n10712) );
  NAND2_X1 U13638 ( .A1(n10712), .A2(n13349), .ZN(n13482) );
  INV_X1 U13639 ( .A(n13482), .ZN(n10738) );
  NOR2_X1 U13640 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21126), .ZN(
        n21291) );
  NAND2_X1 U13641 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10717) );
  NAND2_X1 U13642 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10716) );
  NAND2_X1 U13643 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10715) );
  AOI22_X1 U13644 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10714) );
  INV_X1 U13645 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10722) );
  NAND2_X1 U13646 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11700), .ZN(
        n10718) );
  OAI21_X1 U13647 ( .B1(n11703), .B2(n11865), .A(n10718), .ZN(n10719) );
  AOI21_X1 U13648 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n10719), .ZN(n10721) );
  NAND2_X1 U13649 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10720) );
  OAI211_X1 U13650 ( .C1(n11699), .C2(n10722), .A(n10721), .B(n10720), .ZN(
        n10726) );
  OAI22_X1 U13651 ( .A1(n10724), .A2(n10723), .B1(n11273), .B2(n11873), .ZN(
        n10725) );
  NOR2_X1 U13652 ( .A1(n10726), .A2(n10725), .ZN(n10732) );
  NAND2_X1 U13653 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10730) );
  NAND2_X1 U13654 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10729) );
  NAND2_X1 U13655 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10728) );
  NAND2_X1 U13656 ( .A1(n11755), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10727) );
  MUX2_X1 U13657 ( .A(n10999), .B(n11456), .S(n11423), .Z(n10972) );
  MUX2_X1 U13658 ( .A(n10972), .B(P2_EBX_REG_4__SCAN_IN), .S(n11966), .Z(
        n10734) );
  AND2_X1 U13659 ( .A1(n10734), .A2(n10735), .ZN(n10736) );
  OR2_X1 U13660 ( .A1(n10736), .A2(n10791), .ZN(n10739) );
  INV_X1 U13661 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13675) );
  XNOR2_X1 U13662 ( .A(n10739), .B(n13675), .ZN(n13483) );
  INV_X1 U13663 ( .A(n13483), .ZN(n10737) );
  NAND2_X1 U13664 ( .A1(n10738), .A2(n10737), .ZN(n10741) );
  INV_X1 U13665 ( .A(n10739), .ZN(n19680) );
  NAND2_X1 U13666 ( .A1(n19680), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10740) );
  NAND2_X1 U13667 ( .A1(n10741), .A2(n10740), .ZN(n13667) );
  INV_X1 U13668 ( .A(n11456), .ZN(n10742) );
  INV_X1 U13669 ( .A(n11454), .ZN(n10787) );
  NAND2_X1 U13670 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10746) );
  NAND2_X1 U13671 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10745) );
  NAND2_X1 U13672 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10744) );
  AOI22_X1 U13673 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10743) );
  NAND2_X1 U13674 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10750) );
  NAND2_X1 U13675 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10749) );
  NAND2_X1 U13676 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10748) );
  NAND2_X1 U13677 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10747) );
  AOI22_X1 U13678 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11754), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10756) );
  NAND2_X1 U13679 ( .A1(n11755), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10754) );
  AOI22_X1 U13680 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10753) );
  NAND2_X1 U13681 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10752) );
  NAND2_X1 U13682 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10751) );
  AND4_X1 U13683 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n10755) );
  NAND4_X1 U13684 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n11182) );
  INV_X1 U13685 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11707) );
  INV_X1 U13686 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11310) );
  OAI22_X1 U13687 ( .A1(n11707), .A2(n10759), .B1(n20162), .B2(n11310), .ZN(
        n10763) );
  INV_X1 U13688 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11702) );
  INV_X1 U13689 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10761) );
  OAI22_X1 U13690 ( .A1(n11702), .A2(n10760), .B1(n20136), .B2(n10761), .ZN(
        n10762) );
  NOR2_X1 U13691 ( .A1(n10763), .A2(n10762), .ZN(n10786) );
  INV_X1 U13692 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10766) );
  INV_X1 U13693 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14274) );
  OAI22_X1 U13694 ( .A1(n10766), .A2(n10764), .B1(n10765), .B2(n14274), .ZN(
        n10771) );
  INV_X1 U13695 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10769) );
  INV_X1 U13696 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10768) );
  OAI22_X1 U13697 ( .A1(n10769), .A2(n10767), .B1(n20257), .B2(n10768), .ZN(
        n10770) );
  NOR2_X1 U13698 ( .A1(n10771), .A2(n10770), .ZN(n10785) );
  INV_X1 U13699 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11894) );
  INV_X1 U13700 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11901) );
  OAI22_X1 U13701 ( .A1(n11894), .A2(n19991), .B1(n10772), .B2(n11901), .ZN(
        n10777) );
  INV_X1 U13702 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11316) );
  INV_X1 U13703 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10775) );
  OAI22_X1 U13704 ( .A1(n11316), .A2(n10773), .B1(n13341), .B2(n10775), .ZN(
        n10776) );
  NOR2_X1 U13705 ( .A1(n10777), .A2(n10776), .ZN(n10784) );
  INV_X1 U13706 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11312) );
  INV_X1 U13707 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11698) );
  OAI22_X1 U13708 ( .A1(n11312), .A2(n10778), .B1(n20205), .B2(n11698), .ZN(
        n10782) );
  INV_X1 U13709 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11309) );
  INV_X1 U13710 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10780) );
  OAI22_X1 U13711 ( .A1(n11309), .A2(n10779), .B1(n20100), .B2(n10780), .ZN(
        n10781) );
  NOR2_X1 U13712 ( .A1(n10782), .A2(n10781), .ZN(n10783) );
  NAND2_X1 U13713 ( .A1(n11454), .A2(n10788), .ZN(n10789) );
  INV_X1 U13714 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13309) );
  MUX2_X1 U13715 ( .A(n13309), .B(n11182), .S(n14271), .Z(n10790) );
  OR2_X1 U13716 ( .A1(n10791), .A2(n10790), .ZN(n10792) );
  NAND2_X1 U13717 ( .A1(n10837), .A2(n10792), .ZN(n14458) );
  INV_X1 U13718 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21051) );
  XNOR2_X1 U13719 ( .A(n10793), .B(n21051), .ZN(n13668) );
  NAND2_X1 U13720 ( .A1(n10793), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10794) );
  INV_X1 U13721 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11725) );
  INV_X1 U13722 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11330) );
  OAI22_X1 U13723 ( .A1(n11725), .A2(n10759), .B1(n20162), .B2(n11330), .ZN(
        n10798) );
  INV_X1 U13724 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10796) );
  INV_X1 U13725 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10795) );
  OAI22_X1 U13726 ( .A1(n10796), .A2(n10760), .B1(n10772), .B2(n10795), .ZN(
        n10797) );
  NOR2_X1 U13727 ( .A1(n10798), .A2(n10797), .ZN(n10812) );
  INV_X1 U13728 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11336) );
  INV_X1 U13729 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11733) );
  OAI22_X1 U13730 ( .A1(n11336), .A2(n10773), .B1(n13341), .B2(n11733), .ZN(
        n10802) );
  INV_X1 U13731 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10800) );
  INV_X1 U13732 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10799) );
  OAI22_X1 U13733 ( .A1(n10800), .A2(n20205), .B1(n20257), .B2(n10799), .ZN(
        n10801) );
  NOR2_X1 U13734 ( .A1(n10802), .A2(n10801), .ZN(n10811) );
  INV_X1 U13735 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11720) );
  INV_X1 U13736 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10824) );
  OAI22_X1 U13737 ( .A1(n11720), .A2(n19991), .B1(n20136), .B2(n10824), .ZN(
        n10804) );
  INV_X1 U13738 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11332) );
  INV_X1 U13739 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11917) );
  OAI22_X1 U13740 ( .A1(n11332), .A2(n10778), .B1(n20100), .B2(n11917), .ZN(
        n10803) );
  NOR2_X1 U13741 ( .A1(n10804), .A2(n10803), .ZN(n10810) );
  INV_X1 U13742 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13317) );
  INV_X1 U13743 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10805) );
  OAI22_X1 U13744 ( .A1(n13317), .A2(n10765), .B1(n10764), .B2(n10805), .ZN(
        n10808) );
  INV_X1 U13745 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10806) );
  INV_X1 U13746 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11329) );
  OAI22_X1 U13747 ( .A1(n10806), .A2(n10767), .B1(n10779), .B2(n11329), .ZN(
        n10807) );
  NOR2_X1 U13748 ( .A1(n10808), .A2(n10807), .ZN(n10809) );
  NAND4_X1 U13749 ( .A1(n10812), .A2(n10811), .A3(n10810), .A4(n10809), .ZN(
        n10835) );
  NAND2_X1 U13750 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10816) );
  NAND2_X1 U13751 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10815) );
  NAND2_X1 U13752 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10814) );
  AOI22_X1 U13753 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10813) );
  NAND4_X1 U13754 ( .A1(n10816), .A2(n10815), .A3(n10814), .A4(n10813), .ZN(
        n10822) );
  NAND2_X1 U13755 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10820) );
  NAND2_X1 U13756 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10819) );
  NAND2_X1 U13757 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10818) );
  NAND2_X1 U13758 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10817) );
  NAND4_X1 U13759 ( .A1(n10820), .A2(n10819), .A3(n10818), .A4(n10817), .ZN(
        n10821) );
  NOR2_X1 U13760 ( .A1(n10822), .A2(n10821), .ZN(n10833) );
  NAND2_X1 U13761 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10823) );
  OAI21_X1 U13762 ( .B1(n10824), .B2(n11699), .A(n10823), .ZN(n10831) );
  NAND2_X1 U13763 ( .A1(n11755), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10828) );
  NAND2_X1 U13764 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n11700), .ZN(
        n10825) );
  OAI21_X1 U13765 ( .B1(n11703), .B2(n13317), .A(n10825), .ZN(n10826) );
  AOI21_X1 U13766 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n10826), .ZN(n10827) );
  OAI211_X1 U13767 ( .C1(n11720), .C2(n10829), .A(n10828), .B(n10827), .ZN(
        n10830) );
  NOR2_X1 U13768 ( .A1(n10831), .A2(n10830), .ZN(n10832) );
  NAND2_X1 U13769 ( .A1(n9699), .A2(n11185), .ZN(n10834) );
  MUX2_X1 U13770 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n11185), .S(n14271), .Z(
        n10836) );
  NAND2_X1 U13771 ( .A1(n10837), .A2(n10836), .ZN(n10838) );
  NAND2_X1 U13772 ( .A1(n10844), .A2(n10838), .ZN(n14286) );
  INV_X1 U13773 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11408) );
  NAND2_X1 U13774 ( .A1(n10839), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10840) );
  MUX2_X1 U13775 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n11189), .S(n14271), .Z(
        n10843) );
  XNOR2_X1 U13776 ( .A(n10844), .B(n10110), .ZN(n14481) );
  INV_X1 U13777 ( .A(n14481), .ZN(n10842) );
  INV_X1 U13778 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10841) );
  NAND2_X1 U13779 ( .A1(n10842), .A2(n10841), .ZN(n14292) );
  NAND2_X1 U13780 ( .A1(n11966), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10846) );
  AND2_X2 U13781 ( .A1(n10845), .A2(n10846), .ZN(n10853) );
  NOR2_X1 U13782 ( .A1(n10845), .A2(n10846), .ZN(n10847) );
  OR2_X1 U13783 ( .A1(n10853), .A2(n10847), .ZN(n19653) );
  NOR2_X1 U13784 ( .A1(n19653), .A2(n11189), .ZN(n10848) );
  NAND2_X1 U13785 ( .A1(n10848), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14435) );
  INV_X1 U13786 ( .A(n10848), .ZN(n10850) );
  INV_X1 U13787 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10849) );
  NAND2_X1 U13788 ( .A1(n10850), .A2(n10849), .ZN(n14434) );
  INV_X1 U13789 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13302) );
  NOR2_X1 U13790 ( .A1(n14271), .A2(n13302), .ZN(n10851) );
  XNOR2_X1 U13791 ( .A(n10853), .B(n10851), .ZN(n14470) );
  AOI21_X1 U13792 ( .B1(n14470), .B2(n10880), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16506) );
  INV_X1 U13793 ( .A(n16506), .ZN(n10852) );
  NAND3_X1 U13794 ( .A1(n10857), .A2(P2_EBX_REG_10__SCAN_IN), .A3(n11966), 
        .ZN(n10855) );
  INV_X1 U13795 ( .A(n10845), .ZN(n10854) );
  OAI211_X1 U13796 ( .C1(n10857), .C2(P2_EBX_REG_10__SCAN_IN), .A(n10855), .B(
        n10945), .ZN(n19641) );
  OR2_X1 U13797 ( .A1(n19641), .A2(n11189), .ZN(n10856) );
  INV_X1 U13798 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16492) );
  INV_X1 U13799 ( .A(n10866), .ZN(n10858) );
  INV_X1 U13800 ( .A(n10868), .ZN(n10861) );
  NAND3_X1 U13801 ( .A1(n11966), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10859), 
        .ZN(n10860) );
  NAND2_X1 U13802 ( .A1(n10861), .A2(n10860), .ZN(n19629) );
  NOR2_X1 U13803 ( .A1(n19629), .A2(n11189), .ZN(n10863) );
  INV_X1 U13804 ( .A(n10863), .ZN(n10862) );
  INV_X1 U13805 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16478) );
  AND2_X1 U13806 ( .A1(n10863), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16469) );
  OR3_X1 U13807 ( .A1(n19641), .A2(n11189), .A3(n16492), .ZN(n16485) );
  INV_X1 U13808 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10864) );
  NOR2_X1 U13809 ( .A1(n11189), .A2(n10864), .ZN(n10865) );
  NAND2_X1 U13810 ( .A1(n14470), .A2(n10865), .ZN(n16504) );
  NAND2_X1 U13811 ( .A1(n16485), .A2(n16504), .ZN(n16467) );
  NAND2_X1 U13812 ( .A1(n11966), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10867) );
  OR2_X1 U13813 ( .A1(n10866), .A2(n10867), .ZN(n10869) );
  NAND2_X1 U13814 ( .A1(n10869), .A2(n10872), .ZN(n19619) );
  NOR2_X1 U13815 ( .A1(n19619), .A2(n11189), .ZN(n10870) );
  NAND2_X1 U13816 ( .A1(n10870), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16993) );
  NOR2_X1 U13817 ( .A1(n10870), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16994) );
  INV_X1 U13818 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10871) );
  NOR2_X1 U13819 ( .A1(n14271), .A2(n10871), .ZN(n10902) );
  NAND2_X1 U13820 ( .A1(n11966), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10900) );
  INV_X1 U13821 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10873) );
  NOR2_X1 U13822 ( .A1(n14271), .A2(n10873), .ZN(n10896) );
  OR2_X2 U13823 ( .A1(n10898), .A2(n10896), .ZN(n10891) );
  INV_X1 U13824 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10874) );
  NOR2_X1 U13825 ( .A1(n14271), .A2(n10874), .ZN(n10875) );
  INV_X1 U13826 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10876) );
  NOR2_X1 U13827 ( .A1(n14271), .A2(n10876), .ZN(n10893) );
  NAND2_X1 U13828 ( .A1(n11966), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10881) );
  INV_X1 U13829 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n16969) );
  INV_X1 U13830 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10885) );
  INV_X1 U13831 ( .A(n10925), .ZN(n10878) );
  NAND3_X1 U13832 ( .A1(n10889), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n11966), 
        .ZN(n10877) );
  INV_X1 U13833 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16373) );
  OAI21_X1 U13834 ( .B1(n15972), .B2(n11189), .A(n16373), .ZN(n16240) );
  NAND2_X1 U13835 ( .A1(n11966), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10879) );
  XNOR2_X1 U13836 ( .A(n9749), .B(n10879), .ZN(n15987) );
  NOR2_X1 U13837 ( .A1(n10919), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16263) );
  INV_X1 U13838 ( .A(n10881), .ZN(n10882) );
  NAND2_X1 U13839 ( .A1(n9752), .A2(n10882), .ZN(n10883) );
  AOI21_X1 U13840 ( .B1(n10914), .B2(n10880), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16273) );
  NOR2_X1 U13841 ( .A1(n16263), .A2(n16273), .ZN(n16249) );
  INV_X1 U13842 ( .A(n10884), .ZN(n10887) );
  NOR2_X1 U13843 ( .A1(n14271), .A2(n10885), .ZN(n10886) );
  INV_X1 U13844 ( .A(n10945), .ZN(n10935) );
  AOI21_X1 U13845 ( .B1(n10887), .B2(n10886), .A(n10935), .ZN(n10888) );
  AND2_X1 U13846 ( .A1(n10889), .A2(n10888), .ZN(n10907) );
  AOI21_X1 U13847 ( .B1(n10907), .B2(n10880), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16238) );
  NAND3_X1 U13848 ( .A1(n10891), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n11966), 
        .ZN(n10890) );
  OAI211_X1 U13849 ( .C1(n10891), .C2(P2_EBX_REG_16__SCAN_IN), .A(n10890), .B(
        n10945), .ZN(n19602) );
  OR2_X1 U13850 ( .A1(n19602), .A2(n11189), .ZN(n10892) );
  INV_X1 U13851 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16444) );
  XNOR2_X1 U13852 ( .A(n10892), .B(n16444), .ZN(n16232) );
  NAND2_X1 U13853 ( .A1(n10894), .A2(n10893), .ZN(n10895) );
  NAND2_X1 U13854 ( .A1(n9752), .A2(n10895), .ZN(n16020) );
  INV_X1 U13855 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16441) );
  NAND2_X1 U13856 ( .A1(n10915), .A2(n16441), .ZN(n16235) );
  INV_X1 U13857 ( .A(n10896), .ZN(n10897) );
  XNOR2_X1 U13858 ( .A(n10898), .B(n10897), .ZN(n10911) );
  NAND2_X1 U13859 ( .A1(n10911), .A2(n10880), .ZN(n10899) );
  INV_X1 U13860 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16459) );
  NAND2_X1 U13861 ( .A1(n10899), .A2(n16459), .ZN(n16301) );
  XNOR2_X1 U13862 ( .A(n9718), .B(n10900), .ZN(n19609) );
  NAND2_X1 U13863 ( .A1(n19609), .A2(n10880), .ZN(n10901) );
  INV_X1 U13864 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17059) );
  NAND2_X1 U13865 ( .A1(n10901), .A2(n17059), .ZN(n16980) );
  NAND2_X1 U13866 ( .A1(n10872), .A2(n10902), .ZN(n10903) );
  NAND2_X1 U13867 ( .A1(n9718), .A2(n10903), .ZN(n14499) );
  OR2_X1 U13868 ( .A1(n14499), .A2(n11189), .ZN(n10904) );
  INV_X1 U13869 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17068) );
  NAND2_X1 U13870 ( .A1(n10904), .A2(n17068), .ZN(n16987) );
  NAND4_X1 U13871 ( .A1(n16235), .A2(n16301), .A3(n16980), .A4(n16987), .ZN(
        n10905) );
  NOR3_X1 U13872 ( .A1(n16238), .A2(n16232), .A3(n10905), .ZN(n10906) );
  INV_X1 U13873 ( .A(n10907), .ZN(n15986) );
  INV_X1 U13874 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10908) );
  OR2_X1 U13875 ( .A1(n11189), .A2(n10908), .ZN(n10909) );
  OR2_X1 U13876 ( .A1(n11189), .A2(n16444), .ZN(n10910) );
  OR2_X1 U13877 ( .A1(n19602), .A2(n10910), .ZN(n16233) );
  INV_X1 U13878 ( .A(n10911), .ZN(n14328) );
  NOR2_X1 U13879 ( .A1(n11189), .A2(n17059), .ZN(n10912) );
  NAND2_X1 U13880 ( .A1(n19609), .A2(n10912), .ZN(n16979) );
  OR2_X1 U13881 ( .A1(n11189), .A2(n17068), .ZN(n10913) );
  OR2_X1 U13882 ( .A1(n14499), .A2(n10913), .ZN(n16986) );
  AND4_X1 U13883 ( .A1(n16233), .A2(n16300), .A3(n16979), .A4(n16986), .ZN(
        n10917) );
  INV_X1 U13884 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16420) );
  INV_X1 U13885 ( .A(n10915), .ZN(n10916) );
  NAND2_X1 U13886 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16236) );
  NAND4_X1 U13887 ( .A1(n16247), .A2(n10917), .A3(n16260), .A4(n16236), .ZN(
        n10922) );
  OR2_X1 U13888 ( .A1(n11189), .A2(n16373), .ZN(n10918) );
  INV_X1 U13889 ( .A(n16262), .ZN(n10920) );
  NAND2_X1 U13890 ( .A1(n11966), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10924) );
  INV_X1 U13891 ( .A(n10930), .ZN(n10926) );
  AOI21_X1 U13892 ( .B1(n10115), .B2(n10927), .A(n10926), .ZN(n16607) );
  AOI21_X1 U13893 ( .B1(n16607), .B2(n10880), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16215) );
  NAND3_X1 U13894 ( .A1(n16607), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n10880), .ZN(n16216) );
  INV_X1 U13895 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10928) );
  NOR2_X1 U13896 ( .A1(n14271), .A2(n10928), .ZN(n10929) );
  NAND2_X1 U13897 ( .A1(n10930), .A2(n10929), .ZN(n10931) );
  NAND2_X1 U13898 ( .A1(n10933), .A2(n10880), .ZN(n10932) );
  XNOR2_X1 U13899 ( .A(n10932), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16208) );
  INV_X1 U13900 ( .A(n10933), .ZN(n16947) );
  INV_X1 U13901 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16363) );
  NOR3_X1 U13902 ( .A1(n16947), .A2(n11189), .A3(n16363), .ZN(n10934) );
  NOR2_X1 U13903 ( .A1(n10935), .A2(n11189), .ZN(n16196) );
  INV_X1 U13904 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16195) );
  INV_X1 U13905 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10941) );
  NAND3_X1 U13906 ( .A1(n11966), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10947), 
        .ZN(n10938) );
  INV_X1 U13907 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16327) );
  NOR3_X1 U13908 ( .A1(n10939), .A2(n11189), .A3(n16327), .ZN(n10962) );
  INV_X1 U13909 ( .A(n10939), .ZN(n15944) );
  AOI21_X1 U13910 ( .B1(n15944), .B2(n10880), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10940) );
  NOR2_X1 U13911 ( .A1(n10962), .A2(n10940), .ZN(n16180) );
  NOR2_X1 U13912 ( .A1(n10942), .A2(n10941), .ZN(n10943) );
  NAND2_X1 U13913 ( .A1(n11966), .A2(n10943), .ZN(n10944) );
  AND2_X1 U13914 ( .A1(n10945), .A2(n10944), .ZN(n10946) );
  NAND2_X1 U13915 ( .A1(n10947), .A2(n10946), .ZN(n16929) );
  INV_X1 U13916 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16339) );
  NAND2_X1 U13917 ( .A1(n10960), .A2(n16339), .ZN(n16184) );
  NAND2_X1 U13918 ( .A1(n11966), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10949) );
  INV_X1 U13919 ( .A(n10949), .ZN(n10950) );
  NAND2_X1 U13920 ( .A1(n10950), .A2(n9748), .ZN(n10951) );
  NAND2_X1 U13921 ( .A1(n10956), .A2(n10951), .ZN(n16924) );
  INV_X1 U13922 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16312) );
  INV_X1 U13923 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12405) );
  NAND2_X1 U13924 ( .A1(n11966), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10954) );
  INV_X1 U13925 ( .A(n10954), .ZN(n10955) );
  NAND2_X1 U13926 ( .A1(n10956), .A2(n10955), .ZN(n10957) );
  NAND2_X1 U13927 ( .A1(n10964), .A2(n10957), .ZN(n16912) );
  AOI21_X1 U13928 ( .B1(n12405), .B2(n16312), .A(n11505), .ZN(n10959) );
  INV_X1 U13929 ( .A(n11505), .ZN(n10958) );
  INV_X1 U13930 ( .A(n10960), .ZN(n10961) );
  NOR2_X1 U13931 ( .A1(n16186), .A2(n10962), .ZN(n11499) );
  INV_X1 U13932 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11130) );
  NOR2_X1 U13933 ( .A1(n14271), .A2(n11130), .ZN(n10965) );
  XNOR2_X1 U13934 ( .A(n10964), .B(n10965), .ZN(n10963) );
  INV_X1 U13935 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12406) );
  OAI21_X1 U13936 ( .B1(n10963), .B2(n11189), .A(n12406), .ZN(n12395) );
  INV_X1 U13937 ( .A(n10963), .ZN(n16893) );
  NAND3_X1 U13938 ( .A1(n16893), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10880), .ZN(n12394) );
  NAND2_X1 U13939 ( .A1(n11522), .A2(n12394), .ZN(n10970) );
  NAND2_X1 U13940 ( .A1(n11966), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10966) );
  XNOR2_X1 U13941 ( .A(n11523), .B(n10966), .ZN(n12033) );
  AOI21_X1 U13942 ( .B1(n12033), .B2(n10880), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11521) );
  INV_X1 U13943 ( .A(n11521), .ZN(n10968) );
  INV_X1 U13944 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11556) );
  NOR2_X1 U13945 ( .A1(n11189), .A2(n11556), .ZN(n10967) );
  NAND2_X1 U13946 ( .A1(n10968), .A2(n11518), .ZN(n10969) );
  XNOR2_X1 U13947 ( .A(n10970), .B(n10969), .ZN(n11487) );
  NOR2_X1 U13948 ( .A1(n10972), .A2(n10971), .ZN(n11017) );
  INV_X1 U13949 ( .A(n10973), .ZN(n10974) );
  XNOR2_X1 U13950 ( .A(n10976), .B(n10974), .ZN(n11000) );
  OAI21_X1 U13951 ( .B1(n14265), .B2(n11003), .A(n11000), .ZN(n10975) );
  OAI21_X1 U13952 ( .B1(n14265), .B2(n10978), .A(n10975), .ZN(n10977) );
  NAND2_X1 U13953 ( .A1(n11003), .A2(n10976), .ZN(n11013) );
  AOI22_X1 U13954 ( .A1(n10977), .A2(n11024), .B1(n11423), .B2(n11013), .ZN(
        n10982) );
  NAND2_X1 U13955 ( .A1(n12713), .A2(n14265), .ZN(n10979) );
  INV_X1 U13956 ( .A(n10978), .ZN(n10996) );
  MUX2_X1 U13957 ( .A(n10979), .B(n10694), .S(n10996), .Z(n10980) );
  INV_X1 U13958 ( .A(n10980), .ZN(n10981) );
  NOR2_X1 U13959 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  OAI22_X1 U13960 ( .A1(n11017), .A2(n11423), .B1(n10983), .B2(n10995), .ZN(
        n10986) );
  OAI22_X1 U13961 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21165), .B1(
        n21291), .B2(n10984), .ZN(n11015) );
  INV_X1 U13962 ( .A(n11015), .ZN(n11002) );
  NAND2_X1 U13963 ( .A1(n10999), .A2(n11423), .ZN(n10985) );
  NAND3_X1 U13964 ( .A1(n10986), .A2(n11002), .A3(n10985), .ZN(n10987) );
  MUX2_X1 U13965 ( .A(n10987), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n17100), .Z(n10990) );
  NAND2_X1 U13966 ( .A1(n11015), .A2(n10988), .ZN(n10989) );
  NAND2_X1 U13967 ( .A1(n13219), .A2(n14265), .ZN(n12710) );
  INV_X1 U13968 ( .A(n10990), .ZN(n10991) );
  NAND2_X1 U13969 ( .A1(n12710), .A2(n10991), .ZN(n10992) );
  OAI21_X1 U13970 ( .B1(n11024), .B2(n13219), .A(n10992), .ZN(n10994) );
  NAND2_X1 U13971 ( .A1(n10994), .A2(n10993), .ZN(n11040) );
  INV_X1 U13972 ( .A(n10995), .ZN(n10997) );
  NAND2_X1 U13973 ( .A1(n10997), .A2(n10996), .ZN(n10998) );
  NOR2_X1 U13974 ( .A1(n10999), .A2(n10998), .ZN(n11004) );
  NAND2_X1 U13975 ( .A1(n11004), .A2(n11000), .ZN(n11001) );
  NAND2_X1 U13976 ( .A1(n11002), .A2(n11001), .ZN(n13434) );
  AND2_X1 U13977 ( .A1(n11004), .A2(n11003), .ZN(n11005) );
  OAI21_X1 U13978 ( .B1(n13434), .B2(n11005), .A(n11007), .ZN(n11009) );
  NOR2_X1 U13979 ( .A1(n11007), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(n11008) );
  OAI21_X1 U13980 ( .B1(n11740), .B2(n9812), .A(n11008), .ZN(n20483) );
  AND2_X1 U13981 ( .A1(n11009), .A2(n20483), .ZN(n20502) );
  NOR2_X1 U13982 ( .A1(n11011), .A2(n9699), .ZN(n11012) );
  NAND2_X1 U13983 ( .A1(n20502), .A2(n11012), .ZN(n11019) );
  NAND2_X1 U13984 ( .A1(n11014), .A2(n11013), .ZN(n11016) );
  AOI21_X1 U13985 ( .B1(n11017), .B2(n11016), .A(n11015), .ZN(n20498) );
  INV_X1 U13986 ( .A(n12019), .ZN(n13443) );
  NOR2_X1 U13987 ( .A1(n11011), .A2(n13443), .ZN(n20496) );
  NAND2_X1 U13988 ( .A1(n20498), .A2(n20496), .ZN(n11018) );
  NAND2_X1 U13989 ( .A1(n11019), .A2(n11018), .ZN(n11486) );
  NAND2_X1 U13990 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20373) );
  INV_X1 U13991 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20374) );
  INV_X1 U13992 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20395) );
  NOR2_X1 U13993 ( .A1(n20374), .A2(n20395), .ZN(n20384) );
  NOR2_X1 U13994 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20387) );
  NOR3_X1 U13995 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20384), .A3(n20387), 
        .ZN(n12711) );
  NAND2_X1 U13996 ( .A1(n20373), .A2(n12711), .ZN(n13444) );
  INV_X1 U13997 ( .A(n13444), .ZN(n13432) );
  NAND2_X1 U13998 ( .A1(n11020), .A2(n13432), .ZN(n11021) );
  OR2_X1 U13999 ( .A1(n13434), .A2(n11021), .ZN(n11034) );
  OAI21_X1 U14000 ( .B1(n11023), .B2(n19880), .A(n11022), .ZN(n11032) );
  NAND2_X1 U14001 ( .A1(n9699), .A2(n10993), .ZN(n11409) );
  NAND2_X1 U14002 ( .A1(n11409), .A2(n11024), .ZN(n11025) );
  NAND2_X1 U14003 ( .A1(n11025), .A2(n19905), .ZN(n11027) );
  AOI21_X1 U14004 ( .B1(n11027), .B2(n11026), .A(n10466), .ZN(n11031) );
  NAND2_X1 U14005 ( .A1(n11028), .A2(n19905), .ZN(n11029) );
  NAND2_X1 U14006 ( .A1(n11029), .A2(n12019), .ZN(n11415) );
  NAND2_X1 U14007 ( .A1(n10401), .A2(n10474), .ZN(n11030) );
  NAND4_X1 U14008 ( .A1(n11032), .A2(n11031), .A3(n11415), .A4(n11030), .ZN(
        n11410) );
  INV_X1 U14009 ( .A(n11410), .ZN(n11033) );
  AND2_X1 U14010 ( .A1(n11034), .A2(n11033), .ZN(n12741) );
  MUX2_X1 U14011 ( .A(n11020), .B(n19880), .S(n9699), .Z(n11035) );
  INV_X1 U14012 ( .A(n13434), .ZN(n13424) );
  NAND3_X1 U14013 ( .A1(n11035), .A2(n13424), .A3(n20373), .ZN(n11036) );
  NAND2_X1 U14014 ( .A1(n12741), .A2(n11036), .ZN(n11037) );
  NOR2_X1 U14015 ( .A1(n11486), .A2(n11037), .ZN(n11039) );
  INV_X1 U14016 ( .A(n12710), .ZN(n12740) );
  NAND3_X1 U14017 ( .A1(n12740), .A2(n19880), .A3(n13432), .ZN(n11038) );
  NAND3_X1 U14018 ( .A1(n11040), .A2(n11039), .A3(n11038), .ZN(n11041) );
  OR2_X1 U14019 ( .A1(n19558), .A2(n20312), .ZN(n19561) );
  NOR2_X1 U14020 ( .A1(n11011), .A2(n10694), .ZN(n20495) );
  NAND2_X1 U14021 ( .A1(n11487), .A2(n19866), .ZN(n11485) );
  NAND2_X1 U14022 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11045) );
  AND2_X1 U14023 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11043) );
  AOI21_X1 U14024 ( .B1(n11534), .B2(P2_REIP_REG_10__SCAN_IN), .A(n11043), 
        .ZN(n11044) );
  OAI211_X1 U14025 ( .C1(n11134), .C2(n10104), .A(n11045), .B(n11044), .ZN(
        n13313) );
  NAND2_X1 U14026 ( .A1(n11046), .A2(n11047), .ZN(n11052) );
  INV_X1 U14027 ( .A(n11048), .ZN(n11050) );
  NAND2_X1 U14028 ( .A1(n11050), .A2(n11049), .ZN(n11051) );
  NAND2_X1 U14029 ( .A1(n11052), .A2(n11051), .ZN(n13488) );
  AOI22_X1 U14030 ( .A1(n11534), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11055) );
  NAND2_X1 U14031 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11054) );
  NAND2_X1 U14032 ( .A1(n11536), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14033 ( .A1(n11534), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11060) );
  NAND2_X1 U14034 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11059) );
  NAND2_X1 U14035 ( .A1(n11536), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14036 ( .A1(n11534), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11064) );
  NAND2_X1 U14037 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11063) );
  NAND2_X1 U14038 ( .A1(n11536), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11062) );
  INV_X1 U14039 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U14040 ( .A1(n11534), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11066) );
  NAND2_X1 U14041 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11065) );
  OAI211_X1 U14042 ( .C1(n13325), .C2(n11134), .A(n11066), .B(n11065), .ZN(
        n13319) );
  INV_X1 U14043 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11069) );
  INV_X2 U14044 ( .A(n11100), .ZN(n11534) );
  AOI22_X1 U14045 ( .A1(n11534), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11068) );
  NAND2_X1 U14046 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11067) );
  OAI211_X1 U14047 ( .C1(n11069), .C2(n11134), .A(n11068), .B(n11067), .ZN(
        n13285) );
  AOI22_X1 U14048 ( .A1(n11534), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11072) );
  NAND2_X1 U14049 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11071) );
  NAND2_X1 U14050 ( .A1(n11536), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14051 ( .A1(n11534), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11074) );
  NAND2_X1 U14052 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11073) );
  OAI211_X1 U14053 ( .C1(n11134), .C2(n10102), .A(n11074), .B(n11073), .ZN(
        n13473) );
  AND2_X2 U14054 ( .A1(n13474), .A2(n13473), .ZN(n13476) );
  INV_X1 U14055 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14056 ( .A1(n11534), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11076) );
  NAND2_X1 U14057 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11075) );
  OAI211_X1 U14058 ( .C1(n11134), .C2(n11077), .A(n11076), .B(n11075), .ZN(
        n13468) );
  AOI22_X1 U14059 ( .A1(n11534), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11080) );
  NAND2_X1 U14060 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11079) );
  NAND2_X1 U14061 ( .A1(n11536), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11078) );
  INV_X1 U14062 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U14063 ( .A1(n11534), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11082) );
  NAND2_X1 U14064 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11081) );
  OAI211_X1 U14065 ( .C1(n11134), .C2(n11083), .A(n11082), .B(n11081), .ZN(
        n13664) );
  AOI22_X1 U14066 ( .A1(n11534), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11086) );
  NAND2_X1 U14067 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11085) );
  NAND2_X1 U14068 ( .A1(n11536), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14069 ( .A1(n11534), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11089) );
  NAND2_X1 U14070 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11088) );
  NAND2_X1 U14071 ( .A1(n11536), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U14072 ( .A1(n11534), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11093) );
  NAND2_X1 U14073 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11092) );
  NAND2_X1 U14074 ( .A1(n11536), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11091) );
  INV_X1 U14075 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U14076 ( .A1(n11534), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11095) );
  NAND2_X1 U14077 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11094) );
  OAI211_X1 U14078 ( .C1(n11134), .C2(n11096), .A(n11095), .B(n11094), .ZN(
        n16073) );
  AOI22_X1 U14079 ( .A1(n11534), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11099) );
  NAND2_X1 U14080 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11098) );
  NAND2_X1 U14081 ( .A1(n11536), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14082 ( .A1(n11534), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11103) );
  NAND2_X1 U14083 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11102) );
  NAND2_X1 U14084 ( .A1(n11536), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11101) );
  INV_X1 U14085 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14086 ( .A1(n11534), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11105) );
  NAND2_X1 U14087 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11104) );
  OAI211_X1 U14088 ( .C1(n11134), .C2(n11106), .A(n11105), .B(n11104), .ZN(
        n15965) );
  INV_X1 U14089 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11109) );
  AOI22_X1 U14090 ( .A1(n11534), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11108) );
  NAND2_X1 U14091 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11107) );
  OAI211_X1 U14092 ( .C1(n11134), .C2(n11109), .A(n11108), .B(n11107), .ZN(
        n16063) );
  AOI22_X1 U14093 ( .A1(n11534), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11113) );
  NAND2_X1 U14094 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11112) );
  NAND2_X1 U14095 ( .A1(n11536), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11111) );
  AND3_X1 U14096 ( .A1(n11113), .A2(n11112), .A3(n11111), .ZN(n16055) );
  AOI22_X1 U14097 ( .A1(n11534), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11116) );
  NAND2_X1 U14098 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11115) );
  NAND2_X1 U14099 ( .A1(n11536), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14100 ( .A1(n11534), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11118) );
  NAND2_X1 U14101 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11117) );
  OAI211_X1 U14102 ( .C1(n11134), .C2(n10941), .A(n11118), .B(n11117), .ZN(
        n16048) );
  AOI22_X1 U14103 ( .A1(n11534), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11121) );
  NAND2_X1 U14104 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11120) );
  NAND2_X1 U14105 ( .A1(n11536), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11119) );
  AND3_X1 U14106 ( .A1(n11121), .A2(n11120), .A3(n11119), .ZN(n15931) );
  OR2_X2 U14107 ( .A1(n15930), .A2(n15931), .ZN(n16033) );
  AOI22_X1 U14108 ( .A1(n11534), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11124) );
  NAND2_X1 U14109 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U14110 ( .A1(n11536), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11122) );
  AND3_X1 U14111 ( .A1(n11124), .A2(n11123), .A3(n11122), .ZN(n16032) );
  AOI22_X1 U14112 ( .A1(n11534), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11127) );
  NAND2_X1 U14113 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11126) );
  NAND2_X1 U14114 ( .A1(n11536), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11125) );
  AND3_X1 U14115 ( .A1(n11127), .A2(n11126), .A3(n11125), .ZN(n11507) );
  AOI22_X1 U14116 ( .A1(n11534), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11129) );
  NAND2_X1 U14117 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11128) );
  OAI211_X1 U14118 ( .C1(n11134), .C2(n11130), .A(n11129), .B(n11128), .ZN(
        n12388) );
  INV_X1 U14119 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U14120 ( .A1(n11534), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11132) );
  NAND2_X1 U14121 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11131) );
  OAI211_X1 U14122 ( .C1(n11134), .C2(n11133), .A(n11132), .B(n11131), .ZN(
        n11532) );
  NAND2_X1 U14123 ( .A1(n13413), .A2(n9699), .ZN(n11138) );
  INV_X1 U14124 ( .A(n13384), .ZN(n11137) );
  NAND2_X1 U14125 ( .A1(n11138), .A2(n11137), .ZN(n11139) );
  NAND2_X1 U14126 ( .A1(n11482), .A2(n11139), .ZN(n19870) );
  NAND2_X1 U14127 ( .A1(n11170), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11142) );
  AND2_X2 U14128 ( .A1(n10485), .A2(n20101), .ZN(n11157) );
  AOI22_X1 U14129 ( .A1(n11143), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n11157), .ZN(n11141) );
  AND2_X1 U14130 ( .A1(n11142), .A2(n11141), .ZN(n11402) );
  NAND2_X1 U14131 ( .A1(n11143), .A2(P2_EAX_REG_4__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U14132 ( .A1(n11157), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11144) );
  OAI211_X1 U14133 ( .C1(n11376), .C2(n11456), .A(n11145), .B(n11144), .ZN(
        n11146) );
  INV_X1 U14134 ( .A(n11146), .ZN(n11148) );
  NAND2_X1 U14135 ( .A1(n11170), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11147) );
  MUX2_X1 U14136 ( .A(n19905), .B(n20492), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11150) );
  INV_X1 U14137 ( .A(n11149), .ZN(n11162) );
  NAND2_X1 U14138 ( .A1(n11162), .A2(n11157), .ZN(n11168) );
  AND2_X1 U14139 ( .A1(n11150), .A2(n11168), .ZN(n11151) );
  NAND2_X1 U14140 ( .A1(n11170), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11156) );
  INV_X1 U14141 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19817) );
  NAND2_X1 U14142 ( .A1(n14265), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11153) );
  OAI211_X1 U14143 ( .C1(n19905), .C2(n19817), .A(n20101), .B(n11153), .ZN(
        n11154) );
  INV_X1 U14144 ( .A(n11154), .ZN(n11155) );
  NAND2_X1 U14145 ( .A1(n11156), .A2(n11155), .ZN(n12839) );
  INV_X1 U14146 ( .A(n11161), .ZN(n12842) );
  INV_X1 U14147 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20396) );
  NAND2_X1 U14148 ( .A1(n11170), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11159) );
  AOI22_X1 U14149 ( .A1(n11143), .A2(P2_EAX_REG_1__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11157), .ZN(n11158) );
  NAND2_X1 U14150 ( .A1(n11159), .A2(n11158), .ZN(n11160) );
  NOR2_X1 U14151 ( .A1(n12842), .A2(n11160), .ZN(n11167) );
  OR2_X1 U14152 ( .A1(n11446), .A2(n11376), .ZN(n11165) );
  NAND2_X1 U14153 ( .A1(n11149), .A2(n19905), .ZN(n11163) );
  MUX2_X1 U14154 ( .A(n11163), .B(n20481), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11164) );
  NAND2_X1 U14155 ( .A1(n11165), .A2(n11164), .ZN(n12964) );
  INV_X1 U14156 ( .A(n12964), .ZN(n11166) );
  NAND2_X1 U14157 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11169) );
  OAI211_X1 U14158 ( .C1(n11376), .C2(n11445), .A(n11169), .B(n11168), .ZN(
        n11173) );
  XNOR2_X1 U14159 ( .A(n11174), .B(n11173), .ZN(n12988) );
  NAND2_X1 U14160 ( .A1(n11170), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14161 ( .A1(n11143), .A2(P2_EAX_REG_2__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n11157), .ZN(n11171) );
  NAND2_X1 U14162 ( .A1(n11172), .A2(n11171), .ZN(n12987) );
  NOR2_X1 U14163 ( .A1(n12988), .A2(n12987), .ZN(n12989) );
  NOR2_X1 U14164 ( .A1(n11174), .A2(n11173), .ZN(n11175) );
  NAND2_X1 U14165 ( .A1(n11143), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U14166 ( .A1(n11157), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11176) );
  OAI211_X1 U14167 ( .C1(n11178), .C2(n11376), .A(n11177), .B(n11176), .ZN(
        n11179) );
  INV_X1 U14168 ( .A(n11179), .ZN(n11181) );
  NAND2_X1 U14169 ( .A1(n11170), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11180) );
  NAND2_X1 U14170 ( .A1(n11181), .A2(n11180), .ZN(n13352) );
  AOI22_X1 U14171 ( .A1(n11170), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11143), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U14172 ( .A1(n10218), .A2(n11182), .B1(n11157), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11183) );
  NAND2_X1 U14173 ( .A1(n11184), .A2(n11183), .ZN(n13680) );
  OR2_X1 U14174 ( .A1(n11376), .A2(n11185), .ZN(n11186) );
  NAND2_X1 U14175 ( .A1(n11170), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14176 ( .A1(n11143), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11157), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11187) );
  NAND2_X1 U14177 ( .A1(n11188), .A2(n11187), .ZN(n14091) );
  NAND2_X1 U14178 ( .A1(n14092), .A2(n14091), .ZN(n11191) );
  OR2_X1 U14179 ( .A1(n11376), .A2(n11189), .ZN(n11190) );
  NAND2_X1 U14180 ( .A1(n11170), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U14181 ( .A1(n11143), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11157), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11192) );
  NAND2_X1 U14182 ( .A1(n11193), .A2(n11192), .ZN(n14303) );
  INV_X1 U14183 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11194) );
  INV_X1 U14184 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13660) );
  OAI22_X1 U14185 ( .A1(n11699), .A2(n11194), .B1(n11697), .B2(n13660), .ZN(
        n11202) );
  INV_X1 U14186 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11200) );
  INV_X1 U14187 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11196) );
  NAND2_X1 U14188 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n11700), .ZN(
        n11195) );
  OAI21_X1 U14189 ( .B1(n11703), .B2(n11196), .A(n11195), .ZN(n11197) );
  AOI21_X1 U14190 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n11197), .ZN(n11199) );
  NAND2_X1 U14191 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11198) );
  OAI211_X1 U14192 ( .C1(n11200), .C2(n11726), .A(n11199), .B(n11198), .ZN(
        n11201) );
  NOR2_X1 U14193 ( .A1(n11202), .A2(n11201), .ZN(n11212) );
  NAND2_X1 U14194 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11206) );
  NAND2_X1 U14195 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11205) );
  NAND2_X1 U14196 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11204) );
  AOI22_X1 U14197 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11203) );
  NAND2_X1 U14198 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11210) );
  NAND2_X1 U14199 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11209) );
  NAND2_X1 U14200 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11208) );
  NAND2_X1 U14201 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11207) );
  AND4_X1 U14202 ( .A1(n11210), .A2(n11209), .A3(n11208), .A4(n11207), .ZN(
        n11211) );
  NAND2_X1 U14203 ( .A1(n11170), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11214) );
  AOI22_X1 U14204 ( .A1(n11143), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11157), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11213) );
  OAI211_X1 U14205 ( .C1(n13290), .C2(n11376), .A(n11214), .B(n11213), .ZN(
        n11215) );
  OAI22_X1 U14206 ( .A1(n11217), .A2(n11697), .B1(n11699), .B2(n11216), .ZN(
        n11225) );
  NAND2_X1 U14207 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11700), .ZN(
        n11218) );
  OAI21_X1 U14208 ( .B1(n11703), .B2(n11219), .A(n11218), .ZN(n11220) );
  AOI21_X1 U14209 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n11220), .ZN(n11222) );
  NAND2_X1 U14210 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11221) );
  OAI211_X1 U14211 ( .C1(n11726), .C2(n11223), .A(n11222), .B(n11221), .ZN(
        n11224) );
  NOR2_X1 U14212 ( .A1(n11225), .A2(n11224), .ZN(n11233) );
  NAND2_X1 U14213 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11229) );
  NAND2_X1 U14214 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11228) );
  NAND2_X1 U14215 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11227) );
  AOI22_X1 U14216 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11226) );
  AND4_X1 U14217 ( .A1(n11229), .A2(n11228), .A3(n11227), .A4(n11226), .ZN(
        n11232) );
  AOI22_X1 U14218 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10648), .B1(
        n11747), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14219 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n13391), .B1(
        n11760), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11230) );
  NAND4_X1 U14220 ( .A1(n11233), .A2(n11232), .A3(n11231), .A4(n11230), .ZN(
        n13295) );
  AOI22_X1 U14221 ( .A1(n11170), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n10218), 
        .B2(n13295), .ZN(n11235) );
  AOI22_X1 U14222 ( .A1(n11143), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11157), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11234) );
  NAND2_X1 U14223 ( .A1(n11235), .A2(n11234), .ZN(n14468) );
  INV_X1 U14224 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11237) );
  INV_X1 U14225 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11236) );
  OAI22_X1 U14226 ( .A1(n11237), .A2(n11697), .B1(n11699), .B2(n11236), .ZN(
        n11245) );
  INV_X1 U14227 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11243) );
  INV_X1 U14228 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U14229 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11700), .ZN(
        n11238) );
  OAI21_X1 U14230 ( .B1(n11703), .B2(n11239), .A(n11238), .ZN(n11240) );
  AOI21_X1 U14231 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n11240), .ZN(n11242) );
  NAND2_X1 U14232 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11241) );
  OAI211_X1 U14233 ( .C1(n11726), .C2(n11243), .A(n11242), .B(n11241), .ZN(
        n11244) );
  NOR2_X1 U14234 ( .A1(n11245), .A2(n11244), .ZN(n11256) );
  NAND2_X1 U14235 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11249) );
  NAND2_X1 U14236 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11248) );
  NAND2_X1 U14237 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11247) );
  AOI22_X1 U14238 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11246) );
  AND4_X1 U14239 ( .A1(n11249), .A2(n11248), .A3(n11247), .A4(n11246), .ZN(
        n11255) );
  NAND2_X1 U14240 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11253) );
  NAND2_X1 U14241 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11252) );
  NAND2_X1 U14242 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11251) );
  NAND2_X1 U14243 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11250) );
  AND4_X1 U14244 ( .A1(n11253), .A2(n11252), .A3(n11251), .A4(n11250), .ZN(
        n11254) );
  NAND2_X1 U14245 ( .A1(n11143), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n11258) );
  NAND2_X1 U14246 ( .A1(n11157), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11257) );
  OAI211_X1 U14247 ( .C1(n11376), .C2(n13310), .A(n11258), .B(n11257), .ZN(
        n11259) );
  INV_X1 U14248 ( .A(n11259), .ZN(n11261) );
  NAND2_X1 U14249 ( .A1(n11170), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11260) );
  NAND2_X1 U14250 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11265) );
  NAND2_X1 U14251 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11264) );
  NAND2_X1 U14252 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11263) );
  AOI22_X1 U14253 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11262) );
  AND4_X1 U14254 ( .A1(n11265), .A2(n11264), .A3(n11263), .A4(n11262), .ZN(
        n11283) );
  NAND2_X1 U14255 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11700), .ZN(
        n11266) );
  OAI21_X1 U14256 ( .B1(n11703), .B2(n11267), .A(n11266), .ZN(n11268) );
  AOI21_X1 U14257 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n11268), .ZN(n11270) );
  NAND2_X1 U14258 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11269) );
  OAI211_X1 U14259 ( .C1(n11697), .C2(n11271), .A(n11270), .B(n11269), .ZN(
        n11276) );
  OAI22_X1 U14260 ( .A1(n11699), .A2(n11274), .B1(n11273), .B2(n11272), .ZN(
        n11275) );
  NOR2_X1 U14261 ( .A1(n11276), .A2(n11275), .ZN(n11282) );
  NAND2_X1 U14262 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11280) );
  NAND2_X1 U14263 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11279) );
  NAND2_X1 U14264 ( .A1(n11755), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11278) );
  NAND2_X1 U14265 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11277) );
  AND4_X1 U14266 ( .A1(n11280), .A2(n11279), .A3(n11278), .A4(n11277), .ZN(
        n11281) );
  NAND2_X1 U14267 ( .A1(n11170), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14268 ( .A1(n11143), .A2(P2_EAX_REG_11__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n11157), .ZN(n11284) );
  OAI211_X1 U14269 ( .C1(n13478), .C2(n11376), .A(n11285), .B(n11284), .ZN(
        n16473) );
  INV_X1 U14270 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11287) );
  OAI22_X1 U14271 ( .A1(n11287), .A2(n11697), .B1(n11699), .B2(n11286), .ZN(
        n11295) );
  INV_X1 U14272 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11293) );
  INV_X1 U14273 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11289) );
  NAND2_X1 U14274 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11700), .ZN(
        n11288) );
  OAI21_X1 U14275 ( .B1(n11703), .B2(n11289), .A(n11288), .ZN(n11290) );
  AOI21_X1 U14276 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n11290), .ZN(n11292) );
  NAND2_X1 U14277 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11291) );
  OAI211_X1 U14278 ( .C1(n11726), .C2(n11293), .A(n11292), .B(n11291), .ZN(
        n11294) );
  NOR2_X1 U14279 ( .A1(n11295), .A2(n11294), .ZN(n11303) );
  NAND2_X1 U14280 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11299) );
  NAND2_X1 U14281 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11298) );
  NAND2_X1 U14282 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11297) );
  AOI22_X1 U14283 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11296) );
  AND4_X1 U14284 ( .A1(n11299), .A2(n11298), .A3(n11297), .A4(n11296), .ZN(
        n11302) );
  AOI22_X1 U14285 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10648), .B1(
        n11747), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14286 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13391), .B1(
        n11760), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11300) );
  NAND4_X1 U14287 ( .A1(n11303), .A2(n11302), .A3(n11301), .A4(n11300), .ZN(
        n13467) );
  NAND2_X1 U14288 ( .A1(n11143), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n11305) );
  NAND2_X1 U14289 ( .A1(n11157), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11304) );
  OAI211_X1 U14290 ( .C1(n11376), .C2(n10298), .A(n11305), .B(n11304), .ZN(
        n11306) );
  INV_X1 U14291 ( .A(n11306), .ZN(n11308) );
  NAND2_X1 U14292 ( .A1(n11170), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14293 ( .A1(n11170), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n11157), .ZN(n11328) );
  OAI22_X1 U14294 ( .A1(n11699), .A2(n11310), .B1(n11697), .B2(n11309), .ZN(
        n11318) );
  NAND2_X1 U14295 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n11700), .ZN(
        n11311) );
  OAI21_X1 U14296 ( .B1(n11703), .B2(n11312), .A(n11311), .ZN(n11313) );
  AOI21_X1 U14297 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n11313), .ZN(n11315) );
  NAND2_X1 U14298 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11314) );
  OAI211_X1 U14299 ( .C1(n11316), .C2(n11726), .A(n11315), .B(n11314), .ZN(
        n11317) );
  NOR2_X1 U14300 ( .A1(n11318), .A2(n11317), .ZN(n11326) );
  NAND2_X1 U14301 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11322) );
  NAND2_X1 U14302 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11321) );
  NAND2_X1 U14303 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11320) );
  AOI22_X1 U14304 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11319) );
  AND4_X1 U14305 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(
        n11325) );
  AOI22_X1 U14306 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11747), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14307 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11323) );
  NAND4_X1 U14308 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n13508) );
  AOI22_X1 U14309 ( .A1(n10218), .A2(n13508), .B1(n11143), .B2(
        P2_EAX_REG_13__SCAN_IN), .ZN(n11327) );
  NAND2_X1 U14310 ( .A1(n11328), .A2(n11327), .ZN(n14491) );
  OAI22_X1 U14311 ( .A1(n11699), .A2(n11330), .B1(n11697), .B2(n11329), .ZN(
        n11338) );
  NAND2_X1 U14312 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11700), .ZN(
        n11331) );
  OAI21_X1 U14313 ( .B1(n11703), .B2(n11332), .A(n11331), .ZN(n11333) );
  AOI21_X1 U14314 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n11333), .ZN(n11335) );
  NAND2_X1 U14315 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11334) );
  OAI211_X1 U14316 ( .C1(n11336), .C2(n11726), .A(n11335), .B(n11334), .ZN(
        n11337) );
  NOR2_X1 U14317 ( .A1(n11338), .A2(n11337), .ZN(n11349) );
  NAND2_X1 U14318 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U14319 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11341) );
  NAND2_X1 U14320 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11340) );
  AOI22_X1 U14321 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11339) );
  AND4_X1 U14322 ( .A1(n11342), .A2(n11341), .A3(n11340), .A4(n11339), .ZN(
        n11348) );
  NAND2_X1 U14323 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11346) );
  NAND2_X1 U14324 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11345) );
  NAND2_X1 U14325 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11344) );
  NAND2_X1 U14326 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11343) );
  AND4_X1 U14327 ( .A1(n11346), .A2(n11345), .A3(n11344), .A4(n11343), .ZN(
        n11347) );
  NAND2_X1 U14328 ( .A1(n11170), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14329 ( .A1(n11143), .A2(P2_EAX_REG_14__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n11157), .ZN(n11350) );
  OAI211_X1 U14330 ( .C1(n13661), .C2(n11376), .A(n11351), .B(n11350), .ZN(
        n11352) );
  INV_X1 U14331 ( .A(n11352), .ZN(n17050) );
  INV_X1 U14332 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11354) );
  INV_X1 U14333 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11353) );
  OAI22_X1 U14334 ( .A1(n11699), .A2(n11354), .B1(n11697), .B2(n11353), .ZN(
        n11362) );
  INV_X1 U14335 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11360) );
  INV_X1 U14336 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11356) );
  NAND2_X1 U14337 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11700), .ZN(
        n11355) );
  OAI21_X1 U14338 ( .B1(n11703), .B2(n11356), .A(n11355), .ZN(n11357) );
  AOI21_X1 U14339 ( .B1(n11742), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n11357), .ZN(n11359) );
  NAND2_X1 U14340 ( .A1(n11729), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11358) );
  OAI211_X1 U14341 ( .C1(n11360), .C2(n11726), .A(n11359), .B(n11358), .ZN(
        n11361) );
  NOR2_X1 U14342 ( .A1(n11362), .A2(n11361), .ZN(n11373) );
  NAND2_X1 U14343 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11366) );
  NAND2_X1 U14344 ( .A1(n11747), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11365) );
  NAND2_X1 U14345 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11364) );
  AOI22_X1 U14346 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11363) );
  AND4_X1 U14347 ( .A1(n11366), .A2(n11365), .A3(n11364), .A4(n11363), .ZN(
        n11372) );
  NAND2_X1 U14348 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11370) );
  NAND2_X1 U14349 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11369) );
  NAND2_X1 U14350 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11368) );
  NAND2_X1 U14351 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11367) );
  AND4_X1 U14352 ( .A1(n11370), .A2(n11369), .A3(n11368), .A4(n11367), .ZN(
        n11371) );
  NAND2_X1 U14353 ( .A1(n11170), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14354 ( .A1(n11143), .A2(P2_EAX_REG_15__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n11157), .ZN(n11374) );
  OAI211_X1 U14355 ( .C1(n14175), .C2(n11376), .A(n11375), .B(n11374), .ZN(
        n14320) );
  NAND2_X1 U14356 ( .A1(n11170), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14357 ( .A1(n11143), .A2(P2_EAX_REG_16__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n11157), .ZN(n11377) );
  NAND2_X1 U14358 ( .A1(n11378), .A2(n11377), .ZN(n14179) );
  NAND2_X1 U14359 ( .A1(n11170), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14360 ( .A1(n11143), .A2(P2_EAX_REG_17__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n11157), .ZN(n11379) );
  AND2_X1 U14361 ( .A1(n11380), .A2(n11379), .ZN(n14331) );
  NAND2_X1 U14362 ( .A1(n11170), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14363 ( .A1(n11143), .A2(P2_EAX_REG_18__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n11157), .ZN(n11381) );
  INV_X1 U14364 ( .A(n11170), .ZN(n11400) );
  INV_X1 U14365 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20425) );
  AOI22_X1 U14366 ( .A1(n11143), .A2(P2_EAX_REG_19__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n11157), .ZN(n11383) );
  OAI21_X1 U14367 ( .B1(n11400), .B2(n20425), .A(n11383), .ZN(n15995) );
  NAND2_X1 U14368 ( .A1(n11170), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14369 ( .A1(n11143), .A2(P2_EAX_REG_20__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n11157), .ZN(n11384) );
  AND2_X1 U14370 ( .A1(n11385), .A2(n11384), .ZN(n15981) );
  NAND2_X1 U14371 ( .A1(n11170), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14372 ( .A1(n11143), .A2(P2_EAX_REG_21__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n11157), .ZN(n11386) );
  AND2_X1 U14373 ( .A1(n11387), .A2(n11386), .ZN(n15967) );
  INV_X1 U14374 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16220) );
  AOI22_X1 U14375 ( .A1(n11143), .A2(P2_EAX_REG_22__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n11157), .ZN(n11388) );
  OAI21_X1 U14376 ( .B1(n11400), .B2(n16220), .A(n11388), .ZN(n16117) );
  INV_X1 U14377 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20432) );
  AOI22_X1 U14378 ( .A1(n11143), .A2(P2_EAX_REG_23__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n11157), .ZN(n11389) );
  OAI21_X1 U14379 ( .B1(n11400), .B2(n20432), .A(n11389), .ZN(n16109) );
  NAND2_X1 U14380 ( .A1(n11170), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14381 ( .A1(n11143), .A2(P2_EAX_REG_24__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n11157), .ZN(n11390) );
  AND2_X1 U14382 ( .A1(n11391), .A2(n11390), .ZN(n15952) );
  NAND2_X1 U14383 ( .A1(n11170), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14384 ( .A1(n11143), .A2(P2_EAX_REG_25__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n11157), .ZN(n11392) );
  AND2_X1 U14385 ( .A1(n11393), .A2(n11392), .ZN(n16102) );
  INV_X1 U14386 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20436) );
  AOI22_X1 U14387 ( .A1(n11143), .A2(P2_EAX_REG_26__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n11157), .ZN(n11394) );
  OAI21_X1 U14388 ( .B1(n11400), .B2(n20436), .A(n11394), .ZN(n15938) );
  NAND2_X1 U14389 ( .A1(n11170), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14390 ( .A1(n11143), .A2(P2_EAX_REG_27__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n11157), .ZN(n11395) );
  AND2_X1 U14391 ( .A1(n11396), .A2(n11395), .ZN(n16090) );
  NAND2_X1 U14392 ( .A1(n11170), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14393 ( .A1(n11143), .A2(P2_EAX_REG_28__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n11157), .ZN(n11397) );
  AND2_X1 U14394 ( .A1(n11398), .A2(n11397), .ZN(n11508) );
  INV_X1 U14395 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20442) );
  AOI22_X1 U14396 ( .A1(n11143), .A2(P2_EAX_REG_29__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n11157), .ZN(n11399) );
  OAI21_X1 U14397 ( .B1(n11400), .B2(n20442), .A(n11399), .ZN(n12402) );
  AOI21_X1 U14398 ( .B1(n11402), .B2(n11401), .A(n11554), .ZN(n12015) );
  INV_X1 U14399 ( .A(n11403), .ZN(n11948) );
  AND2_X1 U14400 ( .A1(n11948), .A2(n14265), .ZN(n11404) );
  OR2_X1 U14401 ( .A1(n11404), .A2(n13423), .ZN(n11405) );
  INV_X1 U14402 ( .A(n20133), .ZN(n20458) );
  AND2_X2 U14403 ( .A1(n20458), .A2(n12616), .ZN(n19825) );
  INV_X1 U14404 ( .A(n19825), .ZN(n19856) );
  INV_X1 U14405 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n11406) );
  NOR2_X1 U14406 ( .A1(n19856), .A2(n11406), .ZN(n11493) );
  AOI21_X1 U14407 ( .B1(n12015), .B2(n19854), .A(n11493), .ZN(n11442) );
  AND2_X1 U14408 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16323) );
  NAND2_X1 U14409 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11431) );
  NAND2_X1 U14410 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16427) );
  INV_X1 U14411 ( .A(n16427), .ZN(n11407) );
  NAND2_X1 U14412 ( .A1(n11407), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16416) );
  NAND2_X1 U14413 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11432) );
  INV_X1 U14414 ( .A(n11432), .ZN(n11427) );
  INV_X1 U14415 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13355) );
  NOR3_X1 U14416 ( .A1(n13355), .A2(n21051), .A3(n13675), .ZN(n14087) );
  INV_X1 U14417 ( .A(n14087), .ZN(n14088) );
  NOR2_X1 U14418 ( .A1(n11408), .A2(n14088), .ZN(n14307) );
  NAND2_X1 U14419 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n14307), .ZN(
        n14444) );
  NOR2_X1 U14420 ( .A1(n10849), .A2(n14444), .ZN(n11433) );
  NAND2_X1 U14421 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19852) );
  NAND2_X1 U14422 ( .A1(n11482), .A2(n13427), .ZN(n16431) );
  INV_X1 U14423 ( .A(n19852), .ZN(n19862) );
  NAND2_X1 U14424 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19862), .ZN(
        n11411) );
  AOI22_X1 U14425 ( .A1(n19876), .A2(n19852), .B1(n16431), .B2(n11411), .ZN(
        n13364) );
  INV_X1 U14426 ( .A(n11412), .ZN(n11422) );
  NAND2_X1 U14427 ( .A1(n11414), .A2(n14265), .ZN(n13404) );
  NAND2_X1 U14428 ( .A1(n13404), .A2(n11415), .ZN(n11417) );
  NAND2_X1 U14429 ( .A1(n11417), .A2(n11416), .ZN(n11420) );
  INV_X1 U14430 ( .A(n11947), .ZN(n12606) );
  NAND2_X1 U14431 ( .A1(n10483), .A2(n10474), .ZN(n11418) );
  AOI22_X1 U14432 ( .A1(n12606), .A2(n11418), .B1(n13429), .B2(n19880), .ZN(
        n11419) );
  NAND3_X1 U14433 ( .A1(n11413), .A2(n11420), .A3(n11419), .ZN(n11421) );
  AOI21_X1 U14434 ( .B1(n11422), .B2(n10466), .A(n11421), .ZN(n13410) );
  INV_X1 U14435 ( .A(n10484), .ZN(n11425) );
  AND2_X1 U14436 ( .A1(n10466), .A2(n11423), .ZN(n11424) );
  NAND2_X1 U14437 ( .A1(n11425), .A2(n11424), .ZN(n13382) );
  NAND2_X1 U14438 ( .A1(n13410), .A2(n13382), .ZN(n11426) );
  NAND2_X1 U14439 ( .A1(n13364), .A2(n17054), .ZN(n14443) );
  NAND2_X1 U14440 ( .A1(n11433), .A2(n14306), .ZN(n16509) );
  INV_X1 U14441 ( .A(n16509), .ZN(n16415) );
  NAND2_X1 U14442 ( .A1(n11427), .A2(n16415), .ZN(n11428) );
  NOR2_X1 U14443 ( .A1(n16416), .A2(n11428), .ZN(n11429) );
  NOR2_X1 U14444 ( .A1(n16492), .A2(n16478), .ZN(n17058) );
  AND3_X1 U14445 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n17058), .ZN(n17048) );
  NAND2_X1 U14446 ( .A1(n17048), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16434) );
  NAND2_X1 U14447 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16395) );
  INV_X1 U14448 ( .A(n16395), .ZN(n11430) );
  NAND2_X1 U14449 ( .A1(n16374), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16359) );
  NOR2_X1 U14450 ( .A1(n11431), .A2(n16359), .ZN(n16348) );
  NAND3_X1 U14451 ( .A1(n16323), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16335), .ZN(n12403) );
  NAND2_X1 U14452 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11557) );
  NOR2_X1 U14453 ( .A1(n12403), .A2(n11557), .ZN(n11440) );
  NOR3_X1 U14454 ( .A1(n16434), .A2(n16416), .A3(n11432), .ZN(n11437) );
  OR2_X1 U14455 ( .A1(n16432), .A2(n11433), .ZN(n11436) );
  INV_X1 U14456 ( .A(n19825), .ZN(n19838) );
  NOR2_X1 U14457 ( .A1(n11482), .A2(n19825), .ZN(n19851) );
  AOI21_X1 U14458 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19862), .A(
        n16436), .ZN(n11435) );
  NAND2_X1 U14459 ( .A1(n19876), .A2(n19852), .ZN(n11434) );
  NOR2_X1 U14460 ( .A1(n16431), .A2(n11434), .ZN(n19861) );
  NOR3_X1 U14461 ( .A1(n19851), .A2(n11435), .A3(n19861), .ZN(n14086) );
  AND2_X1 U14462 ( .A1(n11436), .A2(n14086), .ZN(n16508) );
  OAI21_X1 U14463 ( .B1(n16432), .B2(n11437), .A(n16508), .ZN(n16410) );
  INV_X1 U14464 ( .A(n16410), .ZN(n16421) );
  NAND2_X1 U14465 ( .A1(n16421), .A2(n16432), .ZN(n11560) );
  INV_X1 U14466 ( .A(n11560), .ZN(n11439) );
  INV_X1 U14467 ( .A(n11557), .ZN(n12404) );
  NAND3_X1 U14468 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16360) );
  INV_X1 U14469 ( .A(n16360), .ZN(n11438) );
  AOI21_X1 U14470 ( .B1(n16395), .B2(n17054), .A(n16410), .ZN(n16376) );
  OAI211_X1 U14471 ( .C1(n16432), .C2(n11438), .A(n16376), .B(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16347) );
  NAND2_X1 U14472 ( .A1(n16347), .A2(n11560), .ZN(n16340) );
  OAI21_X1 U14473 ( .B1(n16323), .B2(n11439), .A(n16340), .ZN(n16317) );
  AOI21_X1 U14474 ( .B1(n16312), .B2(n11560), .A(n16317), .ZN(n12400) );
  OAI211_X1 U14475 ( .C1(n11439), .C2(n12404), .A(n12400), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11561) );
  OAI21_X1 U14476 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n11440), .A(
        n11561), .ZN(n11441) );
  OAI211_X1 U14477 ( .C1(n9693), .C2(n19870), .A(n11442), .B(n11441), .ZN(
        n11443) );
  XOR2_X1 U14478 ( .A(n11445), .B(n11444), .Z(n19836) );
  NAND2_X1 U14479 ( .A1(n12844), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12843) );
  XNOR2_X1 U14480 ( .A(n11447), .B(n11446), .ZN(n11448) );
  NOR2_X1 U14481 ( .A1(n12843), .A2(n11448), .ZN(n11449) );
  INV_X1 U14482 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21108) );
  XNOR2_X1 U14483 ( .A(n12843), .B(n11448), .ZN(n12733) );
  NOR2_X1 U14484 ( .A1(n21108), .A2(n12733), .ZN(n12732) );
  NOR2_X1 U14485 ( .A1(n11449), .A2(n12732), .ZN(n11450) );
  XOR2_X1 U14486 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11450), .Z(
        n19835) );
  NOR2_X1 U14487 ( .A1(n19836), .A2(n19835), .ZN(n19834) );
  NOR2_X1 U14488 ( .A1(n11450), .A2(n19876), .ZN(n11451) );
  XNOR2_X1 U14489 ( .A(n11452), .B(n13355), .ZN(n13360) );
  NAND2_X1 U14490 ( .A1(n11452), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11453) );
  INV_X1 U14491 ( .A(n11457), .ZN(n11458) );
  OAI21_X1 U14492 ( .B1(n13670), .B2(n13669), .A(n11459), .ZN(n11467) );
  INV_X1 U14493 ( .A(n11466), .ZN(n11465) );
  INV_X1 U14494 ( .A(n11470), .ZN(n11460) );
  NAND2_X1 U14495 ( .A1(n13671), .A2(n11460), .ZN(n11464) );
  INV_X1 U14496 ( .A(n13669), .ZN(n11461) );
  NAND3_X1 U14497 ( .A1(n11462), .A2(n11461), .A3(n11465), .ZN(n11463) );
  NAND2_X1 U14498 ( .A1(n11467), .A2(n11466), .ZN(n11468) );
  INV_X1 U14499 ( .A(n11473), .ZN(n11474) );
  NAND2_X1 U14500 ( .A1(n11472), .A2(n11474), .ZN(n11475) );
  INV_X1 U14501 ( .A(n11478), .ZN(n11479) );
  NAND3_X1 U14502 ( .A1(n11479), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n10880), .ZN(n11480) );
  INV_X1 U14503 ( .A(n16434), .ZN(n11481) );
  INV_X1 U14504 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16375) );
  NAND3_X1 U14505 ( .A1(n11485), .A2(n11484), .A3(n11483), .ZN(P2_U3016) );
  AND2_X1 U14506 ( .A1(n13429), .A2(n13124), .ZN(n12016) );
  NAND2_X1 U14507 ( .A1(n11486), .A2(n12016), .ZN(n19563) );
  NAND2_X1 U14508 ( .A1(n11487), .A2(n19828), .ZN(n11498) );
  NAND2_X1 U14509 ( .A1(n11007), .A2(n20101), .ZN(n20455) );
  NAND2_X1 U14510 ( .A1(n20133), .A2(n20455), .ZN(n20482) );
  NAND2_X1 U14511 ( .A1(n20482), .A2(n17100), .ZN(n11489) );
  AND2_X1 U14512 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20472) );
  INV_X1 U14513 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17006) );
  INV_X1 U14514 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16992) );
  INV_X1 U14515 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16305) );
  NAND2_X1 U14516 ( .A1(n11994), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12007) );
  INV_X1 U14517 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16285) );
  NAND2_X1 U14518 ( .A1(n11992), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11990) );
  INV_X1 U14519 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12008) );
  INV_X1 U14520 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16211) );
  INV_X1 U14521 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16199) );
  INV_X1 U14522 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16188) );
  INV_X1 U14523 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16173) );
  INV_X1 U14524 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16166) );
  XNOR2_X1 U14525 ( .A(n11542), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12012) );
  NAND2_X1 U14526 ( .A1(n17100), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11574) );
  INV_X1 U14527 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21150) );
  NAND2_X1 U14528 ( .A1(n21150), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11491) );
  NAND2_X1 U14529 ( .A1(n11574), .A2(n11491), .ZN(n15261) );
  NOR2_X1 U14530 ( .A1(n12012), .A2(n19840), .ZN(n11492) );
  AOI211_X1 U14531 ( .C1(n19837), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n11493), .B(n11492), .ZN(n11494) );
  OAI21_X1 U14532 ( .B1(n9693), .B2(n16307), .A(n11494), .ZN(n11495) );
  INV_X1 U14533 ( .A(n11495), .ZN(n11496) );
  NAND3_X1 U14534 ( .A1(n11498), .A2(n11497), .A3(n11496), .ZN(P2_U2984) );
  XNOR2_X2 U14535 ( .A(n11502), .B(n11501), .ZN(n16171) );
  INV_X1 U14536 ( .A(n11502), .ZN(n11504) );
  XNOR2_X1 U14537 ( .A(n11505), .B(n12405), .ZN(n11506) );
  NAND2_X1 U14538 ( .A1(n16163), .A2(n19866), .ZN(n11517) );
  OAI21_X1 U14539 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n9719), .ZN(n16170) );
  AOI21_X1 U14540 ( .B1(n11507), .B2(n16035), .A(n12389), .ZN(n16907) );
  AND2_X1 U14541 ( .A1(n9772), .A2(n11508), .ZN(n11509) );
  OR2_X1 U14542 ( .A1(n12401), .A2(n11509), .ZN(n16905) );
  NAND2_X1 U14543 ( .A1(n19825), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n16165) );
  INV_X1 U14544 ( .A(n12403), .ZN(n11510) );
  NAND2_X1 U14545 ( .A1(n11510), .A2(n12405), .ZN(n11511) );
  OAI211_X1 U14546 ( .C1(n16905), .C2(n17070), .A(n16165), .B(n11511), .ZN(
        n11513) );
  NOR2_X1 U14547 ( .A1(n12400), .A2(n12405), .ZN(n11512) );
  AOI211_X1 U14548 ( .C1(n16907), .C2(n17086), .A(n11513), .B(n11512), .ZN(
        n11514) );
  NAND2_X1 U14549 ( .A1(n11517), .A2(n11516), .ZN(P2_U3018) );
  INV_X1 U14550 ( .A(n11518), .ZN(n11520) );
  MUX2_X1 U14551 ( .A(n11525), .B(n11524), .S(n11966), .Z(n16885) );
  NAND2_X1 U14552 ( .A1(n16885), .A2(n10880), .ZN(n11526) );
  XOR2_X1 U14553 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11526), .Z(
        n11527) );
  NAND2_X1 U14554 ( .A1(n11528), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11530) );
  INV_X1 U14555 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11529) );
  NAND2_X1 U14556 ( .A1(n9765), .A2(n11531), .ZN(n11549) );
  AOI22_X1 U14557 ( .A1(n11534), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11539) );
  NAND2_X1 U14558 ( .A1(n11535), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11538) );
  NAND2_X1 U14559 ( .A1(n11536), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11537) );
  AND3_X1 U14560 ( .A1(n11539), .A2(n11538), .A3(n11537), .ZN(n11540) );
  XNOR2_X2 U14561 ( .A(n11541), .B(n11540), .ZN(n16953) );
  NOR2_X1 U14562 ( .A1(n16953), .A2(n16307), .ZN(n11547) );
  NAND2_X1 U14563 ( .A1(n11542), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11544) );
  NAND2_X1 U14564 ( .A1(n19825), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11555) );
  NAND2_X1 U14565 ( .A1(n19837), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11545) );
  OAI211_X1 U14566 ( .C1(n11977), .C2(n19840), .A(n11555), .B(n11545), .ZN(
        n11546) );
  NAND2_X1 U14567 ( .A1(n11550), .A2(n19866), .ZN(n11567) );
  NAND2_X1 U14568 ( .A1(n9765), .A2(n11551), .ZN(n11566) );
  AOI222_X1 U14569 ( .A1(n11170), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11143), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11157), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11553) );
  XNOR2_X1 U14570 ( .A(n11554), .B(n11553), .ZN(n19718) );
  INV_X1 U14571 ( .A(n11555), .ZN(n11559) );
  NOR4_X1 U14572 ( .A1(n12403), .A2(n11557), .A3(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A4(n11556), .ZN(n11558) );
  NAND3_X1 U14573 ( .A1(n11561), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n11560), .ZN(n11562) );
  OAI211_X1 U14574 ( .C1(n16953), .C2(n19870), .A(n11563), .B(n11562), .ZN(
        n11564) );
  NAND3_X1 U14575 ( .A1(n11567), .A2(n11566), .A3(n11565), .ZN(P2_U3015) );
  NAND2_X1 U14576 ( .A1(n19896), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U14577 ( .A1(n11593), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11570) );
  OAI22_X1 U14578 ( .A1(n20481), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B1(
        n20492), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19942) );
  INV_X1 U14579 ( .A(n19942), .ZN(n11569) );
  OR2_X1 U14580 ( .A1(n20133), .A2(n11569), .ZN(n20165) );
  NAND2_X1 U14581 ( .A1(n11570), .A2(n20165), .ZN(n11571) );
  NOR2_X1 U14582 ( .A1(n20133), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11572) );
  AOI21_X1 U14583 ( .B1(n11593), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11572), .ZN(n11573) );
  NAND2_X1 U14584 ( .A1(n11836), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11575) );
  NAND2_X1 U14585 ( .A1(n12969), .A2(n11575), .ZN(n11576) );
  NAND2_X1 U14586 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20203) );
  NAND2_X1 U14587 ( .A1(n20203), .A2(n20470), .ZN(n11578) );
  NOR2_X1 U14588 ( .A1(n20470), .A2(n20481), .ZN(n20311) );
  NAND2_X1 U14589 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20311), .ZN(
        n14257) );
  NAND2_X1 U14590 ( .A1(n11578), .A2(n14257), .ZN(n13336) );
  NOR2_X1 U14591 ( .A1(n13336), .A2(n20133), .ZN(n11579) );
  AOI21_X1 U14592 ( .B1(n11593), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11579), .ZN(n11584) );
  NAND2_X1 U14593 ( .A1(n11836), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11589) );
  NAND2_X1 U14594 ( .A1(n11584), .A2(n11589), .ZN(n11581) );
  INV_X1 U14595 ( .A(n11581), .ZN(n11580) );
  NAND2_X1 U14596 ( .A1(n11582), .A2(n11580), .ZN(n11588) );
  NAND2_X1 U14597 ( .A1(n11577), .A2(n11583), .ZN(n11587) );
  INV_X1 U14598 ( .A(n11584), .ZN(n11590) );
  OAI21_X1 U14599 ( .B1(n11590), .B2(n11596), .A(n11589), .ZN(n11585) );
  OAI21_X1 U14600 ( .B1(n11589), .B2(n11590), .A(n11585), .ZN(n11586) );
  INV_X1 U14601 ( .A(n11589), .ZN(n11591) );
  NAND2_X1 U14602 ( .A1(n11591), .A2(n11590), .ZN(n11592) );
  NAND2_X1 U14603 ( .A1(n11836), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13217) );
  NAND2_X1 U14604 ( .A1(n11593), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11598) );
  NAND2_X1 U14605 ( .A1(n13217), .A2(n11598), .ZN(n11594) );
  NAND2_X1 U14606 ( .A1(n13216), .A2(n11594), .ZN(n11603) );
  NAND2_X1 U14607 ( .A1(n20463), .A2(n20311), .ZN(n20071) );
  NOR2_X1 U14608 ( .A1(n20492), .A2(n20071), .ZN(n20091) );
  AOI21_X1 U14609 ( .B1(n14257), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n20091), .ZN(n11597) );
  OR2_X1 U14610 ( .A1(n20133), .A2(n11597), .ZN(n13344) );
  AND2_X1 U14611 ( .A1(n11598), .A2(n13344), .ZN(n11599) );
  INV_X1 U14612 ( .A(n13217), .ZN(n11601) );
  NOR2_X1 U14613 ( .A1(n19668), .A2(n11865), .ZN(n11604) );
  NAND2_X1 U14614 ( .A1(n13465), .A2(n13508), .ZN(n13507) );
  INV_X1 U14615 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11608) );
  OAI22_X1 U14616 ( .A1(n11699), .A2(n11608), .B1(n11697), .B2(n11607), .ZN(
        n11616) );
  INV_X1 U14617 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11614) );
  INV_X1 U14618 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14619 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n11700), .ZN(
        n11609) );
  OAI21_X1 U14620 ( .B1(n11703), .B2(n11610), .A(n11609), .ZN(n11611) );
  AOI21_X1 U14621 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n11611), .ZN(n11613) );
  NAND2_X1 U14622 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11612) );
  OAI211_X1 U14623 ( .C1(n11614), .C2(n11726), .A(n11613), .B(n11612), .ZN(
        n11615) );
  NOR2_X1 U14624 ( .A1(n11616), .A2(n11615), .ZN(n11624) );
  NAND2_X1 U14625 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11620) );
  NAND2_X1 U14626 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11619) );
  NAND2_X1 U14627 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11618) );
  AOI22_X1 U14628 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11617) );
  AND4_X1 U14629 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11623) );
  AOI22_X1 U14630 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11747), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14631 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11621) );
  NAND4_X1 U14632 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n14082) );
  OAI22_X1 U14633 ( .A1(n11626), .A2(n11699), .B1(n11697), .B2(n11625), .ZN(
        n11634) );
  NAND2_X1 U14634 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11700), .ZN(
        n11627) );
  OAI21_X1 U14635 ( .B1(n11703), .B2(n11628), .A(n11627), .ZN(n11629) );
  AOI21_X1 U14636 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n11629), .ZN(n11631) );
  NAND2_X1 U14637 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11630) );
  OAI211_X1 U14638 ( .C1(n11726), .C2(n11632), .A(n11631), .B(n11630), .ZN(
        n11633) );
  NOR2_X1 U14639 ( .A1(n11634), .A2(n11633), .ZN(n11642) );
  NAND2_X1 U14640 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11638) );
  NAND2_X1 U14641 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11637) );
  NAND2_X1 U14642 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11636) );
  AOI22_X1 U14643 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11635) );
  AND4_X1 U14644 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11641) );
  AOI22_X1 U14645 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11747), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14646 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11760), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11639) );
  AND4_X1 U14647 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n14330) );
  INV_X1 U14648 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11644) );
  INV_X1 U14649 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11643) );
  OAI22_X1 U14650 ( .A1(n11644), .A2(n11699), .B1(n11697), .B2(n11643), .ZN(
        n11652) );
  INV_X1 U14651 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11650) );
  INV_X1 U14652 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11646) );
  NAND2_X1 U14653 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11700), .ZN(
        n11645) );
  OAI21_X1 U14654 ( .B1(n11703), .B2(n11646), .A(n11645), .ZN(n11647) );
  AOI21_X1 U14655 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n11647), .ZN(n11649) );
  NAND2_X1 U14656 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11648) );
  OAI211_X1 U14657 ( .C1(n11726), .C2(n11650), .A(n11649), .B(n11648), .ZN(
        n11651) );
  NOR2_X1 U14658 ( .A1(n11652), .A2(n11651), .ZN(n11660) );
  INV_X1 U14659 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19884) );
  NAND2_X1 U14660 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11656) );
  NAND2_X1 U14661 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11655) );
  NAND2_X1 U14662 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11654) );
  AOI22_X1 U14663 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11653) );
  AND4_X1 U14664 ( .A1(n11656), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(
        n11659) );
  AOI22_X1 U14665 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11747), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14666 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n11760), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11657) );
  NAND4_X1 U14667 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n16072) );
  OAI22_X1 U14668 ( .A1(n11662), .A2(n11699), .B1(n11697), .B2(n11661), .ZN(
        n11670) );
  NAND2_X1 U14669 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11700), .ZN(
        n11663) );
  OAI21_X1 U14670 ( .B1(n11703), .B2(n11664), .A(n11663), .ZN(n11665) );
  AOI21_X1 U14671 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n11665), .ZN(n11667) );
  NAND2_X1 U14672 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11666) );
  OAI211_X1 U14673 ( .C1(n11726), .C2(n11668), .A(n11667), .B(n11666), .ZN(
        n11669) );
  NOR2_X1 U14674 ( .A1(n11670), .A2(n11669), .ZN(n11678) );
  NAND2_X1 U14675 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11674) );
  NAND2_X1 U14676 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11673) );
  NAND2_X1 U14677 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11672) );
  AOI22_X1 U14678 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11671) );
  AND4_X1 U14679 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n11677) );
  AOI22_X1 U14680 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11747), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14681 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n11760), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11675) );
  AND4_X1 U14682 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(
        n16145) );
  NOR2_X2 U14683 ( .A1(n16071), .A2(n16145), .ZN(n16067) );
  OAI22_X1 U14684 ( .A1(n11680), .A2(n11699), .B1(n11697), .B2(n11679), .ZN(
        n11688) );
  NAND2_X1 U14685 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11700), .ZN(
        n11681) );
  OAI21_X1 U14686 ( .B1(n11703), .B2(n11682), .A(n11681), .ZN(n11683) );
  AOI21_X1 U14687 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n11683), .ZN(n11685) );
  NAND2_X1 U14688 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11684) );
  OAI211_X1 U14689 ( .C1(n11726), .C2(n11686), .A(n11685), .B(n11684), .ZN(
        n11687) );
  NOR2_X1 U14690 ( .A1(n11688), .A2(n11687), .ZN(n11696) );
  NAND2_X1 U14691 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11692) );
  NAND2_X1 U14692 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11691) );
  NAND2_X1 U14693 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11690) );
  AOI22_X1 U14694 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11742), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11689) );
  AND4_X1 U14695 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11695) );
  AOI22_X1 U14696 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11747), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14697 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11760), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U14698 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n16069) );
  NAND2_X1 U14699 ( .A1(n16067), .A2(n16069), .ZN(n16068) );
  OAI22_X1 U14700 ( .A1(n11699), .A2(n11698), .B1(n11697), .B2(n11901), .ZN(
        n11709) );
  NAND2_X1 U14701 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n11700), .ZN(
        n11701) );
  OAI21_X1 U14702 ( .B1(n11703), .B2(n11702), .A(n11701), .ZN(n11704) );
  AOI21_X1 U14703 ( .B1(n11718), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n11704), .ZN(n11706) );
  NAND2_X1 U14704 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11705) );
  OAI211_X1 U14705 ( .C1(n11707), .C2(n11726), .A(n11706), .B(n11705), .ZN(
        n11708) );
  NOR2_X1 U14706 ( .A1(n11709), .A2(n11708), .ZN(n11717) );
  NAND2_X1 U14707 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11713) );
  NAND2_X1 U14708 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11712) );
  NAND2_X1 U14709 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11711) );
  AOI22_X1 U14710 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11710) );
  AND4_X1 U14711 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n11716) );
  AOI22_X1 U14712 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11747), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14713 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11714) );
  AND4_X1 U14714 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n16127) );
  NOR2_X2 U14715 ( .A1(n16068), .A2(n16127), .ZN(n16060) );
  AOI22_X1 U14716 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11754), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11724) );
  INV_X1 U14717 ( .A(n11718), .ZN(n11751) );
  AOI22_X1 U14718 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11719) );
  OAI21_X1 U14719 ( .B1(n11751), .B2(n11720), .A(n11719), .ZN(n11721) );
  AOI21_X1 U14720 ( .B1(n11722), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n11721), .ZN(n11723) );
  OAI211_X1 U14721 ( .C1(n11726), .C2(n11725), .A(n11724), .B(n11723), .ZN(
        n11739) );
  AOI22_X1 U14722 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11747), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14723 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11727) );
  NAND2_X1 U14724 ( .A1(n11728), .A2(n11727), .ZN(n11738) );
  INV_X1 U14725 ( .A(n11740), .ZN(n11732) );
  NAND2_X1 U14726 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11731) );
  NAND2_X1 U14727 ( .A1(n11729), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11730) );
  OAI211_X1 U14728 ( .C1(n11732), .C2(n13317), .A(n11731), .B(n11730), .ZN(
        n11737) );
  INV_X1 U14729 ( .A(n10643), .ZN(n11734) );
  OAI22_X1 U14730 ( .A1(n11735), .A2(n11917), .B1(n11734), .B2(n11733), .ZN(
        n11736) );
  NAND2_X1 U14731 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11746) );
  NAND2_X1 U14732 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14733 ( .A1(n10643), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11744) );
  AOI22_X1 U14734 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11729), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11743) );
  AND4_X1 U14735 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(
        n11764) );
  AOI22_X1 U14736 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11747), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11763) );
  INV_X1 U14737 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11930) );
  NAND2_X1 U14738 ( .A1(n11722), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11750) );
  AOI22_X1 U14739 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11749) );
  OAI211_X1 U14740 ( .C1(n11751), .C2(n11930), .A(n11750), .B(n11749), .ZN(
        n11752) );
  INV_X1 U14741 ( .A(n11752), .ZN(n11759) );
  NAND2_X1 U14742 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U14743 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11757) );
  NAND2_X1 U14744 ( .A1(n11755), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11756) );
  AND4_X1 U14745 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11762) );
  AOI22_X1 U14746 ( .A1(n11760), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11761) );
  NAND4_X1 U14747 ( .A1(n11764), .A2(n11763), .A3(n11762), .A4(n11761), .ZN(
        n11787) );
  INV_X1 U14748 ( .A(n10387), .ZN(n11931) );
  AOI22_X1 U14749 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14750 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14751 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11774) );
  INV_X1 U14752 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13234) );
  INV_X1 U14753 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11767) );
  OR2_X1 U14754 ( .A1(n11911), .A2(n11767), .ZN(n11771) );
  INV_X1 U14755 ( .A(n11768), .ZN(n11770) );
  NAND2_X1 U14756 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11769) );
  NAND2_X1 U14757 ( .A1(n11770), .A2(n11769), .ZN(n11935) );
  OAI211_X1 U14758 ( .C1(n11876), .C2(n13234), .A(n11771), .B(n11935), .ZN(
        n11772) );
  INV_X1 U14759 ( .A(n11772), .ZN(n11773) );
  NAND4_X1 U14760 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(
        n11786) );
  AOI22_X1 U14761 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14762 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U14763 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11782) );
  INV_X1 U14764 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11779) );
  INV_X1 U14765 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11777) );
  OR2_X1 U14766 ( .A1(n11911), .A2(n11777), .ZN(n11778) );
  INV_X1 U14767 ( .A(n11935), .ZN(n11927) );
  OAI211_X1 U14768 ( .C1(n11876), .C2(n11779), .A(n11778), .B(n11927), .ZN(
        n11780) );
  INV_X1 U14769 ( .A(n11780), .ZN(n11781) );
  NAND4_X1 U14770 ( .A1(n11784), .A2(n11783), .A3(n11782), .A4(n11781), .ZN(
        n11785) );
  AND2_X1 U14771 ( .A1(n11786), .A2(n11785), .ZN(n11792) );
  AND2_X1 U14772 ( .A1(n11787), .A2(n11792), .ZN(n11812) );
  NAND2_X1 U14773 ( .A1(n11812), .A2(n14265), .ZN(n11791) );
  INV_X1 U14774 ( .A(n11787), .ZN(n11789) );
  NAND2_X1 U14775 ( .A1(n14265), .A2(n11792), .ZN(n11788) );
  NAND2_X1 U14776 ( .A1(n11789), .A2(n11788), .ZN(n11790) );
  NAND2_X1 U14777 ( .A1(n11791), .A2(n11790), .ZN(n11815) );
  INV_X1 U14778 ( .A(n11792), .ZN(n11793) );
  NOR2_X1 U14779 ( .A1(n14265), .A2(n11793), .ZN(n16053) );
  AOI22_X1 U14780 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U14781 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U14782 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U14783 ( .A1(n10592), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11795) );
  OAI211_X1 U14784 ( .C1(n11876), .C2(n11796), .A(n11935), .B(n11795), .ZN(
        n11797) );
  INV_X1 U14785 ( .A(n11797), .ZN(n11798) );
  NAND4_X1 U14786 ( .A1(n11801), .A2(n11800), .A3(n11799), .A4(n11798), .ZN(
        n11810) );
  AOI22_X1 U14787 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11932), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U14788 ( .A1(n11936), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U14789 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11895), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11806) );
  NAND2_X1 U14790 ( .A1(n10592), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11802) );
  OAI211_X1 U14791 ( .C1(n11876), .C2(n11803), .A(n11927), .B(n11802), .ZN(
        n11804) );
  INV_X1 U14792 ( .A(n11804), .ZN(n11805) );
  NAND4_X1 U14793 ( .A1(n11808), .A2(n11807), .A3(n11806), .A4(n11805), .ZN(
        n11809) );
  AND2_X1 U14794 ( .A1(n11810), .A2(n11809), .ZN(n11811) );
  INV_X1 U14795 ( .A(n11811), .ZN(n16955) );
  INV_X1 U14796 ( .A(n11812), .ZN(n11813) );
  AND2_X1 U14797 ( .A1(n11812), .A2(n11811), .ZN(n11816) );
  INV_X1 U14798 ( .A(n16053), .ZN(n11814) );
  INV_X1 U14799 ( .A(n11816), .ZN(n11834) );
  AOI22_X1 U14800 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U14801 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U14802 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11821) );
  INV_X1 U14803 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11818) );
  OR2_X1 U14804 ( .A1(n11911), .A2(n19884), .ZN(n11817) );
  OAI211_X1 U14805 ( .C1(n11876), .C2(n11818), .A(n11817), .B(n11935), .ZN(
        n11819) );
  INV_X1 U14806 ( .A(n11819), .ZN(n11820) );
  NAND4_X1 U14807 ( .A1(n11823), .A2(n11822), .A3(n11821), .A4(n11820), .ZN(
        n11833) );
  AOI22_X1 U14808 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U14809 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14810 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11829) );
  INV_X1 U14811 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11826) );
  INV_X1 U14812 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11824) );
  OR2_X1 U14813 ( .A1(n11911), .A2(n11824), .ZN(n11825) );
  OAI211_X1 U14814 ( .C1(n11876), .C2(n11826), .A(n11825), .B(n11927), .ZN(
        n11827) );
  INV_X1 U14815 ( .A(n11827), .ZN(n11828) );
  NAND4_X1 U14816 ( .A1(n11831), .A2(n11830), .A3(n11829), .A4(n11828), .ZN(
        n11832) );
  NAND2_X1 U14817 ( .A1(n11833), .A2(n11832), .ZN(n11837) );
  NAND2_X1 U14818 ( .A1(n11834), .A2(n11837), .ZN(n11835) );
  NOR2_X1 U14819 ( .A1(n14265), .A2(n11837), .ZN(n16046) );
  INV_X1 U14820 ( .A(n11861), .ZN(n11859) );
  AOI22_X1 U14821 ( .A1(n11936), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14822 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14823 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11847) );
  OR2_X1 U14824 ( .A1(n11911), .A2(n11842), .ZN(n11843) );
  OAI211_X1 U14825 ( .C1(n10387), .C2(n11844), .A(n11843), .B(n11935), .ZN(
        n11845) );
  INV_X1 U14826 ( .A(n11845), .ZN(n11846) );
  NAND4_X1 U14827 ( .A1(n11849), .A2(n11848), .A3(n11847), .A4(n11846), .ZN(
        n11858) );
  AOI22_X1 U14828 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14829 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14830 ( .A1(n11895), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11854) );
  INV_X1 U14831 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n21045) );
  OR2_X1 U14832 ( .A1(n10573), .A2(n21045), .ZN(n11850) );
  OAI211_X1 U14833 ( .C1(n11876), .C2(n11851), .A(n11850), .B(n11927), .ZN(
        n11852) );
  INV_X1 U14834 ( .A(n11852), .ZN(n11853) );
  NAND4_X1 U14835 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11857) );
  AND2_X1 U14836 ( .A1(n11858), .A2(n11857), .ZN(n11860) );
  NAND2_X1 U14837 ( .A1(n11859), .A2(n11860), .ZN(n11884) );
  INV_X1 U14838 ( .A(n11860), .ZN(n11863) );
  AOI21_X1 U14839 ( .B1(n11861), .B2(n11863), .A(n19668), .ZN(n11862) );
  NOR2_X1 U14840 ( .A1(n14265), .A2(n11863), .ZN(n16041) );
  AOI22_X1 U14841 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14842 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14843 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11870) );
  INV_X1 U14844 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11867) );
  OR2_X1 U14845 ( .A1(n11911), .A2(n11865), .ZN(n11866) );
  OAI211_X1 U14846 ( .C1(n11876), .C2(n11867), .A(n11866), .B(n11935), .ZN(
        n11868) );
  INV_X1 U14847 ( .A(n11868), .ZN(n11869) );
  NAND4_X1 U14848 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11883) );
  AOI22_X1 U14849 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U14850 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14851 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11879) );
  INV_X1 U14852 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11875) );
  OR2_X1 U14853 ( .A1(n11911), .A2(n11873), .ZN(n11874) );
  OAI211_X1 U14854 ( .C1(n11876), .C2(n11875), .A(n11874), .B(n11927), .ZN(
        n11877) );
  INV_X1 U14855 ( .A(n11877), .ZN(n11878) );
  NAND4_X1 U14856 ( .A1(n11881), .A2(n11880), .A3(n11879), .A4(n11878), .ZN(
        n11882) );
  NAND2_X1 U14857 ( .A1(n11883), .A2(n11882), .ZN(n11885) );
  AOI21_X1 U14858 ( .B1(n11884), .B2(n11885), .A(n19668), .ZN(n11887) );
  INV_X1 U14859 ( .A(n11884), .ZN(n11886) );
  INV_X1 U14860 ( .A(n11885), .ZN(n11888) );
  NAND2_X1 U14861 ( .A1(n11886), .A2(n11888), .ZN(n16025) );
  NAND2_X1 U14862 ( .A1(n11887), .A2(n16025), .ZN(n11889) );
  NAND2_X1 U14863 ( .A1(n9699), .A2(n11888), .ZN(n16037) );
  NOR2_X2 U14864 ( .A1(n16038), .A2(n16037), .ZN(n16036) );
  AOI22_X1 U14865 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10585), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14866 ( .A1(n11936), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11895), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11890) );
  NAND2_X1 U14867 ( .A1(n11891), .A2(n11890), .ZN(n11905) );
  AOI21_X1 U14868 ( .B1(n11932), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n11927), .ZN(n11893) );
  AOI22_X1 U14869 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11892) );
  OAI211_X1 U14870 ( .C1(n10573), .C2(n11894), .A(n11893), .B(n11892), .ZN(
        n11904) );
  AOI22_X1 U14871 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U14872 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11895), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11896) );
  NAND2_X1 U14873 ( .A1(n11897), .A2(n11896), .ZN(n11903) );
  AOI22_X1 U14874 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11900) );
  AOI21_X1 U14875 ( .B1(n11936), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n11935), .ZN(n11899) );
  OAI211_X1 U14876 ( .C1(n11898), .C2(n11901), .A(n11900), .B(n11899), .ZN(
        n11902) );
  OAI22_X1 U14877 ( .A1(n11905), .A2(n11904), .B1(n11903), .B2(n11902), .ZN(
        n16028) );
  INV_X1 U14878 ( .A(n16028), .ZN(n11906) );
  AOI22_X1 U14879 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U14880 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11907) );
  NAND2_X1 U14881 ( .A1(n11908), .A2(n11907), .ZN(n11921) );
  AOI21_X1 U14882 ( .B1(n9705), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A(n11927), .ZN(n11910) );
  AOI22_X1 U14883 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11909) );
  OAI211_X1 U14884 ( .C1(n11911), .C2(n13317), .A(n11910), .B(n11909), .ZN(
        n11920) );
  AOI22_X1 U14885 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U14886 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11913) );
  NAND2_X1 U14887 ( .A1(n11914), .A2(n11913), .ZN(n11919) );
  AOI22_X1 U14888 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11916) );
  AOI21_X1 U14889 ( .B1(n9705), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n11935), .ZN(n11915) );
  OAI211_X1 U14890 ( .C1(n11911), .C2(n11917), .A(n11916), .B(n11915), .ZN(
        n11918) );
  OAI22_X1 U14891 ( .A1(n11921), .A2(n11920), .B1(n11919), .B2(n11918), .ZN(
        n11923) );
  NOR3_X1 U14892 ( .A1(n16025), .A2(n9699), .A3(n16028), .ZN(n11922) );
  XOR2_X1 U14893 ( .A(n11923), .B(n11922), .Z(n16021) );
  INV_X1 U14894 ( .A(n11922), .ZN(n11924) );
  INV_X1 U14895 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n21174) );
  AOI22_X1 U14896 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11926) );
  NAND2_X1 U14897 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11925) );
  OAI211_X1 U14898 ( .C1(n21174), .C2(n11911), .A(n11926), .B(n11925), .ZN(
        n11943) );
  AOI21_X1 U14899 ( .B1(n9705), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A(n11927), .ZN(n11929) );
  AOI22_X1 U14900 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10592), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11928) );
  OAI211_X1 U14901 ( .C1(n10573), .C2(n11930), .A(n11929), .B(n11928), .ZN(
        n11942) );
  AOI22_X1 U14902 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U14903 ( .A1(n11932), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11933) );
  NAND2_X1 U14904 ( .A1(n11934), .A2(n11933), .ZN(n11941) );
  INV_X1 U14905 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U14906 ( .A1(n11766), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11938) );
  AOI21_X1 U14907 ( .B1(n11936), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n11935), .ZN(n11937) );
  OAI211_X1 U14908 ( .C1(n11911), .C2(n11939), .A(n11938), .B(n11937), .ZN(
        n11940) );
  OAI22_X1 U14909 ( .A1(n11943), .A2(n11942), .B1(n11941), .B2(n11940), .ZN(
        n11944) );
  INV_X1 U14910 ( .A(n11944), .ZN(n11945) );
  XNOR2_X1 U14911 ( .A(n11946), .B(n11945), .ZN(n15268) );
  AND2_X1 U14912 ( .A1(n11947), .A2(n20373), .ZN(n13433) );
  NAND2_X1 U14913 ( .A1(n11948), .A2(n13433), .ZN(n11949) );
  NOR2_X1 U14914 ( .A1(n11949), .A2(n13434), .ZN(n11950) );
  AOI21_X1 U14915 ( .B1(n13219), .B2(n13427), .A(n11950), .ZN(n12742) );
  INV_X1 U14916 ( .A(n11951), .ZN(n11952) );
  NAND2_X1 U14917 ( .A1(n11953), .A2(n11952), .ZN(n11954) );
  NAND2_X1 U14918 ( .A1(n12742), .A2(n11954), .ZN(n11955) );
  AND2_X1 U14919 ( .A1(n19905), .A2(n19896), .ZN(n11956) );
  NOR4_X1 U14920 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n11960) );
  NOR4_X1 U14921 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n11959) );
  NOR4_X1 U14922 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n11958) );
  NOR4_X1 U14923 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n11957) );
  NAND4_X1 U14924 ( .A1(n11960), .A2(n11959), .A3(n11958), .A4(n11957), .ZN(
        n11965) );
  NOR4_X1 U14925 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_14__SCAN_IN), .ZN(n11963) );
  NOR4_X1 U14926 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n11962) );
  NOR4_X1 U14927 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n11961) );
  INV_X1 U14928 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20399) );
  NAND4_X1 U14929 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n20399), .ZN(
        n11964) );
  AOI22_X1 U14930 ( .A1(n12015), .A2(n19772), .B1(BUF1_REG_30__SCAN_IN), .B2(
        n19719), .ZN(n11975) );
  AND2_X1 U14931 ( .A1(n11966), .A2(n19905), .ZN(n11967) );
  NAND2_X1 U14932 ( .A1(n13223), .A2(BUF2_REG_14__SCAN_IN), .ZN(n11970) );
  INV_X1 U14933 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n11968) );
  OR2_X1 U14934 ( .A1(n13223), .A2(n11968), .ZN(n11969) );
  NAND2_X1 U14935 ( .A1(n11970), .A2(n11969), .ZN(n19818) );
  INV_X1 U14936 ( .A(n19818), .ZN(n11972) );
  INV_X1 U14937 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n11971) );
  OAI22_X1 U14938 ( .A1(n16155), .A2(n11972), .B1(n19744), .B2(n11971), .ZN(
        n11973) );
  AOI21_X1 U14939 ( .B1(n19717), .B2(BUF2_REG_30__SCAN_IN), .A(n11973), .ZN(
        n11974) );
  OAI21_X1 U14940 ( .B1(n15268), .B2(n19754), .A(n11976), .ZN(P2_U2889) );
  NOR2_X1 U14941 ( .A1(n11980), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11979) );
  OR2_X1 U14942 ( .A1(n11542), .A2(n11979), .ZN(n12391) );
  INV_X1 U14943 ( .A(n12391), .ZN(n16899) );
  OAI21_X1 U14944 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n9740), .A(
        n10152), .ZN(n16164) );
  INV_X1 U14945 ( .A(n16164), .ZN(n16910) );
  AOI21_X1 U14946 ( .B1(n16173), .B2(n11981), .A(n9740), .ZN(n16922) );
  OAI21_X1 U14947 ( .B1(n11982), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n11981), .ZN(n16182) );
  INV_X1 U14948 ( .A(n16182), .ZN(n15934) );
  AOI21_X1 U14949 ( .B1(n16188), .B2(n11983), .A(n11982), .ZN(n16935) );
  INV_X1 U14950 ( .A(n11983), .ZN(n11984) );
  AOI21_X1 U14951 ( .B1(n16199), .B2(n11986), .A(n11984), .ZN(n16201) );
  INV_X1 U14952 ( .A(n11986), .ZN(n11987) );
  AOI21_X1 U14953 ( .B1(n16211), .B2(n11985), .A(n11987), .ZN(n16945) );
  OAI21_X1 U14954 ( .B1(n11989), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n11985), .ZN(n16222) );
  INV_X1 U14955 ( .A(n16222), .ZN(n16606) );
  NOR2_X1 U14956 ( .A1(n9793), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11988) );
  INV_X1 U14957 ( .A(n12009), .ZN(n11991) );
  AOI21_X1 U14958 ( .B1(n10144), .B2(n11990), .A(n11991), .ZN(n16268) );
  AND2_X1 U14959 ( .A1(n12007), .A2(n16285), .ZN(n11993) );
  NOR2_X1 U14960 ( .A1(n11992), .A2(n11993), .ZN(n16283) );
  AOI21_X1 U14961 ( .B1(n16305), .B2(n12006), .A(n11994), .ZN(n14319) );
  AOI21_X1 U14962 ( .B1(n16992), .B2(n12005), .A(n11995), .ZN(n16985) );
  AOI21_X1 U14963 ( .B1(n17006), .B2(n12004), .A(n11996), .ZN(n19634) );
  AOI21_X1 U14964 ( .B1(n17022), .B2(n11997), .A(n11998), .ZN(n17015) );
  AOI21_X1 U14965 ( .B1(n14295), .B2(n12003), .A(n9750), .ZN(n14480) );
  AOI21_X1 U14966 ( .B1(n17036), .B2(n12002), .A(n11999), .ZN(n17029) );
  AOI21_X1 U14967 ( .B1(n17047), .B2(n12001), .A(n12000), .ZN(n17037) );
  OAI22_X1 U14968 ( .A1(n17100), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n16537) );
  INV_X1 U14969 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19689) );
  OAI22_X1 U14970 ( .A1(n17100), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19689), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16536) );
  AND2_X1 U14971 ( .A1(n16537), .A2(n16536), .ZN(n14378) );
  OAI21_X1 U14972 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12001), .ZN(n19839) );
  NAND2_X1 U14973 ( .A1(n14378), .A2(n19839), .ZN(n14503) );
  NOR2_X1 U14974 ( .A1(n17037), .A2(n14503), .ZN(n19663) );
  OAI21_X1 U14975 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12000), .A(
        n12002), .ZN(n19833) );
  NAND2_X1 U14976 ( .A1(n19663), .A2(n19833), .ZN(n14454) );
  NOR2_X1 U14977 ( .A1(n17029), .A2(n14454), .ZN(n14278) );
  OAI21_X1 U14978 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11999), .A(
        n12003), .ZN(n14279) );
  NAND2_X1 U14979 ( .A1(n14278), .A2(n14279), .ZN(n14478) );
  NOR2_X1 U14980 ( .A1(n14480), .A2(n14478), .ZN(n19655) );
  OAI21_X1 U14981 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n9750), .A(
        n11997), .ZN(n19657) );
  NAND2_X1 U14982 ( .A1(n19655), .A2(n19657), .ZN(n14466) );
  NOR2_X1 U14983 ( .A1(n17015), .A2(n14466), .ZN(n19643) );
  OAI21_X1 U14984 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n11998), .A(
        n12004), .ZN(n19645) );
  NAND2_X1 U14985 ( .A1(n19643), .A2(n19645), .ZN(n19633) );
  NOR2_X1 U14986 ( .A1(n19634), .A2(n19633), .ZN(n19632) );
  OAI21_X1 U14987 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11996), .A(
        n12005), .ZN(n19622) );
  NAND2_X1 U14988 ( .A1(n19632), .A2(n19622), .ZN(n14492) );
  NOR2_X1 U14989 ( .A1(n16985), .A2(n14492), .ZN(n19612) );
  OAI21_X1 U14990 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11995), .A(
        n12006), .ZN(n19613) );
  NAND2_X1 U14991 ( .A1(n19612), .A2(n19613), .ZN(n14318) );
  NOR2_X1 U14992 ( .A1(n14319), .A2(n14318), .ZN(n19598) );
  OAI21_X1 U14993 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11994), .A(
        n12007), .ZN(n19599) );
  NAND2_X1 U14994 ( .A1(n19598), .A2(n19599), .ZN(n16006) );
  NOR2_X1 U14995 ( .A1(n16283), .A2(n16006), .ZN(n19586) );
  OAI21_X1 U14996 ( .B1(n11992), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n11990), .ZN(n19587) );
  NAND2_X1 U14997 ( .A1(n19586), .A2(n19587), .ZN(n15988) );
  NOR2_X1 U14998 ( .A1(n16268), .A2(n15988), .ZN(n15974) );
  AND2_X1 U14999 ( .A1(n12009), .A2(n12008), .ZN(n12010) );
  OR2_X1 U15000 ( .A1(n12010), .A2(n9793), .ZN(n16253) );
  NAND2_X1 U15001 ( .A1(n15974), .A2(n16253), .ZN(n12011) );
  NOR2_X1 U15002 ( .A1(n9783), .A2(n15973), .ZN(n15962) );
  NOR2_X1 U15003 ( .A1(n16606), .A2(n16605), .ZN(n16604) );
  NOR2_X1 U15004 ( .A1(n19656), .A2(n16604), .ZN(n16944) );
  NOR2_X1 U15005 ( .A1(n16935), .A2(n16934), .ZN(n16933) );
  NOR2_X1 U15006 ( .A1(n15934), .A2(n15935), .ZN(n15933) );
  NOR2_X1 U15007 ( .A1(n19656), .A2(n15933), .ZN(n16921) );
  NOR2_X1 U15008 ( .A1(n16922), .A2(n16921), .ZN(n16920) );
  INV_X1 U15009 ( .A(n12012), .ZN(n12013) );
  NAND4_X1 U15010 ( .A1(n20312), .A2(n17100), .A3(n21150), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19704) );
  INV_X1 U15011 ( .A(n12015), .ZN(n12030) );
  NAND2_X1 U15012 ( .A1(n11020), .A2(n12016), .ZN(n12017) );
  INV_X1 U15013 ( .A(n11022), .ZN(n12018) );
  NAND2_X1 U15014 ( .A1(n12018), .A2(n13124), .ZN(n12709) );
  NAND2_X1 U15015 ( .A1(n12629), .A2(n19688), .ZN(n19557) );
  NOR2_X1 U15016 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13444), .ZN(n12024) );
  AND2_X1 U15017 ( .A1(n12019), .A2(n12024), .ZN(n12020) );
  NOR2_X1 U15018 ( .A1(n20101), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20070) );
  INV_X1 U15019 ( .A(n20070), .ZN(n13460) );
  NOR2_X1 U15020 ( .A1(n19558), .A2(n13460), .ZN(n17092) );
  INV_X1 U15021 ( .A(n17092), .ZN(n12021) );
  NAND2_X1 U15022 ( .A1(n19704), .A2(n12021), .ZN(n12022) );
  OR2_X1 U15023 ( .A1(n19825), .A2(n12022), .ZN(n12023) );
  NAND2_X1 U15024 ( .A1(n19676), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19690) );
  NAND2_X1 U15025 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19672), .ZN(
        n12029) );
  NOR2_X2 U15026 ( .A1(n12629), .A2(n14265), .ZN(n19821) );
  INV_X1 U15027 ( .A(n12024), .ZN(n12025) );
  NAND2_X1 U15028 ( .A1(n19821), .A2(n12025), .ZN(n16886) );
  AND2_X1 U15029 ( .A1(n20373), .A2(n21150), .ZN(n12026) );
  NOR2_X1 U15030 ( .A1(n12629), .A2(n12026), .ZN(n12032) );
  INV_X1 U15031 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16952) );
  NAND2_X1 U15032 ( .A1(n12032), .A2(n16952), .ZN(n12027) );
  NAND2_X2 U15033 ( .A1(n16886), .A2(n12027), .ZN(n19678) );
  AOI22_X1 U15034 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19678), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19697), .ZN(n12028) );
  OAI211_X1 U15035 ( .C1(n12030), .C2(n19703), .A(n12029), .B(n12028), .ZN(
        n12034) );
  AND2_X1 U15036 ( .A1(n14265), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12031) );
  NAND2_X1 U15037 ( .A1(n14265), .A2(n20373), .ZN(n12035) );
  OAI21_X1 U15038 ( .B1(n16890), .B2(n12039), .A(n12038), .ZN(P2_U2825) );
  NOR2_X2 U15039 ( .A1(n12045), .A2(n17603), .ZN(n12175) );
  AOI22_X1 U15040 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12055) );
  INV_X2 U15041 ( .A(n10339), .ZN(n17797) );
  AOI22_X1 U15042 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12054) );
  NOR2_X1 U15043 ( .A1(n12046), .A2(n12041), .ZN(n12177) );
  INV_X1 U15044 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n21187) );
  AOI22_X1 U15045 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12040) );
  OAI21_X1 U15046 ( .B1(n12215), .B2(n21187), .A(n12040), .ZN(n12052) );
  AOI22_X1 U15047 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17820), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12050) );
  NOR2_X2 U15048 ( .A1(n12042), .A2(n12043), .ZN(n12093) );
  CLKBUF_X3 U15049 ( .A(n12093), .Z(n17856) );
  AOI22_X1 U15050 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15051 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12048) );
  NOR2_X2 U15052 ( .A1(n12046), .A2(n12045), .ZN(n12128) );
  AOI22_X1 U15053 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12130), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15054 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12051) );
  AOI211_X1 U15055 ( .C1(n17859), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n12052), .B(n12051), .ZN(n12053) );
  NAND3_X1 U15056 ( .A1(n12055), .A2(n12054), .A3(n12053), .ZN(n18036) );
  AOI22_X1 U15057 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12065) );
  INV_X2 U15058 ( .A(n10339), .ZN(n17758) );
  AOI22_X1 U15059 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12064) );
  INV_X1 U15060 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n21193) );
  AOI22_X1 U15061 ( .A1(n12130), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12056) );
  OAI21_X1 U15062 ( .B1(n9754), .B2(n21193), .A(n12056), .ZN(n12062) );
  AOI22_X1 U15063 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12060) );
  INV_X2 U15064 ( .A(n12215), .ZN(n17880) );
  AOI22_X1 U15065 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17856), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15066 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15067 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12057) );
  NAND4_X1 U15068 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n12057), .ZN(
        n12061) );
  AOI211_X1 U15069 ( .C1(n12175), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n12062), .B(n12061), .ZN(n12063) );
  NAND3_X1 U15070 ( .A1(n12065), .A2(n12064), .A3(n12063), .ZN(n12250) );
  AOI22_X1 U15071 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15072 ( .A1(n12105), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12074) );
  INV_X1 U15073 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n21181) );
  AOI22_X1 U15074 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12066) );
  OAI21_X1 U15075 ( .B1(n10339), .B2(n21181), .A(n12066), .ZN(n12072) );
  AOI22_X1 U15076 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17820), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15077 ( .A1(n12175), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12091), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15078 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15079 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12067) );
  NAND4_X1 U15080 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12071) );
  AOI211_X1 U15081 ( .C1(n17855), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n12072), .B(n12071), .ZN(n12073) );
  AOI22_X1 U15082 ( .A1(n12105), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15083 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15084 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15085 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12130), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12076) );
  NAND4_X1 U15086 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(
        n12085) );
  AOI22_X1 U15087 ( .A1(n17857), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12086), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12083) );
  INV_X2 U15088 ( .A(n16558), .ZN(n17875) );
  AOI22_X1 U15089 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12175), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15090 ( .A1(n12093), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12091), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15091 ( .A1(n12128), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12080) );
  NAND4_X1 U15092 ( .A1(n12083), .A2(n12082), .A3(n12081), .A4(n12080), .ZN(
        n12084) );
  INV_X2 U15093 ( .A(n9754), .ZN(n17857) );
  AOI22_X1 U15094 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17797), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17857), .ZN(n12090) );
  AOI22_X1 U15095 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n12216), .ZN(n12089) );
  AOI22_X1 U15096 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n12130), .ZN(n12088) );
  AOI22_X1 U15097 ( .A1(n12128), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12086), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15098 ( .A1(n12105), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n16556), .ZN(n12100) );
  INV_X1 U15099 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n21120) );
  AOI22_X1 U15100 ( .A1(n12093), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12092), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12094) );
  OAI21_X1 U15101 ( .B1(n21120), .B2(n17745), .A(n12094), .ZN(n12097) );
  AOI22_X1 U15102 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12175), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15103 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15104 ( .A1(n17857), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15105 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9695), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15106 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12101) );
  NAND4_X1 U15107 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12111) );
  INV_X2 U15108 ( .A(n9746), .ZN(n17873) );
  AOI22_X1 U15109 ( .A1(n12175), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15110 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15111 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17763), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15112 ( .A1(n17844), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12106) );
  NAND4_X1 U15113 ( .A1(n12109), .A2(n12108), .A3(n12107), .A4(n12106), .ZN(
        n12110) );
  AOI22_X1 U15114 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15115 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15116 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15117 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12112) );
  NAND4_X1 U15118 ( .A1(n12115), .A2(n12114), .A3(n12113), .A4(n12112), .ZN(
        n12121) );
  AOI22_X1 U15119 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15120 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15121 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15122 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12116) );
  NAND4_X1 U15123 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(
        n12120) );
  INV_X1 U15124 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18205) );
  INV_X1 U15125 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18692) );
  AOI21_X1 U15126 ( .B1(n17116), .B2(n12122), .A(n18463), .ZN(n12148) );
  INV_X1 U15127 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18817) );
  XOR2_X1 U15128 ( .A(n18044), .B(n12123), .Z(n18499) );
  NAND2_X1 U15129 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12126), .ZN(
        n12143) );
  XOR2_X1 U15130 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12126), .Z(
        n18513) );
  INV_X1 U15131 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18842) );
  OR2_X1 U15132 ( .A1(n18842), .A2(n12127), .ZN(n12139) );
  XOR2_X1 U15133 ( .A(n18842), .B(n12127), .Z(n18536) );
  INV_X1 U15134 ( .A(n18066), .ZN(n12256) );
  NAND2_X1 U15135 ( .A1(n12256), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12138) );
  XNOR2_X1 U15136 ( .A(n18066), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18545) );
  AOI22_X1 U15137 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15138 ( .A1(n17857), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12136) );
  INV_X1 U15139 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18897) );
  AOI22_X1 U15140 ( .A1(n12175), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12129) );
  OAI21_X1 U15141 ( .B1(n12221), .B2(n18897), .A(n12129), .ZN(n12135) );
  AOI22_X1 U15142 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12091), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15143 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15144 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15145 ( .A1(n12086), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12130), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12131) );
  INV_X1 U15146 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19519) );
  NOR2_X1 U15147 ( .A1(n18553), .A2(n19519), .ZN(n18552) );
  NAND2_X1 U15148 ( .A1(n18545), .A2(n18552), .ZN(n18544) );
  NAND2_X1 U15149 ( .A1(n12138), .A2(n18544), .ZN(n18535) );
  NAND2_X1 U15150 ( .A1(n18536), .A2(n18535), .ZN(n18534) );
  NAND2_X1 U15151 ( .A1(n12139), .A2(n18534), .ZN(n18523) );
  XNOR2_X1 U15152 ( .A(n12252), .B(n12140), .ZN(n12141) );
  XOR2_X1 U15153 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12141), .Z(
        n18524) );
  NAND2_X1 U15154 ( .A1(n18523), .A2(n18524), .ZN(n18522) );
  NAND2_X1 U15155 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12141), .ZN(
        n12142) );
  NAND2_X1 U15156 ( .A1(n18522), .A2(n12142), .ZN(n18512) );
  XOR2_X1 U15157 ( .A(n12145), .B(n12144), .Z(n12146) );
  XOR2_X1 U15158 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12146), .Z(
        n18483) );
  NAND2_X1 U15159 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12146), .ZN(
        n12147) );
  NAND2_X1 U15160 ( .A1(n12148), .A2(n12149), .ZN(n12150) );
  OR2_X2 U15161 ( .A1(n12151), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18423) );
  NAND2_X1 U15163 ( .A1(n18423), .A2(n18461), .ZN(n18379) );
  INV_X1 U15164 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18699) );
  INV_X1 U15165 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18721) );
  INV_X1 U15166 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18776) );
  INV_X1 U15167 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18424) );
  NOR2_X1 U15168 ( .A1(n18776), .A2(n18424), .ZN(n18756) );
  NAND2_X1 U15169 ( .A1(n18756), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18736) );
  INV_X1 U15170 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18749) );
  NOR2_X1 U15171 ( .A1(n18736), .A2(n18749), .ZN(n18732) );
  NAND2_X1 U15172 ( .A1(n18732), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18718) );
  NOR2_X1 U15173 ( .A1(n18721), .A2(n18718), .ZN(n18689) );
  INV_X1 U15174 ( .A(n18689), .ZN(n18700) );
  NOR2_X1 U15175 ( .A1(n18699), .A2(n18700), .ZN(n18345) );
  INV_X1 U15176 ( .A(n18345), .ZN(n18671) );
  NOR2_X1 U15177 ( .A1(n18379), .A2(n18671), .ZN(n12154) );
  NOR2_X1 U15178 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18435) );
  INV_X1 U15179 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18413) );
  NAND2_X1 U15180 ( .A1(n12152), .A2(n18382), .ZN(n12153) );
  INV_X1 U15181 ( .A(n12153), .ZN(n12155) );
  NAND2_X1 U15182 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18662) );
  NAND2_X1 U15183 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18290) );
  INV_X1 U15184 ( .A(n18290), .ZN(n18642) );
  NAND2_X1 U15185 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18642), .ZN(
        n18629) );
  INV_X1 U15186 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18636) );
  OR2_X1 U15187 ( .A1(n18629), .A2(n18636), .ZN(n12156) );
  INV_X1 U15188 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18321) );
  NOR2_X1 U15189 ( .A1(n18662), .A2(n18321), .ZN(n18638) );
  INV_X1 U15190 ( .A(n18638), .ZN(n18309) );
  NOR2_X1 U15191 ( .A1(n18309), .A2(n12156), .ZN(n12349) );
  NAND2_X1 U15192 ( .A1(n12349), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18246) );
  NAND2_X1 U15193 ( .A1(n18321), .A2(n18382), .ZN(n18320) );
  NOR2_X1 U15194 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18320), .ZN(
        n12157) );
  INV_X1 U15195 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18306) );
  NAND2_X1 U15196 ( .A1(n12157), .A2(n18306), .ZN(n18282) );
  NOR2_X1 U15197 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18282), .ZN(
        n18275) );
  INV_X1 U15198 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21089) );
  NAND3_X1 U15199 ( .A1(n18275), .A2(n18636), .A3(n21089), .ZN(n12158) );
  INV_X1 U15200 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18609) );
  NAND2_X1 U15201 ( .A1(n18248), .A2(n18609), .ZN(n18247) );
  NAND3_X1 U15202 ( .A1(n18252), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n18247), .ZN(n12163) );
  NAND2_X1 U15203 ( .A1(n12163), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12162) );
  INV_X1 U15204 ( .A(n18247), .ZN(n18231) );
  INV_X1 U15205 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18588) );
  INV_X1 U15206 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18585) );
  NAND2_X1 U15207 ( .A1(n18463), .A2(n12163), .ZN(n18230) );
  NOR2_X1 U15208 ( .A1(n18588), .A2(n18585), .ZN(n12303) );
  INV_X1 U15209 ( .A(n18201), .ZN(n12345) );
  AOI21_X1 U15210 ( .B1(n18463), .B2(n18200), .A(n12345), .ZN(n18183) );
  NOR2_X1 U15211 ( .A1(n18382), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16593) );
  AOI21_X1 U15212 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18382), .A(
        n16593), .ZN(n18182) );
  NOR2_X1 U15213 ( .A1(n18183), .A2(n18182), .ZN(n18181) );
  AOI22_X1 U15214 ( .A1(n17879), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15215 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9698), .B1(
        n17826), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15216 ( .A1(n16556), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12166) );
  INV_X2 U15217 ( .A(n17745), .ZN(n16555) );
  AOI22_X1 U15218 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12165) );
  NAND4_X1 U15219 ( .A1(n12168), .A2(n12167), .A3(n12166), .A4(n12165), .ZN(
        n12174) );
  AOI22_X1 U15220 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17763), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12172) );
  INV_X2 U15221 ( .A(n12215), .ZN(n17839) );
  AOI22_X1 U15222 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17839), .ZN(n12171) );
  AOI22_X1 U15223 ( .A1(n17758), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15224 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17855), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12169) );
  NAND4_X1 U15225 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(
        n12173) );
  AOI22_X1 U15226 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15227 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12185) );
  INV_X1 U15228 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n21247) );
  AOI22_X1 U15229 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12176) );
  OAI21_X1 U15230 ( .B1(n9746), .B2(n21247), .A(n12176), .ZN(n12183) );
  AOI22_X1 U15231 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15232 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17763), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15233 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15234 ( .A1(n12130), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12178) );
  NAND4_X1 U15235 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12182) );
  NOR2_X1 U15236 ( .A1(n19539), .A2(n12326), .ZN(n12328) );
  AOI22_X1 U15237 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17797), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15238 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12193) );
  INV_X1 U15239 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18925) );
  AOI22_X1 U15240 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12187) );
  OAI21_X1 U15241 ( .B1(n17745), .B2(n18925), .A(n12187), .ZN(n12192) );
  AOI22_X1 U15242 ( .A1(n17857), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15243 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15244 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12175), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15245 ( .A1(n17820), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12188) );
  NAND2_X1 U15246 ( .A1(n12328), .A2(n17926), .ZN(n12337) );
  AOI22_X1 U15247 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12198) );
  INV_X1 U15248 ( .A(n16558), .ZN(n17820) );
  AOI22_X1 U15249 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17820), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15250 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15251 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12195) );
  NAND4_X1 U15252 ( .A1(n12198), .A2(n12197), .A3(n12196), .A4(n12195), .ZN(
        n12204) );
  AOI22_X1 U15253 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15254 ( .A1(n9698), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U15255 ( .A1(n17857), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15256 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17763), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12199) );
  NAND4_X1 U15257 ( .A1(n12202), .A2(n12201), .A3(n12200), .A4(n12199), .ZN(
        n12203) );
  AOI22_X1 U15258 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15259 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15260 ( .A1(n9698), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17826), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15261 ( .A1(n17857), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12130), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12205) );
  NAND4_X1 U15262 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12214) );
  AOI22_X1 U15263 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15264 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15265 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15266 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12209) );
  NAND4_X1 U15267 ( .A1(n12212), .A2(n12211), .A3(n12210), .A4(n12209), .ZN(
        n12213) );
  NOR2_X1 U15268 ( .A1(n18917), .A2(n17926), .ZN(n19359) );
  AOI22_X1 U15269 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15270 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15271 ( .A1(n17857), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15272 ( .A1(n12130), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12217) );
  NAND4_X1 U15273 ( .A1(n12220), .A2(n12219), .A3(n12218), .A4(n12217), .ZN(
        n12227) );
  AOI22_X1 U15274 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17855), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15275 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15276 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15277 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12222) );
  NAND4_X1 U15278 ( .A1(n12225), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        n12226) );
  AOI22_X1 U15279 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15280 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15281 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15282 ( .A1(n17758), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12228) );
  NAND4_X1 U15283 ( .A1(n12231), .A2(n12230), .A3(n12229), .A4(n12228), .ZN(
        n12237) );
  AOI22_X1 U15284 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15285 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15286 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15287 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12232) );
  NAND4_X1 U15288 ( .A1(n12235), .A2(n12234), .A3(n12233), .A4(n12232), .ZN(
        n12236) );
  AOI22_X1 U15289 ( .A1(n9698), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17857), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15290 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17797), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15291 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12238) );
  OAI21_X1 U15292 ( .B1(n17745), .B2(n18897), .A(n12238), .ZN(n12244) );
  AOI22_X1 U15293 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15294 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17856), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15295 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15296 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12239) );
  NAND4_X1 U15297 ( .A1(n12242), .A2(n12241), .A3(n12240), .A4(n12239), .ZN(
        n12243) );
  NOR2_X1 U15298 ( .A1(n17562), .A2(n19539), .ZN(n12291) );
  OR2_X1 U15299 ( .A1(n12326), .A2(n12291), .ZN(n12289) );
  NOR2_X1 U15300 ( .A1(n12280), .A2(n12289), .ZN(n12248) );
  OAI211_X1 U15301 ( .C1(n18914), .C2(n19359), .A(n12300), .B(n12248), .ZN(
        n12331) );
  NOR2_X1 U15302 ( .A1(n12337), .A2(n12331), .ZN(n17109) );
  INV_X1 U15303 ( .A(n17109), .ZN(n19326) );
  NOR4_X1 U15304 ( .A1(n16595), .A2(n17116), .A3(n18181), .A4(n19326), .ZN(
        n12343) );
  NAND2_X1 U15305 ( .A1(n16683), .A2(n18066), .ZN(n12254) );
  NAND2_X1 U15306 ( .A1(n12249), .A2(n12254), .ZN(n12253) );
  NAND2_X1 U15307 ( .A1(n12253), .A2(n12252), .ZN(n12262) );
  NOR2_X1 U15308 ( .A1(n18047), .A2(n12262), .ZN(n12251) );
  NAND2_X1 U15309 ( .A1(n12251), .A2(n12250), .ZN(n12268) );
  NOR2_X1 U15310 ( .A1(n18041), .A2(n12268), .ZN(n12272) );
  NAND2_X1 U15311 ( .A1(n12272), .A2(n18036), .ZN(n12273) );
  XOR2_X1 U15312 ( .A(n12251), .B(n12250), .Z(n12266) );
  INV_X1 U15313 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18840) );
  XNOR2_X1 U15314 ( .A(n12253), .B(n12252), .ZN(n12260) );
  NOR2_X1 U15315 ( .A1(n18840), .A2(n12260), .ZN(n12261) );
  XNOR2_X1 U15316 ( .A(n18056), .B(n12254), .ZN(n12258) );
  NOR2_X1 U15317 ( .A1(n12258), .A2(n18842), .ZN(n12259) );
  NOR2_X1 U15318 ( .A1(n12256), .A2(n19519), .ZN(n12257) );
  NAND3_X1 U15319 ( .A1(n18553), .A2(n12256), .A3(n19519), .ZN(n12255) );
  OAI221_X1 U15320 ( .B1(n12257), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18553), .C2(n12256), .A(n12255), .ZN(n18533) );
  XOR2_X1 U15321 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12258), .Z(
        n18532) );
  NOR2_X1 U15322 ( .A1(n18533), .A2(n18532), .ZN(n18531) );
  NOR2_X1 U15323 ( .A1(n12259), .A2(n18531), .ZN(n18521) );
  XOR2_X1 U15324 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12260), .Z(
        n18520) );
  NOR2_X1 U15325 ( .A1(n18521), .A2(n18520), .ZN(n18519) );
  NOR2_X1 U15326 ( .A1(n12261), .A2(n18519), .ZN(n12263) );
  XNOR2_X1 U15327 ( .A(n12262), .B(n18047), .ZN(n12264) );
  NOR2_X1 U15328 ( .A1(n12263), .A2(n12264), .ZN(n12265) );
  INV_X1 U15329 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18811) );
  XNOR2_X1 U15330 ( .A(n12264), .B(n12263), .ZN(n18508) );
  XOR2_X1 U15331 ( .A(n18817), .B(n12266), .Z(n18495) );
  XNOR2_X1 U15332 ( .A(n12268), .B(n18041), .ZN(n12270) );
  NOR2_X1 U15333 ( .A1(n12269), .A2(n12270), .ZN(n12271) );
  XNOR2_X1 U15334 ( .A(n12270), .B(n12269), .ZN(n18488) );
  INV_X1 U15335 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18808) );
  XOR2_X1 U15336 ( .A(n12272), .B(n17116), .Z(n12275) );
  NAND2_X1 U15337 ( .A1(n12274), .A2(n12275), .ZN(n18472) );
  INV_X1 U15338 ( .A(n12273), .ZN(n12278) );
  OR2_X1 U15339 ( .A1(n12275), .A2(n12274), .ZN(n18473) );
  OAI21_X1 U15340 ( .B1(n12278), .B2(n12277), .A(n18473), .ZN(n12276) );
  INV_X1 U15341 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21202) );
  NOR2_X2 U15342 ( .A1(n18460), .A2(n21202), .ZN(n18459) );
  NAND2_X1 U15343 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18566) );
  INV_X1 U15344 ( .A(n18566), .ZN(n12301) );
  NAND2_X1 U15345 ( .A1(n12349), .A2(n12301), .ZN(n18587) );
  OR2_X2 U15346 ( .A1(n18623), .A2(n18587), .ZN(n18229) );
  INV_X1 U15347 ( .A(n12303), .ZN(n18568) );
  NOR2_X2 U15348 ( .A1(n18229), .A2(n18568), .ZN(n18570) );
  INV_X1 U15349 ( .A(n18570), .ZN(n18195) );
  NAND2_X1 U15350 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17142) );
  NOR2_X1 U15351 ( .A1(n18195), .A2(n17142), .ZN(n17147) );
  INV_X1 U15352 ( .A(n19542), .ZN(n19550) );
  NOR2_X1 U15353 ( .A1(n18914), .A2(n17926), .ZN(n19337) );
  NAND3_X1 U15354 ( .A1(n12300), .A2(n12329), .A3(n19337), .ZN(n14658) );
  INV_X1 U15355 ( .A(n18909), .ZN(n12296) );
  NAND2_X1 U15356 ( .A1(n18914), .A2(n18922), .ZN(n12287) );
  NOR2_X1 U15357 ( .A1(n12326), .A2(n12287), .ZN(n12284) );
  NAND4_X1 U15358 ( .A1(n12300), .A2(n18917), .A3(n12284), .A4(n17562), .ZN(
        n18124) );
  INV_X1 U15359 ( .A(n18124), .ZN(n18122) );
  INV_X1 U15360 ( .A(n12326), .ZN(n18904) );
  NOR2_X1 U15361 ( .A1(n18929), .A2(n17562), .ZN(n12281) );
  NAND4_X1 U15362 ( .A1(n18909), .A2(n18914), .A3(n12285), .A4(n12281), .ZN(
        n12282) );
  INV_X1 U15363 ( .A(n12282), .ZN(n12297) );
  OAI21_X1 U15364 ( .B1(n18929), .B2(n19359), .A(n12283), .ZN(n12332) );
  OAI21_X1 U15365 ( .B1(n12329), .B2(n12284), .A(n12332), .ZN(n12295) );
  NOR2_X1 U15366 ( .A1(n18929), .A2(n12285), .ZN(n12294) );
  INV_X1 U15367 ( .A(n12285), .ZN(n12325) );
  AOI21_X1 U15368 ( .B1(n18904), .B2(n18893), .A(n19359), .ZN(n12286) );
  AOI21_X1 U15369 ( .B1(n12287), .B2(n12325), .A(n12286), .ZN(n12288) );
  AOI21_X1 U15370 ( .B1(n12325), .B2(n12289), .A(n12288), .ZN(n12293) );
  OR3_X1 U15371 ( .A1(n12296), .A2(n12291), .A3(n12290), .ZN(n12292) );
  OAI211_X1 U15372 ( .C1(n18914), .C2(n12294), .A(n12293), .B(n12292), .ZN(
        n12330) );
  AOI21_X1 U15373 ( .B1(n12296), .B2(n12295), .A(n12330), .ZN(n12298) );
  NAND2_X1 U15374 ( .A1(n12297), .A2(n12298), .ZN(n12372) );
  NAND2_X1 U15375 ( .A1(n19343), .A2(n12372), .ZN(n19331) );
  NAND2_X1 U15376 ( .A1(n18125), .A2(n19343), .ZN(n12299) );
  OAI21_X1 U15377 ( .B1(n12300), .B2(n12299), .A(n12298), .ZN(n19335) );
  NOR2_X4 U15378 ( .A1(n18763), .A2(n19358), .ZN(n18783) );
  OR2_X1 U15379 ( .A1(n17147), .A2(n18601), .ZN(n12341) );
  NOR2_X1 U15380 ( .A1(n18587), .A2(n18697), .ZN(n18228) );
  NAND2_X1 U15381 ( .A1(n12303), .A2(n18228), .ZN(n18572) );
  OR2_X1 U15382 ( .A1(n17142), .A2(n18572), .ZN(n12339) );
  NOR2_X1 U15383 ( .A1(n19326), .A2(n18036), .ZN(n18730) );
  INV_X1 U15384 ( .A(n18763), .ZN(n18758) );
  INV_X1 U15385 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21225) );
  NOR3_X1 U15386 ( .A1(n21225), .A2(n18808), .A3(n21202), .ZN(n18669) );
  NAND3_X1 U15387 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18668) );
  NAND2_X1 U15388 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18820) );
  NOR2_X1 U15389 ( .A1(n18668), .A2(n18820), .ZN(n18778) );
  NAND2_X1 U15390 ( .A1(n18669), .A2(n18778), .ZN(n18684) );
  NOR2_X1 U15391 ( .A1(n18671), .A2(n18684), .ZN(n18661) );
  NOR2_X1 U15392 ( .A1(n18587), .A2(n18568), .ZN(n17125) );
  NAND2_X1 U15393 ( .A1(n18661), .A2(n17125), .ZN(n12305) );
  NOR2_X1 U15394 ( .A1(n19519), .A2(n18684), .ZN(n18712) );
  INV_X1 U15395 ( .A(n18712), .ZN(n18771) );
  NOR2_X1 U15396 ( .A1(n18671), .A2(n18771), .ZN(n18686) );
  NAND2_X1 U15397 ( .A1(n12349), .A2(n18686), .ZN(n18563) );
  INV_X1 U15398 ( .A(n18563), .ZN(n12302) );
  NAND2_X1 U15399 ( .A1(n12301), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18580) );
  INV_X1 U15400 ( .A(n18580), .ZN(n18221) );
  NAND2_X1 U15401 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18221), .ZN(
        n18562) );
  NOR2_X1 U15402 ( .A1(n18205), .A2(n18562), .ZN(n12350) );
  AOI21_X1 U15403 ( .B1(n12302), .B2(n12350), .A(n19345), .ZN(n12304) );
  AOI21_X1 U15404 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18844) );
  NOR2_X1 U15405 ( .A1(n18844), .A2(n18668), .ZN(n18779) );
  NAND2_X1 U15406 ( .A1(n18779), .A2(n18669), .ZN(n18685) );
  NOR2_X1 U15407 ( .A1(n18671), .A2(n18685), .ZN(n18627) );
  NAND2_X1 U15408 ( .A1(n12349), .A2(n18627), .ZN(n18607) );
  OAI21_X1 U15409 ( .B1(n18566), .B2(n18607), .A(n19334), .ZN(n18590) );
  OAI21_X1 U15410 ( .B1(n12303), .B2(n19353), .A(n18590), .ZN(n18567) );
  AOI211_X1 U15411 ( .C1(n19331), .C2(n12305), .A(n12304), .B(n18567), .ZN(
        n16659) );
  NAND2_X1 U15412 ( .A1(n19503), .A2(n19492), .ZN(n19497) );
  NOR2_X1 U15413 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19497), .ZN(n19552) );
  INV_X1 U15414 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n17110) );
  INV_X2 U15415 ( .A(n18833), .ZN(n18828) );
  NAND2_X1 U15416 ( .A1(n19364), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12313) );
  OAI22_X1 U15417 ( .A1(n12306), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19371), .B2(n19350), .ZN(n12311) );
  OAI22_X1 U15418 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19375), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12308), .ZN(n12315) );
  NOR2_X1 U15419 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19375), .ZN(
        n12309) );
  NAND2_X1 U15420 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12308), .ZN(
        n12314) );
  AOI22_X1 U15421 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12315), .B1(
        n12309), .B2(n12314), .ZN(n12324) );
  OAI21_X1 U15422 ( .B1(n12312), .B2(n12311), .A(n12324), .ZN(n12310) );
  INV_X1 U15423 ( .A(n12322), .ZN(n12318) );
  OAI21_X1 U15424 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19364), .A(
        n12313), .ZN(n12319) );
  XOR2_X1 U15425 ( .A(n12313), .B(n12320), .Z(n12317) );
  INV_X1 U15426 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19330) );
  AND2_X1 U15427 ( .A1(n12314), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12316) );
  OAI22_X1 U15428 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19330), .B1(
        n12316), .B2(n12315), .ZN(n12321) );
  OAI21_X1 U15429 ( .B1(n12318), .B2(n12319), .A(n19324), .ZN(n17108) );
  NOR2_X1 U15430 ( .A1(n12320), .A2(n12319), .ZN(n12323) );
  OAI21_X1 U15431 ( .B1(n12326), .B2(n12325), .A(n18914), .ZN(n12336) );
  INV_X1 U15432 ( .A(n19324), .ZN(n17257) );
  NAND2_X1 U15433 ( .A1(n19419), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19548) );
  INV_X2 U15434 ( .A(n19548), .ZN(n19484) );
  NAND2_X1 U15435 ( .A1(n19484), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19480) );
  OAI211_X1 U15436 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19419), .B(n19474), .ZN(n19537) );
  OAI21_X1 U15437 ( .B1(n18904), .B2(n18125), .A(n19537), .ZN(n12327) );
  NAND2_X1 U15438 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19540) );
  OAI21_X1 U15439 ( .B1(n12328), .B2(n12327), .A(n19540), .ZN(n17256) );
  NOR3_X1 U15440 ( .A1(n12329), .A2(n17257), .A3(n17256), .ZN(n12335) );
  NOR2_X1 U15441 ( .A1(n12331), .A2(n12330), .ZN(n12334) );
  OAI21_X1 U15442 ( .B1(n12334), .B2(n12333), .A(n12332), .ZN(n16580) );
  AOI211_X1 U15443 ( .C1(n19321), .C2(n12336), .A(n12335), .B(n16580), .ZN(
        n12338) );
  NAND2_X1 U15444 ( .A1(n19503), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19396) );
  NOR2_X1 U15445 ( .A1(n19396), .A2(n19393), .ZN(n19535) );
  INV_X1 U15446 ( .A(n19535), .ZN(n19391) );
  AOI221_X4 U15447 ( .B1(n17108), .B2(n12338), .C1(n12337), .C2(n12338), .A(
        n19391), .ZN(n18854) );
  OAI211_X1 U15448 ( .C1(n18758), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16659), .B(n18841), .ZN(n16592) );
  NAND2_X1 U15449 ( .A1(n12341), .A2(n12340), .ZN(n12342) );
  INV_X1 U15450 ( .A(n18833), .ZN(n18869) );
  AND2_X1 U15451 ( .A1(n12344), .A2(n18833), .ZN(n12348) );
  NAND2_X1 U15452 ( .A1(n18036), .A2(n18868), .ZN(n18740) );
  AND3_X1 U15453 ( .A1(n12345), .A2(n18788), .A3(n18182), .ZN(n12347) );
  AND3_X1 U15454 ( .A1(n16593), .A2(n18868), .A3(n18183), .ZN(n12346) );
  AOI211_X1 U15455 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n12348), .A(
        n12347), .B(n12346), .ZN(n12352) );
  NAND2_X1 U15456 ( .A1(n18869), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n18188) );
  INV_X1 U15457 ( .A(n18730), .ZN(n18603) );
  OAI22_X1 U15458 ( .A1(n18731), .A2(n18601), .B1(n18729), .B2(n18603), .ZN(
        n18667) );
  INV_X1 U15459 ( .A(n18627), .ZN(n18663) );
  AOI21_X1 U15460 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19358), .A(
        n19331), .ZN(n18852) );
  INV_X1 U15461 ( .A(n18661), .ZN(n18625) );
  OAI22_X1 U15462 ( .A1(n19353), .A2(n18663), .B1(n18852), .B2(n18625), .ZN(
        n18586) );
  AOI21_X1 U15463 ( .B1(n18345), .B2(n18667), .A(n18586), .ZN(n18561) );
  NOR2_X1 U15464 ( .A1(n18561), .A2(n18871), .ZN(n18656) );
  NAND2_X1 U15465 ( .A1(n12349), .A2(n18656), .ZN(n18615) );
  INV_X1 U15466 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16591) );
  NAND2_X1 U15467 ( .A1(n12350), .A2(n16591), .ZN(n18199) );
  NAND3_X1 U15468 ( .A1(n12352), .A2(n18188), .A3(n12351), .ZN(P3_U2834) );
  INV_X1 U15469 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17328) );
  INV_X1 U15470 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18337) );
  NAND2_X1 U15471 ( .A1(n12357), .A2(n10330), .ZN(n18295) );
  INV_X1 U15472 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21230) );
  NAND3_X1 U15473 ( .A1(n18269), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12355) );
  NAND2_X1 U15474 ( .A1(n18234), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12353) );
  INV_X1 U15475 ( .A(n12353), .ZN(n12365) );
  NAND2_X1 U15476 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12365), .ZN(
        n12354) );
  INV_X1 U15477 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18244) );
  NOR3_X1 U15478 ( .A1(n18244), .A2(n17328), .A3(n12353), .ZN(n12366) );
  AOI21_X1 U15479 ( .B1(n17328), .B2(n12354), .A(n12366), .ZN(n18227) );
  XNOR2_X1 U15480 ( .A(n18244), .B(n12365), .ZN(n18240) );
  INV_X1 U15481 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18270) );
  INV_X1 U15482 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18286) );
  INV_X1 U15483 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18548) );
  NOR2_X1 U15484 ( .A1(n18295), .A2(n18548), .ZN(n18267) );
  NAND2_X1 U15485 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18267), .ZN(
        n12363) );
  OR2_X1 U15486 ( .A1(n18286), .A2(n12363), .ZN(n12356) );
  NOR2_X1 U15487 ( .A1(n12355), .A2(n18548), .ZN(n12364) );
  AOI21_X1 U15488 ( .B1(n18270), .B2(n12356), .A(n12364), .ZN(n18273) );
  XOR2_X1 U15489 ( .A(n18286), .B(n12363), .Z(n18289) );
  INV_X1 U15490 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n21075) );
  INV_X1 U15491 ( .A(n12357), .ZN(n18316) );
  NOR2_X1 U15492 ( .A1(n18316), .A2(n18548), .ZN(n18307) );
  NAND2_X1 U15493 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18307), .ZN(
        n12358) );
  AOI21_X1 U15494 ( .B1(n21075), .B2(n12358), .A(n18267), .ZN(n18308) );
  NOR2_X1 U15495 ( .A1(n18336), .A2(n18548), .ZN(n12360) );
  INV_X1 U15496 ( .A(n12360), .ZN(n12359) );
  AOI21_X1 U15497 ( .B1(n18337), .B2(n12359), .A(n18307), .ZN(n18339) );
  NOR2_X1 U15498 ( .A1(n18349), .A2(n18548), .ZN(n18347) );
  NAND2_X1 U15499 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18347), .ZN(
        n17426) );
  AOI21_X1 U15500 ( .B1(n18350), .B2(n17426), .A(n12360), .ZN(n18348) );
  INV_X1 U15501 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18213) );
  INV_X1 U15502 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18184) );
  NAND2_X1 U15503 ( .A1(n17149), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17111) );
  NAND2_X1 U15504 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n12371), .ZN(
        n17126) );
  INV_X1 U15505 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17276) );
  NOR2_X1 U15506 ( .A1(n18348), .A2(n10325), .ZN(n17418) );
  NOR2_X1 U15507 ( .A1(n17418), .A2(n10186), .ZN(n17409) );
  NOR2_X1 U15508 ( .A1(n18339), .A2(n17409), .ZN(n17408) );
  NOR2_X1 U15509 ( .A1(n17408), .A2(n10186), .ZN(n17402) );
  INV_X1 U15510 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18327) );
  XOR2_X1 U15511 ( .A(n18327), .B(n18307), .Z(n18324) );
  INV_X1 U15512 ( .A(n18324), .ZN(n17403) );
  OAI21_X1 U15514 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18267), .A(
        n12363), .ZN(n18297) );
  INV_X1 U15515 ( .A(n18297), .ZN(n17381) );
  NOR2_X1 U15516 ( .A1(n17379), .A2(n10186), .ZN(n17366) );
  NOR2_X1 U15518 ( .A1(n17365), .A2(n10186), .ZN(n17358) );
  INV_X1 U15520 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17348) );
  INV_X1 U15521 ( .A(n12364), .ZN(n18226) );
  AOI21_X1 U15522 ( .B1(n17348), .B2(n18226), .A(n12365), .ZN(n18257) );
  NOR2_X1 U15523 ( .A1(n17339), .A2(n10186), .ZN(n17327) );
  NOR2_X1 U15524 ( .A1(n17326), .A2(n10186), .ZN(n17319) );
  INV_X1 U15525 ( .A(n12366), .ZN(n18187) );
  NOR2_X1 U15526 ( .A1(n10179), .A2(n18548), .ZN(n12367) );
  AOI21_X1 U15527 ( .B1(n18213), .B2(n18187), .A(n12367), .ZN(n18217) );
  NOR2_X1 U15528 ( .A1(n17318), .A2(n10186), .ZN(n17309) );
  NAND2_X1 U15529 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n12367), .ZN(
        n12369) );
  OAI21_X1 U15530 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n12367), .A(
        n12369), .ZN(n12368) );
  INV_X1 U15531 ( .A(n12368), .ZN(n18203) );
  NOR2_X1 U15533 ( .A1(n17308), .A2(n10186), .ZN(n17301) );
  NOR2_X1 U15534 ( .A1(n18184), .A2(n12369), .ZN(n12370) );
  AOI21_X1 U15535 ( .B1(n18184), .B2(n12369), .A(n12370), .ZN(n18194) );
  INV_X1 U15536 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12377) );
  INV_X1 U15537 ( .A(n12370), .ZN(n17112) );
  AOI21_X1 U15538 ( .B1(n12377), .B2(n17112), .A(n12371), .ZN(n17139) );
  INV_X1 U15539 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19538) );
  NAND3_X1 U15540 ( .A1(n17110), .A2(n19393), .A3(n19538), .ZN(n19401) );
  NOR2_X1 U15541 ( .A1(n19503), .A2(n19401), .ZN(n17591) );
  AOI211_X1 U15542 ( .C1(n9776), .C2(n17139), .A(n17284), .B(n19399), .ZN(
        n12386) );
  NOR3_X1 U15543 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17587) );
  NAND2_X1 U15544 ( .A1(n17587), .A2(n17906), .ZN(n17582) );
  NOR2_X1 U15545 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17582), .ZN(n17561) );
  INV_X1 U15546 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17553) );
  NAND2_X1 U15547 ( .A1(n17561), .A2(n17553), .ZN(n17552) );
  NOR2_X1 U15548 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17552), .ZN(n17533) );
  INV_X1 U15549 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17530) );
  NAND2_X1 U15550 ( .A1(n17533), .A2(n17530), .ZN(n17529) );
  NOR2_X1 U15551 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17529), .ZN(n17502) );
  INV_X1 U15552 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17854) );
  NAND2_X1 U15553 ( .A1(n17502), .A2(n17854), .ZN(n17491) );
  NOR2_X1 U15554 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17491), .ZN(n17490) );
  INV_X1 U15555 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17481) );
  NAND2_X1 U15556 ( .A1(n17490), .A2(n17481), .ZN(n17480) );
  NOR2_X1 U15557 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17480), .ZN(n17467) );
  INV_X1 U15558 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17454) );
  NAND2_X1 U15559 ( .A1(n17467), .A2(n17454), .ZN(n17452) );
  NOR2_X1 U15560 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17452), .ZN(n17438) );
  INV_X1 U15561 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17431) );
  NAND2_X1 U15562 ( .A1(n17438), .A2(n17431), .ZN(n17430) );
  NOR2_X1 U15563 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17430), .ZN(n17419) );
  INV_X1 U15564 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17412) );
  NAND2_X1 U15565 ( .A1(n17419), .A2(n17412), .ZN(n17410) );
  NOR2_X1 U15566 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17410), .ZN(n17399) );
  INV_X1 U15567 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17393) );
  NAND2_X1 U15568 ( .A1(n17399), .A2(n17393), .ZN(n17391) );
  NOR2_X1 U15569 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17391), .ZN(n17374) );
  INV_X1 U15570 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17703) );
  NAND2_X1 U15571 ( .A1(n17374), .A2(n17703), .ZN(n17369) );
  NOR2_X1 U15572 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17369), .ZN(n17356) );
  INV_X1 U15573 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17626) );
  NAND2_X1 U15574 ( .A1(n17356), .A2(n17626), .ZN(n17351) );
  NOR2_X1 U15575 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17351), .ZN(n17338) );
  INV_X1 U15576 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17624) );
  NAND2_X1 U15577 ( .A1(n17338), .A2(n17624), .ZN(n17332) );
  NOR2_X1 U15578 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17332), .ZN(n17317) );
  INV_X1 U15579 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17671) );
  NAND2_X1 U15580 ( .A1(n17317), .A2(n17671), .ZN(n17313) );
  NOR2_X1 U15581 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17313), .ZN(n17299) );
  INV_X1 U15582 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17659) );
  NOR2_X1 U15583 ( .A1(n17299), .A2(n17659), .ZN(n12374) );
  NAND2_X1 U15584 ( .A1(n19535), .A2(n19324), .ZN(n18123) );
  NAND2_X1 U15585 ( .A1(n19555), .A2(n17562), .ZN(n19553) );
  NAND2_X1 U15586 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18125), .ZN(n12373) );
  AOI211_X4 U15587 ( .C1(n19538), .C2(n19540), .A(n19553), .B(n12373), .ZN(
        n17616) );
  NAND2_X1 U15588 ( .A1(n17299), .A2(n17659), .ZN(n17274) );
  NAND2_X1 U15589 ( .A1(n17616), .A2(n17274), .ZN(n17296) );
  OR2_X1 U15590 ( .A1(n12374), .A2(n17296), .ZN(n12384) );
  NAND2_X1 U15591 ( .A1(n19393), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19259) );
  OR2_X1 U15592 ( .A1(n19396), .A2(n19259), .ZN(n19389) );
  NOR2_X2 U15593 ( .A1(n19492), .A2(n17604), .ZN(n17598) );
  INV_X1 U15594 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19475) );
  NAND3_X1 U15595 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(P3_REIP_REG_28__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n12376) );
  INV_X1 U15596 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19468) );
  INV_X1 U15597 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19465) );
  INV_X1 U15598 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19459) );
  INV_X1 U15599 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n21324) );
  INV_X1 U15600 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19445) );
  INV_X1 U15601 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n21135) );
  INV_X1 U15602 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19426) );
  INV_X1 U15603 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19423) );
  INV_X1 U15604 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19424) );
  NOR2_X1 U15605 ( .A1(n19423), .A2(n19424), .ZN(n17576) );
  INV_X1 U15606 ( .A(n17576), .ZN(n17599) );
  NOR2_X1 U15607 ( .A1(n19426), .A2(n17599), .ZN(n17573) );
  NAND3_X1 U15608 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .A3(n17573), .ZN(n17485) );
  NAND3_X1 U15609 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n17486) );
  INV_X1 U15610 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19439) );
  INV_X1 U15611 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19437) );
  NOR2_X1 U15612 ( .A1(n19439), .A2(n19437), .ZN(n17472) );
  INV_X1 U15613 ( .A(n17472), .ZN(n17496) );
  NOR4_X1 U15614 ( .A1(n21135), .A2(n17485), .A3(n17486), .A4(n17496), .ZN(
        n17448) );
  NAND2_X1 U15615 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17448), .ZN(n17440) );
  NOR3_X1 U15616 ( .A1(n21324), .A2(n19445), .A3(n17440), .ZN(n17376) );
  NAND3_X1 U15617 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(P3_REIP_REG_17__SCAN_IN), 
        .A3(P3_REIP_REG_16__SCAN_IN), .ZN(n17377) );
  INV_X1 U15618 ( .A(n17377), .ZN(n12375) );
  INV_X1 U15619 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19455) );
  INV_X1 U15620 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19453) );
  INV_X1 U15621 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19451) );
  NOR3_X1 U15622 ( .A1(n19455), .A2(n19453), .A3(n19451), .ZN(n17378) );
  NAND4_X1 U15623 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n17376), .A3(n12375), 
        .A4(n17378), .ZN(n17359) );
  NOR2_X1 U15624 ( .A1(n19459), .A2(n17359), .ZN(n17345) );
  AND2_X1 U15625 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17345), .ZN(n17337) );
  NAND2_X1 U15626 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17337), .ZN(n17316) );
  NOR3_X1 U15627 ( .A1(n19468), .A2(n19465), .A3(n17316), .ZN(n12378) );
  NAND2_X1 U15628 ( .A1(n12378), .A2(n17620), .ZN(n17297) );
  INV_X1 U15629 ( .A(n19540), .ZN(n19411) );
  AOI211_X1 U15630 ( .C1(n19539), .C2(n19537), .A(n19411), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n12379) );
  INV_X1 U15631 ( .A(n12379), .ZN(n19385) );
  NOR2_X1 U15632 ( .A1(n17600), .A2(n17604), .ZN(n17388) );
  OAI21_X1 U15633 ( .B1(n12376), .B2(n17297), .A(n17619), .ZN(n17287) );
  OAI22_X1 U15634 ( .A1(n12377), .A2(n17605), .B1(n19475), .B2(n17287), .ZN(
        n12383) );
  AND2_X1 U15635 ( .A1(n17600), .A2(n12378), .ZN(n17298) );
  NAND4_X1 U15636 ( .A1(n17298), .A2(P3_REIP_REG_28__SCAN_IN), .A3(
        P3_REIP_REG_27__SCAN_IN), .A4(n19475), .ZN(n12381) );
  AOI211_X4 U15637 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18125), .A(n12379), .B(
        n19553), .ZN(n17617) );
  NAND2_X1 U15638 ( .A1(n17617), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n12380) );
  NAND2_X1 U15639 ( .A1(n12381), .A2(n12380), .ZN(n12382) );
  AOI21_X1 U15640 ( .B1(n12406), .B2(n9719), .A(n11528), .ZN(n12413) );
  OAI21_X2 U15641 ( .B1(n12389), .B2(n12388), .A(n12387), .ZN(n16894) );
  NOR2_X1 U15642 ( .A1(n16894), .A2(n16307), .ZN(n12393) );
  NAND2_X1 U15643 ( .A1(n19825), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12407) );
  NAND2_X1 U15644 ( .A1(n19837), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12390) );
  OAI211_X1 U15645 ( .C1(n12391), .C2(n19840), .A(n12407), .B(n12390), .ZN(
        n12392) );
  AOI211_X1 U15646 ( .C1(n12413), .C2(n11531), .A(n12393), .B(n12392), .ZN(
        n12399) );
  NAND2_X1 U15647 ( .A1(n12395), .A2(n12394), .ZN(n12397) );
  NAND2_X1 U15648 ( .A1(n12399), .A2(n12398), .ZN(P2_U2985) );
  NOR2_X1 U15649 ( .A1(n12400), .A2(n12406), .ZN(n12412) );
  XOR2_X1 U15650 ( .A(n12402), .B(n12401), .Z(n16895) );
  AOI211_X1 U15651 ( .C1(n12406), .C2(n12405), .A(n12404), .B(n12403), .ZN(
        n12409) );
  INV_X1 U15652 ( .A(n12407), .ZN(n12408) );
  AOI211_X1 U15653 ( .C1(n16895), .C2(n19854), .A(n12409), .B(n12408), .ZN(
        n12410) );
  OAI21_X1 U15654 ( .B1(n16894), .B2(n19870), .A(n12410), .ZN(n12411) );
  AOI211_X1 U15655 ( .C1(n12413), .C2(n11551), .A(n12412), .B(n12411), .ZN(
        n12415) );
  NAND2_X1 U15656 ( .A1(n12415), .A2(n12414), .ZN(P2_U3017) );
  NOR4_X1 U15657 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12419) );
  NOR4_X1 U15658 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12418) );
  NOR4_X1 U15659 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12417) );
  NOR4_X1 U15660 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12416) );
  AND4_X1 U15661 ( .A1(n12419), .A2(n12418), .A3(n12417), .A4(n12416), .ZN(
        n12424) );
  NOR4_X1 U15662 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12422) );
  NOR4_X1 U15663 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12421) );
  NOR4_X1 U15664 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12420) );
  INV_X1 U15665 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20954) );
  AND4_X1 U15666 ( .A1(n12422), .A2(n12421), .A3(n12420), .A4(n20954), .ZN(
        n12423) );
  NAND2_X1 U15667 ( .A1(n12424), .A2(n12423), .ZN(n12425) );
  AND2_X2 U15668 ( .A1(n12425), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15109)
         );
  INV_X1 U15669 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21064) );
  NOR3_X1 U15670 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21064), .ZN(n12427) );
  NOR4_X1 U15671 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12426) );
  NAND4_X1 U15672 ( .A1(n15109), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12427), .A4(
        n12426), .ZN(U214) );
  INV_X1 U15673 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20493) );
  NOR2_X1 U15674 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n20493), .ZN(n12429) );
  NOR4_X1 U15675 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12428) );
  INV_X1 U15676 ( .A(P2_BE_N_REG_2__SCAN_IN), .ZN(n21240) );
  NAND4_X1 U15677 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n12429), .A3(n12428), .A4(
        n21240), .ZN(n12430) );
  NOR2_X1 U15678 ( .A1(n13223), .A2(n12430), .ZN(n17167) );
  NAND2_X1 U15679 ( .A1(n17167), .A2(U214), .ZN(U212) );
  NOR2_X1 U15680 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12430), .ZN(n17239)
         );
  NOR2_X1 U15681 ( .A1(n9712), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12431) );
  NAND2_X1 U15682 ( .A1(n16622), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12433) );
  XNOR2_X1 U15683 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12528) );
  INV_X1 U15684 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12829) );
  AOI222_X1 U15685 ( .A1(n12526), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n12526), .B2(n12829), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n12829), .ZN(n12612) );
  AND2_X4 U15686 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14740) );
  AND2_X2 U15687 ( .A1(n12441), .A2(n14740), .ZN(n15015) );
  AND2_X2 U15688 ( .A1(n12441), .A2(n12440), .ZN(n14908) );
  AOI22_X1 U15689 ( .A1(n15015), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14908), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12438) );
  AND2_X2 U15690 ( .A1(n12439), .A2(n13533), .ZN(n14948) );
  AOI22_X1 U15691 ( .A1(n9708), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14948), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12437) );
  AND2_X2 U15692 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12870) );
  AND2_X4 U15693 ( .A1(n12870), .A2(n14740), .ZN(n15075) );
  AOI22_X1 U15694 ( .A1(n14929), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15696 ( .A1(n12892), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13960), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12445) );
  AND2_X2 U15697 ( .A1(n12869), .A2(n13533), .ZN(n13700) );
  AOI22_X1 U15698 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13700), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15699 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12443) );
  NAND2_X1 U15700 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12449) );
  NAND2_X1 U15701 ( .A1(n14908), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12448) );
  NAND2_X1 U15702 ( .A1(n12555), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12447) );
  NAND2_X1 U15703 ( .A1(n9710), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12446) );
  NAND2_X1 U15704 ( .A1(n15040), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12453) );
  NAND2_X1 U15705 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12452) );
  NAND2_X1 U15706 ( .A1(n14948), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12451) );
  NAND2_X1 U15707 ( .A1(n14930), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12450) );
  NAND2_X1 U15708 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12457) );
  NAND2_X1 U15709 ( .A1(n15073), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12455) );
  NAND2_X1 U15710 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12454) );
  NAND2_X1 U15711 ( .A1(n15075), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12460) );
  NAND2_X1 U15712 ( .A1(n14929), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12459) );
  NAND3_X1 U15713 ( .A1(n12460), .A2(n12459), .A3(n12458), .ZN(n12461) );
  NAND4_X4 U15714 ( .A1(n12465), .A2(n12464), .A3(n12463), .A4(n12462), .ZN(
        n13832) );
  NAND2_X1 U15715 ( .A1(n13547), .A2(n13832), .ZN(n12486) );
  NAND2_X1 U15716 ( .A1(n12612), .A2(n13972), .ZN(n12540) );
  NAND2_X1 U15717 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12469) );
  NAND2_X1 U15718 ( .A1(n14908), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12468) );
  INV_X1 U15719 ( .A(n12555), .ZN(n14344) );
  NAND2_X1 U15720 ( .A1(n12555), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12467) );
  NAND2_X1 U15721 ( .A1(n13960), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12466) );
  NAND2_X1 U15722 ( .A1(n15082), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12473) );
  NAND2_X1 U15723 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12472) );
  NAND2_X1 U15724 ( .A1(n14948), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12471) );
  NAND2_X1 U15725 ( .A1(n14930), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12470) );
  NAND2_X1 U15726 ( .A1(n12892), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12477) );
  NAND2_X1 U15727 ( .A1(n15059), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12476) );
  NAND2_X1 U15728 ( .A1(n15053), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12475) );
  NAND2_X1 U15729 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12474) );
  NAND2_X1 U15730 ( .A1(n14947), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12481) );
  NAND2_X1 U15731 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12480) );
  NAND2_X1 U15732 ( .A1(n14929), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12479) );
  NAND2_X1 U15733 ( .A1(n15075), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12478) );
  NAND4_X4 U15734 ( .A1(n12485), .A2(n12484), .A3(n12483), .A4(n12482), .ZN(
        n13587) );
  NAND2_X1 U15735 ( .A1(n12486), .A2(n13587), .ZN(n12497) );
  AOI22_X1 U15736 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9710), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15737 ( .A1(n14908), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15738 ( .A1(n12892), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15059), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15739 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12487) );
  NAND4_X1 U15740 ( .A1(n12490), .A2(n12489), .A3(n12488), .A4(n12487), .ZN(
        n12496) );
  AOI22_X1 U15741 ( .A1(n15015), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12573), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U15742 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15743 ( .A1(n14948), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13700), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15744 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9701), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12491) );
  NAND4_X1 U15745 ( .A1(n12494), .A2(n12493), .A3(n12492), .A4(n12491), .ZN(
        n12495) );
  NAND2_X1 U15746 ( .A1(n12497), .A2(n15107), .ZN(n12498) );
  NAND2_X1 U15747 ( .A1(n12498), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12501) );
  NAND2_X1 U15748 ( .A1(n12501), .A2(n13587), .ZN(n12534) );
  XNOR2_X1 U15749 ( .A(n12499), .B(n12504), .ZN(n12609) );
  NAND2_X1 U15750 ( .A1(n12534), .A2(n12609), .ZN(n12512) );
  NAND2_X1 U15751 ( .A1(n13971), .A2(n12609), .ZN(n12500) );
  NAND2_X1 U15752 ( .A1(n12501), .A2(n12500), .ZN(n12511) );
  NOR2_X1 U15753 ( .A1(n12853), .A2(n12975), .ZN(n12505) );
  NAND2_X1 U15754 ( .A1(n12764), .A2(n15107), .ZN(n12502) );
  NAND2_X1 U15755 ( .A1(n15286), .A2(n12502), .ZN(n12522) );
  AND2_X1 U15756 ( .A1(n12777), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12503) );
  NOR2_X1 U15757 ( .A1(n12504), .A2(n12503), .ZN(n12506) );
  OAI211_X1 U15758 ( .C1(n12505), .C2(n12522), .A(n13972), .B(n12506), .ZN(
        n12509) );
  INV_X1 U15759 ( .A(n12506), .ZN(n12507) );
  NAND3_X1 U15760 ( .A1(n13971), .A2(n14530), .A3(n12507), .ZN(n12508) );
  NAND2_X1 U15761 ( .A1(n12509), .A2(n12508), .ZN(n12510) );
  OAI21_X1 U15762 ( .B1(n12512), .B2(n12511), .A(n12510), .ZN(n12514) );
  NAND2_X1 U15763 ( .A1(n12512), .A2(n12511), .ZN(n12513) );
  NAND2_X1 U15764 ( .A1(n12514), .A2(n12513), .ZN(n12520) );
  XNOR2_X1 U15765 ( .A(n12434), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12515) );
  XNOR2_X1 U15766 ( .A(n12516), .B(n12515), .ZN(n12610) );
  INV_X1 U15767 ( .A(n12610), .ZN(n12518) );
  NAND2_X1 U15768 ( .A1(n13972), .A2(n12518), .ZN(n12521) );
  INV_X1 U15769 ( .A(n12522), .ZN(n12517) );
  OAI211_X1 U15770 ( .C1(n12518), .C2(n14103), .A(n12521), .B(n12517), .ZN(
        n12519) );
  NAND2_X1 U15771 ( .A1(n12520), .A2(n12519), .ZN(n12525) );
  INV_X1 U15772 ( .A(n12521), .ZN(n12523) );
  NAND2_X1 U15773 ( .A1(n12523), .A2(n12522), .ZN(n12524) );
  NAND2_X1 U15774 ( .A1(n12525), .A2(n12524), .ZN(n12536) );
  AND2_X1 U15775 ( .A1(n12829), .A2(n12526), .ZN(n12527) );
  NAND2_X1 U15776 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12527), .ZN(
        n12611) );
  NOR2_X1 U15777 ( .A1(n12529), .A2(n12528), .ZN(n12530) );
  OR2_X1 U15778 ( .A1(n12531), .A2(n12530), .ZN(n12608) );
  INV_X1 U15779 ( .A(n12608), .ZN(n12533) );
  AND2_X1 U15780 ( .A1(n12611), .A2(n12533), .ZN(n12532) );
  AOI22_X1 U15781 ( .A1(n12536), .A2(n12532), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n9922), .ZN(n12538) );
  OAI22_X1 U15782 ( .A1(n12611), .A2(n12534), .B1(n12533), .B2(n14401), .ZN(
        n12535) );
  OAI21_X1 U15783 ( .B1(n12536), .B2(n12535), .A(n13971), .ZN(n12537) );
  NOR2_X1 U15784 ( .A1(n14103), .A2(n14401), .ZN(n12541) );
  NAND2_X1 U15785 ( .A1(n12612), .A2(n12541), .ZN(n12542) );
  AOI22_X1 U15786 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9709), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15787 ( .A1(n14908), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15788 ( .A1(n14948), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U15789 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U15790 ( .A1(n12892), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15791 ( .A1(n15015), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15059), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15792 ( .A1(n12573), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13700), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15793 ( .A1(n14947), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9702), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12548) );
  NAND2_X2 U15794 ( .A1(n12554), .A2(n12780), .ZN(n12759) );
  INV_X1 U15795 ( .A(n12759), .ZN(n12553) );
  NAND2_X1 U15796 ( .A1(n12772), .A2(n12590), .ZN(n12918) );
  AOI22_X1 U15797 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14908), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U15798 ( .A1(n9707), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14948), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15799 ( .A1(n12555), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15800 ( .A1(n15015), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12556) );
  NAND4_X1 U15801 ( .A1(n12559), .A2(n12558), .A3(n12557), .A4(n12556), .ZN(
        n12566) );
  AOI22_X1 U15802 ( .A1(n12892), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15059), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15803 ( .A1(n13960), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15804 ( .A1(n14947), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12583), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U15805 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12561) );
  NAND4_X1 U15806 ( .A1(n12564), .A2(n12563), .A3(n12562), .A4(n12561), .ZN(
        n12565) );
  OR2_X4 U15807 ( .A1(n12566), .A2(n12565), .ZN(n13577) );
  NAND2_X1 U15808 ( .A1(n12918), .A2(n13577), .ZN(n12758) );
  INV_X1 U15809 ( .A(n12758), .ZN(n12567) );
  AOI22_X1 U15810 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14908), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15811 ( .A1(n12892), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13960), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12571) );
  AOI22_X1 U15812 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U15813 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15814 ( .A1(n15015), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15040), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U15815 ( .A1(n14929), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U15816 ( .A1(n14948), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U15817 ( .A1(n12892), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15059), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U15818 ( .A1(n14908), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15819 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13960), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15820 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12579) );
  NAND4_X1 U15821 ( .A1(n12582), .A2(n12581), .A3(n12580), .A4(n12579), .ZN(
        n12589) );
  AOI22_X1 U15822 ( .A1(n15015), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9708), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12587) );
  CLKBUF_X3 U15823 ( .A(n12583), .Z(n15087) );
  AOI22_X1 U15824 ( .A1(n14947), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15825 ( .A1(n14948), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15826 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12584) );
  NAND4_X1 U15827 ( .A1(n12587), .A2(n12586), .A3(n12585), .A4(n12584), .ZN(
        n12588) );
  INV_X1 U15828 ( .A(n13077), .ZN(n20508) );
  NOR2_X1 U15829 ( .A1(n12767), .A2(n20508), .ZN(n12592) );
  INV_X1 U15830 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20951) );
  NAND2_X1 U15831 ( .A1(n20951), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20942) );
  INV_X1 U15832 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n12593) );
  NAND2_X1 U15833 ( .A1(n12593), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n12594) );
  AND2_X1 U15834 ( .A1(n20942), .A2(n12594), .ZN(n12754) );
  OR2_X1 U15835 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n12754), .ZN(n16666) );
  OR3_X1 U15836 ( .A1(n12831), .A2(n13587), .A3(n16666), .ZN(n12603) );
  NAND2_X1 U15837 ( .A1(n15107), .A2(n13564), .ZN(n12595) );
  OR2_X4 U15838 ( .A1(n12759), .A2(n12596), .ZN(n12761) );
  AOI21_X2 U15839 ( .B1(n12761), .B2(n13571), .A(n12597), .ZN(n12598) );
  NOR2_X1 U15840 ( .A1(n12766), .A2(n12764), .ZN(n14742) );
  INV_X1 U15841 ( .A(n16666), .ZN(n13068) );
  AND2_X1 U15842 ( .A1(n14742), .A2(n13068), .ZN(n12601) );
  NAND2_X1 U15843 ( .A1(n16614), .A2(n12601), .ZN(n12821) );
  OR2_X1 U15844 ( .A1(n12821), .A2(n20508), .ZN(n12602) );
  NAND2_X1 U15845 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16878) );
  NOR2_X1 U15846 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16878), .ZN(n20647) );
  AND2_X1 U15847 ( .A1(n20646), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OAI21_X1 U15848 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n20133), .A(n12629), 
        .ZN(n12605) );
  AOI21_X1 U15849 ( .B1(P2_MEMORYFETCH_REG_SCAN_IN), .B2(n19688), .A(n12605), 
        .ZN(n12604) );
  INV_X1 U15850 ( .A(n12604), .ZN(P2_U2814) );
  NOR2_X1 U15851 ( .A1(P2_READREQUEST_REG_SCAN_IN), .A2(n12605), .ZN(n12607)
         );
  AOI22_X1 U15852 ( .A1(n12607), .A2(n19688), .B1(n12606), .B2(n19557), .ZN(
        P2_U3612) );
  NOR3_X1 U15853 ( .A1(n12610), .A2(n12609), .A3(n12608), .ZN(n12613) );
  OAI21_X1 U15854 ( .B1(n12613), .B2(n12612), .A(n12611), .ZN(n15281) );
  INV_X1 U15855 ( .A(n12766), .ZN(n12614) );
  NAND2_X1 U15856 ( .A1(n15282), .A2(n13077), .ZN(n12668) );
  NOR2_X1 U15857 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20866) );
  NAND2_X1 U15858 ( .A1(n15926), .A2(n21133), .ZN(n20511) );
  INV_X1 U15859 ( .A(n20511), .ZN(n12669) );
  AOI21_X1 U15860 ( .B1(n12668), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n12669), 
        .ZN(n12615) );
  NAND2_X1 U15861 ( .A1(n12831), .A2(n12615), .ZN(P1_U2801) );
  OR2_X1 U15862 ( .A1(n12616), .A2(n20312), .ZN(n13446) );
  INV_X1 U15863 ( .A(n20373), .ZN(n20385) );
  NAND2_X1 U15864 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20484) );
  OR2_X1 U15865 ( .A1(n20484), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19793) );
  INV_X1 U15866 ( .A(n19557), .ZN(n12617) );
  OAI21_X1 U15867 ( .B1(n20385), .B2(n19793), .A(n12617), .ZN(n12618) );
  AOI21_X1 U15868 ( .B1(n20101), .B2(n13446), .A(n12618), .ZN(n12627) );
  NOR2_X1 U15869 ( .A1(n12711), .A2(n13429), .ZN(n12621) );
  AOI21_X1 U15870 ( .B1(n20312), .B2(n11007), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n17096) );
  AOI21_X1 U15871 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20373), .A(n17096), 
        .ZN(n12619) );
  AOI21_X1 U15872 ( .B1(n12621), .B2(n12620), .A(n12619), .ZN(n12625) );
  INV_X1 U15873 ( .A(n12711), .ZN(n20380) );
  INV_X1 U15874 ( .A(n12622), .ZN(n12623) );
  OAI21_X1 U15875 ( .B1(n20380), .B2(n21150), .A(n12623), .ZN(n12624) );
  AOI21_X1 U15876 ( .B1(n12625), .B2(n12624), .A(n12627), .ZN(n12626) );
  AOI21_X1 U15877 ( .B1(n12627), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .A(n12626), .ZN(n12628) );
  INV_X1 U15878 ( .A(n12628), .ZN(P2_U3610) );
  INV_X1 U15879 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n12633) );
  INV_X1 U15880 ( .A(n12629), .ZN(n12630) );
  AOI21_X2 U15881 ( .B1(n12630), .B2(n20373), .A(n19821), .ZN(n19822) );
  NAND2_X1 U15882 ( .A1(n19822), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U15883 ( .A1(n13225), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n12694), .ZN(n19735) );
  INV_X1 U15884 ( .A(n19735), .ZN(n12631) );
  NAND2_X1 U15885 ( .A1(n19819), .A2(n12631), .ZN(n12650) );
  OAI211_X1 U15886 ( .C1(n12708), .C2(n12633), .A(n12632), .B(n12650), .ZN(
        P2_U2977) );
  INV_X1 U15887 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n12636) );
  NAND2_X1 U15888 ( .A1(n19822), .A2(P2_LWORD_REG_3__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U15889 ( .A1(n13225), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13223), .ZN(n19886) );
  INV_X1 U15890 ( .A(n19886), .ZN(n12634) );
  NAND2_X1 U15891 ( .A1(n19819), .A2(n12634), .ZN(n12660) );
  OAI211_X1 U15892 ( .C1(n12636), .C2(n12708), .A(n12635), .B(n12660), .ZN(
        P2_U2970) );
  INV_X1 U15893 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16111) );
  NAND2_X1 U15894 ( .A1(n19822), .A2(P2_UWORD_REG_7__SCAN_IN), .ZN(n12638) );
  AOI22_X1 U15895 ( .A1(n13225), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n12694), .ZN(n19908) );
  INV_X1 U15896 ( .A(n19908), .ZN(n12637) );
  NAND2_X1 U15897 ( .A1(n19819), .A2(n12637), .ZN(n12663) );
  OAI211_X1 U15898 ( .C1(n12708), .C2(n16111), .A(n12638), .B(n12663), .ZN(
        P2_U2959) );
  INV_X1 U15899 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n12725) );
  NAND2_X1 U15900 ( .A1(n19822), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12639) );
  INV_X1 U15901 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17204) );
  INV_X1 U15902 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n18162) );
  AOI22_X1 U15903 ( .A1(n13225), .A2(n17204), .B1(n18162), .B2(n13223), .ZN(
        n19740) );
  NAND2_X1 U15904 ( .A1(n19819), .A2(n19740), .ZN(n12645) );
  OAI211_X1 U15905 ( .C1(n12725), .C2(n12708), .A(n12639), .B(n12645), .ZN(
        P2_U2960) );
  INV_X1 U15906 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19795) );
  NAND2_X1 U15907 ( .A1(n19822), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12642) );
  NAND2_X1 U15908 ( .A1(n13223), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12641) );
  INV_X1 U15909 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n17198) );
  OR2_X1 U15910 ( .A1(n13223), .A2(n17198), .ZN(n12640) );
  NAND2_X1 U15911 ( .A1(n12641), .A2(n12640), .ZN(n19730) );
  NAND2_X1 U15912 ( .A1(n19819), .A2(n19730), .ZN(n12643) );
  OAI211_X1 U15913 ( .C1(n19795), .C2(n12708), .A(n12642), .B(n12643), .ZN(
        P2_U2979) );
  INV_X1 U15914 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n12715) );
  NAND2_X1 U15915 ( .A1(n19822), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12644) );
  OAI211_X1 U15916 ( .C1(n12715), .C2(n12708), .A(n12644), .B(n12643), .ZN(
        P2_U2964) );
  INV_X1 U15917 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19801) );
  NAND2_X1 U15918 ( .A1(n19822), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12646) );
  OAI211_X1 U15919 ( .C1(n19801), .C2(n12708), .A(n12646), .B(n12645), .ZN(
        P2_U2975) );
  INV_X1 U15920 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n12649) );
  NAND2_X1 U15921 ( .A1(n19822), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15922 ( .A1(n13225), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n12694), .ZN(n19891) );
  INV_X1 U15923 ( .A(n19891), .ZN(n12647) );
  NAND2_X1 U15924 ( .A1(n19819), .A2(n12647), .ZN(n12652) );
  OAI211_X1 U15925 ( .C1(n12649), .C2(n12708), .A(n12648), .B(n12652), .ZN(
        P2_U2971) );
  INV_X1 U15926 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n16096) );
  NAND2_X1 U15927 ( .A1(n19822), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12651) );
  OAI211_X1 U15928 ( .C1(n12708), .C2(n16096), .A(n12651), .B(n12650), .ZN(
        P2_U2962) );
  INV_X1 U15929 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U15930 ( .A1(n19822), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n12653) );
  OAI211_X1 U15931 ( .C1(n12708), .C2(n12654), .A(n12653), .B(n12652), .ZN(
        P2_U2956) );
  INV_X1 U15932 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n12657) );
  NAND2_X1 U15933 ( .A1(n19822), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U15934 ( .A1(n13225), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n13223), .ZN(n19733) );
  INV_X1 U15935 ( .A(n19733), .ZN(n12655) );
  NAND2_X1 U15936 ( .A1(n19819), .A2(n12655), .ZN(n12666) );
  OAI211_X1 U15937 ( .C1(n12708), .C2(n12657), .A(n12656), .B(n12666), .ZN(
        P2_U2978) );
  INV_X1 U15938 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n16077) );
  NAND2_X1 U15939 ( .A1(n19822), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U15940 ( .A1(n13225), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n12694), .ZN(n19727) );
  INV_X1 U15941 ( .A(n19727), .ZN(n12658) );
  NAND2_X1 U15942 ( .A1(n19819), .A2(n12658), .ZN(n12704) );
  OAI211_X1 U15943 ( .C1(n12708), .C2(n16077), .A(n12659), .B(n12704), .ZN(
        P2_U2965) );
  INV_X1 U15944 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n12662) );
  NAND2_X1 U15945 ( .A1(n19822), .A2(P2_UWORD_REG_3__SCAN_IN), .ZN(n12661) );
  OAI211_X1 U15946 ( .C1(n12708), .C2(n12662), .A(n12661), .B(n12660), .ZN(
        P2_U2955) );
  INV_X1 U15947 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n12665) );
  NAND2_X1 U15948 ( .A1(n19822), .A2(P2_LWORD_REG_7__SCAN_IN), .ZN(n12664) );
  OAI211_X1 U15949 ( .C1(n12708), .C2(n12665), .A(n12664), .B(n12663), .ZN(
        P2_U2974) );
  INV_X1 U15950 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n21132) );
  NAND2_X1 U15951 ( .A1(n19822), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12667) );
  OAI211_X1 U15952 ( .C1(n12708), .C2(n21132), .A(n12667), .B(n12666), .ZN(
        P2_U2963) );
  NAND2_X2 U15953 ( .A1(n13587), .A2(n13571), .ZN(n15147) );
  AND2_X1 U15954 ( .A1(n15286), .A2(n15129), .ZN(n12784) );
  INV_X1 U15955 ( .A(n21026), .ZN(n12671) );
  OAI21_X1 U15956 ( .B1(n12669), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n12671), 
        .ZN(n12670) );
  OAI21_X1 U15957 ( .B1(n12784), .B2(n12671), .A(n12670), .ZN(P1_U3487) );
  INV_X1 U15958 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n12673) );
  INV_X1 U15959 ( .A(n19819), .ZN(n12706) );
  AOI22_X1 U15960 ( .A1(n13225), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n13223), .ZN(n19737) );
  NOR2_X1 U15961 ( .A1(n12706), .A2(n19737), .ZN(n12674) );
  AOI21_X1 U15962 ( .B1(n19821), .B2(P2_EAX_REG_25__SCAN_IN), .A(n12674), .ZN(
        n12672) );
  OAI21_X1 U15963 ( .B1(n12707), .B2(n12673), .A(n12672), .ZN(P2_U2961) );
  INV_X1 U15964 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n12676) );
  AOI21_X1 U15965 ( .B1(n19821), .B2(P2_EAX_REG_9__SCAN_IN), .A(n12674), .ZN(
        n12675) );
  OAI21_X1 U15966 ( .B1(n12707), .B2(n12676), .A(n12675), .ZN(P2_U2976) );
  INV_X1 U15967 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n12678) );
  AOI22_X1 U15968 ( .A1(n13225), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n12694), .ZN(n14335) );
  NOR2_X1 U15969 ( .A1(n12706), .A2(n14335), .ZN(n12683) );
  AOI21_X1 U15970 ( .B1(n19821), .B2(P2_EAX_REG_1__SCAN_IN), .A(n12683), .ZN(
        n12677) );
  OAI21_X1 U15971 ( .B1(n12707), .B2(n12678), .A(n12677), .ZN(P2_U2968) );
  INV_X1 U15972 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U15973 ( .A1(n13225), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13223), .ZN(n19881) );
  NOR2_X1 U15974 ( .A1(n12706), .A2(n19881), .ZN(n12691) );
  AOI21_X1 U15975 ( .B1(n19821), .B2(P2_EAX_REG_18__SCAN_IN), .A(n12691), .ZN(
        n12679) );
  OAI21_X1 U15976 ( .B1(n12707), .B2(n12680), .A(n12679), .ZN(P2_U2954) );
  INV_X1 U15977 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U15978 ( .A1(n13225), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n12694), .ZN(n19897) );
  NOR2_X1 U15979 ( .A1(n12706), .A2(n19897), .ZN(n12688) );
  AOI21_X1 U15980 ( .B1(n19821), .B2(P2_EAX_REG_22__SCAN_IN), .A(n12688), .ZN(
        n12681) );
  OAI21_X1 U15981 ( .B1(n12707), .B2(n12682), .A(n12681), .ZN(P2_U2958) );
  INV_X1 U15982 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n12685) );
  AOI21_X1 U15983 ( .B1(n19821), .B2(P2_EAX_REG_17__SCAN_IN), .A(n12683), .ZN(
        n12684) );
  OAI21_X1 U15984 ( .B1(n12707), .B2(n12685), .A(n12684), .ZN(P2_U2953) );
  INV_X1 U15985 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n12687) );
  INV_X1 U15986 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n21094) );
  INV_X1 U15987 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21293) );
  OAI22_X1 U15988 ( .A1(n12694), .A2(n21094), .B1(n21293), .B2(n13225), .ZN(
        n19747) );
  INV_X1 U15989 ( .A(n19747), .ZN(n16132) );
  NOR2_X1 U15990 ( .A1(n12706), .A2(n16132), .ZN(n12697) );
  AOI21_X1 U15991 ( .B1(n19821), .B2(P2_EAX_REG_5__SCAN_IN), .A(n12697), .ZN(
        n12686) );
  OAI21_X1 U15992 ( .B1(n12707), .B2(n12687), .A(n12686), .ZN(P2_U2972) );
  INV_X1 U15993 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n12690) );
  AOI21_X1 U15994 ( .B1(n19821), .B2(P2_EAX_REG_6__SCAN_IN), .A(n12688), .ZN(
        n12689) );
  OAI21_X1 U15995 ( .B1(n12707), .B2(n12690), .A(n12689), .ZN(P2_U2973) );
  INV_X1 U15996 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n12693) );
  AOI21_X1 U15997 ( .B1(n19821), .B2(P2_EAX_REG_2__SCAN_IN), .A(n12691), .ZN(
        n12692) );
  OAI21_X1 U15998 ( .B1(n12707), .B2(n12693), .A(n12692), .ZN(P2_U2969) );
  INV_X1 U15999 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U16000 ( .A1(n13225), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n12694), .ZN(n19780) );
  NOR2_X1 U16001 ( .A1(n12706), .A2(n19780), .ZN(n12700) );
  AOI21_X1 U16002 ( .B1(n19821), .B2(P2_EAX_REG_16__SCAN_IN), .A(n12700), .ZN(
        n12695) );
  OAI21_X1 U16003 ( .B1(n12707), .B2(n12696), .A(n12695), .ZN(P2_U2952) );
  INV_X1 U16004 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n12699) );
  AOI21_X1 U16005 ( .B1(n19821), .B2(P2_EAX_REG_21__SCAN_IN), .A(n12697), .ZN(
        n12698) );
  OAI21_X1 U16006 ( .B1(n12707), .B2(n12699), .A(n12698), .ZN(P2_U2957) );
  INV_X1 U16007 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12702) );
  AOI21_X1 U16008 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n19821), .A(n12700), .ZN(
        n12701) );
  OAI21_X1 U16009 ( .B1(n12707), .B2(n12702), .A(n12701), .ZN(P2_U2967) );
  INV_X1 U16010 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n12705) );
  NAND2_X1 U16011 ( .A1(n19821), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n12703) );
  OAI211_X1 U16012 ( .C1(n12707), .C2(n12705), .A(n12704), .B(n12703), .ZN(
        P2_U2980) );
  INV_X1 U16013 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19787) );
  INV_X1 U16014 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n19786) );
  AOI22_X1 U16015 ( .A1(n13225), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13223), .ZN(n19722) );
  OAI222_X1 U16016 ( .A1(n12708), .A2(n19787), .B1(n12707), .B2(n19786), .C1(
        n12706), .C2(n19722), .ZN(P2_U2982) );
  OAI21_X1 U16017 ( .B1(n12710), .B2(n12709), .A(n12708), .ZN(n12712) );
  OR2_X1 U16018 ( .A1(n19816), .A2(n12713), .ZN(n19782) );
  INV_X2 U16019 ( .A(n19793), .ZN(n19814) );
  NAND2_X1 U16020 ( .A1(n19816), .A2(n19793), .ZN(n19791) );
  INV_X2 U16021 ( .A(n19791), .ZN(n19813) );
  AOI22_X1 U16022 ( .A1(n19814), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12714) );
  OAI21_X1 U16023 ( .B1(n12715), .B2(n19782), .A(n12714), .ZN(P2_U2923) );
  INV_X1 U16024 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14181) );
  AOI22_X1 U16025 ( .A1(n19814), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12716) );
  OAI21_X1 U16026 ( .B1(n14181), .B2(n19782), .A(n12716), .ZN(P2_U2935) );
  INV_X1 U16027 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14334) );
  AOI22_X1 U16028 ( .A1(n19814), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12717) );
  OAI21_X1 U16029 ( .B1(n14334), .B2(n19782), .A(n12717), .ZN(P2_U2934) );
  AOI22_X1 U16030 ( .A1(n19814), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12718) );
  OAI21_X1 U16031 ( .B1(n12654), .B2(n19782), .A(n12718), .ZN(P2_U2931) );
  AOI22_X1 U16032 ( .A1(n19814), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12719) );
  OAI21_X1 U16033 ( .B1(n12662), .B2(n19782), .A(n12719), .ZN(P2_U2932) );
  INV_X1 U16034 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n21238) );
  AOI22_X1 U16035 ( .A1(n19814), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12720) );
  OAI21_X1 U16036 ( .B1(n21238), .B2(n19782), .A(n12720), .ZN(P2_U2933) );
  AOI22_X1 U16037 ( .A1(n19814), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12721) );
  OAI21_X1 U16038 ( .B1(n16077), .B2(n19782), .A(n12721), .ZN(P2_U2922) );
  AOI22_X1 U16039 ( .A1(n19814), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12722) );
  OAI21_X1 U16040 ( .B1(n16096), .B2(n19782), .A(n12722), .ZN(P2_U2925) );
  AOI22_X1 U16041 ( .A1(n19814), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12723) );
  OAI21_X1 U16042 ( .B1(n21132), .B2(n19782), .A(n12723), .ZN(P2_U2924) );
  AOI22_X1 U16043 ( .A1(n19814), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12724) );
  OAI21_X1 U16044 ( .B1(n12725), .B2(n19782), .A(n12724), .ZN(P2_U2927) );
  INV_X1 U16045 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n16104) );
  AOI22_X1 U16046 ( .A1(n19814), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12726) );
  OAI21_X1 U16047 ( .B1(n16104), .B2(n19782), .A(n12726), .ZN(P2_U2926) );
  INV_X1 U16048 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n16131) );
  AOI22_X1 U16049 ( .A1(n19814), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12727) );
  OAI21_X1 U16050 ( .B1(n16131), .B2(n19782), .A(n12727), .ZN(P2_U2930) );
  AOI22_X1 U16051 ( .A1(n19814), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12728) );
  OAI21_X1 U16052 ( .B1(n16111), .B2(n19782), .A(n12728), .ZN(P2_U2928) );
  INV_X1 U16053 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n16121) );
  AOI22_X1 U16054 ( .A1(n19814), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12729) );
  OAI21_X1 U16055 ( .B1(n16121), .B2(n19782), .A(n12729), .ZN(P2_U2929) );
  INV_X1 U16056 ( .A(n9706), .ZN(n12738) );
  OAI21_X1 U16057 ( .B1(n19691), .B2(n12837), .A(n12730), .ZN(n12731) );
  XOR2_X1 U16058 ( .A(n12731), .B(n21108), .Z(n16524) );
  AOI21_X1 U16059 ( .B1(n21108), .B2(n12733), .A(n12732), .ZN(n16523) );
  AND2_X1 U16060 ( .A1(n19825), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n16522) );
  AOI21_X1 U16061 ( .B1(n11531), .B2(n16523), .A(n16522), .ZN(n12735) );
  NAND2_X1 U16062 ( .A1(n17038), .A2(n19689), .ZN(n12734) );
  OAI211_X1 U16063 ( .C1(n17046), .C2(n19689), .A(n12735), .B(n12734), .ZN(
        n12736) );
  AOI21_X1 U16064 ( .B1(n19828), .B2(n16524), .A(n12736), .ZN(n12737) );
  OAI21_X1 U16065 ( .B1(n12738), .B2(n16307), .A(n12737), .ZN(P2_U3013) );
  NOR2_X1 U16066 ( .A1(n17100), .A2(n20484), .ZN(n17094) );
  NOR2_X1 U16067 ( .A1(n11022), .A2(n13444), .ZN(n12739) );
  NAND2_X1 U16068 ( .A1(n12740), .A2(n12739), .ZN(n12743) );
  INV_X1 U16069 ( .A(n13219), .ZN(n13428) );
  NAND2_X1 U16070 ( .A1(n13428), .A2(n13423), .ZN(n13123) );
  NAND4_X1 U16071 ( .A1(n12743), .A2(n12742), .A3(n12741), .A4(n13123), .ZN(
        n13437) );
  INV_X1 U16072 ( .A(n13437), .ZN(n13402) );
  OAI22_X1 U16073 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20101), .B1(n13402), 
        .B2(n19561), .ZN(n12744) );
  AOI21_X1 U16074 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17094), .A(n12744), .ZN(
        n16553) );
  INV_X1 U16075 ( .A(n16553), .ZN(n12746) );
  NOR2_X1 U16076 ( .A1(n11022), .A2(n14265), .ZN(n13431) );
  INV_X1 U16077 ( .A(n20455), .ZN(n16547) );
  NAND4_X1 U16078 ( .A1(n12746), .A2(n13431), .A3(n9812), .A4(n16547), .ZN(
        n12745) );
  OAI21_X1 U16079 ( .B1(n12746), .B2(n21165), .A(n12745), .ZN(P2_U3595) );
  INV_X1 U16080 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n21320) );
  NAND2_X1 U16081 ( .A1(n20619), .A2(n13832), .ZN(n13066) );
  AOI22_X1 U16082 ( .A1(n21029), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20644), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12747) );
  OAI21_X1 U16083 ( .B1(n21320), .B2(n13066), .A(n12747), .ZN(P1_U2906) );
  INV_X1 U16084 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U16085 ( .A1(n20647), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20644), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12748) );
  OAI21_X1 U16086 ( .B1(n12940), .B2(n13066), .A(n12748), .ZN(P1_U2912) );
  INV_X1 U16087 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U16088 ( .A1(n20647), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20644), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12749) );
  OAI21_X1 U16089 ( .B1(n12943), .B2(n13066), .A(n12749), .ZN(P1_U2907) );
  INV_X1 U16090 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U16091 ( .A1(n20647), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20644), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12750) );
  OAI21_X1 U16092 ( .B1(n12937), .B2(n13066), .A(n12750), .ZN(P1_U2908) );
  INV_X1 U16093 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U16094 ( .A1(n20647), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20644), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12751) );
  OAI21_X1 U16095 ( .B1(n12930), .B2(n13066), .A(n12751), .ZN(P1_U2909) );
  INV_X1 U16096 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U16097 ( .A1(n20647), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20644), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12752) );
  OAI21_X1 U16098 ( .B1(n12953), .B2(n13066), .A(n12752), .ZN(P1_U2910) );
  INV_X1 U16099 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12950) );
  AOI22_X1 U16100 ( .A1(n20647), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20644), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12753) );
  OAI21_X1 U16101 ( .B1(n12950), .B2(n13066), .A(n12753), .ZN(P1_U2911) );
  NAND2_X1 U16102 ( .A1(n12756), .A2(n12755), .ZN(n12773) );
  INV_X1 U16103 ( .A(n13571), .ZN(n12763) );
  NAND2_X1 U16104 ( .A1(n12763), .A2(n13097), .ZN(n12854) );
  NAND2_X1 U16105 ( .A1(n12854), .A2(n12764), .ZN(n12757) );
  OAI21_X1 U16106 ( .B1(n12778), .B2(n12757), .A(n12975), .ZN(n12762) );
  NAND2_X1 U16107 ( .A1(n12759), .A2(n13079), .ZN(n12760) );
  NAND2_X1 U16108 ( .A1(n12763), .A2(n13832), .ZN(n13271) );
  NAND2_X2 U16109 ( .A1(n13271), .A2(n15147), .ZN(n15218) );
  NAND2_X1 U16110 ( .A1(n13558), .A2(n13832), .ZN(n12858) );
  INV_X1 U16111 ( .A(n16646), .ZN(n16639) );
  NAND2_X1 U16112 ( .A1(n16639), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12788) );
  NOR2_X1 U16113 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21003) );
  NAND2_X1 U16114 ( .A1(n21003), .A2(n9922), .ZN(n12981) );
  NAND2_X1 U16115 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12795) );
  OAI21_X1 U16116 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n12795), .ZN(n20701) );
  OR2_X1 U16117 ( .A1(n12981), .A2(n20701), .ZN(n12770) );
  AND2_X1 U16118 ( .A1(n12788), .A2(n12770), .ZN(n12771) );
  NAND3_X1 U16119 ( .A1(n13082), .A2(n12773), .A3(n13107), .ZN(n12774) );
  XNOR2_X2 U16120 ( .A(n12775), .B(n12790), .ZN(n13718) );
  MUX2_X1 U16121 ( .A(n12981), .B(n16646), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n12776) );
  NAND2_X1 U16122 ( .A1(n12778), .A2(n12779), .ZN(n12862) );
  NAND2_X1 U16123 ( .A1(n13519), .A2(n12780), .ZN(n13101) );
  NAND2_X1 U16124 ( .A1(n12975), .A2(n13587), .ZN(n13838) );
  NAND4_X1 U16125 ( .A1(n13101), .A2(n21003), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n13838), .ZN(n12781) );
  NOR2_X1 U16126 ( .A1(n12782), .A2(n12781), .ZN(n12787) );
  NAND2_X1 U16127 ( .A1(n12759), .A2(n13571), .ZN(n12783) );
  AOI22_X1 U16128 ( .A1(n12784), .A2(n12783), .B1(n12758), .B2(n14536), .ZN(
        n12786) );
  NAND3_X1 U16129 ( .A1(n12815), .A2(n12761), .A3(n13587), .ZN(n12785) );
  NAND4_X1 U16130 ( .A1(n12862), .A2(n12787), .A3(n12786), .A4(n12785), .ZN(
        n12880) );
  NAND2_X1 U16131 ( .A1(n12788), .A2(n9712), .ZN(n12789) );
  INV_X1 U16133 ( .A(n12981), .ZN(n12797) );
  INV_X1 U16134 ( .A(n12795), .ZN(n12794) );
  NAND2_X1 U16135 ( .A1(n12794), .A2(n16622), .ZN(n13765) );
  NAND2_X1 U16136 ( .A1(n12795), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12796) );
  NAND2_X1 U16137 ( .A1(n13765), .A2(n12796), .ZN(n14049) );
  AOI22_X1 U16138 ( .A1(n12797), .A2(n14049), .B1(n16639), .B2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12798) );
  INV_X1 U16139 ( .A(n12793), .ZN(n12799) );
  NAND2_X1 U16140 ( .A1(n12799), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12803) );
  NAND2_X1 U16141 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10340), .ZN(
        n13747) );
  NAND2_X1 U16142 ( .A1(n20737), .A2(n13747), .ZN(n12800) );
  NOR3_X1 U16143 ( .A1(n20737), .A2(n16622), .A3(n20698), .ZN(n14556) );
  NAND2_X1 U16144 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14556), .ZN(
        n14548) );
  NAND2_X1 U16145 ( .A1(n12800), .A2(n14548), .ZN(n14190) );
  OAI22_X1 U16146 ( .A1(n12981), .A2(n14190), .B1(n16646), .B2(n20737), .ZN(
        n12801) );
  INV_X1 U16147 ( .A(n12801), .ZN(n12802) );
  INV_X1 U16148 ( .A(n13544), .ZN(n13983) );
  OR2_X1 U16149 ( .A1(n13173), .A2(n13983), .ZN(n12804) );
  XNOR2_X1 U16150 ( .A(n12804), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20574) );
  NOR2_X1 U16151 ( .A1(n12766), .A2(n13587), .ZN(n12852) );
  NAND2_X1 U16152 ( .A1(n20574), .A2(n12852), .ZN(n13511) );
  NAND2_X1 U16153 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21028) );
  NAND2_X1 U16154 ( .A1(n13587), .A2(n21028), .ZN(n12806) );
  INV_X1 U16155 ( .A(n12761), .ZN(n12954) );
  NOR2_X1 U16156 ( .A1(n12818), .A2(n15286), .ZN(n12805) );
  NAND2_X1 U16157 ( .A1(n12954), .A2(n12805), .ZN(n15275) );
  OAI21_X1 U16158 ( .B1(n12767), .B2(n12806), .A(n15275), .ZN(n12807) );
  NAND2_X1 U16159 ( .A1(n16614), .A2(n12807), .ZN(n12809) );
  NAND3_X1 U16160 ( .A1(n15282), .A2(n12764), .A3(n21028), .ZN(n12808) );
  NAND2_X1 U16161 ( .A1(n12809), .A2(n12808), .ZN(n12917) );
  INV_X1 U16162 ( .A(n21028), .ZN(n20943) );
  NOR2_X1 U16163 ( .A1(n16666), .A2(n20943), .ZN(n12811) );
  AND2_X1 U16164 ( .A1(n12810), .A2(n12811), .ZN(n12812) );
  AND2_X1 U16165 ( .A1(n16614), .A2(n12812), .ZN(n16640) );
  OR2_X1 U16166 ( .A1(n12917), .A2(n16640), .ZN(n12823) );
  NAND2_X1 U16167 ( .A1(n12761), .A2(n12975), .ZN(n12813) );
  AND2_X1 U16168 ( .A1(n12814), .A2(n12813), .ZN(n12979) );
  OAI211_X1 U16169 ( .C1(n12764), .C2(n12759), .A(n12815), .B(n13832), .ZN(
        n12860) );
  NAND2_X1 U16170 ( .A1(n12979), .A2(n12860), .ZN(n12816) );
  NAND2_X1 U16171 ( .A1(n12816), .A2(n12766), .ZN(n13075) );
  OR2_X1 U16172 ( .A1(n13838), .A2(n13558), .ZN(n12817) );
  AND2_X1 U16173 ( .A1(n13075), .A2(n12817), .ZN(n12820) );
  NOR2_X1 U16174 ( .A1(n15287), .A2(n12818), .ZN(n12819) );
  NAND2_X1 U16175 ( .A1(n12954), .A2(n12819), .ZN(n13105) );
  OR2_X1 U16176 ( .A1(n16614), .A2(n13105), .ZN(n13050) );
  OAI211_X1 U16177 ( .C1(n12821), .C2(n20943), .A(n12820), .B(n13050), .ZN(
        n12822) );
  NAND2_X1 U16178 ( .A1(n16616), .A2(n13077), .ZN(n12825) );
  INV_X1 U16179 ( .A(n16878), .ZN(n21290) );
  NAND2_X1 U16180 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21290), .ZN(n16883) );
  INV_X1 U16181 ( .A(n16883), .ZN(n13536) );
  NAND2_X1 U16182 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13536), .ZN(n12824) );
  NAND2_X1 U16183 ( .A1(n12825), .A2(n12824), .ZN(n12828) );
  NAND2_X1 U16184 ( .A1(n12828), .A2(n21003), .ZN(n14745) );
  INV_X1 U16185 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n12826) );
  NOR2_X1 U16186 ( .A1(n12826), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12827) );
  NOR2_X1 U16187 ( .A1(n12828), .A2(n12827), .ZN(n21012) );
  INV_X1 U16188 ( .A(n21012), .ZN(n21014) );
  OAI22_X1 U16189 ( .A1(n13511), .A2(n14745), .B1(n12829), .B2(n21014), .ZN(
        P1_U3468) );
  AND2_X1 U16190 ( .A1(n16636), .A2(n20943), .ZN(n12830) );
  INV_X2 U16191 ( .A(n12931), .ZN(n13015) );
  INV_X1 U16192 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20621) );
  OR2_X1 U16193 ( .A1(n13015), .A2(n12764), .ZN(n12926) );
  INV_X1 U16194 ( .A(DATAI_15_), .ZN(n12833) );
  INV_X1 U16195 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12832) );
  MUX2_X1 U16196 ( .A(n12833), .B(n12832), .S(n15109), .Z(n15603) );
  INV_X1 U16197 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n12834) );
  OAI222_X1 U16198 ( .A1(n13001), .A2(n20621), .B1(n12926), .B2(n15603), .C1(
        n12931), .C2(n12834), .ZN(P1_U2967) );
  INV_X1 U16199 ( .A(n14515), .ZN(n12836) );
  INV_X1 U16200 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12835) );
  NAND2_X1 U16201 ( .A1(n12836), .A2(n12835), .ZN(n12838) );
  AND2_X1 U16202 ( .A1(n12838), .A2(n12837), .ZN(n15260) );
  NAND2_X1 U16203 ( .A1(n19825), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n15256) );
  OAI21_X1 U16204 ( .B1(n19870), .B2(n15264), .A(n15256), .ZN(n12847) );
  NOR2_X1 U16205 ( .A1(n12840), .A2(n12839), .ZN(n12841) );
  NOR2_X1 U16206 ( .A1(n12842), .A2(n12841), .ZN(n19775) );
  INV_X1 U16207 ( .A(n19775), .ZN(n12845) );
  OAI21_X1 U16208 ( .B1(n12844), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12843), .ZN(n15257) );
  OAI22_X1 U16209 ( .A1(n17070), .A2(n12845), .B1(n19859), .B2(n15257), .ZN(
        n12846) );
  AOI211_X1 U16210 ( .C1(n19866), .C2(n15260), .A(n12847), .B(n12846), .ZN(
        n12849) );
  INV_X1 U16211 ( .A(n19851), .ZN(n16520) );
  MUX2_X1 U16212 ( .A(n16432), .B(n16520), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n12848) );
  NAND2_X1 U16213 ( .A1(n12849), .A2(n12848), .ZN(P2_U3046) );
  INV_X1 U16214 ( .A(n14740), .ZN(n12850) );
  OAI21_X1 U16215 ( .B1(n12850), .B2(n12434), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12851) );
  NAND2_X1 U16216 ( .A1(n14344), .A2(n12851), .ZN(n12874) );
  INV_X1 U16217 ( .A(n12874), .ZN(n12879) );
  OR2_X1 U16218 ( .A1(n21012), .A2(n21010), .ZN(n12878) );
  INV_X1 U16219 ( .A(n13908), .ZN(n20600) );
  INV_X1 U16220 ( .A(n12852), .ZN(n12867) );
  NAND2_X1 U16221 ( .A1(n12853), .A2(n12975), .ZN(n12855) );
  NAND2_X1 U16222 ( .A1(n12855), .A2(n12854), .ZN(n12856) );
  INV_X1 U16223 ( .A(n12857), .ZN(n12859) );
  AND4_X1 U16224 ( .A1(n12861), .A2(n12860), .A3(n12859), .A4(n12858), .ZN(
        n12863) );
  AND2_X1 U16225 ( .A1(n12863), .A2(n12862), .ZN(n13102) );
  NAND2_X1 U16226 ( .A1(n12864), .A2(n13103), .ZN(n12865) );
  NOR2_X1 U16227 ( .A1(n12810), .A2(n12865), .ZN(n12866) );
  XNOR2_X1 U16228 ( .A(n12868), .B(n13262), .ZN(n12873) );
  MUX2_X1 U16229 ( .A(n12869), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14740), .Z(n12871) );
  NOR2_X1 U16230 ( .A1(n12871), .A2(n12870), .ZN(n12872) );
  NAND2_X1 U16231 ( .A1(n13105), .A2(n15275), .ZN(n13516) );
  AOI22_X1 U16232 ( .A1(n14742), .A2(n12873), .B1(n12872), .B2(n13516), .ZN(
        n12876) );
  NAND3_X1 U16233 ( .A1(n14744), .A2(n13519), .A3(n12874), .ZN(n12875) );
  OAI211_X1 U16234 ( .C1(n20600), .C2(n14744), .A(n12876), .B(n12875), .ZN(
        n13527) );
  INV_X1 U16235 ( .A(n13527), .ZN(n12877) );
  OAI222_X1 U16236 ( .A1(n21014), .A2(n13262), .B1(n12879), .B2(n12878), .C1(
        n14745), .C2(n12877), .ZN(P1_U3469) );
  INV_X1 U16237 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12904) );
  AOI22_X1 U16238 ( .A1(n15015), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15081), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12884) );
  AOI22_X1 U16239 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13960), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12883) );
  AOI22_X1 U16240 ( .A1(n15040), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12882) );
  AOI22_X1 U16241 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12881) );
  NAND4_X1 U16242 ( .A1(n12884), .A2(n12883), .A3(n12882), .A4(n12881), .ZN(
        n12891) );
  AOI22_X1 U16243 ( .A1(n12892), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16244 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U16245 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U16246 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12886) );
  NAND4_X1 U16247 ( .A1(n12889), .A2(n12888), .A3(n12887), .A4(n12886), .ZN(
        n12890) );
  AOI21_X1 U16248 ( .B1(n12975), .B2(n13194), .A(n9922), .ZN(n12903) );
  AOI22_X1 U16249 ( .A1(n12892), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12896) );
  AOI22_X1 U16250 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U16251 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9710), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U16252 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12893) );
  NAND4_X1 U16253 ( .A1(n12896), .A2(n12895), .A3(n12894), .A4(n12893), .ZN(
        n12902) );
  AOI22_X1 U16254 ( .A1(n15015), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15082), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U16255 ( .A1(n14947), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U16256 ( .A1(n14948), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U16257 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12897) );
  NAND4_X1 U16258 ( .A1(n12900), .A2(n12899), .A3(n12898), .A4(n12897), .ZN(
        n12901) );
  NAND2_X1 U16259 ( .A1(n13079), .A2(n14535), .ZN(n12905) );
  OAI211_X1 U16260 ( .C1(n14103), .C2(n12904), .A(n12903), .B(n12905), .ZN(
        n13140) );
  NAND2_X1 U16261 ( .A1(n13139), .A2(n13140), .ZN(n12909) );
  NOR2_X1 U16262 ( .A1(n13547), .A2(n9922), .ZN(n13185) );
  INV_X1 U16263 ( .A(n14535), .ZN(n14104) );
  NAND2_X1 U16264 ( .A1(n13185), .A2(n14104), .ZN(n13137) );
  INV_X1 U16265 ( .A(n13137), .ZN(n12907) );
  INV_X1 U16266 ( .A(n13194), .ZN(n12906) );
  MUX2_X1 U16267 ( .A(n12907), .B(n14531), .S(n12906), .Z(n13138) );
  NAND2_X1 U16268 ( .A1(n13138), .A2(n13140), .ZN(n12910) );
  AOI21_X1 U16269 ( .B1(n13721), .B2(n12780), .A(n14046), .ZN(n12916) );
  INV_X1 U16270 ( .A(n12911), .ZN(n15925) );
  NAND2_X1 U16271 ( .A1(n12780), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14797) );
  NAND2_X1 U16272 ( .A1(n15925), .A2(n14780), .ZN(n12915) );
  NAND2_X1 U16273 ( .A1(n9937), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13263) );
  INV_X1 U16274 ( .A(n13263), .ZN(n13615) );
  NAND2_X1 U16275 ( .A1(n13615), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12913) );
  INV_X1 U16276 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n14046) );
  AOI22_X1 U16277 ( .A1(n15246), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n14046), .ZN(n12912) );
  AND2_X1 U16278 ( .A1(n12913), .A2(n12912), .ZN(n12914) );
  NAND2_X1 U16279 ( .A1(n12915), .A2(n12914), .ZN(n13151) );
  NAND2_X1 U16280 ( .A1(n12916), .A2(n13151), .ZN(n13154) );
  OAI21_X1 U16281 ( .B1(n12916), .B2(n13151), .A(n13154), .ZN(n15483) );
  NAND2_X1 U16282 ( .A1(n12917), .A2(n13077), .ZN(n12922) );
  INV_X1 U16283 ( .A(n12918), .ZN(n12920) );
  INV_X1 U16284 ( .A(n13577), .ZN(n15533) );
  NOR2_X1 U16285 ( .A1(n13547), .A2(n20508), .ZN(n12919) );
  AND4_X1 U16286 ( .A1(n12920), .A2(n15533), .A3(n13519), .A4(n12919), .ZN(
        n13051) );
  NAND2_X1 U16287 ( .A1(n13051), .A2(n12779), .ZN(n12921) );
  NAND2_X1 U16288 ( .A1(n12759), .A2(n13577), .ZN(n12923) );
  NAND2_X2 U16289 ( .A1(n15606), .A2(n12923), .ZN(n15614) );
  INV_X1 U16290 ( .A(n15109), .ZN(n15105) );
  NAND2_X1 U16291 ( .A1(n15105), .A2(DATAI_0_), .ZN(n12925) );
  NAND2_X1 U16292 ( .A1(n15109), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12924) );
  AND2_X1 U16293 ( .A1(n12925), .A2(n12924), .ZN(n15596) );
  INV_X1 U16294 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20650) );
  OAI222_X1 U16295 ( .A1(n15483), .A2(n15614), .B1(n15608), .B2(n15596), .C1(
        n15606), .C2(n20650), .ZN(P1_U2904) );
  INV_X1 U16296 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15593) );
  INV_X1 U16297 ( .A(n15596), .ZN(n12927) );
  NAND2_X1 U16298 ( .A1(n13030), .A2(n12927), .ZN(n13038) );
  NAND2_X1 U16299 ( .A1(n13015), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n12928) );
  OAI211_X1 U16300 ( .C1(n15593), .C2(n13001), .A(n13038), .B(n12928), .ZN(
        P1_U2937) );
  MUX2_X1 U16301 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n15109), .Z(
        n15545) );
  NAND2_X1 U16302 ( .A1(n13030), .A2(n15545), .ZN(n12947) );
  NAND2_X1 U16303 ( .A1(n13015), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n12929) );
  OAI211_X1 U16304 ( .C1(n12930), .C2(n13001), .A(n12947), .B(n12929), .ZN(
        P1_U2948) );
  INV_X1 U16305 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20632) );
  MUX2_X1 U16306 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n15109), .Z(
        n15552) );
  NAND2_X1 U16307 ( .A1(n13030), .A2(n15552), .ZN(n12949) );
  NAND2_X1 U16308 ( .A1(n13015), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n12932) );
  OAI211_X1 U16309 ( .C1(n20632), .C2(n13001), .A(n12949), .B(n12932), .ZN(
        P1_U2961) );
  INV_X1 U16310 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20634) );
  MUX2_X1 U16311 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n15109), .Z(
        n15556) );
  NAND2_X1 U16312 ( .A1(n13030), .A2(n15556), .ZN(n12939) );
  NAND2_X1 U16313 ( .A1(n13015), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n12933) );
  OAI211_X1 U16314 ( .C1(n20634), .C2(n13001), .A(n12939), .B(n12933), .ZN(
        P1_U2960) );
  INV_X1 U16315 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20626) );
  MUX2_X1 U16316 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n15109), .Z(
        n15541) );
  NAND2_X1 U16317 ( .A1(n13030), .A2(n15541), .ZN(n12936) );
  NAND2_X1 U16318 ( .A1(n13015), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n12934) );
  OAI211_X1 U16319 ( .C1(n20626), .C2(n13001), .A(n12936), .B(n12934), .ZN(
        P1_U2964) );
  NAND2_X1 U16320 ( .A1(n13015), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n12935) );
  OAI211_X1 U16321 ( .C1(n12937), .C2(n13001), .A(n12936), .B(n12935), .ZN(
        P1_U2949) );
  NAND2_X1 U16322 ( .A1(n13015), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n12938) );
  OAI211_X1 U16323 ( .C1(n12940), .C2(n13001), .A(n12939), .B(n12938), .ZN(
        P1_U2945) );
  INV_X1 U16324 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20630) );
  MUX2_X1 U16325 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n15109), .Z(
        n15549) );
  NAND2_X1 U16326 ( .A1(n13030), .A2(n15549), .ZN(n12952) );
  NAND2_X1 U16327 ( .A1(n13015), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n12941) );
  OAI211_X1 U16328 ( .C1(n20630), .C2(n13001), .A(n12952), .B(n12941), .ZN(
        P1_U2962) );
  MUX2_X1 U16329 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n15109), .Z(
        n15611) );
  NAND2_X1 U16330 ( .A1(n13030), .A2(n15611), .ZN(n12945) );
  NAND2_X1 U16331 ( .A1(n13015), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n12942) );
  OAI211_X1 U16332 ( .C1(n12943), .C2(n13001), .A(n12945), .B(n12942), .ZN(
        P1_U2950) );
  INV_X1 U16333 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20624) );
  NAND2_X1 U16334 ( .A1(n13015), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n12944) );
  OAI211_X1 U16335 ( .C1(n20624), .C2(n13001), .A(n12945), .B(n12944), .ZN(
        P1_U2965) );
  INV_X1 U16336 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20628) );
  NAND2_X1 U16337 ( .A1(n13015), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n12946) );
  OAI211_X1 U16338 ( .C1(n20628), .C2(n13001), .A(n12947), .B(n12946), .ZN(
        P1_U2963) );
  NAND2_X1 U16339 ( .A1(n13015), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n12948) );
  OAI211_X1 U16340 ( .C1(n12950), .C2(n13001), .A(n12949), .B(n12948), .ZN(
        P1_U2946) );
  NAND2_X1 U16341 ( .A1(n13015), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n12951) );
  OAI211_X1 U16342 ( .C1(n12953), .C2(n13001), .A(n12952), .B(n12951), .ZN(
        P1_U2947) );
  INV_X1 U16343 ( .A(n14744), .ZN(n12956) );
  MUX2_X1 U16344 ( .A(n12954), .B(n14742), .S(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n12955) );
  AOI21_X1 U16345 ( .B1(n15925), .B2(n12956), .A(n12955), .ZN(n16618) );
  OAI22_X1 U16346 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21010), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21133), .ZN(n12957) );
  AOI22_X1 U16347 ( .A1(n21012), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n12957), .B2(n21014), .ZN(n12958) );
  OAI21_X1 U16348 ( .B1(n16618), .B2(n14745), .A(n12958), .ZN(P1_U3474) );
  INV_X1 U16349 ( .A(n16155), .ZN(n16973) );
  OR2_X1 U16350 ( .A1(n12962), .A2(n12961), .ZN(n12963) );
  XNOR2_X1 U16351 ( .A(n12965), .B(n12964), .ZN(n19702) );
  XNOR2_X1 U16352 ( .A(n20478), .B(n19702), .ZN(n12970) );
  NAND2_X1 U16353 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12966) );
  NAND4_X1 U16354 ( .A1(n12967), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12966), 
        .A4(n20101), .ZN(n12968) );
  NAND2_X1 U16355 ( .A1(n19776), .A2(n19775), .ZN(n19774) );
  NAND2_X1 U16356 ( .A1(n12970), .A2(n19774), .ZN(n12993) );
  OAI21_X1 U16357 ( .B1(n12970), .B2(n19774), .A(n12993), .ZN(n12971) );
  NAND2_X1 U16358 ( .A1(n12971), .A2(n19773), .ZN(n12973) );
  INV_X1 U16359 ( .A(n19702), .ZN(n20474) );
  INV_X1 U16360 ( .A(n19744), .ZN(n19771) );
  AOI22_X1 U16361 ( .A1(n19772), .A2(n20474), .B1(n19771), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n12972) );
  OAI211_X1 U16362 ( .C1(n14335), .C2(n19779), .A(n12973), .B(n12972), .ZN(
        P2_U2918) );
  NAND3_X1 U16363 ( .A1(n9922), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16876) );
  INV_X1 U16364 ( .A(n16876), .ZN(n12974) );
  INV_X1 U16365 ( .A(n16764), .ZN(n16770) );
  NAND2_X1 U16366 ( .A1(n12975), .A2(n13571), .ZN(n13198) );
  OAI21_X1 U16367 ( .B1(n16636), .B2(n13194), .A(n13198), .ZN(n12976) );
  OAI21_X1 U16368 ( .B1(n12977), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13163), .ZN(n20654) );
  AND2_X1 U16369 ( .A1(n12979), .A2(n12978), .ZN(n15274) );
  NAND2_X1 U16370 ( .A1(n16614), .A2(n15274), .ZN(n16628) );
  OR2_X2 U16371 ( .A1(n12981), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16808) );
  INV_X1 U16372 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n12980) );
  OR2_X1 U16373 ( .A1(n16808), .A2(n12980), .ZN(n20660) );
  INV_X1 U16374 ( .A(n20866), .ZN(n20807) );
  NAND2_X1 U16375 ( .A1(n20807), .A2(n12981), .ZN(n21027) );
  NAND2_X1 U16376 ( .A1(n21027), .A2(n9922), .ZN(n12982) );
  NAND2_X1 U16377 ( .A1(n9922), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16637) );
  INV_X1 U16378 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20514) );
  NAND2_X1 U16379 ( .A1(n20514), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12983) );
  NAND2_X1 U16380 ( .A1(n16637), .A2(n12983), .ZN(n13158) );
  OAI21_X1 U16381 ( .B1(n16759), .B2(n13158), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12984) );
  OAI211_X1 U16382 ( .C1(n20654), .C2(n20516), .A(n20660), .B(n12984), .ZN(
        n12985) );
  INV_X1 U16383 ( .A(n12985), .ZN(n12986) );
  OAI21_X1 U16384 ( .B1(n16770), .B2(n15483), .A(n12986), .ZN(P1_U2999) );
  NAND2_X1 U16385 ( .A1(n12988), .A2(n12987), .ZN(n12990) );
  NAND2_X1 U16386 ( .A1(n12990), .A2(n10225), .ZN(n20468) );
  INV_X1 U16387 ( .A(n20468), .ZN(n19750) );
  INV_X1 U16388 ( .A(n19772), .ZN(n16085) );
  XNOR2_X1 U16389 ( .A(n20466), .B(n20468), .ZN(n12996) );
  NAND2_X1 U16390 ( .A1(n14255), .A2(n19702), .ZN(n12994) );
  NAND2_X1 U16391 ( .A1(n12994), .A2(n12993), .ZN(n12995) );
  NAND2_X1 U16392 ( .A1(n12996), .A2(n12995), .ZN(n19751) );
  OAI21_X1 U16393 ( .B1(n12996), .B2(n12995), .A(n19751), .ZN(n12997) );
  NAND2_X1 U16394 ( .A1(n12997), .A2(n19773), .ZN(n13000) );
  INV_X1 U16395 ( .A(n19881), .ZN(n12998) );
  AOI22_X1 U16396 ( .A1(n19746), .A2(n12998), .B1(n19771), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n12999) );
  OAI211_X1 U16397 ( .C1(n19750), .C2(n16085), .A(n13000), .B(n12999), .ZN(
        P2_U2917) );
  AOI22_X1 U16398 ( .A1(n13042), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n13015), .ZN(n13004) );
  NAND2_X1 U16399 ( .A1(n15105), .A2(DATAI_2_), .ZN(n13003) );
  NAND2_X1 U16400 ( .A1(n15109), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13002) );
  AND2_X1 U16401 ( .A1(n13003), .A2(n13002), .ZN(n13557) );
  INV_X1 U16402 ( .A(n13557), .ZN(n15583) );
  NAND2_X1 U16403 ( .A1(n13030), .A2(n15583), .ZN(n13019) );
  NAND2_X1 U16404 ( .A1(n13004), .A2(n13019), .ZN(P1_U2939) );
  AOI22_X1 U16405 ( .A1(n13042), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n13015), .ZN(n13007) );
  INV_X1 U16406 ( .A(DATAI_7_), .ZN(n13006) );
  NAND2_X1 U16407 ( .A1(n15109), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13005) );
  OAI21_X1 U16408 ( .B1(n15109), .B2(n13006), .A(n13005), .ZN(n15560) );
  NAND2_X1 U16409 ( .A1(n13030), .A2(n15560), .ZN(n13023) );
  NAND2_X1 U16410 ( .A1(n13007), .A2(n13023), .ZN(P1_U2944) );
  AOI22_X1 U16411 ( .A1(n13042), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n13015), .ZN(n13008) );
  MUX2_X1 U16412 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n15109), .Z(
        n15605) );
  NAND2_X1 U16413 ( .A1(n13030), .A2(n15605), .ZN(n13032) );
  NAND2_X1 U16414 ( .A1(n13008), .A2(n13032), .ZN(P1_U2966) );
  AOI22_X1 U16415 ( .A1(n13042), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n13015), .ZN(n13011) );
  INV_X1 U16416 ( .A(DATAI_5_), .ZN(n13010) );
  NAND2_X1 U16417 ( .A1(n15109), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13009) );
  OAI21_X1 U16418 ( .B1(n15109), .B2(n13010), .A(n13009), .ZN(n15570) );
  NAND2_X1 U16419 ( .A1(n13030), .A2(n15570), .ZN(n13040) );
  NAND2_X1 U16420 ( .A1(n13011), .A2(n13040), .ZN(P1_U2942) );
  AOI22_X1 U16421 ( .A1(n13042), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n13015), .ZN(n13014) );
  INV_X1 U16422 ( .A(DATAI_4_), .ZN(n13013) );
  NAND2_X1 U16423 ( .A1(n15109), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13012) );
  OAI21_X1 U16424 ( .B1(n15109), .B2(n13013), .A(n13012), .ZN(n15575) );
  NAND2_X1 U16425 ( .A1(n13030), .A2(n15575), .ZN(n13036) );
  NAND2_X1 U16426 ( .A1(n13014), .A2(n13036), .ZN(P1_U2941) );
  AOI22_X1 U16427 ( .A1(n13042), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n13015), .ZN(n13018) );
  INV_X1 U16428 ( .A(DATAI_6_), .ZN(n13017) );
  NAND2_X1 U16429 ( .A1(n15109), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13016) );
  OAI21_X1 U16430 ( .B1(n15109), .B2(n13017), .A(n13016), .ZN(n15566) );
  NAND2_X1 U16431 ( .A1(n13030), .A2(n15566), .ZN(n13021) );
  NAND2_X1 U16432 ( .A1(n13018), .A2(n13021), .ZN(P1_U2943) );
  AOI22_X1 U16433 ( .A1(n13042), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n13015), .ZN(n13020) );
  NAND2_X1 U16434 ( .A1(n13020), .A2(n13019), .ZN(P1_U2954) );
  AOI22_X1 U16435 ( .A1(n13042), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n13015), .ZN(n13022) );
  NAND2_X1 U16436 ( .A1(n13022), .A2(n13021), .ZN(P1_U2958) );
  AOI22_X1 U16437 ( .A1(n13042), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n13015), .ZN(n13024) );
  NAND2_X1 U16438 ( .A1(n13024), .A2(n13023), .ZN(P1_U2959) );
  AOI22_X1 U16439 ( .A1(n13042), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n13015), .ZN(n13027) );
  NAND2_X1 U16440 ( .A1(n15105), .A2(DATAI_1_), .ZN(n13026) );
  NAND2_X1 U16441 ( .A1(n15109), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13025) );
  AND2_X1 U16442 ( .A1(n13026), .A2(n13025), .ZN(n13586) );
  INV_X1 U16443 ( .A(n13586), .ZN(n15588) );
  NAND2_X1 U16444 ( .A1(n13030), .A2(n15588), .ZN(n13034) );
  NAND2_X1 U16445 ( .A1(n13027), .A2(n13034), .ZN(P1_U2953) );
  AOI22_X1 U16446 ( .A1(n13042), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n13015), .ZN(n13031) );
  NAND2_X1 U16447 ( .A1(n15105), .A2(DATAI_3_), .ZN(n13029) );
  NAND2_X1 U16448 ( .A1(n15109), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13028) );
  AND2_X1 U16449 ( .A1(n13029), .A2(n13028), .ZN(n13570) );
  INV_X1 U16450 ( .A(n13570), .ZN(n15579) );
  NAND2_X1 U16451 ( .A1(n13030), .A2(n15579), .ZN(n13043) );
  NAND2_X1 U16452 ( .A1(n13031), .A2(n13043), .ZN(P1_U2955) );
  AOI22_X1 U16453 ( .A1(n13042), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n13015), .ZN(n13033) );
  NAND2_X1 U16454 ( .A1(n13033), .A2(n13032), .ZN(P1_U2951) );
  AOI22_X1 U16455 ( .A1(n13042), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n13015), .ZN(n13035) );
  NAND2_X1 U16456 ( .A1(n13035), .A2(n13034), .ZN(P1_U2938) );
  AOI22_X1 U16457 ( .A1(n13042), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n13015), .ZN(n13037) );
  NAND2_X1 U16458 ( .A1(n13037), .A2(n13036), .ZN(P1_U2956) );
  AOI22_X1 U16459 ( .A1(n13042), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n13015), .ZN(n13039) );
  NAND2_X1 U16460 ( .A1(n13039), .A2(n13038), .ZN(P1_U2952) );
  AOI22_X1 U16461 ( .A1(n13042), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n13015), .ZN(n13041) );
  NAND2_X1 U16462 ( .A1(n13041), .A2(n13040), .ZN(P1_U2957) );
  AOI22_X1 U16463 ( .A1(n13042), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n13015), .ZN(n13044) );
  NAND2_X1 U16464 ( .A1(n13044), .A2(n13043), .ZN(P1_U2940) );
  INV_X1 U16465 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13045) );
  OR2_X1 U16466 ( .A1(n15149), .A2(n13045), .ZN(n13047) );
  NAND2_X1 U16467 ( .A1(n12765), .A2(n13045), .ZN(n13046) );
  NAND2_X1 U16468 ( .A1(n13047), .A2(n13046), .ZN(n13112) );
  INV_X1 U16469 ( .A(n13112), .ZN(n13049) );
  OR2_X1 U16470 ( .A1(n15218), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13048) );
  NAND2_X1 U16471 ( .A1(n13049), .A2(n13048), .ZN(n20651) );
  NAND2_X1 U16472 ( .A1(n13051), .A2(n15162), .ZN(n13052) );
  NAND2_X1 U16473 ( .A1(n20618), .A2(n13577), .ZN(n15529) );
  OAI222_X1 U16474 ( .A1(n20651), .A2(n16730), .B1(n20618), .B2(n13045), .C1(
        n15483), .C2(n15513), .ZN(P1_U2872) );
  INV_X1 U16475 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15573) );
  AOI22_X1 U16476 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20647), .B1(n20646), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13054) );
  OAI21_X1 U16477 ( .B1(n15573), .B2(n13066), .A(n13054), .ZN(P1_U2916) );
  INV_X1 U16478 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15564) );
  AOI22_X1 U16479 ( .A1(n20647), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13055) );
  OAI21_X1 U16480 ( .B1(n15564), .B2(n13066), .A(n13055), .ZN(P1_U2914) );
  INV_X1 U16481 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U16482 ( .A1(n21029), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13056) );
  OAI21_X1 U16483 ( .B1(n13057), .B2(n13066), .A(n13056), .ZN(P1_U2917) );
  INV_X1 U16484 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U16485 ( .A1(n21029), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13058) );
  OAI21_X1 U16486 ( .B1(n13059), .B2(n13066), .A(n13058), .ZN(P1_U2915) );
  INV_X1 U16487 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n21327) );
  AOI22_X1 U16488 ( .A1(n21029), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13060) );
  OAI21_X1 U16489 ( .B1(n21327), .B2(n13066), .A(n13060), .ZN(P1_U2919) );
  INV_X1 U16490 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U16491 ( .A1(n21029), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13061) );
  OAI21_X1 U16492 ( .B1(n13062), .B2(n13066), .A(n13061), .ZN(P1_U2918) );
  INV_X1 U16493 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16494 ( .A1(n21029), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13063) );
  OAI21_X1 U16495 ( .B1(n13064), .B2(n13066), .A(n13063), .ZN(P1_U2913) );
  AOI22_X1 U16496 ( .A1(n21029), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13065) );
  OAI21_X1 U16497 ( .B1(n15593), .B2(n13066), .A(n13065), .ZN(P1_U2920) );
  AOI21_X1 U16498 ( .B1(n13587), .B2(n16666), .A(n20943), .ZN(n13067) );
  NAND2_X1 U16499 ( .A1(n15281), .A2(n13067), .ZN(n13073) );
  OAI21_X1 U16500 ( .B1(n13587), .B2(n13068), .A(n21028), .ZN(n13833) );
  INV_X1 U16501 ( .A(n13833), .ZN(n13069) );
  NAND2_X1 U16502 ( .A1(n12810), .A2(n13069), .ZN(n13070) );
  NAND3_X1 U16503 ( .A1(n13070), .A2(n13832), .A3(n15108), .ZN(n13071) );
  NAND2_X1 U16504 ( .A1(n16614), .A2(n13071), .ZN(n13072) );
  MUX2_X1 U16505 ( .A(n13073), .B(n13072), .S(n13097), .Z(n13076) );
  OR3_X1 U16506 ( .A1(n16614), .A2(n12764), .A3(n12761), .ZN(n13074) );
  NAND3_X1 U16507 ( .A1(n13076), .A2(n13075), .A3(n13074), .ZN(n13078) );
  INV_X1 U16508 ( .A(n13117), .ZN(n13084) );
  OAI21_X1 U16509 ( .B1(n13107), .B2(n13079), .A(n15275), .ZN(n13080) );
  NOR2_X1 U16510 ( .A1(n15274), .A2(n13080), .ZN(n13081) );
  AND2_X1 U16511 ( .A1(n13082), .A2(n13081), .ZN(n13083) );
  AOI22_X1 U16512 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16513 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U16514 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9710), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U16515 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13087) );
  NAND4_X1 U16516 ( .A1(n13090), .A2(n13089), .A3(n13088), .A4(n13087), .ZN(
        n13096) );
  AOI22_X1 U16517 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15082), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U16518 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16519 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16520 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13091) );
  NAND4_X1 U16521 ( .A1(n13094), .A2(n13093), .A3(n13092), .A4(n13091), .ZN(
        n13095) );
  XNOR2_X1 U16522 ( .A(n13195), .B(n13194), .ZN(n13098) );
  OAI211_X1 U16523 ( .C1(n13098), .C2(n16636), .A(n13097), .B(n15107), .ZN(
        n13099) );
  INV_X1 U16524 ( .A(n13099), .ZN(n13100) );
  NAND2_X1 U16525 ( .A1(n10328), .A2(n13100), .ZN(n13164) );
  XOR2_X1 U16526 ( .A(n13162), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n13157) );
  OAI211_X1 U16527 ( .C1(n13103), .C2(n13832), .A(n13102), .B(n13101), .ZN(
        n13104) );
  INV_X1 U16528 ( .A(n13105), .ZN(n15278) );
  INV_X1 U16529 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14736) );
  NAND2_X1 U16530 ( .A1(n13210), .A2(n14736), .ZN(n13115) );
  NAND2_X1 U16531 ( .A1(n12810), .A2(n14536), .ZN(n13106) );
  OAI21_X1 U16532 ( .B1(n13107), .B2(n13547), .A(n13106), .ZN(n13108) );
  INV_X1 U16533 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n20617) );
  NAND2_X1 U16534 ( .A1(n15146), .A2(n20617), .ZN(n13111) );
  NAND2_X1 U16535 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13109) );
  OAI211_X1 U16536 ( .C1(n9691), .C2(P1_EBX_REG_1__SCAN_IN), .A(n15149), .B(
        n13109), .ZN(n13110) );
  NAND2_X1 U16537 ( .A1(n13111), .A2(n13110), .ZN(n13203) );
  XNOR2_X1 U16538 ( .A(n13203), .B(n13112), .ZN(n13849) );
  XNOR2_X1 U16539 ( .A(n13849), .B(n15162), .ZN(n20614) );
  INV_X1 U16540 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21016) );
  NOR2_X1 U16541 ( .A1(n16808), .A2(n21016), .ZN(n13113) );
  AOI21_X1 U16542 ( .B1(n16857), .B2(n20614), .A(n13113), .ZN(n13114) );
  OAI21_X1 U16543 ( .B1(n15871), .B2(n13115), .A(n13114), .ZN(n13121) );
  NAND2_X1 U16544 ( .A1(n20656), .A2(n10008), .ZN(n13119) );
  OR2_X1 U16545 ( .A1(n13117), .A2(n13116), .ZN(n13118) );
  NAND2_X1 U16546 ( .A1(n15914), .A2(n10008), .ZN(n20661) );
  AOI21_X1 U16547 ( .B1(n15228), .B2(n20661), .A(n14736), .ZN(n13120) );
  AOI211_X1 U16548 ( .C1(n16861), .C2(n13157), .A(n13121), .B(n13120), .ZN(
        n13122) );
  INV_X1 U16549 ( .A(n13122), .ZN(P1_U3030) );
  NAND2_X1 U16550 ( .A1(n13123), .A2(n13382), .ZN(n13125) );
  AND2_X2 U16551 ( .A1(n13125), .A2(n13124), .ZN(n19712) );
  NAND2_X1 U16552 ( .A1(n19712), .A2(n19905), .ZN(n19713) );
  INV_X1 U16553 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n21322) );
  MUX2_X1 U16554 ( .A(n21322), .B(n15264), .S(n19712), .Z(n13126) );
  OAI21_X1 U16555 ( .B1(n20487), .B2(n19713), .A(n13126), .ZN(P2_U2887) );
  XOR2_X1 U16556 ( .A(n13127), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .Z(n13132)
         );
  AND2_X1 U16557 ( .A1(n13306), .A2(n13128), .ZN(n13129) );
  OR2_X1 U16558 ( .A1(n13129), .A2(n13320), .ZN(n14282) );
  NOR2_X1 U16559 ( .A1(n14282), .A2(n19716), .ZN(n13130) );
  AOI21_X1 U16560 ( .B1(P2_EBX_REG_6__SCAN_IN), .B2(n19716), .A(n13130), .ZN(
        n13131) );
  OAI21_X1 U16561 ( .B1(n13132), .B2(n19713), .A(n13131), .ZN(P2_U2881) );
  INV_X1 U16562 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13133) );
  MUX2_X1 U16563 ( .A(n13133), .B(n19869), .S(n19712), .Z(n13134) );
  OAI21_X1 U16564 ( .B1(n20466), .B2(n19713), .A(n13134), .ZN(P2_U2885) );
  NAND2_X1 U16565 ( .A1(n13971), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13136) );
  NOR2_X1 U16566 ( .A1(n13832), .A2(n9922), .ZN(n13187) );
  NAND2_X1 U16567 ( .A1(n13187), .A2(n13195), .ZN(n13135) );
  XNOR2_X1 U16568 ( .A(n13170), .B(n13168), .ZN(n13142) );
  NAND2_X1 U16569 ( .A1(n13139), .A2(n12908), .ZN(n13141) );
  INV_X1 U16570 ( .A(n13142), .ZN(n13145) );
  INV_X1 U16571 ( .A(n13143), .ZN(n13144) );
  NAND2_X1 U16572 ( .A1(n13145), .A2(n13144), .ZN(n13146) );
  NAND2_X1 U16573 ( .A1(n13540), .A2(n14780), .ZN(n13150) );
  AOI22_X1 U16574 ( .A1(n15246), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n14046), .ZN(n13147) );
  AND2_X1 U16575 ( .A1(n13148), .A2(n13147), .ZN(n13149) );
  INV_X1 U16576 ( .A(n13151), .ZN(n13152) );
  NAND2_X1 U16577 ( .A1(n14046), .A2(n20514), .ZN(n15101) );
  NAND2_X1 U16578 ( .A1(n13152), .A2(n14983), .ZN(n13153) );
  NAND2_X1 U16579 ( .A1(n13154), .A2(n13153), .ZN(n13155) );
  NAND2_X1 U16580 ( .A1(n13156), .A2(n13155), .ZN(n13330) );
  OAI21_X1 U16581 ( .B1(n13156), .B2(n13155), .A(n13330), .ZN(n20613) );
  NAND2_X1 U16582 ( .A1(n13157), .A2(n16772), .ZN(n13161) );
  INV_X1 U16583 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13842) );
  OAI22_X1 U16584 ( .A1(n16774), .A2(n13842), .B1(n16808), .B2(n21016), .ZN(
        n13159) );
  AOI21_X1 U16585 ( .B1(n16742), .B2(n13842), .A(n13159), .ZN(n13160) );
  OAI211_X1 U16586 ( .C1(n16770), .C2(n20613), .A(n13161), .B(n13160), .ZN(
        P1_U2998) );
  INV_X1 U16587 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n21256) );
  OAI222_X1 U16588 ( .A1(n20613), .A2(n15614), .B1(n15608), .B2(n13586), .C1(
        n15606), .C2(n21256), .ZN(P1_U2903) );
  NAND2_X1 U16589 ( .A1(n13162), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13167) );
  INV_X1 U16590 ( .A(n13163), .ZN(n13165) );
  NAND2_X1 U16591 ( .A1(n13165), .A2(n13164), .ZN(n13166) );
  INV_X1 U16592 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13211) );
  INV_X1 U16593 ( .A(n13168), .ZN(n13169) );
  AOI22_X1 U16594 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13178) );
  AOI22_X1 U16595 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13177) );
  AOI22_X1 U16596 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9710), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13176) );
  AOI22_X1 U16597 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13175) );
  NAND4_X1 U16598 ( .A1(n13178), .A2(n13177), .A3(n13176), .A4(n13175), .ZN(
        n13184) );
  AOI22_X1 U16599 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15040), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U16600 ( .A1(n14947), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U16601 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U16602 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13179) );
  NAND4_X1 U16603 ( .A1(n13182), .A2(n13181), .A3(n13180), .A4(n13179), .ZN(
        n13183) );
  INV_X1 U16604 ( .A(n13185), .ZN(n13186) );
  INV_X1 U16605 ( .A(n13187), .ZN(n13189) );
  INV_X1 U16606 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13188) );
  OAI22_X1 U16607 ( .A1(n13189), .A2(n13197), .B1(n14103), .B2(n13188), .ZN(
        n13190) );
  NAND2_X1 U16608 ( .A1(n13195), .A2(n13194), .ZN(n13196) );
  NAND2_X1 U16609 ( .A1(n13196), .A2(n13197), .ZN(n13814) );
  OAI21_X1 U16610 ( .B1(n13197), .B2(n13196), .A(n13814), .ZN(n13200) );
  INV_X1 U16611 ( .A(n13198), .ZN(n13199) );
  AOI21_X1 U16612 ( .B1(n13200), .B2(n14536), .A(n13199), .ZN(n13201) );
  NAND2_X1 U16613 ( .A1(n13202), .A2(n13201), .ZN(n13450) );
  XNOR2_X1 U16614 ( .A(n13449), .B(n13450), .ZN(n13335) );
  INV_X1 U16615 ( .A(n15224), .ZN(n15909) );
  OAI21_X1 U16616 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n15909), .A(
        n15228), .ZN(n13209) );
  NAND2_X1 U16617 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15222) );
  NOR3_X1 U16618 ( .A1(n10008), .A2(n15222), .A3(n15863), .ZN(n13208) );
  AOI21_X1 U16619 ( .B1(n13849), .B2(n15162), .A(n13203), .ZN(n13270) );
  MUX2_X1 U16620 ( .A(n15159), .B(n15147), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13204) );
  OAI21_X1 U16621 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n15218), .A(
        n13204), .ZN(n13205) );
  INV_X1 U16622 ( .A(n13205), .ZN(n13269) );
  XNOR2_X1 U16623 ( .A(n13270), .B(n13269), .ZN(n13945) );
  NAND2_X1 U16624 ( .A1(n13116), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13206) );
  AOI21_X1 U16625 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14425) );
  NAND2_X1 U16626 ( .A1(n15914), .A2(n14425), .ZN(n13455) );
  OAI211_X1 U16627 ( .C1(n20652), .C2(n13945), .A(n13206), .B(n13455), .ZN(
        n13207) );
  AOI211_X1 U16628 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n13209), .A(
        n13208), .B(n13207), .ZN(n13214) );
  NAND2_X1 U16629 ( .A1(n15224), .A2(n13210), .ZN(n15846) );
  INV_X1 U16630 ( .A(n15846), .ZN(n13212) );
  NAND3_X1 U16631 ( .A1(n13212), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13211), .ZN(n13213) );
  OAI211_X1 U16632 ( .C1(n13335), .C2(n20653), .A(n13214), .B(n13213), .ZN(
        P1_U3029) );
  NAND2_X1 U16633 ( .A1(n19749), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20072) );
  OAI21_X1 U16634 ( .B1(n20072), .B2(n20260), .A(n20458), .ZN(n13230) );
  NAND3_X1 U16635 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20463), .A3(
        n20481), .ZN(n19992) );
  INV_X1 U16636 ( .A(n19992), .ZN(n13222) );
  NAND2_X1 U16637 ( .A1(n16542), .A2(n17100), .ZN(n17095) );
  NAND2_X1 U16638 ( .A1(n17096), .A2(n20484), .ZN(n13220) );
  NOR2_X1 U16639 ( .A1(n20492), .A2(n19992), .ZN(n20044) );
  INV_X1 U16640 ( .A(n20044), .ZN(n13226) );
  OAI211_X1 U16641 ( .C1(n10764), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n13226), 
        .B(n20133), .ZN(n13221) );
  OAI211_X1 U16642 ( .C1(n13230), .C2(n13222), .A(n20320), .B(n13221), .ZN(
        n20035) );
  INV_X1 U16643 ( .A(n20035), .ZN(n13235) );
  NOR2_X1 U16644 ( .A1(n20133), .A2(n21150), .ZN(n20471) );
  AOI22_X1 U16645 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19909), .ZN(n20176) );
  AOI22_X1 U16646 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19909), .ZN(n20325) );
  NAND2_X1 U16647 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20320), .ZN(n19890) );
  INV_X1 U16648 ( .A(n20314), .ZN(n13651) );
  OAI22_X1 U16649 ( .A1(n20325), .A2(n20066), .B1(n13651), .B2(n13226), .ZN(
        n13227) );
  AOI21_X1 U16650 ( .B1(n20322), .B2(n20022), .A(n13227), .ZN(n13233) );
  INV_X1 U16651 ( .A(n10764), .ZN(n13228) );
  OAI21_X1 U16652 ( .B1(n13228), .B2(n20044), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13229) );
  OAI21_X1 U16653 ( .B1(n13230), .B2(n19992), .A(n13229), .ZN(n20034) );
  NAND2_X1 U16654 ( .A1(n20034), .A2(n13231), .ZN(n13232) );
  OAI211_X1 U16655 ( .C1(n13235), .C2(n13234), .A(n13233), .B(n13232), .ZN(
        P2_U3088) );
  INV_X1 U16656 ( .A(n13330), .ZN(n13240) );
  XNOR2_X1 U16657 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13943) );
  AOI21_X1 U16658 ( .B1(n14983), .B2(n13943), .A(n15245), .ZN(n13237) );
  NAND2_X1 U16659 ( .A1(n15246), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n13236) );
  OAI211_X1 U16660 ( .C1(n13263), .C2(n12434), .A(n13237), .B(n13236), .ZN(
        n13238) );
  INV_X1 U16661 ( .A(n13238), .ZN(n13239) );
  OAI21_X2 U16662 ( .B1(n13539), .B2(n14797), .A(n13239), .ZN(n13327) );
  NAND2_X1 U16663 ( .A1(n13240), .A2(n13327), .ZN(n13328) );
  NAND2_X1 U16664 ( .A1(n15245), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13326) );
  AOI22_X1 U16665 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14908), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U16666 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U16667 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16668 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13241) );
  NAND4_X1 U16669 ( .A1(n13244), .A2(n13243), .A3(n13242), .A4(n13241), .ZN(
        n13250) );
  AOI22_X1 U16670 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U16671 ( .A1(n15083), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16672 ( .A1(n15082), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U16673 ( .A1(n9710), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13245) );
  NAND4_X1 U16674 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        n13249) );
  AOI22_X1 U16675 ( .A1(n13972), .A2(n13813), .B1(n13971), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13251) );
  NAND2_X1 U16676 ( .A1(n13254), .A2(n13640), .ZN(n13255) );
  INV_X1 U16677 ( .A(n13256), .ZN(n13259) );
  INV_X1 U16678 ( .A(n13618), .ZN(n13258) );
  OAI21_X1 U16679 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13259), .A(
        n13258), .ZN(n20603) );
  AOI22_X1 U16680 ( .A1(n14983), .A2(n20603), .B1(n15245), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13261) );
  NAND2_X1 U16681 ( .A1(n15246), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n13260) );
  OAI211_X1 U16682 ( .C1(n13263), .C2(n13262), .A(n13261), .B(n13260), .ZN(
        n13264) );
  INV_X1 U16683 ( .A(n13264), .ZN(n13265) );
  OAI21_X2 U16684 ( .B1(n13637), .B2(n14797), .A(n13265), .ZN(n13267) );
  NAND2_X1 U16685 ( .A1(n13268), .A2(n13267), .ZN(n13623) );
  OAI21_X1 U16686 ( .B1(n13268), .B2(n13267), .A(n13266), .ZN(n13498) );
  OR2_X1 U16687 ( .A1(n15165), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n13276) );
  INV_X1 U16688 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13852) );
  NAND2_X1 U16689 ( .A1(n15149), .A2(n13852), .ZN(n13274) );
  INV_X1 U16690 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13272) );
  NAND2_X1 U16691 ( .A1(n15162), .A2(n13272), .ZN(n13273) );
  NAND3_X1 U16692 ( .A1(n13274), .A2(n15129), .A3(n13273), .ZN(n13275) );
  NAND2_X1 U16693 ( .A1(n13276), .A2(n13275), .ZN(n13277) );
  NAND2_X1 U16694 ( .A1(n13278), .A2(n13277), .ZN(n13633) );
  OR2_X1 U16695 ( .A1(n13278), .A2(n13277), .ZN(n13279) );
  NAND2_X1 U16696 ( .A1(n13633), .A2(n13279), .ZN(n13456) );
  INV_X1 U16697 ( .A(n13456), .ZN(n20594) );
  AOI22_X1 U16698 ( .A1(n21040), .A2(n20594), .B1(n21041), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13280) );
  OAI21_X1 U16699 ( .B1(n13498), .B2(n15513), .A(n13280), .ZN(P1_U2869) );
  INV_X1 U16700 ( .A(n19749), .ZN(n20460) );
  AOI21_X1 U16701 ( .B1(n20460), .B2(n16970), .A(n13281), .ZN(n13282) );
  INV_X1 U16702 ( .A(n13282), .ZN(P2_U2884) );
  NAND2_X1 U16703 ( .A1(n20478), .A2(n16970), .ZN(n13284) );
  NAND2_X1 U16704 ( .A1(n9706), .A2(n19712), .ZN(n13283) );
  OAI211_X1 U16705 ( .C1(n19712), .C2(n19693), .A(n13284), .B(n13283), .ZN(
        P2_U2886) );
  INV_X1 U16706 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20641) );
  OAI222_X1 U16707 ( .A1(n13498), .A2(n15614), .B1(n15608), .B2(n13570), .C1(
        n15606), .C2(n20641), .ZN(P1_U2901) );
  OR2_X1 U16708 ( .A1(n13322), .A2(n13285), .ZN(n13286) );
  NAND2_X1 U16709 ( .A1(n13286), .A2(n13296), .ZN(n19662) );
  INV_X1 U16710 ( .A(n19662), .ZN(n17025) );
  NOR2_X1 U16711 ( .A1(n19712), .A2(n11069), .ZN(n13292) );
  AOI211_X1 U16712 ( .C1(n13290), .C2(n13288), .A(n19713), .B(n13289), .ZN(
        n13291) );
  AOI211_X1 U16713 ( .C1(n17025), .C2(n19712), .A(n13292), .B(n13291), .ZN(
        n13293) );
  INV_X1 U16714 ( .A(n13293), .ZN(P2_U2879) );
  OAI211_X1 U16715 ( .C1(n13289), .C2(n13295), .A(n13294), .B(n16970), .ZN(
        n13301) );
  NAND2_X1 U16716 ( .A1(n13297), .A2(n13296), .ZN(n13299) );
  INV_X1 U16717 ( .A(n13312), .ZN(n13298) );
  AND2_X1 U16718 ( .A1(n13299), .A2(n13298), .ZN(n17019) );
  NAND2_X1 U16719 ( .A1(n19712), .A2(n17019), .ZN(n13300) );
  OAI211_X1 U16720 ( .C1(n19712), .C2(n13302), .A(n13301), .B(n13300), .ZN(
        P2_U2878) );
  OAI211_X1 U16721 ( .C1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .C2(n19665), .A(
        n13127), .B(n16970), .ZN(n13308) );
  NAND2_X1 U16722 ( .A1(n13303), .A2(n13304), .ZN(n13305) );
  AND2_X1 U16723 ( .A1(n13306), .A2(n13305), .ZN(n17033) );
  NAND2_X1 U16724 ( .A1(n17033), .A2(n19712), .ZN(n13307) );
  OAI211_X1 U16725 ( .C1(n19712), .C2(n13309), .A(n13308), .B(n13307), .ZN(
        P2_U2882) );
  OAI211_X1 U16726 ( .C1(n11606), .C2(n11605), .A(n16970), .B(n13311), .ZN(
        n13316) );
  NOR2_X1 U16727 ( .A1(n13313), .A2(n13312), .ZN(n13314) );
  NOR2_X1 U16728 ( .A1(n13314), .A2(n13474), .ZN(n19646) );
  NAND2_X1 U16729 ( .A1(n19712), .A2(n19646), .ZN(n13315) );
  OAI211_X1 U16730 ( .C1(n19712), .C2(n10104), .A(n13316), .B(n13315), .ZN(
        P2_U2877) );
  NOR2_X1 U16731 ( .A1(n13127), .A2(n13317), .ZN(n13318) );
  OAI211_X1 U16732 ( .C1(n13318), .C2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n16970), .B(n13288), .ZN(n13324) );
  NOR2_X1 U16733 ( .A1(n13320), .A2(n13319), .ZN(n13321) );
  OR2_X1 U16734 ( .A1(n13322), .A2(n13321), .ZN(n14298) );
  INV_X1 U16735 ( .A(n14298), .ZN(n14484) );
  NAND2_X1 U16736 ( .A1(n14484), .A2(n19712), .ZN(n13323) );
  OAI211_X1 U16737 ( .C1(n19712), .C2(n13325), .A(n13324), .B(n13323), .ZN(
        P2_U2880) );
  NAND2_X1 U16738 ( .A1(n13327), .A2(n13326), .ZN(n13331) );
  INV_X1 U16739 ( .A(n13328), .ZN(n13329) );
  AOI21_X1 U16740 ( .B1(n13331), .B2(n13330), .A(n13329), .ZN(n13956) );
  AOI22_X1 U16741 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13332) );
  OAI21_X1 U16742 ( .B1(n13943), .B2(n16769), .A(n13332), .ZN(n13333) );
  AOI21_X1 U16743 ( .B1(n13956), .B2(n16764), .A(n13333), .ZN(n13334) );
  OAI21_X1 U16744 ( .B1(n20516), .B2(n13335), .A(n13334), .ZN(P1_U2997) );
  NOR2_X2 U16745 ( .A1(n20166), .A2(n20260), .ZN(n20280) );
  OAI21_X1 U16746 ( .B1(n20280), .B2(n20250), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13340) );
  NOR2_X1 U16747 ( .A1(n13336), .A2(n19942), .ZN(n19990) );
  NAND2_X1 U16748 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19990), .ZN(
        n13339) );
  AOI21_X1 U16749 ( .B1(n13341), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13337) );
  NAND3_X1 U16750 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20481), .ZN(n20259) );
  NOR2_X1 U16751 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20259), .ZN(
        n20248) );
  OAI21_X1 U16752 ( .B1(n13337), .B2(n20248), .A(n20320), .ZN(n13338) );
  INV_X1 U16753 ( .A(n20325), .ZN(n20173) );
  AOI22_X1 U16754 ( .A1(n20280), .A2(n20173), .B1(n20250), .B2(n20322), .ZN(
        n13346) );
  INV_X1 U16755 ( .A(n19990), .ZN(n13343) );
  OAI21_X1 U16756 ( .B1(n10601), .B2(n20248), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13342) );
  OAI21_X1 U16757 ( .B1(n13344), .B2(n13343), .A(n13342), .ZN(n20249) );
  AOI22_X1 U16758 ( .A1(n20249), .A2(n13231), .B1(n20314), .B2(n20248), .ZN(
        n13345) );
  OAI211_X1 U16759 ( .C1(n20254), .C2(n13347), .A(n13346), .B(n13345), .ZN(
        P2_U3144) );
  INV_X1 U16760 ( .A(n13956), .ZN(n13471) );
  INV_X1 U16761 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20643) );
  OAI222_X1 U16762 ( .A1(n13471), .A2(n15614), .B1(n15608), .B2(n13557), .C1(
        n15606), .C2(n20643), .ZN(P1_U2902) );
  NAND2_X1 U16763 ( .A1(n13349), .A2(n13348), .ZN(n13351) );
  XNOR2_X1 U16764 ( .A(n13351), .B(n13350), .ZN(n17042) );
  NOR2_X1 U16765 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16432), .ZN(
        n13365) );
  OR2_X1 U16766 ( .A1(n13353), .A2(n13352), .ZN(n13354) );
  NAND2_X1 U16767 ( .A1(n13354), .A2(n13490), .ZN(n19748) );
  INV_X1 U16768 ( .A(n19748), .ZN(n20459) );
  OAI22_X1 U16769 ( .A1(n19856), .A2(n13356), .B1(n14086), .B2(n13355), .ZN(
        n13357) );
  AOI21_X1 U16770 ( .B1(n20459), .B2(n19854), .A(n13357), .ZN(n13358) );
  OAI21_X1 U16771 ( .B1(n13359), .B2(n19870), .A(n13358), .ZN(n13363) );
  NOR2_X1 U16772 ( .A1(n9797), .A2(n13360), .ZN(n17041) );
  INV_X1 U16773 ( .A(n13361), .ZN(n17040) );
  NOR3_X1 U16774 ( .A1(n17041), .A2(n17040), .A3(n19859), .ZN(n13362) );
  AOI211_X1 U16775 ( .C1(n13365), .C2(n13364), .A(n13363), .B(n13362), .ZN(
        n13366) );
  OAI21_X1 U16776 ( .B1(n17042), .B2(n16500), .A(n13366), .ZN(P2_U3043) );
  OR2_X1 U16777 ( .A1(n20072), .A2(n20209), .ZN(n13367) );
  AND2_X1 U16778 ( .A1(n13367), .A2(n20458), .ZN(n13373) );
  NOR2_X1 U16779 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19941) );
  NAND2_X1 U16780 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19941), .ZN(
        n13377) );
  NAND2_X1 U16781 ( .A1(n13373), .A2(n13377), .ZN(n13371) );
  INV_X1 U16782 ( .A(n20203), .ZN(n13368) );
  NAND2_X1 U16783 ( .A1(n13368), .A2(n19941), .ZN(n13374) );
  OAI211_X1 U16784 ( .C1(n10767), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n13374), 
        .B(n20133), .ZN(n13369) );
  AND2_X1 U16785 ( .A1(n13369), .A2(n20320), .ZN(n13370) );
  NAND2_X1 U16786 ( .A1(n13371), .A2(n13370), .ZN(n19986) );
  INV_X1 U16787 ( .A(n19986), .ZN(n19974) );
  INV_X1 U16788 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13381) );
  OAI22_X1 U16789 ( .A1(n20325), .A2(n20019), .B1(n13651), .B2(n13374), .ZN(
        n13372) );
  AOI21_X1 U16790 ( .B1(n20322), .B2(n19981), .A(n13372), .ZN(n13380) );
  INV_X1 U16791 ( .A(n13373), .ZN(n13378) );
  INV_X1 U16792 ( .A(n10767), .ZN(n13375) );
  INV_X1 U16793 ( .A(n13374), .ZN(n19984) );
  OAI21_X1 U16794 ( .B1(n13375), .B2(n19984), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13376) );
  OAI21_X1 U16795 ( .B1(n13378), .B2(n13377), .A(n13376), .ZN(n19985) );
  NAND2_X1 U16796 ( .A1(n19985), .A2(n13231), .ZN(n13379) );
  OAI211_X1 U16797 ( .C1(n19974), .C2(n13381), .A(n13380), .B(n13379), .ZN(
        P2_U3072) );
  INV_X1 U16798 ( .A(n13410), .ZN(n13409) );
  INV_X1 U16799 ( .A(n13382), .ZN(n13383) );
  NOR2_X1 U16800 ( .A1(n13384), .A2(n13383), .ZN(n13397) );
  NAND2_X1 U16801 ( .A1(n13413), .A2(n9973), .ZN(n13407) );
  NOR2_X1 U16802 ( .A1(n10578), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13392) );
  AOI21_X1 U16803 ( .B1(n13413), .B2(n10346), .A(n13392), .ZN(n13385) );
  OAI211_X1 U16804 ( .C1(n10449), .C2(n13397), .A(n13407), .B(n13385), .ZN(
        n13389) );
  NOR2_X1 U16805 ( .A1(n13427), .A2(n13423), .ZN(n13396) );
  NAND3_X1 U16806 ( .A1(n13413), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13386) );
  OAI21_X1 U16807 ( .B1(n13396), .B2(n13392), .A(n13386), .ZN(n13388) );
  MUX2_X1 U16808 ( .A(n13389), .B(n13388), .S(n13387), .Z(n13390) );
  MUX2_X1 U16809 ( .A(n13387), .B(n16551), .S(n13437), .Z(n13439) );
  INV_X1 U16810 ( .A(n13392), .ZN(n13394) );
  NAND2_X1 U16811 ( .A1(n13394), .A2(n13393), .ZN(n13395) );
  MUX2_X1 U16812 ( .A(n13397), .B(n13396), .S(n13395), .Z(n13400) );
  NAND2_X1 U16813 ( .A1(n13413), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13398) );
  MUX2_X1 U16814 ( .A(n13407), .B(n13398), .S(n10346), .Z(n13399) );
  OAI211_X1 U16815 ( .C1(n19869), .C2(n13410), .A(n13400), .B(n13399), .ZN(
        n16548) );
  NAND2_X1 U16816 ( .A1(n13402), .A2(n10346), .ZN(n13401) );
  OAI21_X1 U16817 ( .B1(n16548), .B2(n13402), .A(n13401), .ZN(n13438) );
  NOR2_X1 U16818 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13438), .ZN(
        n13421) );
  NAND2_X1 U16819 ( .A1(n13404), .A2(n13403), .ZN(n13412) );
  NOR2_X1 U16820 ( .A1(n10586), .A2(n10578), .ZN(n13405) );
  NAND2_X1 U16821 ( .A1(n13412), .A2(n13405), .ZN(n13406) );
  NAND2_X1 U16822 ( .A1(n13407), .A2(n13406), .ZN(n13408) );
  AOI21_X1 U16823 ( .B1(n9706), .B2(n13409), .A(n13408), .ZN(n16540) );
  INV_X1 U16824 ( .A(n16540), .ZN(n13417) );
  OR2_X1 U16825 ( .A1(n15264), .A2(n13410), .ZN(n13416) );
  MUX2_X1 U16826 ( .A(n13413), .B(n13412), .S(n13411), .Z(n13414) );
  INV_X1 U16827 ( .A(n13414), .ZN(n13415) );
  NAND2_X1 U16828 ( .A1(n13416), .A2(n13415), .ZN(n16530) );
  AOI211_X1 U16829 ( .C1(n13417), .C2(n20481), .A(n20492), .B(n16530), .ZN(
        n13419) );
  OAI21_X1 U16830 ( .B1(n13417), .B2(n20481), .A(n13437), .ZN(n13418) );
  AOI211_X1 U16831 ( .C1(n16551), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n13419), .B(n13418), .ZN(n13420) );
  AOI222_X1 U16832 ( .A1(n13421), .A2(n13420), .B1(n13421), .B2(n20470), .C1(
        n13420), .C2(n20470), .ZN(n13422) );
  OAI21_X1 U16833 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13439), .A(
        n13422), .ZN(n13442) );
  INV_X1 U16834 ( .A(n13423), .ZN(n13425) );
  OAI22_X1 U16835 ( .A1(n13428), .A2(n13425), .B1(n11403), .B2(n13424), .ZN(
        n13426) );
  AOI21_X1 U16836 ( .B1(n13428), .B2(n13427), .A(n13426), .ZN(n20500) );
  INV_X1 U16837 ( .A(n11011), .ZN(n13430) );
  AOI22_X1 U16838 ( .A1(n13431), .A2(n9812), .B1(n13430), .B2(n13429), .ZN(
        n13436) );
  NOR4_X1 U16839 ( .A1(n11403), .A2(n13434), .A3(n13433), .A4(n13432), .ZN(
        n19562) );
  OAI21_X1 U16840 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19562), .ZN(n13435) );
  NAND3_X1 U16841 ( .A1(n20500), .A2(n13436), .A3(n13435), .ZN(n13441) );
  OAI22_X1 U16842 ( .A1(n13439), .A2(n13438), .B1(n21165), .B2(n13437), .ZN(
        n13440) );
  AOI211_X1 U16843 ( .C1(n21126), .C2(n13442), .A(n13441), .B(n13440), .ZN(
        n17106) );
  AOI21_X1 U16844 ( .B1(n17106), .B2(n11007), .A(n17100), .ZN(n13448) );
  NOR4_X1 U16845 ( .A1(n13445), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n13444), 
        .A4(n13443), .ZN(n13447) );
  NOR2_X1 U16846 ( .A1(n17101), .A2(n17100), .ZN(n17099) );
  INV_X1 U16847 ( .A(n17094), .ZN(n16678) );
  OAI21_X1 U16848 ( .B1(n17099), .B2(n20101), .A(n16678), .ZN(P2_U3593) );
  NAND2_X1 U16849 ( .A1(n13450), .A2(n13449), .ZN(n13453) );
  NAND2_X1 U16850 ( .A1(n13451), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13452) );
  XNOR2_X1 U16851 ( .A(n13814), .B(n13813), .ZN(n13454) );
  OAI22_X1 U16852 ( .A1(n13637), .A2(n14401), .B1(n16636), .B2(n13454), .ZN(
        n13807) );
  XNOR2_X1 U16853 ( .A(n13808), .B(n13807), .ZN(n13502) );
  NOR2_X1 U16854 ( .A1(n15234), .A2(n15914), .ZN(n15896) );
  NOR2_X1 U16855 ( .A1(n14425), .A2(n15896), .ZN(n16872) );
  AOI21_X1 U16856 ( .B1(n15222), .B2(n15224), .A(n20658), .ZN(n16822) );
  NAND2_X1 U16857 ( .A1(n16822), .A2(n13455), .ZN(n13855) );
  INV_X1 U16858 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20955) );
  OAI22_X1 U16859 ( .A1(n16808), .A2(n20955), .B1(n20652), .B2(n13456), .ZN(
        n13457) );
  AOI221_X1 U16860 ( .B1(n16872), .B2(n13852), .C1(n13855), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n13457), .ZN(n13458) );
  OAI21_X1 U16861 ( .B1(n20653), .B2(n13502), .A(n13458), .ZN(P1_U3028) );
  NOR3_X1 U16862 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n17100), .A3(n20373), 
        .ZN(n17093) );
  AOI21_X1 U16863 ( .B1(n17101), .B2(n20385), .A(n17093), .ZN(n13463) );
  INV_X1 U16864 ( .A(n17101), .ZN(n13461) );
  OAI21_X1 U16865 ( .B1(n20385), .B2(n19558), .A(n19561), .ZN(n13459) );
  NAND3_X1 U16866 ( .A1(n13461), .A2(n13460), .A3(n13459), .ZN(n13462) );
  OAI211_X1 U16867 ( .C1(n13463), .C2(n11007), .A(n19704), .B(n13462), .ZN(
        P2_U3177) );
  INV_X1 U16868 ( .A(n13465), .ZN(n13466) );
  OAI211_X1 U16869 ( .C1(n13464), .C2(n13467), .A(n13466), .B(n16970), .ZN(
        n13470) );
  OAI21_X1 U16870 ( .B1(n13476), .B2(n13468), .A(n13504), .ZN(n19627) );
  INV_X1 U16871 ( .A(n19627), .ZN(n17085) );
  NAND2_X1 U16872 ( .A1(n19712), .A2(n17085), .ZN(n13469) );
  OAI211_X1 U16873 ( .C1(n19712), .C2(n11077), .A(n13470), .B(n13469), .ZN(
        P2_U2875) );
  INV_X1 U16874 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13472) );
  OAI222_X1 U16875 ( .A1(n13945), .A2(n16730), .B1(n20618), .B2(n13472), .C1(
        n15513), .C2(n13471), .ZN(P1_U2870) );
  NOR2_X1 U16876 ( .A1(n13474), .A2(n13473), .ZN(n13475) );
  NOR2_X1 U16877 ( .A1(n13476), .A2(n13475), .ZN(n19637) );
  INV_X1 U16878 ( .A(n19637), .ZN(n13477) );
  NOR2_X1 U16879 ( .A1(n19716), .A2(n13477), .ZN(n13480) );
  AOI211_X1 U16880 ( .C1(n13478), .C2(n13311), .A(n19713), .B(n13464), .ZN(
        n13479) );
  AOI211_X1 U16881 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n19716), .A(n13480), .B(
        n13479), .ZN(n13481) );
  INV_X1 U16882 ( .A(n13481), .ZN(P2_U2876) );
  XOR2_X1 U16883 ( .A(n13482), .B(n13483), .Z(n19827) );
  INV_X1 U16884 ( .A(n19827), .ZN(n13497) );
  XNOR2_X1 U16885 ( .A(n13485), .B(n13675), .ZN(n13486) );
  XNOR2_X1 U16886 ( .A(n13484), .B(n13486), .ZN(n19830) );
  NAND2_X1 U16887 ( .A1(n13488), .A2(n13487), .ZN(n13489) );
  NAND2_X1 U16888 ( .A1(n13303), .A2(n13489), .ZN(n19826) );
  OAI21_X1 U16889 ( .B1(n16432), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n14086), .ZN(n13678) );
  NAND2_X1 U16890 ( .A1(n13678), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13494) );
  AOI21_X1 U16891 ( .B1(n13491), .B2(n13490), .A(n13681), .ZN(n19759) );
  INV_X1 U16892 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20400) );
  NAND2_X1 U16893 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14306), .ZN(
        n13674) );
  OAI22_X1 U16894 ( .A1(n19856), .A2(n20400), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13674), .ZN(n13492) );
  AOI21_X1 U16895 ( .B1(n19854), .B2(n19759), .A(n13492), .ZN(n13493) );
  OAI211_X1 U16896 ( .C1(n19826), .C2(n19870), .A(n13494), .B(n13493), .ZN(
        n13495) );
  AOI21_X1 U16897 ( .B1(n19830), .B2(n11551), .A(n13495), .ZN(n13496) );
  OAI21_X1 U16898 ( .B1(n13497), .B2(n16500), .A(n13496), .ZN(P2_U3042) );
  INV_X1 U16899 ( .A(n13498), .ZN(n20607) );
  AOI22_X1 U16900 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13499) );
  OAI21_X1 U16901 ( .B1(n20603), .B2(n16769), .A(n13499), .ZN(n13500) );
  AOI21_X1 U16902 ( .B1(n20607), .B2(n16764), .A(n13500), .ZN(n13501) );
  OAI21_X1 U16903 ( .B1(n13502), .B2(n20516), .A(n13501), .ZN(P1_U2996) );
  AND2_X1 U16904 ( .A1(n13504), .A2(n13503), .ZN(n13506) );
  OR2_X1 U16905 ( .A1(n13506), .A2(n13505), .ZN(n14494) );
  INV_X2 U16906 ( .A(n19712), .ZN(n19716) );
  OAI211_X1 U16907 ( .C1(n13465), .C2(n13508), .A(n13507), .B(n16970), .ZN(
        n13510) );
  NAND2_X1 U16908 ( .A1(n19716), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13509) );
  OAI211_X1 U16909 ( .C1(n14494), .C2(n19716), .A(n13510), .B(n13509), .ZN(
        P2_U2874) );
  NAND2_X1 U16910 ( .A1(n13511), .A2(n16616), .ZN(n13512) );
  NOR2_X1 U16911 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21133), .ZN(n13528) );
  AOI21_X1 U16912 ( .B1(n13512), .B2(n21133), .A(n13528), .ZN(n13514) );
  AOI21_X1 U16913 ( .B1(n16616), .B2(n21133), .A(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13513) );
  XNOR2_X1 U16914 ( .A(n9712), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13517) );
  XNOR2_X1 U16915 ( .A(n14740), .B(n12434), .ZN(n13518) );
  INV_X1 U16916 ( .A(n13518), .ZN(n21011) );
  AOI22_X1 U16917 ( .A1(n14742), .A2(n13517), .B1(n21011), .B2(n13516), .ZN(
        n13521) );
  NAND3_X1 U16918 ( .A1(n14744), .A2(n13519), .A3(n13518), .ZN(n13520) );
  OAI211_X1 U16919 ( .C1(n13515), .C2(n14744), .A(n13521), .B(n13520), .ZN(
        n21004) );
  NAND2_X1 U16920 ( .A1(n21004), .A2(n16616), .ZN(n13524) );
  INV_X1 U16921 ( .A(n16616), .ZN(n13522) );
  NAND2_X1 U16922 ( .A1(n13522), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13523) );
  NAND2_X1 U16923 ( .A1(n13524), .A2(n13523), .ZN(n16623) );
  NAND2_X1 U16924 ( .A1(n16623), .A2(n21133), .ZN(n13526) );
  NAND2_X1 U16925 ( .A1(n13528), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13525) );
  NAND2_X1 U16926 ( .A1(n13526), .A2(n13525), .ZN(n13531) );
  MUX2_X1 U16927 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13527), .S(
        n16616), .Z(n16627) );
  AOI22_X1 U16928 ( .A1(n13528), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16627), .B2(n21133), .ZN(n13529) );
  INV_X1 U16929 ( .A(n13529), .ZN(n13530) );
  NAND2_X1 U16930 ( .A1(n13531), .A2(n13530), .ZN(n13532) );
  NAND2_X1 U16931 ( .A1(n13534), .A2(n13532), .ZN(n16631) );
  NAND2_X1 U16932 ( .A1(n13534), .A2(n14739), .ZN(n13535) );
  NAND2_X1 U16933 ( .A1(n16631), .A2(n13535), .ZN(n15923) );
  INV_X1 U16934 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20517) );
  NAND2_X1 U16935 ( .A1(n15923), .A2(n20517), .ZN(n13537) );
  NAND2_X1 U16936 ( .A1(n13537), .A2(n13536), .ZN(n13538) );
  NAND2_X1 U16937 ( .A1(n14046), .A2(n21133), .ZN(n16879) );
  INV_X1 U16938 ( .A(n16879), .ZN(n21033) );
  INV_X1 U16939 ( .A(n20663), .ZN(n13643) );
  NAND2_X1 U16940 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n12826), .ZN(n15924) );
  NAND2_X1 U16941 ( .A1(n13643), .A2(n15924), .ZN(n15273) );
  AND2_X1 U16942 ( .A1(n13540), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20733) );
  AOI21_X1 U16943 ( .B1(n13639), .B2(n20733), .A(n20807), .ZN(n14554) );
  OAI21_X1 U16944 ( .B1(n13639), .B2(n20733), .A(n14554), .ZN(n13762) );
  MUX2_X1 U16945 ( .A(n13762), .B(n16622), .S(n20663), .Z(n13541) );
  OAI21_X1 U16946 ( .B1(n15273), .B2(n13515), .A(n13541), .ZN(P1_U3476) );
  INV_X1 U16947 ( .A(n13721), .ZN(n15927) );
  INV_X1 U16948 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19889) );
  INV_X1 U16949 ( .A(DATAI_28_), .ZN(n13542) );
  NAND2_X1 U16950 ( .A1(n16764), .A2(n15105), .ZN(n13593) );
  OAI22_X1 U16951 ( .A1(n19889), .A2(n13592), .B1(n13542), .B2(n13593), .ZN(
        n20906) );
  INV_X1 U16952 ( .A(n20906), .ZN(n20842) );
  INV_X1 U16953 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n21269) );
  INV_X1 U16954 ( .A(DATAI_20_), .ZN(n13543) );
  NOR2_X1 U16955 ( .A1(n13515), .A2(n13544), .ZN(n20776) );
  INV_X1 U16956 ( .A(n13984), .ZN(n13910) );
  NOR3_X1 U16957 ( .A1(n16622), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13552) );
  INV_X1 U16958 ( .A(n13552), .ZN(n14188) );
  NOR2_X1 U16959 ( .A1(n20779), .A2(n14188), .ZN(n13548) );
  AOI21_X1 U16960 ( .B1(n20776), .B2(n13910), .A(n13548), .ZN(n13550) );
  OAI22_X1 U16961 ( .A1(n13550), .A2(n20807), .B1(n14188), .B2(n14046), .ZN(
        n13545) );
  INV_X1 U16962 ( .A(n13545), .ZN(n13598) );
  INV_X1 U16963 ( .A(n15575), .ZN(n13636) );
  NOR2_X1 U16964 ( .A1(n14128), .A2(n13636), .ZN(n13992) );
  NAND2_X1 U16965 ( .A1(n13596), .A2(n13547), .ZN(n20841) );
  INV_X1 U16966 ( .A(n13548), .ZN(n13597) );
  OAI22_X1 U16967 ( .A1(n13598), .A2(n20909), .B1(n20841), .B2(n13597), .ZN(
        n13549) );
  AOI21_X1 U16968 ( .B1(n20801), .B2(n20905), .A(n13549), .ZN(n13554) );
  OR2_X1 U16969 ( .A1(n13540), .A2(n20514), .ZN(n15270) );
  OAI211_X1 U16970 ( .C1(n13722), .C2(n15270), .A(n15926), .B(n13550), .ZN(
        n13551) );
  OAI211_X1 U16971 ( .C1(n15926), .C2(n13552), .A(n13551), .B(n20744), .ZN(
        n13600) );
  NAND2_X1 U16972 ( .A1(n13600), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n13553) );
  OAI211_X1 U16973 ( .C1(n13603), .C2(n20842), .A(n13554), .B(n13553), .ZN(
        P1_U3077) );
  INV_X1 U16974 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n17174) );
  INV_X1 U16975 ( .A(DATAI_26_), .ZN(n13555) );
  OAI22_X1 U16976 ( .A1(n17174), .A2(n13592), .B1(n13555), .B2(n13593), .ZN(
        n20894) );
  INV_X1 U16977 ( .A(n20894), .ZN(n20832) );
  INV_X1 U16978 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n17189) );
  INV_X1 U16979 ( .A(DATAI_18_), .ZN(n13556) );
  NOR2_X1 U16980 ( .A1(n14128), .A2(n13557), .ZN(n14016) );
  NAND2_X1 U16981 ( .A1(n13596), .A2(n13558), .ZN(n20831) );
  OAI22_X1 U16982 ( .A1(n13598), .A2(n20897), .B1(n20831), .B2(n13597), .ZN(
        n13559) );
  AOI21_X1 U16983 ( .B1(n20801), .B2(n20893), .A(n13559), .ZN(n13561) );
  NAND2_X1 U16984 ( .A1(n13600), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n13560) );
  OAI211_X1 U16985 ( .C1(n13603), .C2(n20832), .A(n13561), .B(n13560), .ZN(
        P1_U3075) );
  INV_X1 U16986 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19895) );
  INV_X1 U16987 ( .A(DATAI_30_), .ZN(n13562) );
  OAI22_X1 U16988 ( .A1(n19895), .A2(n13592), .B1(n13562), .B2(n13593), .ZN(
        n20918) );
  INV_X1 U16989 ( .A(n20918), .ZN(n20852) );
  INV_X1 U16990 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n17182) );
  INV_X1 U16991 ( .A(DATAI_22_), .ZN(n13563) );
  INV_X1 U16992 ( .A(n15566), .ZN(n13981) );
  NOR2_X1 U16993 ( .A1(n14128), .A2(n13981), .ZN(n14012) );
  NAND2_X1 U16994 ( .A1(n13596), .A2(n13564), .ZN(n20851) );
  OAI22_X1 U16995 ( .A1(n13598), .A2(n20921), .B1(n20851), .B2(n13597), .ZN(
        n13565) );
  AOI21_X1 U16996 ( .B1(n20801), .B2(n20917), .A(n13565), .ZN(n13567) );
  NAND2_X1 U16997 ( .A1(n13600), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13566) );
  OAI211_X1 U16998 ( .C1(n13603), .C2(n20852), .A(n13567), .B(n13566), .ZN(
        P1_U3079) );
  INV_X1 U16999 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19885) );
  INV_X1 U17000 ( .A(DATAI_27_), .ZN(n13568) );
  OAI22_X1 U17001 ( .A1(n19885), .A2(n13592), .B1(n13568), .B2(n13593), .ZN(
        n20900) );
  INV_X1 U17002 ( .A(n20900), .ZN(n20837) );
  INV_X1 U17003 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n17187) );
  INV_X1 U17004 ( .A(DATAI_19_), .ZN(n13569) );
  NOR2_X1 U17005 ( .A1(n14128), .A2(n13570), .ZN(n14002) );
  NAND2_X1 U17006 ( .A1(n13596), .A2(n13571), .ZN(n20836) );
  OAI22_X1 U17007 ( .A1(n13598), .A2(n20903), .B1(n20836), .B2(n13597), .ZN(
        n13572) );
  AOI21_X1 U17008 ( .B1(n20801), .B2(n20899), .A(n13572), .ZN(n13574) );
  NAND2_X1 U17009 ( .A1(n13600), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n13573) );
  OAI211_X1 U17010 ( .C1(n13603), .C2(n20837), .A(n13574), .B(n13573), .ZN(
        P1_U3076) );
  INV_X1 U17011 ( .A(DATAI_31_), .ZN(n13575) );
  INV_X1 U17012 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19903) );
  OAI22_X1 U17013 ( .A1(n13575), .A2(n13593), .B1(n19903), .B2(n13592), .ZN(
        n20927) );
  INV_X1 U17014 ( .A(n20927), .ZN(n20858) );
  INV_X1 U17015 ( .A(DATAI_23_), .ZN(n13576) );
  INV_X1 U17016 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n17180) );
  INV_X1 U17017 ( .A(n15560), .ZN(n14123) );
  NOR2_X1 U17018 ( .A1(n14128), .A2(n14123), .ZN(n14021) );
  NAND2_X1 U17019 ( .A1(n13596), .A2(n13577), .ZN(n20857) );
  OAI22_X1 U17020 ( .A1(n13598), .A2(n20931), .B1(n20857), .B2(n13597), .ZN(
        n13578) );
  AOI21_X1 U17021 ( .B1(n20801), .B2(n20924), .A(n13578), .ZN(n13580) );
  NAND2_X1 U17022 ( .A1(n13600), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13579) );
  OAI211_X1 U17023 ( .C1(n13603), .C2(n20858), .A(n13580), .B(n13579), .ZN(
        P1_U3080) );
  INV_X1 U17024 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17178) );
  INV_X1 U17025 ( .A(DATAI_24_), .ZN(n13581) );
  OAI22_X1 U17026 ( .A1(n17178), .A2(n13592), .B1(n13581), .B2(n13593), .ZN(
        n20882) );
  INV_X1 U17027 ( .A(n20882), .ZN(n20816) );
  INV_X1 U17028 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n21227) );
  INV_X1 U17029 ( .A(DATAI_16_), .ZN(n21176) );
  NOR2_X1 U17030 ( .A1(n14128), .A2(n15596), .ZN(n14007) );
  NAND2_X1 U17031 ( .A1(n13596), .A2(n13832), .ZN(n20815) );
  OAI22_X1 U17032 ( .A1(n13598), .A2(n20885), .B1(n20815), .B2(n13597), .ZN(
        n13582) );
  AOI21_X1 U17033 ( .B1(n20801), .B2(n20875), .A(n13582), .ZN(n13584) );
  NAND2_X1 U17034 ( .A1(n13600), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13583) );
  OAI211_X1 U17035 ( .C1(n13603), .C2(n20816), .A(n13584), .B(n13583), .ZN(
        P1_U3073) );
  INV_X1 U17036 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n17176) );
  INV_X1 U17037 ( .A(DATAI_25_), .ZN(n21259) );
  OAI22_X1 U17038 ( .A1(n17176), .A2(n13592), .B1(n21259), .B2(n13593), .ZN(
        n20888) );
  INV_X1 U17039 ( .A(n20888), .ZN(n20827) );
  INV_X1 U17040 ( .A(DATAI_17_), .ZN(n13585) );
  INV_X1 U17041 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n17191) );
  NOR2_X1 U17042 ( .A1(n14128), .A2(n13586), .ZN(n13997) );
  NAND2_X1 U17043 ( .A1(n13596), .A2(n13587), .ZN(n20826) );
  OAI22_X1 U17044 ( .A1(n13598), .A2(n20891), .B1(n20826), .B2(n13597), .ZN(
        n13588) );
  AOI21_X1 U17045 ( .B1(n20801), .B2(n20887), .A(n13588), .ZN(n13590) );
  NAND2_X1 U17046 ( .A1(n13600), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13589) );
  OAI211_X1 U17047 ( .C1(n13603), .C2(n20827), .A(n13590), .B(n13589), .ZN(
        P1_U3074) );
  INV_X1 U17048 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n17170) );
  INV_X1 U17049 ( .A(DATAI_29_), .ZN(n13591) );
  OAI22_X1 U17050 ( .A1(n17170), .A2(n13592), .B1(n13591), .B2(n13593), .ZN(
        n20912) );
  INV_X1 U17051 ( .A(n20912), .ZN(n20847) );
  INV_X1 U17052 ( .A(DATAI_21_), .ZN(n13594) );
  INV_X1 U17053 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17184) );
  INV_X1 U17054 ( .A(n15570), .ZN(n13595) );
  NOR2_X1 U17055 ( .A1(n14128), .A2(n13595), .ZN(n14027) );
  NAND2_X1 U17056 ( .A1(n13596), .A2(n15107), .ZN(n20846) );
  OAI22_X1 U17057 ( .A1(n13598), .A2(n20915), .B1(n20846), .B2(n13597), .ZN(
        n13599) );
  AOI21_X1 U17058 ( .B1(n20801), .B2(n20911), .A(n13599), .ZN(n13602) );
  NAND2_X1 U17059 ( .A1(n13600), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13601) );
  OAI211_X1 U17060 ( .C1(n13603), .C2(n20847), .A(n13602), .B(n13601), .ZN(
        P1_U3078) );
  INV_X1 U17061 ( .A(n13972), .ZN(n14105) );
  AOI22_X1 U17062 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n15071), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13607) );
  AOI22_X1 U17063 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13606) );
  AOI22_X1 U17064 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13960), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13605) );
  AOI22_X1 U17065 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13604) );
  NAND4_X1 U17066 ( .A1(n13607), .A2(n13606), .A3(n13605), .A4(n13604), .ZN(
        n13613) );
  INV_X1 U17067 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n21076) );
  AOI22_X1 U17068 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15040), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13611) );
  AOI22_X1 U17069 ( .A1(n14947), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13610) );
  AOI22_X1 U17070 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n15081), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13609) );
  AOI22_X1 U17071 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13608) );
  NAND4_X1 U17072 ( .A1(n13611), .A2(n13610), .A3(n13609), .A4(n13608), .ZN(
        n13612) );
  NOR2_X1 U17073 ( .A1(n13613), .A2(n13612), .ZN(n13815) );
  INV_X1 U17074 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13614) );
  OAI22_X1 U17075 ( .A1(n14105), .A2(n13815), .B1(n14103), .B2(n13614), .ZN(
        n13693) );
  XNOR2_X1 U17076 ( .A(n13695), .B(n13693), .ZN(n13812) );
  NAND2_X1 U17077 ( .A1(n13615), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13621) );
  INV_X1 U17078 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20582) );
  AOI21_X1 U17079 ( .B1(n20582), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13617) );
  AOI21_X1 U17080 ( .B1(n15246), .B2(P1_EAX_REG_4__SCAN_IN), .A(n13617), .ZN(
        n13620) );
  OAI21_X1 U17081 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13618), .A(
        n13688), .ZN(n20584) );
  NOR2_X1 U17082 ( .A1(n20584), .A2(n15101), .ZN(n13619) );
  AOI21_X1 U17083 ( .B1(n13621), .B2(n13620), .A(n13619), .ZN(n13622) );
  INV_X1 U17084 ( .A(n13623), .ZN(n13626) );
  NAND2_X1 U17085 ( .A1(n13626), .A2(n13625), .ZN(n13715) );
  INV_X1 U17086 ( .A(n13715), .ZN(n13627) );
  AOI21_X1 U17087 ( .B1(n13624), .B2(n13266), .A(n13627), .ZN(n13822) );
  INV_X1 U17088 ( .A(n13822), .ZN(n20586) );
  NAND2_X1 U17089 ( .A1(n15147), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13628) );
  OAI211_X1 U17090 ( .C1(n15287), .C2(P1_EBX_REG_4__SCAN_IN), .A(n15149), .B(
        n13628), .ZN(n13629) );
  OAI21_X1 U17091 ( .B1(n15159), .B2(P1_EBX_REG_4__SCAN_IN), .A(n13629), .ZN(
        n13632) );
  INV_X1 U17092 ( .A(n13632), .ZN(n13630) );
  NAND2_X1 U17093 ( .A1(n13633), .A2(n13632), .ZN(n13634) );
  NAND2_X1 U17094 ( .A1(n13758), .A2(n13634), .ZN(n20579) );
  INV_X1 U17095 ( .A(n20579), .ZN(n13857) );
  AOI22_X1 U17096 ( .A1(n21040), .A2(n13857), .B1(n21041), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13635) );
  OAI21_X1 U17097 ( .B1(n20586), .B2(n15513), .A(n13635), .ZN(P1_U2868) );
  INV_X1 U17098 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21197) );
  OAI222_X1 U17099 ( .A1(n20586), .A2(n15614), .B1(n15608), .B2(n13636), .C1(
        n21197), .C2(n15606), .ZN(P1_U2900) );
  INV_X1 U17100 ( .A(n13722), .ZN(n13638) );
  NAND2_X1 U17101 ( .A1(n13638), .A2(n20733), .ZN(n13719) );
  OAI21_X1 U17102 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n13637), .A(n13719), 
        .ZN(n13641) );
  OR2_X1 U17103 ( .A1(n13539), .A2(n13640), .ZN(n14547) );
  NOR2_X1 U17104 ( .A1(n14547), .A2(n15270), .ZN(n13985) );
  NOR3_X1 U17105 ( .A1(n13641), .A2(n13865), .A3(n13985), .ZN(n13642) );
  NOR2_X1 U17106 ( .A1(n13642), .A2(n20807), .ZN(n14553) );
  NAND2_X1 U17107 ( .A1(n14553), .A2(n13643), .ZN(n13645) );
  NAND2_X1 U17108 ( .A1(n20663), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13644) );
  OAI211_X1 U17109 ( .C1(n20600), .C2(n15273), .A(n13645), .B(n13644), .ZN(
        P1_U3475) );
  OAI21_X1 U17110 ( .B1(n20305), .B2(n20366), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13647) );
  NAND2_X1 U17111 ( .A1(n13647), .A2(n20458), .ZN(n13657) );
  INV_X1 U17112 ( .A(n13657), .ZN(n13649) );
  AND3_X1 U17113 ( .A1(n20492), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n20311), .ZN(n20303) );
  NOR2_X1 U17114 ( .A1(n20492), .A2(n20259), .ZN(n20278) );
  NOR2_X1 U17115 ( .A1(n20303), .A2(n20278), .ZN(n13656) );
  INV_X1 U17116 ( .A(n10779), .ZN(n13654) );
  AOI211_X1 U17117 ( .C1(n13654), .C2(n20101), .A(n20303), .B(n20458), .ZN(
        n13648) );
  AOI211_X2 U17118 ( .C1(n13649), .C2(n13656), .A(n20074), .B(n13648), .ZN(
        n20309) );
  INV_X1 U17119 ( .A(n20366), .ZN(n13652) );
  INV_X1 U17120 ( .A(n20303), .ZN(n13650) );
  OAI22_X1 U17121 ( .A1(n13652), .A2(n20325), .B1(n13651), .B2(n13650), .ZN(
        n13653) );
  AOI21_X1 U17122 ( .B1(n20305), .B2(n20322), .A(n13653), .ZN(n13659) );
  OAI21_X1 U17123 ( .B1(n13654), .B2(n20303), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13655) );
  NAND2_X1 U17124 ( .A1(n20306), .A2(n13231), .ZN(n13658) );
  OAI211_X1 U17125 ( .C1(n20309), .C2(n13660), .A(n13659), .B(n13658), .ZN(
        P2_U3160) );
  INV_X1 U17126 ( .A(n13661), .ZN(n13663) );
  OAI211_X1 U17127 ( .C1(n9872), .C2(n13663), .A(n16970), .B(n13662), .ZN(
        n13666) );
  OAI21_X1 U17128 ( .B1(n13505), .B2(n13664), .A(n14172), .ZN(n19618) );
  INV_X1 U17129 ( .A(n19618), .ZN(n17062) );
  NAND2_X1 U17130 ( .A1(n17062), .A2(n19712), .ZN(n13665) );
  OAI211_X1 U17131 ( .C1(n19712), .C2(n11083), .A(n13666), .B(n13665), .ZN(
        P2_U2873) );
  XNOR2_X1 U17132 ( .A(n13667), .B(n13668), .ZN(n17031) );
  OR2_X1 U17133 ( .A1(n13669), .A2(n13670), .ZN(n13673) );
  OAI21_X1 U17134 ( .B1(n13671), .B2(n13669), .A(n13670), .ZN(n13672) );
  OAI21_X1 U17135 ( .B1(n13673), .B2(n13671), .A(n13672), .ZN(n17030) );
  AOI221_X1 U17136 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n21051), .C2(n13675), .A(
        n13674), .ZN(n13677) );
  INV_X1 U17137 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n21260) );
  NOR2_X1 U17138 ( .A1(n21260), .A2(n19856), .ZN(n13676) );
  AOI211_X1 U17139 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n13678), .A(
        n13677), .B(n13676), .ZN(n13685) );
  OAI21_X1 U17140 ( .B1(n13681), .B2(n13680), .A(n13679), .ZN(n19757) );
  INV_X1 U17141 ( .A(n17033), .ZN(n13682) );
  OAI22_X1 U17142 ( .A1(n19757), .A2(n17070), .B1(n19870), .B2(n13682), .ZN(
        n13683) );
  INV_X1 U17143 ( .A(n13683), .ZN(n13684) );
  OAI211_X1 U17144 ( .C1(n17030), .C2(n19859), .A(n13685), .B(n13684), .ZN(
        n13686) );
  INV_X1 U17145 ( .A(n13686), .ZN(n13687) );
  OAI21_X1 U17146 ( .B1(n17031), .B2(n16500), .A(n13687), .ZN(P2_U3041) );
  INV_X1 U17147 ( .A(n15245), .ZN(n14830) );
  INV_X1 U17148 ( .A(n13688), .ZN(n13690) );
  INV_X1 U17149 ( .A(n13974), .ZN(n13689) );
  OAI21_X1 U17150 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13690), .A(
        n13689), .ZN(n20572) );
  NAND2_X1 U17151 ( .A1(n14983), .A2(n20572), .ZN(n13691) );
  OAI21_X1 U17152 ( .B1(n20559), .B2(n14830), .A(n13691), .ZN(n13692) );
  AOI21_X1 U17153 ( .B1(n15246), .B2(P1_EAX_REG_5__SCAN_IN), .A(n13692), .ZN(
        n13710) );
  INV_X1 U17154 ( .A(n13693), .ZN(n13694) );
  AOI22_X1 U17155 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U17156 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9710), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13698) );
  AOI22_X1 U17157 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U17158 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13696) );
  NAND4_X1 U17159 ( .A1(n13699), .A2(n13698), .A3(n13697), .A4(n13696), .ZN(
        n13706) );
  AOI22_X1 U17160 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15082), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13704) );
  AOI22_X1 U17161 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13703) );
  AOI22_X1 U17162 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U17163 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13701) );
  NAND4_X1 U17164 ( .A1(n13704), .A2(n13703), .A3(n13702), .A4(n13701), .ZN(
        n13705) );
  INV_X1 U17165 ( .A(n14408), .ZN(n13708) );
  INV_X1 U17166 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13707) );
  OAI22_X1 U17167 ( .A1(n14105), .A2(n13708), .B1(n14103), .B2(n13707), .ZN(
        n14101) );
  INV_X1 U17168 ( .A(n14101), .ZN(n14399) );
  AND2_X1 U17169 ( .A1(n14399), .A2(n13710), .ZN(n13711) );
  NAND2_X1 U17170 ( .A1(n14400), .A2(n13711), .ZN(n13712) );
  AND2_X1 U17171 ( .A1(n13715), .A2(n13714), .ZN(n13716) );
  NOR2_X2 U17172 ( .A1(n13715), .A2(n13714), .ZN(n13978) );
  OR2_X1 U17173 ( .A1(n13716), .A2(n13978), .ZN(n20568) );
  AOI22_X1 U17174 ( .A1(n15612), .A2(n15570), .B1(P1_EAX_REG_5__SCAN_IN), .B2(
        n15610), .ZN(n13717) );
  OAI21_X1 U17175 ( .B1(n20568), .B2(n15614), .A(n13717), .ZN(P1_U2899) );
  INV_X1 U17176 ( .A(n20924), .ZN(n14137) );
  OR2_X1 U17177 ( .A1(n12911), .A2(n13718), .ZN(n20735) );
  INV_X1 U17178 ( .A(n20735), .ZN(n14549) );
  NAND2_X1 U17179 ( .A1(n20776), .A2(n14549), .ZN(n13723) );
  NAND4_X1 U17180 ( .A1(n13719), .A2(n15926), .A3(n13747), .A4(n13723), .ZN(
        n13720) );
  OAI211_X1 U17181 ( .C1(n15926), .C2(n10340), .A(n13720), .B(n20744), .ZN(
        n13746) );
  NAND2_X1 U17182 ( .A1(n13746), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13727) );
  AOI21_X1 U17183 ( .B1(n13723), .B2(n13747), .A(n20807), .ZN(n13724) );
  AOI21_X1 U17184 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n10340), .A(n13724), 
        .ZN(n13748) );
  OAI22_X1 U17185 ( .A1(n13748), .A2(n20931), .B1(n13747), .B2(n20857), .ZN(
        n13725) );
  AOI21_X1 U17186 ( .B1(n20927), .B2(n20802), .A(n13725), .ZN(n13726) );
  OAI211_X1 U17187 ( .C1(n13752), .C2(n14137), .A(n13727), .B(n13726), .ZN(
        P1_U3096) );
  INV_X1 U17188 ( .A(n20893), .ZN(n14141) );
  NAND2_X1 U17189 ( .A1(n13746), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13730) );
  OAI22_X1 U17190 ( .A1(n13748), .A2(n20897), .B1(n13747), .B2(n20831), .ZN(
        n13728) );
  AOI21_X1 U17191 ( .B1(n20894), .B2(n20802), .A(n13728), .ZN(n13729) );
  OAI211_X1 U17192 ( .C1(n13752), .C2(n14141), .A(n13730), .B(n13729), .ZN(
        P1_U3091) );
  INV_X1 U17193 ( .A(n20917), .ZN(n14157) );
  NAND2_X1 U17194 ( .A1(n13746), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n13733) );
  OAI22_X1 U17195 ( .A1(n13748), .A2(n20921), .B1(n13747), .B2(n20851), .ZN(
        n13731) );
  AOI21_X1 U17196 ( .B1(n20918), .B2(n20802), .A(n13731), .ZN(n13732) );
  OAI211_X1 U17197 ( .C1(n13752), .C2(n14157), .A(n13733), .B(n13732), .ZN(
        P1_U3095) );
  INV_X1 U17198 ( .A(n20875), .ZN(n14149) );
  NAND2_X1 U17199 ( .A1(n13746), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13736) );
  OAI22_X1 U17200 ( .A1(n13748), .A2(n20885), .B1(n13747), .B2(n20815), .ZN(
        n13734) );
  AOI21_X1 U17201 ( .B1(n20882), .B2(n20802), .A(n13734), .ZN(n13735) );
  OAI211_X1 U17202 ( .C1(n13752), .C2(n14149), .A(n13736), .B(n13735), .ZN(
        P1_U3089) );
  INV_X1 U17203 ( .A(n20899), .ZN(n14161) );
  NAND2_X1 U17204 ( .A1(n13746), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13739) );
  OAI22_X1 U17205 ( .A1(n13748), .A2(n20903), .B1(n13747), .B2(n20836), .ZN(
        n13737) );
  AOI21_X1 U17206 ( .B1(n20900), .B2(n20802), .A(n13737), .ZN(n13738) );
  OAI211_X1 U17207 ( .C1(n13752), .C2(n14161), .A(n13739), .B(n13738), .ZN(
        P1_U3092) );
  INV_X1 U17208 ( .A(n20887), .ZN(n14145) );
  NAND2_X1 U17209 ( .A1(n13746), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13742) );
  OAI22_X1 U17210 ( .A1(n13748), .A2(n20891), .B1(n13747), .B2(n20826), .ZN(
        n13740) );
  AOI21_X1 U17211 ( .B1(n20888), .B2(n20802), .A(n13740), .ZN(n13741) );
  OAI211_X1 U17212 ( .C1(n13752), .C2(n14145), .A(n13742), .B(n13741), .ZN(
        P1_U3090) );
  INV_X1 U17213 ( .A(n20905), .ZN(n14169) );
  NAND2_X1 U17214 ( .A1(n13746), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13745) );
  OAI22_X1 U17215 ( .A1(n13748), .A2(n20909), .B1(n13747), .B2(n20841), .ZN(
        n13743) );
  AOI21_X1 U17216 ( .B1(n20906), .B2(n20802), .A(n13743), .ZN(n13744) );
  OAI211_X1 U17217 ( .C1(n13752), .C2(n14169), .A(n13745), .B(n13744), .ZN(
        P1_U3093) );
  INV_X1 U17218 ( .A(n20911), .ZN(n14153) );
  NAND2_X1 U17219 ( .A1(n13746), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13751) );
  OAI22_X1 U17220 ( .A1(n13748), .A2(n20915), .B1(n13747), .B2(n20846), .ZN(
        n13749) );
  AOI21_X1 U17221 ( .B1(n20912), .B2(n20802), .A(n13749), .ZN(n13750) );
  OAI211_X1 U17222 ( .C1(n13752), .C2(n14153), .A(n13751), .B(n13750), .ZN(
        P1_U3094) );
  INV_X1 U17223 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13760) );
  OR2_X1 U17224 ( .A1(n15165), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n13756) );
  NAND2_X1 U17225 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13753) );
  NAND2_X1 U17226 ( .A1(n15149), .A2(n13753), .ZN(n13754) );
  OAI21_X1 U17227 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(n15287), .A(n13754), .ZN(
        n13755) );
  AND2_X1 U17228 ( .A1(n13758), .A2(n13757), .ZN(n13759) );
  OR2_X1 U17229 ( .A1(n13759), .A2(n16854), .ZN(n20560) );
  OAI222_X1 U17230 ( .A1(n20568), .A2(n15513), .B1(n20618), .B2(n13760), .C1(
        n16730), .C2(n20560), .ZN(P1_U2867) );
  INV_X1 U17231 ( .A(n13865), .ZN(n13861) );
  NAND3_X1 U17232 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n16622), .ZN(n20814) );
  OAI21_X1 U17233 ( .B1(n13762), .B2(n13861), .A(n20814), .ZN(n13763) );
  NAND2_X1 U17234 ( .A1(n13763), .A2(n20744), .ZN(n13799) );
  NAND2_X1 U17235 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13774) );
  INV_X1 U17236 ( .A(n13765), .ZN(n20738) );
  NAND2_X1 U17237 ( .A1(n20738), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13802) );
  AND2_X1 U17238 ( .A1(n13908), .A2(n13515), .ZN(n20810) );
  NAND2_X1 U17239 ( .A1(n20810), .A2(n14549), .ZN(n13766) );
  NAND2_X1 U17240 ( .A1(n13766), .A2(n13802), .ZN(n13767) );
  NAND2_X1 U17241 ( .A1(n13767), .A2(n20866), .ZN(n13770) );
  INV_X1 U17242 ( .A(n20814), .ZN(n13768) );
  NAND2_X1 U17243 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13768), .ZN(n13769) );
  NAND2_X1 U17244 ( .A1(n13770), .A2(n13769), .ZN(n13800) );
  NAND2_X1 U17245 ( .A1(n13800), .A2(n14002), .ZN(n13771) );
  OAI21_X1 U17246 ( .B1(n13802), .B2(n20836), .A(n13771), .ZN(n13772) );
  AOI21_X1 U17247 ( .B1(n20926), .B2(n20899), .A(n13772), .ZN(n13773) );
  OAI211_X1 U17248 ( .C1(n13806), .C2(n20837), .A(n13774), .B(n13773), .ZN(
        P1_U3124) );
  NAND2_X1 U17249 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13778) );
  NAND2_X1 U17250 ( .A1(n13800), .A2(n14016), .ZN(n13775) );
  OAI21_X1 U17251 ( .B1(n13802), .B2(n20831), .A(n13775), .ZN(n13776) );
  AOI21_X1 U17252 ( .B1(n20926), .B2(n20893), .A(n13776), .ZN(n13777) );
  OAI211_X1 U17253 ( .C1(n13806), .C2(n20832), .A(n13778), .B(n13777), .ZN(
        P1_U3123) );
  NAND2_X1 U17254 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13782) );
  NAND2_X1 U17255 ( .A1(n13800), .A2(n14007), .ZN(n13779) );
  OAI21_X1 U17256 ( .B1(n13802), .B2(n20815), .A(n13779), .ZN(n13780) );
  AOI21_X1 U17257 ( .B1(n20926), .B2(n20875), .A(n13780), .ZN(n13781) );
  OAI211_X1 U17258 ( .C1(n13806), .C2(n20816), .A(n13782), .B(n13781), .ZN(
        P1_U3121) );
  NAND2_X1 U17259 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13786) );
  NAND2_X1 U17260 ( .A1(n13800), .A2(n14021), .ZN(n13783) );
  OAI21_X1 U17261 ( .B1(n13802), .B2(n20857), .A(n13783), .ZN(n13784) );
  AOI21_X1 U17262 ( .B1(n20926), .B2(n20924), .A(n13784), .ZN(n13785) );
  OAI211_X1 U17263 ( .C1(n13806), .C2(n20858), .A(n13786), .B(n13785), .ZN(
        P1_U3128) );
  NAND2_X1 U17264 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13790) );
  NAND2_X1 U17265 ( .A1(n13800), .A2(n13992), .ZN(n13787) );
  OAI21_X1 U17266 ( .B1(n13802), .B2(n20841), .A(n13787), .ZN(n13788) );
  AOI21_X1 U17267 ( .B1(n20926), .B2(n20905), .A(n13788), .ZN(n13789) );
  OAI211_X1 U17268 ( .C1(n13806), .C2(n20842), .A(n13790), .B(n13789), .ZN(
        P1_U3125) );
  NAND2_X1 U17269 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13794) );
  NAND2_X1 U17270 ( .A1(n13800), .A2(n14027), .ZN(n13791) );
  OAI21_X1 U17271 ( .B1(n13802), .B2(n20846), .A(n13791), .ZN(n13792) );
  AOI21_X1 U17272 ( .B1(n20926), .B2(n20911), .A(n13792), .ZN(n13793) );
  OAI211_X1 U17273 ( .C1(n13806), .C2(n20847), .A(n13794), .B(n13793), .ZN(
        P1_U3126) );
  NAND2_X1 U17274 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13798) );
  NAND2_X1 U17275 ( .A1(n13800), .A2(n14012), .ZN(n13795) );
  OAI21_X1 U17276 ( .B1(n13802), .B2(n20851), .A(n13795), .ZN(n13796) );
  AOI21_X1 U17277 ( .B1(n20926), .B2(n20917), .A(n13796), .ZN(n13797) );
  OAI211_X1 U17278 ( .C1(n13806), .C2(n20852), .A(n13798), .B(n13797), .ZN(
        P1_U3127) );
  NAND2_X1 U17279 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13805) );
  NAND2_X1 U17280 ( .A1(n13800), .A2(n13997), .ZN(n13801) );
  OAI21_X1 U17281 ( .B1(n13802), .B2(n20826), .A(n13801), .ZN(n13803) );
  AOI21_X1 U17282 ( .B1(n20926), .B2(n20887), .A(n13803), .ZN(n13804) );
  OAI211_X1 U17283 ( .C1(n13806), .C2(n20827), .A(n13805), .B(n13804), .ZN(
        P1_U3122) );
  NAND2_X1 U17284 ( .A1(n13808), .A2(n13807), .ZN(n13811) );
  NAND2_X1 U17285 ( .A1(n13809), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13810) );
  NAND2_X2 U17286 ( .A1(n13811), .A2(n13810), .ZN(n14396) );
  INV_X1 U17287 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13853) );
  NAND2_X1 U17288 ( .A1(n13812), .A2(n14530), .ZN(n13819) );
  NAND2_X1 U17289 ( .A1(n13814), .A2(n13813), .ZN(n13816) );
  OR2_X1 U17290 ( .A1(n13816), .A2(n13815), .ZN(n14407) );
  NAND2_X1 U17291 ( .A1(n13816), .A2(n13815), .ZN(n13817) );
  NAND3_X1 U17292 ( .A1(n14407), .A2(n14536), .A3(n13817), .ZN(n13818) );
  NAND2_X1 U17293 ( .A1(n13819), .A2(n13818), .ZN(n14394) );
  XNOR2_X1 U17294 ( .A(n14395), .B(n14394), .ZN(n13860) );
  INV_X1 U17295 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20957) );
  NOR2_X1 U17296 ( .A1(n16808), .A2(n20957), .ZN(n13856) );
  AOI21_X1 U17297 ( .B1(n16759), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13856), .ZN(n13820) );
  OAI21_X1 U17298 ( .B1(n20584), .B2(n16769), .A(n13820), .ZN(n13821) );
  AOI21_X1 U17299 ( .B1(n13822), .B2(n16764), .A(n13821), .ZN(n13823) );
  OAI21_X1 U17300 ( .B1(n13860), .B2(n20516), .A(n13823), .ZN(P1_U2995) );
  NAND2_X1 U17301 ( .A1(n21026), .A2(n12779), .ZN(n13831) );
  NAND2_X1 U17302 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21033), .ZN(n16642) );
  NAND2_X1 U17303 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n9922), .ZN(n13824) );
  OAI22_X1 U17304 ( .A1(n9922), .A2(n16642), .B1(n13824), .B2(n15101), .ZN(
        n13825) );
  INV_X1 U17305 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14645) );
  INV_X1 U17306 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16704) );
  INV_X1 U17307 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14854) );
  INV_X1 U17308 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15667) );
  INV_X1 U17309 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15344) );
  INV_X1 U17310 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15652) );
  INV_X1 U17311 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15633) );
  INV_X1 U17312 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15187) );
  NOR2_X1 U17313 ( .A1(n15252), .A2(n21133), .ZN(n13830) );
  NAND2_X1 U17314 ( .A1(n21026), .A2(n13832), .ZN(n13846) );
  OR2_X1 U17315 ( .A1(n13833), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13845) );
  NAND2_X1 U17316 ( .A1(n15162), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13836) );
  NAND2_X1 U17317 ( .A1(n13845), .A2(n13836), .ZN(n13834) );
  INV_X1 U17318 ( .A(n15180), .ZN(n20565) );
  AOI22_X1 U17319 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n20602), .B1(n20565), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13851) );
  AND2_X1 U17320 ( .A1(n21028), .A2(n20514), .ZN(n13835) );
  NOR2_X1 U17321 ( .A1(n13836), .A2(n13835), .ZN(n13837) );
  INV_X1 U17322 ( .A(n13838), .ZN(n13839) );
  NAND2_X1 U17323 ( .A1(n21026), .A2(n13839), .ZN(n20599) );
  AND2_X1 U17324 ( .A1(n15252), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13841) );
  NAND2_X1 U17325 ( .A1(n20604), .A2(n13842), .ZN(n13844) );
  NAND2_X1 U17326 ( .A1(n20593), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13843) );
  OAI211_X1 U17327 ( .C1(n20599), .C2(n13840), .A(n13844), .B(n13843), .ZN(
        n13848) );
  NOR2_X1 U17328 ( .A1(n20578), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13847) );
  AOI211_X1 U17329 ( .C1(n20595), .C2(n13849), .A(n13848), .B(n13847), .ZN(
        n13850) );
  OAI211_X1 U17330 ( .C1(n20585), .C2(n20613), .A(n13851), .B(n13850), .ZN(
        P1_U2839) );
  NAND2_X1 U17331 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14422) );
  INV_X1 U17332 ( .A(n14422), .ZN(n14424) );
  AOI21_X1 U17333 ( .B1(n13853), .B2(n13852), .A(n14424), .ZN(n13854) );
  AOI22_X1 U17334 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13855), .B1(
        n16872), .B2(n13854), .ZN(n13859) );
  AOI21_X1 U17335 ( .B1(n16857), .B2(n13857), .A(n13856), .ZN(n13858) );
  OAI211_X1 U17336 ( .C1(n13860), .C2(n20653), .A(n13859), .B(n13858), .ZN(
        P1_U3027) );
  NOR3_X1 U17337 ( .A1(n20737), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13868) );
  INV_X1 U17338 ( .A(n13868), .ZN(n14125) );
  NOR2_X1 U17339 ( .A1(n20779), .A2(n14125), .ZN(n13899) );
  AOI21_X1 U17340 ( .B1(n20810), .B2(n13910), .A(n13899), .ZN(n13866) );
  OAI211_X1 U17341 ( .C1(n13861), .C2(n15270), .A(n15926), .B(n13866), .ZN(
        n13862) );
  OAI211_X1 U17342 ( .C1(n15926), .C2(n13868), .A(n13862), .B(n20744), .ZN(
        n13863) );
  INV_X1 U17343 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13874) );
  INV_X1 U17344 ( .A(n13989), .ZN(n13864) );
  INV_X1 U17345 ( .A(n13866), .ZN(n13867) );
  NAND2_X1 U17346 ( .A1(n13867), .A2(n20866), .ZN(n13870) );
  NAND2_X1 U17347 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13868), .ZN(n13869) );
  NAND2_X1 U17348 ( .A1(n13870), .A2(n13869), .ZN(n13900) );
  INV_X1 U17349 ( .A(n20857), .ZN(n20923) );
  AOI22_X1 U17350 ( .A1(n13900), .A2(n14021), .B1(n20923), .B2(n13899), .ZN(
        n13871) );
  OAI21_X1 U17351 ( .B1(n20859), .B2(n14137), .A(n13871), .ZN(n13872) );
  AOI21_X1 U17352 ( .B1(n20927), .B2(n14126), .A(n13872), .ZN(n13873) );
  OAI21_X1 U17353 ( .B1(n13905), .B2(n13874), .A(n13873), .ZN(P1_U3112) );
  INV_X1 U17354 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13878) );
  INV_X1 U17355 ( .A(n20815), .ZN(n20874) );
  AOI22_X1 U17356 ( .A1(n13900), .A2(n14007), .B1(n20874), .B2(n13899), .ZN(
        n13875) );
  OAI21_X1 U17357 ( .B1(n20859), .B2(n14149), .A(n13875), .ZN(n13876) );
  AOI21_X1 U17358 ( .B1(n20882), .B2(n14126), .A(n13876), .ZN(n13877) );
  OAI21_X1 U17359 ( .B1(n13905), .B2(n13878), .A(n13877), .ZN(P1_U3105) );
  INV_X1 U17360 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13882) );
  INV_X1 U17361 ( .A(n20826), .ZN(n20886) );
  AOI22_X1 U17362 ( .A1(n13900), .A2(n13997), .B1(n20886), .B2(n13899), .ZN(
        n13879) );
  OAI21_X1 U17363 ( .B1(n20859), .B2(n14145), .A(n13879), .ZN(n13880) );
  AOI21_X1 U17364 ( .B1(n20888), .B2(n14126), .A(n13880), .ZN(n13881) );
  OAI21_X1 U17365 ( .B1(n13905), .B2(n13882), .A(n13881), .ZN(P1_U3106) );
  INV_X1 U17366 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13886) );
  INV_X1 U17367 ( .A(n20836), .ZN(n20898) );
  AOI22_X1 U17368 ( .A1(n13900), .A2(n14002), .B1(n20898), .B2(n13899), .ZN(
        n13883) );
  OAI21_X1 U17369 ( .B1(n20859), .B2(n14161), .A(n13883), .ZN(n13884) );
  AOI21_X1 U17370 ( .B1(n20900), .B2(n14126), .A(n13884), .ZN(n13885) );
  OAI21_X1 U17371 ( .B1(n13905), .B2(n13886), .A(n13885), .ZN(P1_U3108) );
  INV_X1 U17372 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13890) );
  INV_X1 U17373 ( .A(n20831), .ZN(n20892) );
  AOI22_X1 U17374 ( .A1(n13900), .A2(n14016), .B1(n20892), .B2(n13899), .ZN(
        n13887) );
  OAI21_X1 U17375 ( .B1(n20859), .B2(n14141), .A(n13887), .ZN(n13888) );
  AOI21_X1 U17376 ( .B1(n20894), .B2(n14126), .A(n13888), .ZN(n13889) );
  OAI21_X1 U17377 ( .B1(n13905), .B2(n13890), .A(n13889), .ZN(P1_U3107) );
  INV_X1 U17378 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13894) );
  INV_X1 U17379 ( .A(n20846), .ZN(n20910) );
  AOI22_X1 U17380 ( .A1(n13900), .A2(n14027), .B1(n20910), .B2(n13899), .ZN(
        n13891) );
  OAI21_X1 U17381 ( .B1(n20859), .B2(n14153), .A(n13891), .ZN(n13892) );
  AOI21_X1 U17382 ( .B1(n20912), .B2(n14126), .A(n13892), .ZN(n13893) );
  OAI21_X1 U17383 ( .B1(n13905), .B2(n13894), .A(n13893), .ZN(P1_U3110) );
  INV_X1 U17384 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13898) );
  INV_X1 U17385 ( .A(n20841), .ZN(n20904) );
  AOI22_X1 U17386 ( .A1(n13900), .A2(n13992), .B1(n20904), .B2(n13899), .ZN(
        n13895) );
  OAI21_X1 U17387 ( .B1(n20859), .B2(n14169), .A(n13895), .ZN(n13896) );
  AOI21_X1 U17388 ( .B1(n20906), .B2(n14126), .A(n13896), .ZN(n13897) );
  OAI21_X1 U17389 ( .B1(n13905), .B2(n13898), .A(n13897), .ZN(P1_U3109) );
  INV_X1 U17390 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13904) );
  INV_X1 U17391 ( .A(n20851), .ZN(n20916) );
  AOI22_X1 U17392 ( .A1(n13900), .A2(n14012), .B1(n20916), .B2(n13899), .ZN(
        n13901) );
  OAI21_X1 U17393 ( .B1(n20859), .B2(n14157), .A(n13901), .ZN(n13902) );
  AOI21_X1 U17394 ( .B1(n20918), .B2(n14126), .A(n13902), .ZN(n13903) );
  OAI21_X1 U17395 ( .B1(n13905), .B2(n13904), .A(n13903), .ZN(P1_U3111) );
  INV_X1 U17396 ( .A(n20695), .ZN(n20734) );
  NOR3_X1 U17397 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20667) );
  INV_X1 U17398 ( .A(n13515), .ZN(n13907) );
  OR2_X1 U17399 ( .A1(n13908), .A2(n13907), .ZN(n20736) );
  INV_X1 U17400 ( .A(n20736), .ZN(n13911) );
  INV_X1 U17401 ( .A(n20667), .ZN(n13909) );
  NOR2_X1 U17402 ( .A1(n20779), .A2(n13909), .ZN(n13915) );
  AOI21_X1 U17403 ( .B1(n13911), .B2(n13910), .A(n13915), .ZN(n13913) );
  OAI211_X1 U17404 ( .C1(n20695), .C2(n15270), .A(n15926), .B(n13913), .ZN(
        n13912) );
  OAI211_X1 U17405 ( .C1(n15926), .C2(n20667), .A(n13912), .B(n20744), .ZN(
        n13937) );
  NAND2_X1 U17406 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13918) );
  INV_X1 U17407 ( .A(n13913), .ZN(n13914) );
  AOI22_X1 U17408 ( .A1(n13914), .A2(n20866), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20667), .ZN(n13939) );
  INV_X1 U17409 ( .A(n13915), .ZN(n13938) );
  OAI22_X1 U17410 ( .A1(n13939), .A2(n20931), .B1(n20857), .B2(n13938), .ZN(
        n13916) );
  AOI21_X1 U17411 ( .B1(n20689), .B2(n20927), .A(n13916), .ZN(n13917) );
  OAI211_X1 U17412 ( .C1(n20727), .C2(n14137), .A(n13918), .B(n13917), .ZN(
        P1_U3048) );
  NAND2_X1 U17413 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13921) );
  OAI22_X1 U17414 ( .A1(n13939), .A2(n20915), .B1(n20846), .B2(n13938), .ZN(
        n13919) );
  AOI21_X1 U17415 ( .B1(n20689), .B2(n20912), .A(n13919), .ZN(n13920) );
  OAI211_X1 U17416 ( .C1(n20727), .C2(n14153), .A(n13921), .B(n13920), .ZN(
        P1_U3046) );
  NAND2_X1 U17417 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n13924) );
  OAI22_X1 U17418 ( .A1(n13939), .A2(n20921), .B1(n20851), .B2(n13938), .ZN(
        n13922) );
  AOI21_X1 U17419 ( .B1(n20689), .B2(n20918), .A(n13922), .ZN(n13923) );
  OAI211_X1 U17420 ( .C1(n20727), .C2(n14157), .A(n13924), .B(n13923), .ZN(
        P1_U3047) );
  NAND2_X1 U17421 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13927) );
  OAI22_X1 U17422 ( .A1(n13939), .A2(n20909), .B1(n20841), .B2(n13938), .ZN(
        n13925) );
  AOI21_X1 U17423 ( .B1(n20689), .B2(n20906), .A(n13925), .ZN(n13926) );
  OAI211_X1 U17424 ( .C1(n20727), .C2(n14169), .A(n13927), .B(n13926), .ZN(
        P1_U3045) );
  NAND2_X1 U17425 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13930) );
  OAI22_X1 U17426 ( .A1(n13939), .A2(n20903), .B1(n20836), .B2(n13938), .ZN(
        n13928) );
  AOI21_X1 U17427 ( .B1(n20689), .B2(n20900), .A(n13928), .ZN(n13929) );
  OAI211_X1 U17428 ( .C1(n20727), .C2(n14161), .A(n13930), .B(n13929), .ZN(
        P1_U3044) );
  NAND2_X1 U17429 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13933) );
  OAI22_X1 U17430 ( .A1(n13939), .A2(n20897), .B1(n20831), .B2(n13938), .ZN(
        n13931) );
  AOI21_X1 U17431 ( .B1(n20689), .B2(n20894), .A(n13931), .ZN(n13932) );
  OAI211_X1 U17432 ( .C1(n20727), .C2(n14141), .A(n13933), .B(n13932), .ZN(
        P1_U3043) );
  NAND2_X1 U17433 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13936) );
  OAI22_X1 U17434 ( .A1(n13939), .A2(n20891), .B1(n20826), .B2(n13938), .ZN(
        n13934) );
  AOI21_X1 U17435 ( .B1(n20689), .B2(n20888), .A(n13934), .ZN(n13935) );
  OAI211_X1 U17436 ( .C1(n20727), .C2(n14145), .A(n13936), .B(n13935), .ZN(
        P1_U3042) );
  NAND2_X1 U17437 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13942) );
  OAI22_X1 U17438 ( .A1(n13939), .A2(n20885), .B1(n20815), .B2(n13938), .ZN(
        n13940) );
  AOI21_X1 U17439 ( .B1(n20689), .B2(n20882), .A(n13940), .ZN(n13941) );
  OAI211_X1 U17440 ( .C1(n20727), .C2(n14149), .A(n13942), .B(n13941), .ZN(
        P1_U3041) );
  INV_X1 U17441 ( .A(n20585), .ZN(n20606) );
  NOR2_X1 U17442 ( .A1(n13515), .A2(n20599), .ZN(n13955) );
  INV_X1 U17443 ( .A(n13943), .ZN(n13952) );
  INV_X1 U17444 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13950) );
  AOI21_X1 U17445 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_2__SCAN_IN), 
        .A(n20578), .ZN(n13944) );
  NOR2_X1 U17446 ( .A1(n20565), .A2(n13944), .ZN(n20610) );
  NAND2_X1 U17447 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n13944), .ZN(n13949) );
  INV_X1 U17448 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13946) );
  OAI22_X1 U17449 ( .A1(n13946), .A2(n20581), .B1(n20580), .B2(n13945), .ZN(
        n13947) );
  INV_X1 U17450 ( .A(n13947), .ZN(n13948) );
  OAI211_X1 U17451 ( .C1(n13950), .C2(n20610), .A(n13949), .B(n13948), .ZN(
        n13951) );
  AOI21_X1 U17452 ( .B1(n20604), .B2(n13952), .A(n13951), .ZN(n13953) );
  OAI21_X1 U17453 ( .B1(n20592), .B2(n13472), .A(n13953), .ZN(n13954) );
  AOI211_X1 U17454 ( .C1(n13956), .C2(n20606), .A(n13955), .B(n13954), .ZN(
        n13957) );
  INV_X1 U17455 ( .A(n13957), .ZN(P1_U2838) );
  INV_X1 U17456 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13977) );
  AOI22_X1 U17457 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13964) );
  AOI22_X1 U17458 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13963) );
  AOI22_X1 U17459 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9710), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13962) );
  AOI22_X1 U17460 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13961) );
  NAND4_X1 U17461 ( .A1(n13964), .A2(n13963), .A3(n13962), .A4(n13961), .ZN(
        n13970) );
  AOI22_X1 U17462 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15082), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13968) );
  INV_X1 U17463 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n21081) );
  AOI22_X1 U17464 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13967) );
  AOI22_X1 U17465 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13966) );
  AOI22_X1 U17466 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13965) );
  NAND4_X1 U17467 ( .A1(n13968), .A2(n13967), .A3(n13966), .A4(n13965), .ZN(
        n13969) );
  AOI22_X1 U17468 ( .A1(n13972), .A2(n14416), .B1(n13971), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14099) );
  NAND2_X1 U17469 ( .A1(n13959), .A2(n14099), .ZN(n14406) );
  NAND2_X1 U17470 ( .A1(n14406), .A2(n14780), .ZN(n13976) );
  OAI21_X1 U17471 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13974), .A(
        n13973), .ZN(n20551) );
  AOI22_X1 U17472 ( .A1(n14983), .A2(n20551), .B1(n15245), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13975) );
  NAND2_X1 U17473 ( .A1(n13978), .A2(n13979), .ZN(n14098) );
  OR2_X1 U17474 ( .A1(n13978), .A2(n13979), .ZN(n13980) );
  AND2_X1 U17475 ( .A1(n14098), .A2(n13980), .ZN(n20611) );
  INV_X1 U17476 ( .A(n20611), .ZN(n13982) );
  OAI222_X1 U17477 ( .A1(n13982), .A2(n15614), .B1(n15608), .B2(n13981), .C1(
        n15606), .C2(n13977), .ZN(P1_U2898) );
  OR3_X1 U17478 ( .A1(n16622), .A2(n20737), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20873) );
  INV_X1 U17479 ( .A(n20744), .ZN(n13987) );
  NOR2_X1 U17480 ( .A1(n20869), .A2(n13984), .ZN(n13990) );
  NOR2_X1 U17481 ( .A1(n20779), .A2(n20873), .ZN(n14026) );
  NOR4_X1 U17482 ( .A1(n13985), .A2(n13990), .A3(n14026), .A4(n20807), .ZN(
        n13986) );
  AOI211_X2 U17483 ( .C1(n20807), .C2(n20873), .A(n13987), .B(n13986), .ZN(
        n14034) );
  INV_X1 U17484 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13996) );
  NOR2_X2 U17485 ( .A1(n14547), .A2(n13988), .ZN(n14078) );
  INV_X1 U17486 ( .A(n20925), .ZN(n14030) );
  OAI21_X1 U17487 ( .B1(n13990), .B2(n14026), .A(n15926), .ZN(n13991) );
  OAI21_X1 U17488 ( .B1(n20873), .B2(n14046), .A(n13991), .ZN(n14028) );
  AOI22_X1 U17489 ( .A1(n14028), .A2(n13992), .B1(n20904), .B2(n14026), .ZN(
        n13993) );
  OAI21_X1 U17490 ( .B1(n14030), .B2(n20842), .A(n13993), .ZN(n13994) );
  AOI21_X1 U17491 ( .B1(n20905), .B2(n14078), .A(n13994), .ZN(n13995) );
  OAI21_X1 U17492 ( .B1(n14034), .B2(n13996), .A(n13995), .ZN(P1_U3141) );
  INV_X1 U17493 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14001) );
  AOI22_X1 U17494 ( .A1(n14028), .A2(n13997), .B1(n20886), .B2(n14026), .ZN(
        n13998) );
  OAI21_X1 U17495 ( .B1(n14030), .B2(n20827), .A(n13998), .ZN(n13999) );
  AOI21_X1 U17496 ( .B1(n20887), .B2(n14078), .A(n13999), .ZN(n14000) );
  OAI21_X1 U17497 ( .B1(n14034), .B2(n14001), .A(n14000), .ZN(P1_U3138) );
  INV_X1 U17498 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U17499 ( .A1(n14028), .A2(n14002), .B1(n20898), .B2(n14026), .ZN(
        n14003) );
  OAI21_X1 U17500 ( .B1(n14030), .B2(n20837), .A(n14003), .ZN(n14004) );
  AOI21_X1 U17501 ( .B1(n20899), .B2(n14078), .A(n14004), .ZN(n14005) );
  OAI21_X1 U17502 ( .B1(n14034), .B2(n14006), .A(n14005), .ZN(P1_U3140) );
  INV_X1 U17503 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14011) );
  AOI22_X1 U17504 ( .A1(n14028), .A2(n14007), .B1(n20874), .B2(n14026), .ZN(
        n14008) );
  OAI21_X1 U17505 ( .B1(n14030), .B2(n20816), .A(n14008), .ZN(n14009) );
  AOI21_X1 U17506 ( .B1(n20875), .B2(n14078), .A(n14009), .ZN(n14010) );
  OAI21_X1 U17507 ( .B1(n14034), .B2(n14011), .A(n14010), .ZN(P1_U3137) );
  AOI22_X1 U17508 ( .A1(n14028), .A2(n14012), .B1(n20916), .B2(n14026), .ZN(
        n14013) );
  OAI21_X1 U17509 ( .B1(n14030), .B2(n20852), .A(n14013), .ZN(n14014) );
  AOI21_X1 U17510 ( .B1(n20917), .B2(n14078), .A(n14014), .ZN(n14015) );
  OAI21_X1 U17511 ( .B1(n14034), .B2(n21081), .A(n14015), .ZN(P1_U3143) );
  INV_X1 U17512 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14020) );
  AOI22_X1 U17513 ( .A1(n14028), .A2(n14016), .B1(n20892), .B2(n14026), .ZN(
        n14017) );
  OAI21_X1 U17514 ( .B1(n14030), .B2(n20832), .A(n14017), .ZN(n14018) );
  AOI21_X1 U17515 ( .B1(n20893), .B2(n14078), .A(n14018), .ZN(n14019) );
  OAI21_X1 U17516 ( .B1(n14034), .B2(n14020), .A(n14019), .ZN(P1_U3139) );
  INV_X1 U17517 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14025) );
  AOI22_X1 U17518 ( .A1(n14028), .A2(n14021), .B1(n20923), .B2(n14026), .ZN(
        n14022) );
  OAI21_X1 U17519 ( .B1(n14030), .B2(n20858), .A(n14022), .ZN(n14023) );
  AOI21_X1 U17520 ( .B1(n20924), .B2(n14078), .A(n14023), .ZN(n14024) );
  OAI21_X1 U17521 ( .B1(n14034), .B2(n14025), .A(n14024), .ZN(P1_U3144) );
  INV_X1 U17522 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14033) );
  AOI22_X1 U17523 ( .A1(n14028), .A2(n14027), .B1(n20910), .B2(n14026), .ZN(
        n14029) );
  OAI21_X1 U17524 ( .B1(n14030), .B2(n20847), .A(n14029), .ZN(n14031) );
  AOI21_X1 U17525 ( .B1(n20911), .B2(n14078), .A(n14031), .ZN(n14032) );
  OAI21_X1 U17526 ( .B1(n14034), .B2(n14033), .A(n14032), .ZN(P1_U3142) );
  XNOR2_X1 U17527 ( .A(n14035), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14097) );
  XOR2_X1 U17528 ( .A(n14037), .B(n14036), .Z(n14095) );
  INV_X1 U17529 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20403) );
  OAI22_X1 U17530 ( .A1(n20403), .A2(n19856), .B1(n19840), .B2(n14279), .ZN(
        n14039) );
  NOR2_X1 U17531 ( .A1(n17046), .A2(n10155), .ZN(n14038) );
  NOR2_X1 U17532 ( .A1(n14039), .A2(n14038), .ZN(n14040) );
  OAI21_X1 U17533 ( .B1(n14282), .B2(n16307), .A(n14040), .ZN(n14041) );
  AOI21_X1 U17534 ( .B1(n14095), .B2(n19828), .A(n14041), .ZN(n14042) );
  OAI21_X1 U17535 ( .B1(n14097), .B2(n17039), .A(n14042), .ZN(P2_U3008) );
  OAI21_X1 U17536 ( .B1(n14078), .B2(n14043), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14044) );
  INV_X1 U17537 ( .A(n20869), .ZN(n14550) );
  INV_X1 U17538 ( .A(n13840), .ZN(n20868) );
  NAND2_X1 U17539 ( .A1(n14550), .A2(n20868), .ZN(n14048) );
  AOI21_X1 U17540 ( .B1(n14044), .B2(n14048), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n14047) );
  INV_X1 U17541 ( .A(n14556), .ZN(n14045) );
  NOR2_X1 U17542 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14045), .ZN(
        n14052) );
  OAI21_X1 U17543 ( .B1(n20737), .B2(n20701), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20818) );
  NOR2_X1 U17544 ( .A1(n14049), .A2(n14046), .ZN(n20811) );
  NOR2_X1 U17545 ( .A1(n20811), .A2(n14128), .ZN(n20876) );
  NAND2_X1 U17546 ( .A1(n14074), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n14055) );
  INV_X1 U17547 ( .A(n14048), .ZN(n14051) );
  INV_X1 U17548 ( .A(n14049), .ZN(n14050) );
  NOR2_X1 U17549 ( .A1(n14050), .A2(n14046), .ZN(n20871) );
  NOR2_X1 U17550 ( .A1(n20701), .A2(n20737), .ZN(n20812) );
  AOI22_X1 U17551 ( .A1(n14051), .A2(n20866), .B1(n20871), .B2(n20812), .ZN(
        n14076) );
  INV_X1 U17552 ( .A(n14052), .ZN(n14075) );
  OAI22_X1 U17553 ( .A1(n20915), .A2(n14076), .B1(n20846), .B2(n14075), .ZN(
        n14053) );
  AOI21_X1 U17554 ( .B1(n14078), .B2(n20912), .A(n14053), .ZN(n14054) );
  OAI211_X1 U17555 ( .C1(n14584), .C2(n14153), .A(n14055), .B(n14054), .ZN(
        P1_U3150) );
  NAND2_X1 U17556 ( .A1(n14074), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14058) );
  OAI22_X1 U17557 ( .A1(n20909), .A2(n14076), .B1(n20841), .B2(n14075), .ZN(
        n14056) );
  AOI21_X1 U17558 ( .B1(n14078), .B2(n20906), .A(n14056), .ZN(n14057) );
  OAI211_X1 U17559 ( .C1(n14584), .C2(n14169), .A(n14058), .B(n14057), .ZN(
        P1_U3149) );
  NAND2_X1 U17560 ( .A1(n14074), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14061) );
  OAI22_X1 U17561 ( .A1(n14076), .A2(n20897), .B1(n20831), .B2(n14075), .ZN(
        n14059) );
  AOI21_X1 U17562 ( .B1(n14078), .B2(n20894), .A(n14059), .ZN(n14060) );
  OAI211_X1 U17563 ( .C1(n14584), .C2(n14141), .A(n14061), .B(n14060), .ZN(
        P1_U3147) );
  NAND2_X1 U17564 ( .A1(n14074), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14064) );
  OAI22_X1 U17565 ( .A1(n14076), .A2(n20885), .B1(n20815), .B2(n14075), .ZN(
        n14062) );
  AOI21_X1 U17566 ( .B1(n14078), .B2(n20882), .A(n14062), .ZN(n14063) );
  OAI211_X1 U17567 ( .C1(n14584), .C2(n14149), .A(n14064), .B(n14063), .ZN(
        P1_U3145) );
  NAND2_X1 U17568 ( .A1(n14074), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n14067) );
  OAI22_X1 U17569 ( .A1(n14076), .A2(n20903), .B1(n20836), .B2(n14075), .ZN(
        n14065) );
  AOI21_X1 U17570 ( .B1(n14078), .B2(n20900), .A(n14065), .ZN(n14066) );
  OAI211_X1 U17571 ( .C1(n14584), .C2(n14161), .A(n14067), .B(n14066), .ZN(
        P1_U3148) );
  NAND2_X1 U17572 ( .A1(n14074), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14070) );
  OAI22_X1 U17573 ( .A1(n20921), .A2(n14076), .B1(n20851), .B2(n14075), .ZN(
        n14068) );
  AOI21_X1 U17574 ( .B1(n14078), .B2(n20918), .A(n14068), .ZN(n14069) );
  OAI211_X1 U17575 ( .C1(n14584), .C2(n14157), .A(n14070), .B(n14069), .ZN(
        P1_U3151) );
  NAND2_X1 U17576 ( .A1(n14074), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n14073) );
  OAI22_X1 U17577 ( .A1(n14076), .A2(n20891), .B1(n20826), .B2(n14075), .ZN(
        n14071) );
  AOI21_X1 U17578 ( .B1(n14078), .B2(n20888), .A(n14071), .ZN(n14072) );
  OAI211_X1 U17579 ( .C1(n14584), .C2(n14145), .A(n14073), .B(n14072), .ZN(
        P1_U3146) );
  NAND2_X1 U17580 ( .A1(n14074), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n14080) );
  OAI22_X1 U17581 ( .A1(n20931), .A2(n14076), .B1(n20857), .B2(n14075), .ZN(
        n14077) );
  AOI21_X1 U17582 ( .B1(n14078), .B2(n20927), .A(n14077), .ZN(n14079) );
  OAI211_X1 U17583 ( .C1(n14584), .C2(n14137), .A(n14080), .B(n14079), .ZN(
        P1_U3152) );
  OAI21_X1 U17584 ( .B1(n14081), .B2(n14082), .A(n9715), .ZN(n14185) );
  NAND2_X1 U17585 ( .A1(n19716), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n14085) );
  AOI21_X1 U17586 ( .B1(n14083), .B2(n14174), .A(n11090), .ZN(n19605) );
  NAND2_X1 U17587 ( .A1(n19605), .A2(n19712), .ZN(n14084) );
  OAI211_X1 U17588 ( .C1(n14185), .C2(n19713), .A(n14085), .B(n14084), .ZN(
        P2_U2871) );
  OAI21_X1 U17589 ( .B1(n16432), .B2(n14087), .A(n14086), .ZN(n14301) );
  NOR3_X1 U17590 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14088), .A3(
        n14443), .ZN(n14302) );
  NOR2_X1 U17591 ( .A1(n20403), .A2(n19856), .ZN(n14089) );
  AOI211_X1 U17592 ( .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n14301), .A(
        n14302), .B(n14089), .ZN(n14090) );
  INV_X1 U17593 ( .A(n14090), .ZN(n14094) );
  XNOR2_X1 U17594 ( .A(n14092), .B(n14091), .ZN(n19745) );
  OAI22_X1 U17595 ( .A1(n19745), .A2(n17070), .B1(n19870), .B2(n14282), .ZN(
        n14093) );
  AOI211_X1 U17596 ( .C1(n14095), .C2(n19866), .A(n14094), .B(n14093), .ZN(
        n14096) );
  OAI21_X1 U17597 ( .B1(n14097), .B2(n19859), .A(n14096), .ZN(P2_U3040) );
  INV_X1 U17598 ( .A(n14099), .ZN(n14100) );
  INV_X1 U17599 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14102) );
  OAI22_X1 U17600 ( .A1(n14105), .A2(n14104), .B1(n14103), .B2(n14102), .ZN(
        n14106) );
  INV_X1 U17601 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n14122) );
  OAI21_X1 U17602 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n14107), .A(
        n14223), .ZN(n20545) );
  AOI22_X1 U17603 ( .A1(n14983), .A2(n20545), .B1(n15245), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14108) );
  OAI21_X1 U17604 ( .B1(n13616), .B2(n14122), .A(n14108), .ZN(n14109) );
  NAND2_X1 U17605 ( .A1(n14098), .A2(n14110), .ZN(n14111) );
  AND2_X1 U17606 ( .A1(n14222), .A2(n14111), .ZN(n20547) );
  INV_X1 U17607 ( .A(n20547), .ZN(n14124) );
  INV_X1 U17608 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14121) );
  INV_X1 U17609 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21295) );
  NAND2_X1 U17610 ( .A1(n15146), .A2(n21295), .ZN(n14114) );
  NAND2_X1 U17611 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14112) );
  OAI211_X1 U17612 ( .C1(n15287), .C2(P1_EBX_REG_6__SCAN_IN), .A(n15149), .B(
        n14112), .ZN(n14113) );
  OR2_X1 U17613 ( .A1(n15165), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n14118) );
  NAND2_X1 U17614 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14115) );
  NAND2_X1 U17615 ( .A1(n15149), .A2(n14115), .ZN(n14116) );
  OAI21_X1 U17616 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n15287), .A(n14116), .ZN(
        n14117) );
  NAND2_X1 U17617 ( .A1(n14118), .A2(n14117), .ZN(n14119) );
  OR2_X1 U17618 ( .A1(n16856), .A2(n14119), .ZN(n14120) );
  NAND2_X1 U17619 ( .A1(n14241), .A2(n14120), .ZN(n20550) );
  OAI222_X1 U17620 ( .A1(n14124), .A2(n15513), .B1(n20618), .B2(n14121), .C1(
        n16730), .C2(n20550), .ZN(P1_U2865) );
  OAI222_X1 U17621 ( .A1(n14124), .A2(n15614), .B1(n15608), .B2(n14123), .C1(
        n14122), .C2(n15606), .ZN(P1_U2897) );
  NOR2_X1 U17622 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14125), .ZN(
        n14133) );
  OAI21_X1 U17623 ( .B1(n14126), .B2(n14166), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14127) );
  AOI21_X1 U17624 ( .B1(n20810), .B2(n13840), .A(n14133), .ZN(n14130) );
  NAND2_X1 U17625 ( .A1(n14127), .A2(n14130), .ZN(n14129) );
  NOR2_X1 U17626 ( .A1(n20871), .A2(n14128), .ZN(n20700) );
  NAND2_X1 U17627 ( .A1(n14162), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n14136) );
  INV_X1 U17628 ( .A(n14130), .ZN(n14132) );
  INV_X1 U17629 ( .A(n14190), .ZN(n14131) );
  NAND2_X1 U17630 ( .A1(n14131), .A2(n20701), .ZN(n20878) );
  INV_X1 U17631 ( .A(n20878), .ZN(n20870) );
  AOI22_X1 U17632 ( .A1(n14132), .A2(n20866), .B1(n20870), .B2(n20811), .ZN(
        n14164) );
  INV_X1 U17633 ( .A(n14133), .ZN(n14163) );
  OAI22_X1 U17634 ( .A1(n14164), .A2(n20931), .B1(n20857), .B2(n14163), .ZN(
        n14134) );
  AOI21_X1 U17635 ( .B1(n14166), .B2(n20927), .A(n14134), .ZN(n14135) );
  OAI211_X1 U17636 ( .C1(n14170), .C2(n14137), .A(n14136), .B(n14135), .ZN(
        P1_U3104) );
  NAND2_X1 U17637 ( .A1(n14162), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14140) );
  OAI22_X1 U17638 ( .A1(n14164), .A2(n20897), .B1(n20831), .B2(n14163), .ZN(
        n14138) );
  AOI21_X1 U17639 ( .B1(n14166), .B2(n20894), .A(n14138), .ZN(n14139) );
  OAI211_X1 U17640 ( .C1(n14170), .C2(n14141), .A(n14140), .B(n14139), .ZN(
        P1_U3099) );
  NAND2_X1 U17641 ( .A1(n14162), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14144) );
  OAI22_X1 U17642 ( .A1(n14164), .A2(n20891), .B1(n20826), .B2(n14163), .ZN(
        n14142) );
  AOI21_X1 U17643 ( .B1(n14166), .B2(n20888), .A(n14142), .ZN(n14143) );
  OAI211_X1 U17644 ( .C1(n14170), .C2(n14145), .A(n14144), .B(n14143), .ZN(
        P1_U3098) );
  NAND2_X1 U17645 ( .A1(n14162), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14148) );
  OAI22_X1 U17646 ( .A1(n14164), .A2(n20885), .B1(n20815), .B2(n14163), .ZN(
        n14146) );
  AOI21_X1 U17647 ( .B1(n14166), .B2(n20882), .A(n14146), .ZN(n14147) );
  OAI211_X1 U17648 ( .C1(n14170), .C2(n14149), .A(n14148), .B(n14147), .ZN(
        P1_U3097) );
  NAND2_X1 U17649 ( .A1(n14162), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14152) );
  OAI22_X1 U17650 ( .A1(n14164), .A2(n20915), .B1(n20846), .B2(n14163), .ZN(
        n14150) );
  AOI21_X1 U17651 ( .B1(n14166), .B2(n20912), .A(n14150), .ZN(n14151) );
  OAI211_X1 U17652 ( .C1(n14170), .C2(n14153), .A(n14152), .B(n14151), .ZN(
        P1_U3102) );
  NAND2_X1 U17653 ( .A1(n14162), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14156) );
  OAI22_X1 U17654 ( .A1(n14164), .A2(n20921), .B1(n20851), .B2(n14163), .ZN(
        n14154) );
  AOI21_X1 U17655 ( .B1(n14166), .B2(n20918), .A(n14154), .ZN(n14155) );
  OAI211_X1 U17656 ( .C1(n14170), .C2(n14157), .A(n14156), .B(n14155), .ZN(
        P1_U3103) );
  NAND2_X1 U17657 ( .A1(n14162), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14160) );
  OAI22_X1 U17658 ( .A1(n14164), .A2(n20903), .B1(n20836), .B2(n14163), .ZN(
        n14158) );
  AOI21_X1 U17659 ( .B1(n14166), .B2(n20900), .A(n14158), .ZN(n14159) );
  OAI211_X1 U17660 ( .C1(n14170), .C2(n14161), .A(n14160), .B(n14159), .ZN(
        P1_U3100) );
  NAND2_X1 U17661 ( .A1(n14162), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14168) );
  OAI22_X1 U17662 ( .A1(n14164), .A2(n20909), .B1(n20841), .B2(n14163), .ZN(
        n14165) );
  AOI21_X1 U17663 ( .B1(n14166), .B2(n20906), .A(n14165), .ZN(n14167) );
  OAI211_X1 U17664 ( .C1(n14170), .C2(n14169), .A(n14168), .B(n14167), .ZN(
        P1_U3101) );
  NAND2_X1 U17665 ( .A1(n14172), .A2(n14171), .ZN(n14173) );
  NAND2_X1 U17666 ( .A1(n14174), .A2(n14173), .ZN(n16454) );
  NOR2_X1 U17667 ( .A1(n16454), .A2(n19716), .ZN(n14177) );
  AOI211_X1 U17668 ( .C1(n14175), .C2(n13662), .A(n19713), .B(n14081), .ZN(
        n14176) );
  AOI211_X1 U17669 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19716), .A(n14177), .B(
        n14176), .ZN(n14178) );
  INV_X1 U17670 ( .A(n14178), .ZN(P2_U2872) );
  OR2_X1 U17671 ( .A1(n14179), .A2(n14321), .ZN(n14180) );
  NAND2_X1 U17672 ( .A1(n14332), .A2(n14180), .ZN(n16448) );
  INV_X1 U17673 ( .A(n16448), .ZN(n19604) );
  OAI22_X1 U17674 ( .A1(n16155), .A2(n19780), .B1(n19744), .B2(n14181), .ZN(
        n14183) );
  INV_X1 U17675 ( .A(n19717), .ZN(n16158) );
  OAI22_X1 U17676 ( .A1(n16158), .A2(n18894), .B1(n16156), .B2(n21227), .ZN(
        n14182) );
  AOI211_X1 U17677 ( .C1(n19772), .C2(n19604), .A(n14183), .B(n14182), .ZN(
        n14184) );
  OAI21_X1 U17678 ( .B1(n14185), .B2(n19754), .A(n14184), .ZN(P2_U2903) );
  OAI21_X1 U17679 ( .B1(n20769), .B2(n14218), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14187) );
  NAND2_X1 U17680 ( .A1(n20776), .A2(n13840), .ZN(n14186) );
  AOI21_X1 U17681 ( .B1(n14187), .B2(n14186), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n14189) );
  NOR2_X1 U17682 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14188), .ZN(
        n14192) );
  NAND2_X1 U17683 ( .A1(n14214), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n14195) );
  NOR2_X1 U17684 ( .A1(n20868), .A2(n20807), .ZN(n14191) );
  NAND2_X1 U17685 ( .A1(n20701), .A2(n14190), .ZN(n20669) );
  INV_X1 U17686 ( .A(n20669), .ZN(n20665) );
  AOI22_X1 U17687 ( .A1(n20776), .A2(n14191), .B1(n20871), .B2(n20665), .ZN(
        n14216) );
  INV_X1 U17688 ( .A(n14192), .ZN(n14215) );
  OAI22_X1 U17689 ( .A1(n14216), .A2(n20897), .B1(n20831), .B2(n14215), .ZN(
        n14193) );
  AOI21_X1 U17690 ( .B1(n14218), .B2(n20893), .A(n14193), .ZN(n14194) );
  OAI211_X1 U17691 ( .C1(n14221), .C2(n20832), .A(n14195), .B(n14194), .ZN(
        P1_U3067) );
  NAND2_X1 U17692 ( .A1(n14214), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n14198) );
  OAI22_X1 U17693 ( .A1(n14216), .A2(n20885), .B1(n20815), .B2(n14215), .ZN(
        n14196) );
  AOI21_X1 U17694 ( .B1(n14218), .B2(n20875), .A(n14196), .ZN(n14197) );
  OAI211_X1 U17695 ( .C1(n14221), .C2(n20816), .A(n14198), .B(n14197), .ZN(
        P1_U3065) );
  NAND2_X1 U17696 ( .A1(n14214), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n14201) );
  OAI22_X1 U17697 ( .A1(n20931), .A2(n14216), .B1(n14215), .B2(n20857), .ZN(
        n14199) );
  AOI21_X1 U17698 ( .B1(n14218), .B2(n20924), .A(n14199), .ZN(n14200) );
  OAI211_X1 U17699 ( .C1(n14221), .C2(n20858), .A(n14201), .B(n14200), .ZN(
        P1_U3072) );
  NAND2_X1 U17700 ( .A1(n14214), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n14204) );
  OAI22_X1 U17701 ( .A1(n20921), .A2(n14216), .B1(n14215), .B2(n20851), .ZN(
        n14202) );
  AOI21_X1 U17702 ( .B1(n14218), .B2(n20917), .A(n14202), .ZN(n14203) );
  OAI211_X1 U17703 ( .C1(n14221), .C2(n20852), .A(n14204), .B(n14203), .ZN(
        P1_U3071) );
  NAND2_X1 U17704 ( .A1(n14214), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n14207) );
  OAI22_X1 U17705 ( .A1(n20915), .A2(n14216), .B1(n14215), .B2(n20846), .ZN(
        n14205) );
  AOI21_X1 U17706 ( .B1(n14218), .B2(n20911), .A(n14205), .ZN(n14206) );
  OAI211_X1 U17707 ( .C1(n14221), .C2(n20847), .A(n14207), .B(n14206), .ZN(
        P1_U3070) );
  NAND2_X1 U17708 ( .A1(n14214), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14210) );
  OAI22_X1 U17709 ( .A1(n20909), .A2(n14216), .B1(n14215), .B2(n20841), .ZN(
        n14208) );
  AOI21_X1 U17710 ( .B1(n14218), .B2(n20905), .A(n14208), .ZN(n14209) );
  OAI211_X1 U17711 ( .C1(n14221), .C2(n20842), .A(n14210), .B(n14209), .ZN(
        P1_U3069) );
  NAND2_X1 U17712 ( .A1(n14214), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n14213) );
  OAI22_X1 U17713 ( .A1(n14216), .A2(n20903), .B1(n20836), .B2(n14215), .ZN(
        n14211) );
  AOI21_X1 U17714 ( .B1(n14218), .B2(n20899), .A(n14211), .ZN(n14212) );
  OAI211_X1 U17715 ( .C1(n14221), .C2(n20837), .A(n14213), .B(n14212), .ZN(
        P1_U3068) );
  NAND2_X1 U17716 ( .A1(n14214), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n14220) );
  OAI22_X1 U17717 ( .A1(n14216), .A2(n20891), .B1(n20826), .B2(n14215), .ZN(
        n14217) );
  AOI21_X1 U17718 ( .B1(n14218), .B2(n20887), .A(n14217), .ZN(n14219) );
  OAI211_X1 U17719 ( .C1(n14221), .C2(n20827), .A(n14220), .B(n14219), .ZN(
        P1_U3066) );
  AOI21_X1 U17720 ( .B1(n21296), .B2(n14223), .A(n14351), .ZN(n14542) );
  OAI22_X1 U17721 ( .A1(n14542), .A2(n15101), .B1(n14830), .B2(n21296), .ZN(
        n14224) );
  AOI21_X1 U17722 ( .B1(n15246), .B2(P1_EAX_REG_8__SCAN_IN), .A(n14224), .ZN(
        n14236) );
  AOI22_X1 U17723 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14228) );
  AOI22_X1 U17724 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U17725 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14226) );
  AOI22_X1 U17726 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14225) );
  NAND4_X1 U17727 ( .A1(n14228), .A2(n14227), .A3(n14226), .A4(n14225), .ZN(
        n14234) );
  AOI22_X1 U17728 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14232) );
  AOI22_X1 U17729 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9710), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14231) );
  AOI22_X1 U17730 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14230) );
  AOI22_X1 U17731 ( .A1(n15040), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14229) );
  NAND4_X1 U17732 ( .A1(n14232), .A2(n14231), .A3(n14230), .A4(n14229), .ZN(
        n14233) );
  OAI21_X1 U17733 ( .B1(n14234), .B2(n14233), .A(n14780), .ZN(n14235) );
  OAI21_X1 U17734 ( .B1(n14237), .B2(n9733), .A(n14355), .ZN(n14545) );
  INV_X1 U17735 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20962) );
  NAND3_X1 U17736 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20577) );
  NOR2_X1 U17737 ( .A1(n20957), .A2(n20577), .ZN(n20564) );
  NAND3_X1 U17738 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n20564), .ZN(n20544) );
  NOR2_X1 U17739 ( .A1(n20962), .A2(n20544), .ZN(n14387) );
  NAND2_X1 U17740 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14387), .ZN(n15173) );
  NAND2_X1 U17741 ( .A1(n20578), .A2(n15180), .ZN(n16694) );
  OAI21_X1 U17742 ( .B1(n15173), .B2(n20565), .A(n16694), .ZN(n14238) );
  INV_X1 U17743 ( .A(n14238), .ZN(n20536) );
  NAND2_X1 U17744 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14239) );
  OAI211_X1 U17745 ( .C1(n15287), .C2(P1_EBX_REG_8__SCAN_IN), .A(n15149), .B(
        n14239), .ZN(n14240) );
  OAI21_X1 U17746 ( .B1(n15159), .B2(P1_EBX_REG_8__SCAN_IN), .A(n14240), .ZN(
        n14242) );
  AOI21_X1 U17747 ( .B1(n14242), .B2(n14241), .A(n10161), .ZN(n16845) );
  INV_X1 U17748 ( .A(n16845), .ZN(n14245) );
  OAI21_X1 U17749 ( .B1(n20581), .B2(n21296), .A(n16808), .ZN(n14243) );
  AOI21_X1 U17750 ( .B1(n20604), .B2(n14542), .A(n14243), .ZN(n14244) );
  OAI21_X1 U17751 ( .B1(n14245), .B2(n20580), .A(n14244), .ZN(n14249) );
  NAND2_X1 U17752 ( .A1(n20596), .A2(n14387), .ZN(n14247) );
  INV_X1 U17753 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14246) );
  OAI22_X1 U17754 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14247), .B1(n14246), 
        .B2(n20592), .ZN(n14248) );
  AOI211_X1 U17755 ( .C1(n20536), .C2(P1_REIP_REG_8__SCAN_IN), .A(n14249), .B(
        n14248), .ZN(n14250) );
  OAI21_X1 U17756 ( .B1(n14545), .B2(n15476), .A(n14250), .ZN(P1_U2832) );
  AOI22_X1 U17757 ( .A1(n15612), .A2(n15556), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15610), .ZN(n14251) );
  OAI21_X1 U17758 ( .B1(n14545), .B2(n15614), .A(n14251), .ZN(P1_U2896) );
  AOI22_X1 U17759 ( .A1(n16845), .A2(n21040), .B1(n21041), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n14252) );
  OAI21_X1 U17760 ( .B1(n14545), .B2(n15529), .A(n14252), .ZN(P1_U2864) );
  OAI21_X1 U17761 ( .B1(n19907), .B2(n19937), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14256) );
  NAND2_X1 U17762 ( .A1(n14256), .A2(n20458), .ZN(n14260) );
  INV_X1 U17763 ( .A(n14257), .ZN(n14258) );
  AND2_X1 U17764 ( .A1(n14258), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20361) );
  NAND2_X1 U17765 ( .A1(n19941), .A2(n20481), .ZN(n19917) );
  NOR2_X1 U17766 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19917), .ZN(
        n19906) );
  NOR2_X1 U17767 ( .A1(n20361), .A2(n19906), .ZN(n14263) );
  INV_X1 U17768 ( .A(n10765), .ZN(n14261) );
  OAI21_X1 U17769 ( .B1(n14261), .B2(n19906), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14259) );
  INV_X1 U17770 ( .A(n14260), .ZN(n14264) );
  AOI211_X1 U17771 ( .C1(n14261), .C2(n20101), .A(n19906), .B(n20458), .ZN(
        n14262) );
  AOI211_X2 U17772 ( .C1(n14264), .C2(n14263), .A(n20074), .B(n14262), .ZN(
        n19914) );
  AOI22_X1 U17773 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19909), .ZN(n20330) );
  AOI22_X1 U17774 ( .A1(n20285), .A2(n19937), .B1(n19906), .B2(n20326), .ZN(
        n14267) );
  AOI22_X1 U17775 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19909), .ZN(n20179) );
  NAND2_X1 U17776 ( .A1(n19907), .A2(n20327), .ZN(n14266) );
  OAI211_X1 U17777 ( .C1(n19914), .C2(n14268), .A(n14267), .B(n14266), .ZN(
        n14269) );
  AOI21_X1 U17778 ( .B1(n14253), .B2(n19911), .A(n14269), .ZN(n14270) );
  INV_X1 U17779 ( .A(n14270), .ZN(P2_U3049) );
  NOR2_X2 U17780 ( .A1(n16132), .A2(n20074), .ZN(n20350) );
  AOI22_X1 U17781 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19909), .ZN(n20354) );
  INV_X1 U17782 ( .A(n20354), .ZN(n20297) );
  AOI22_X1 U17783 ( .A1(n20297), .A2(n19937), .B1(n19906), .B2(n20349), .ZN(
        n14273) );
  AOI22_X1 U17784 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19909), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19910), .ZN(n20191) );
  NAND2_X1 U17785 ( .A1(n19907), .A2(n20351), .ZN(n14272) );
  OAI211_X1 U17786 ( .C1(n19914), .C2(n14274), .A(n14273), .B(n14272), .ZN(
        n14275) );
  AOI21_X1 U17787 ( .B1(n20350), .B2(n19911), .A(n14275), .ZN(n14276) );
  INV_X1 U17788 ( .A(n14276), .ZN(P2_U3053) );
  NOR2_X1 U17789 ( .A1(n19656), .A2(n14278), .ZN(n14280) );
  XNOR2_X1 U17790 ( .A(n14280), .B(n14279), .ZN(n14281) );
  INV_X1 U17791 ( .A(n19704), .ZN(n19684) );
  NAND2_X1 U17792 ( .A1(n14281), .A2(n19684), .ZN(n14290) );
  INV_X1 U17793 ( .A(n14282), .ZN(n14288) );
  OAI21_X1 U17794 ( .B1(n20403), .B2(n19676), .A(n19856), .ZN(n14284) );
  NOR2_X1 U17795 ( .A1(n10155), .A2(n19690), .ZN(n14283) );
  AOI211_X1 U17796 ( .C1(n19678), .C2(P2_EBX_REG_6__SCAN_IN), .A(n14284), .B(
        n14283), .ZN(n14285) );
  OAI21_X1 U17797 ( .B1(n14286), .B2(n19692), .A(n14285), .ZN(n14287) );
  AOI21_X1 U17798 ( .B1(n14288), .B2(n19698), .A(n14287), .ZN(n14289) );
  OAI211_X1 U17799 ( .C1(n19745), .C2(n19703), .A(n14290), .B(n14289), .ZN(
        P2_U2849) );
  XNOR2_X1 U17800 ( .A(n14291), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14314) );
  NAND2_X1 U17801 ( .A1(n9826), .A2(n14292), .ZN(n14293) );
  XNOR2_X1 U17802 ( .A(n14294), .B(n14293), .ZN(n14312) );
  INV_X1 U17803 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20405) );
  OAI22_X1 U17804 ( .A1(n17046), .A2(n14295), .B1(n20405), .B2(n19856), .ZN(
        n14296) );
  AOI21_X1 U17805 ( .B1(n17038), .B2(n14480), .A(n14296), .ZN(n14297) );
  OAI21_X1 U17806 ( .B1(n14298), .B2(n16307), .A(n14297), .ZN(n14299) );
  AOI21_X1 U17807 ( .B1(n14312), .B2(n19828), .A(n14299), .ZN(n14300) );
  OAI21_X1 U17808 ( .B1(n14314), .B2(n17039), .A(n14300), .ZN(P2_U3007) );
  NOR2_X1 U17809 ( .A1(n14302), .A2(n14301), .ZN(n14440) );
  OR2_X1 U17810 ( .A1(n14304), .A2(n14303), .ZN(n14305) );
  NAND2_X1 U17811 ( .A1(n14305), .A2(n14441), .ZN(n19743) );
  NAND3_X1 U17812 ( .A1(n14307), .A2(n14306), .A3(n10841), .ZN(n14439) );
  NAND2_X1 U17813 ( .A1(n19825), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n14308) );
  OAI211_X1 U17814 ( .C1(n19743), .C2(n17070), .A(n14439), .B(n14308), .ZN(
        n14309) );
  AOI21_X1 U17815 ( .B1(n17086), .B2(n14484), .A(n14309), .ZN(n14310) );
  OAI21_X1 U17816 ( .B1(n14440), .B2(n10841), .A(n14310), .ZN(n14311) );
  AOI21_X1 U17817 ( .B1(n14312), .B2(n19866), .A(n14311), .ZN(n14313) );
  OAI21_X1 U17818 ( .B1(n14314), .B2(n19859), .A(n14313), .ZN(P2_U3039) );
  INV_X1 U17819 ( .A(n14319), .ZN(n16304) );
  NAND2_X1 U17820 ( .A1(n19656), .A2(n19684), .ZN(n19710) );
  AOI21_X1 U17821 ( .B1(P2_REIP_REG_15__SCAN_IN), .B2(n19697), .A(n19825), 
        .ZN(n14316) );
  AOI22_X1 U17822 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n19678), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19672), .ZN(n14315) );
  OAI211_X1 U17823 ( .C1(n16304), .C2(n19710), .A(n14316), .B(n14315), .ZN(
        n14317) );
  INV_X1 U17824 ( .A(n14317), .ZN(n14327) );
  NOR2_X1 U17825 ( .A1(n19656), .A2(n19704), .ZN(n19636) );
  AOI21_X1 U17826 ( .B1(n14319), .B2(n14318), .A(n19598), .ZN(n14325) );
  OR2_X1 U17827 ( .A1(n14320), .A2(n17049), .ZN(n14323) );
  INV_X1 U17828 ( .A(n14321), .ZN(n14322) );
  NAND2_X1 U17829 ( .A1(n14323), .A2(n14322), .ZN(n19723) );
  OAI22_X1 U17830 ( .A1(n16454), .A2(n19687), .B1(n19723), .B2(n19703), .ZN(
        n14324) );
  AOI21_X1 U17831 ( .B1(n19636), .B2(n14325), .A(n14324), .ZN(n14326) );
  OAI211_X1 U17832 ( .C1(n14328), .C2(n19692), .A(n14327), .B(n14326), .ZN(
        P2_U2840) );
  AOI21_X1 U17833 ( .B1(n14330), .B2(n9715), .A(n14329), .ZN(n16971) );
  INV_X1 U17834 ( .A(n16971), .ZN(n14339) );
  NAND2_X1 U17835 ( .A1(n14332), .A2(n14331), .ZN(n14333) );
  NAND2_X1 U17836 ( .A1(n16153), .A2(n14333), .ZN(n16430) );
  INV_X1 U17837 ( .A(n16430), .ZN(n16015) );
  OAI22_X1 U17838 ( .A1(n16155), .A2(n14335), .B1(n19744), .B2(n14334), .ZN(
        n14336) );
  AOI21_X1 U17839 ( .B1(n19772), .B2(n16015), .A(n14336), .ZN(n14338) );
  AOI22_X1 U17840 ( .A1(n19717), .A2(BUF2_REG_17__SCAN_IN), .B1(n19719), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14337) );
  OAI211_X1 U17841 ( .C1(n14339), .C2(n19754), .A(n14338), .B(n14337), .ZN(
        P2_U2902) );
  AOI22_X1 U17842 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14343) );
  AOI22_X1 U17843 ( .A1(n15082), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14342) );
  AOI22_X1 U17844 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U17845 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14340) );
  NAND4_X1 U17846 ( .A1(n14343), .A2(n14342), .A3(n14341), .A4(n14340), .ZN(
        n14350) );
  AOI22_X1 U17847 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15072), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14348) );
  INV_X2 U17848 ( .A(n14344), .ZN(n15076) );
  AOI22_X1 U17849 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14347) );
  AOI22_X1 U17850 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14346) );
  AOI22_X1 U17851 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14345) );
  NAND4_X1 U17852 ( .A1(n14348), .A2(n14347), .A3(n14346), .A4(n14345), .ZN(
        n14349) );
  OAI21_X1 U17853 ( .B1(n14350), .B2(n14349), .A(n14780), .ZN(n14354) );
  XOR2_X1 U17854 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n14351), .Z(n20537) );
  INV_X1 U17855 ( .A(n20537), .ZN(n14590) );
  AOI22_X1 U17856 ( .A1(n14983), .A2(n14590), .B1(n15245), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14353) );
  NAND2_X1 U17857 ( .A1(n13958), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n14352) );
  NOR2_X2 U17858 ( .A1(n14355), .A2(n14451), .ZN(n14594) );
  AOI22_X1 U17859 ( .A1(n15083), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9710), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14359) );
  AOI22_X1 U17860 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15072), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14358) );
  AOI22_X1 U17861 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14357) );
  AOI22_X1 U17862 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14356) );
  NAND4_X1 U17863 ( .A1(n14359), .A2(n14358), .A3(n14357), .A4(n14356), .ZN(
        n14365) );
  AOI22_X1 U17864 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9708), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14363) );
  AOI22_X1 U17865 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14362) );
  AOI22_X1 U17866 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14361) );
  AOI22_X1 U17867 ( .A1(n14930), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14360) );
  NAND4_X1 U17868 ( .A1(n14363), .A2(n14362), .A3(n14361), .A4(n14360), .ZN(
        n14364) );
  OR2_X1 U17869 ( .A1(n14365), .A2(n14364), .ZN(n14366) );
  NAND2_X1 U17870 ( .A1(n14780), .A2(n14366), .ZN(n14370) );
  XNOR2_X1 U17871 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B(n14367), .ZN(
        n15787) );
  OAI22_X1 U17872 ( .A1(n15787), .A2(n15101), .B1(n14830), .B2(n15785), .ZN(
        n14368) );
  INV_X1 U17873 ( .A(n14368), .ZN(n14369) );
  OAI211_X1 U17874 ( .C1(n13616), .C2(n20630), .A(n14370), .B(n14369), .ZN(
        n14593) );
  XNOR2_X1 U17875 ( .A(n14450), .B(n14593), .ZN(n15790) );
  MUX2_X1 U17876 ( .A(n15159), .B(n15129), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n14371) );
  OAI21_X1 U17877 ( .B1(n15218), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n14371), .ZN(n14376) );
  OR2_X1 U17878 ( .A1(n15165), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n14375) );
  NAND2_X1 U17879 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14372) );
  NAND2_X1 U17880 ( .A1(n15149), .A2(n14372), .ZN(n14373) );
  OAI21_X1 U17881 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n15287), .A(n14373), .ZN(
        n14374) );
  AOI21_X1 U17882 ( .B1(n14376), .B2(n16835), .A(n14620), .ZN(n16826) );
  AOI22_X1 U17883 ( .A1(n16826), .A2(n21040), .B1(n21041), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n14377) );
  OAI21_X1 U17884 ( .B1(n15790), .B2(n15513), .A(n14377), .ZN(P1_U2862) );
  NOR2_X1 U17885 ( .A1(n19656), .A2(n14378), .ZN(n16535) );
  XNOR2_X1 U17886 ( .A(n16535), .B(n19839), .ZN(n14379) );
  NAND2_X1 U17887 ( .A1(n14379), .A2(n19684), .ZN(n14386) );
  NOR2_X1 U17888 ( .A1(n19869), .A2(n19687), .ZN(n14384) );
  AOI22_X1 U17889 ( .A1(n19697), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19672), .ZN(n14381) );
  NAND2_X1 U17890 ( .A1(n19678), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n14380) );
  OAI211_X1 U17891 ( .C1(n19692), .C2(n14382), .A(n14381), .B(n14380), .ZN(
        n14383) );
  AOI211_X1 U17892 ( .C1(n20468), .C2(n19671), .A(n14384), .B(n14383), .ZN(
        n14385) );
  OAI211_X1 U17893 ( .C1(n20466), .C2(n19688), .A(n14386), .B(n14385), .ZN(
        P2_U2853) );
  NAND2_X1 U17894 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15172) );
  AOI21_X1 U17895 ( .B1(n15172), .B2(n16694), .A(n20536), .ZN(n16727) );
  INV_X1 U17896 ( .A(n16727), .ZN(n14389) );
  INV_X1 U17897 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20964) );
  NAND3_X1 U17898 ( .A1(n20596), .A2(P1_REIP_REG_8__SCAN_IN), .A3(n14387), 
        .ZN(n20540) );
  NOR2_X1 U17899 ( .A1(n20964), .A2(n20540), .ZN(n14643) );
  INV_X1 U17900 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U17901 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n14389), .B1(n14643), 
        .B2(n14388), .ZN(n14393) );
  AOI22_X1 U17902 ( .A1(n15787), .A2(n20604), .B1(n20595), .B2(n16826), .ZN(
        n14390) );
  OAI211_X1 U17903 ( .C1(n20581), .C2(n15785), .A(n14390), .B(n16808), .ZN(
        n14391) );
  AOI21_X1 U17904 ( .B1(n20602), .B2(P1_EBX_REG_10__SCAN_IN), .A(n14391), .ZN(
        n14392) );
  OAI211_X1 U17905 ( .C1(n15790), .C2(n15476), .A(n14393), .B(n14392), .ZN(
        P1_U2830) );
  NAND2_X1 U17906 ( .A1(n14395), .A2(n14394), .ZN(n14398) );
  NAND2_X1 U17907 ( .A1(n14396), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14397) );
  NAND2_X1 U17908 ( .A1(n14398), .A2(n14397), .ZN(n16767) );
  XNOR2_X1 U17909 ( .A(n14407), .B(n14408), .ZN(n14402) );
  NAND2_X1 U17910 ( .A1(n14402), .A2(n14536), .ZN(n14403) );
  XNOR2_X1 U17911 ( .A(n14404), .B(n16868), .ZN(n16768) );
  NAND2_X1 U17912 ( .A1(n14404), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14405) );
  NAND3_X1 U17913 ( .A1(n14533), .A2(n14406), .A3(n14530), .ZN(n14412) );
  INV_X1 U17914 ( .A(n14407), .ZN(n14409) );
  NAND2_X1 U17915 ( .A1(n14409), .A2(n14408), .ZN(n14415) );
  XNOR2_X1 U17916 ( .A(n14415), .B(n14416), .ZN(n14410) );
  NAND2_X1 U17917 ( .A1(n14410), .A2(n14536), .ZN(n14411) );
  INV_X1 U17918 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21163) );
  NAND2_X1 U17919 ( .A1(n14413), .A2(n21163), .ZN(n16762) );
  INV_X1 U17920 ( .A(n14413), .ZN(n14414) );
  NAND2_X1 U17921 ( .A1(n14414), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16761) );
  INV_X1 U17922 ( .A(n14415), .ZN(n14417) );
  NAND2_X1 U17923 ( .A1(n14417), .A2(n14416), .ZN(n14534) );
  XNOR2_X1 U17924 ( .A(n14534), .B(n14535), .ZN(n14418) );
  AND2_X1 U17925 ( .A1(n14418), .A2(n14536), .ZN(n14419) );
  AOI21_X1 U17926 ( .B1(n14420), .B2(n14530), .A(n14419), .ZN(n14526) );
  INV_X1 U17927 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14523) );
  XNOR2_X1 U17928 ( .A(n14526), .B(n14523), .ZN(n14421) );
  XNOR2_X1 U17929 ( .A(n14525), .B(n14421), .ZN(n16756) );
  INV_X1 U17930 ( .A(n16756), .ZN(n14430) );
  INV_X1 U17931 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16868) );
  NOR2_X1 U17932 ( .A1(n16868), .A2(n14422), .ZN(n15233) );
  NAND2_X1 U17933 ( .A1(n15233), .A2(n16872), .ZN(n16859) );
  NOR2_X1 U17934 ( .A1(n21163), .A2(n16859), .ZN(n16848) );
  NOR2_X1 U17935 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14422), .ZN(
        n16871) );
  INV_X1 U17936 ( .A(n15222), .ZN(n14423) );
  NAND2_X1 U17937 ( .A1(n14424), .A2(n14423), .ZN(n14426) );
  INV_X1 U17938 ( .A(n15233), .ZN(n15221) );
  NOR2_X1 U17939 ( .A1(n14425), .A2(n15221), .ZN(n16823) );
  OAI21_X1 U17940 ( .B1(n16823), .B2(n15863), .A(n15228), .ZN(n15912) );
  AOI21_X1 U17941 ( .B1(n15224), .B2(n14426), .A(n15912), .ZN(n16867) );
  INV_X1 U17942 ( .A(n16867), .ZN(n14427) );
  AOI21_X1 U17943 ( .B1(n15234), .B2(n16871), .A(n14427), .ZN(n16865) );
  OAI21_X1 U17944 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15871), .A(
        n16865), .ZN(n16846) );
  OAI22_X1 U17945 ( .A1(n16808), .A2(n20962), .B1(n20652), .B2(n20550), .ZN(
        n14428) );
  AOI221_X1 U17946 ( .B1(n16848), .B2(n14523), .C1(n16846), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n14428), .ZN(n14429) );
  OAI21_X1 U17947 ( .B1(n14430), .B2(n20653), .A(n14429), .ZN(P1_U3024) );
  XNOR2_X1 U17948 ( .A(n14432), .B(n14433), .ZN(n17023) );
  NAND2_X1 U17949 ( .A1(n14435), .A2(n14434), .ZN(n14437) );
  XOR2_X1 U17950 ( .A(n14437), .B(n14436), .Z(n17024) );
  NAND2_X1 U17951 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19825), .ZN(n14438) );
  OAI221_X1 U17952 ( .B1(n10849), .B2(n14440), .C1(n10849), .C2(n14439), .A(
        n14438), .ZN(n14448) );
  AOI21_X1 U17953 ( .B1(n14442), .B2(n14441), .A(n14469), .ZN(n19739) );
  NOR3_X1 U17954 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n14444), .A3(
        n14443), .ZN(n14445) );
  AOI21_X1 U17955 ( .B1(n19854), .B2(n19739), .A(n14445), .ZN(n14446) );
  OAI21_X1 U17956 ( .B1(n19870), .B2(n19662), .A(n14446), .ZN(n14447) );
  AOI211_X1 U17957 ( .C1(n17024), .C2(n19866), .A(n14448), .B(n14447), .ZN(
        n14449) );
  OAI21_X1 U17958 ( .B1(n17023), .B2(n19859), .A(n14449), .ZN(P2_U3038) );
  AOI21_X1 U17959 ( .B1(n14451), .B2(n14355), .A(n14450), .ZN(n21043) );
  INV_X1 U17960 ( .A(n21043), .ZN(n14453) );
  AOI22_X1 U17961 ( .A1(n15612), .A2(n15552), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15610), .ZN(n14452) );
  OAI21_X1 U17962 ( .B1(n14453), .B2(n15614), .A(n14452), .ZN(P1_U2895) );
  NAND2_X1 U17963 ( .A1(n16007), .A2(n14454), .ZN(n14455) );
  XNOR2_X1 U17964 ( .A(n17029), .B(n14455), .ZN(n14464) );
  OAI21_X1 U17965 ( .B1(n21260), .B2(n19676), .A(n19838), .ZN(n14460) );
  NOR2_X1 U17966 ( .A1(n19690), .A2(n17036), .ZN(n14456) );
  AOI21_X1 U17967 ( .B1(n19678), .B2(P2_EBX_REG_5__SCAN_IN), .A(n14456), .ZN(
        n14457) );
  OAI21_X1 U17968 ( .B1(n14458), .B2(n19692), .A(n14457), .ZN(n14459) );
  NOR2_X1 U17969 ( .A1(n14460), .A2(n14459), .ZN(n14462) );
  NAND2_X1 U17970 ( .A1(n17033), .A2(n19698), .ZN(n14461) );
  OAI211_X1 U17971 ( .C1(n19757), .C2(n19703), .A(n14462), .B(n14461), .ZN(
        n14463) );
  AOI21_X1 U17972 ( .B1(n14464), .B2(n19684), .A(n14463), .ZN(n14465) );
  INV_X1 U17973 ( .A(n14465), .ZN(P2_U2850) );
  NAND2_X1 U17974 ( .A1(n16007), .A2(n14466), .ZN(n14467) );
  XNOR2_X1 U17975 ( .A(n17015), .B(n14467), .ZN(n14476) );
  OAI21_X1 U17976 ( .B1(n14469), .B2(n14468), .A(n16495), .ZN(n19738) );
  INV_X1 U17977 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20409) );
  AOI22_X1 U17978 ( .A1(n14470), .A2(n19679), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19672), .ZN(n14471) );
  OAI211_X1 U17979 ( .C1(n20409), .C2(n19676), .A(n14471), .B(n19856), .ZN(
        n14472) );
  AOI21_X1 U17980 ( .B1(P2_EBX_REG_9__SCAN_IN), .B2(n19678), .A(n14472), .ZN(
        n14474) );
  NAND2_X1 U17981 ( .A1(n17019), .A2(n19698), .ZN(n14473) );
  OAI211_X1 U17982 ( .C1(n19738), .C2(n19703), .A(n14474), .B(n14473), .ZN(
        n14475) );
  AOI21_X1 U17983 ( .B1(n14476), .B2(n19684), .A(n14475), .ZN(n14477) );
  INV_X1 U17984 ( .A(n14477), .ZN(P2_U2846) );
  NAND2_X1 U17985 ( .A1(n16007), .A2(n14478), .ZN(n14479) );
  XNOR2_X1 U17986 ( .A(n14480), .B(n14479), .ZN(n14488) );
  AOI22_X1 U17987 ( .A1(n14481), .A2(n19679), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19672), .ZN(n14482) );
  OAI211_X1 U17988 ( .C1(n20405), .C2(n19676), .A(n14482), .B(n19856), .ZN(
        n14483) );
  AOI21_X1 U17989 ( .B1(P2_EBX_REG_7__SCAN_IN), .B2(n19678), .A(n14483), .ZN(
        n14486) );
  NAND2_X1 U17990 ( .A1(n14484), .A2(n19698), .ZN(n14485) );
  OAI211_X1 U17991 ( .C1(n19743), .C2(n19703), .A(n14486), .B(n14485), .ZN(
        n14487) );
  AOI21_X1 U17992 ( .B1(n14488), .B2(n19684), .A(n14487), .ZN(n14489) );
  INV_X1 U17993 ( .A(n14489), .ZN(P2_U2848) );
  INV_X1 U17994 ( .A(n15549), .ZN(n14490) );
  OAI222_X1 U17995 ( .A1(n15606), .A2(n20630), .B1(n15608), .B2(n14490), .C1(
        n15614), .C2(n15790), .ZN(P1_U2894) );
  OAI21_X1 U17996 ( .B1(n17078), .B2(n14491), .A(n17051), .ZN(n19728) );
  NAND2_X1 U17997 ( .A1(n16007), .A2(n14492), .ZN(n14493) );
  XNOR2_X1 U17998 ( .A(n16985), .B(n14493), .ZN(n14501) );
  INV_X1 U17999 ( .A(n14494), .ZN(n17072) );
  INV_X1 U18000 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U18001 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n19678), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19672), .ZN(n14495) );
  OAI211_X1 U18002 ( .C1(n19676), .C2(n14496), .A(n14495), .B(n19856), .ZN(
        n14497) );
  AOI21_X1 U18003 ( .B1(n17072), .B2(n19698), .A(n14497), .ZN(n14498) );
  OAI21_X1 U18004 ( .B1(n14499), .B2(n19692), .A(n14498), .ZN(n14500) );
  AOI21_X1 U18005 ( .B1(n14501), .B2(n19684), .A(n14500), .ZN(n14502) );
  OAI21_X1 U18006 ( .B1(n19728), .B2(n19703), .A(n14502), .ZN(P2_U2842) );
  NAND2_X1 U18007 ( .A1(n16007), .A2(n14503), .ZN(n14504) );
  XNOR2_X1 U18008 ( .A(n17037), .B(n14504), .ZN(n14511) );
  OAI22_X1 U18009 ( .A1(n19676), .A2(n13356), .B1(n19690), .B2(n17047), .ZN(
        n14507) );
  NOR2_X1 U18010 ( .A1(n19692), .A2(n14505), .ZN(n14506) );
  AOI211_X1 U18011 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19678), .A(n14507), .B(
        n14506), .ZN(n14509) );
  OAI211_X1 U18012 ( .C1(n19748), .C2(n19703), .A(n14509), .B(n14508), .ZN(
        n14510) );
  AOI21_X1 U18013 ( .B1(n14511), .B2(n19684), .A(n14510), .ZN(n14512) );
  OAI21_X1 U18014 ( .B1(n19688), .B2(n19749), .A(n14512), .ZN(P2_U2852) );
  AOI21_X1 U18015 ( .B1(n19690), .B2(n19710), .A(n14513), .ZN(n14514) );
  INV_X1 U18016 ( .A(n14514), .ZN(n14522) );
  INV_X1 U18017 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n14518) );
  AOI22_X1 U18018 ( .A1(n19678), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n19679), .B2(
        n14515), .ZN(n14517) );
  INV_X1 U18019 ( .A(n16537), .ZN(n16529) );
  AOI22_X1 U18020 ( .A1(n19671), .A2(n19775), .B1(n19636), .B2(n16529), .ZN(
        n14516) );
  OAI211_X1 U18021 ( .C1(n14518), .C2(n19676), .A(n14517), .B(n14516), .ZN(
        n14519) );
  AOI21_X1 U18022 ( .B1(n14520), .B2(n19698), .A(n14519), .ZN(n14521) );
  OAI211_X1 U18023 ( .C1(n20487), .C2(n19688), .A(n14522), .B(n14521), .ZN(
        P2_U2855) );
  NAND2_X1 U18024 ( .A1(n14526), .A2(n14523), .ZN(n14524) );
  NAND2_X1 U18025 ( .A1(n14525), .A2(n14524), .ZN(n14529) );
  INV_X1 U18026 ( .A(n14526), .ZN(n14527) );
  NAND2_X1 U18027 ( .A1(n14527), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14528) );
  AND2_X1 U18028 ( .A1(n14531), .A2(n14530), .ZN(n14532) );
  INV_X1 U18029 ( .A(n14534), .ZN(n14537) );
  NAND3_X1 U18030 ( .A1(n14537), .A2(n14536), .A3(n14535), .ZN(n14538) );
  XNOR2_X1 U18031 ( .A(n14585), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14539) );
  NAND2_X1 U18032 ( .A1(n16847), .A2(n16772), .ZN(n14544) );
  INV_X1 U18033 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n14540) );
  OAI22_X1 U18034 ( .A1(n16774), .A2(n21296), .B1(n16808), .B2(n14540), .ZN(
        n14541) );
  AOI21_X1 U18035 ( .B1(n16742), .B2(n14542), .A(n14541), .ZN(n14543) );
  OAI211_X1 U18036 ( .C1(n16770), .C2(n14545), .A(n14544), .B(n14543), .ZN(
        P1_U2991) );
  INV_X1 U18037 ( .A(n14548), .ZN(n14579) );
  AOI21_X1 U18038 ( .B1(n14550), .B2(n14549), .A(n14579), .ZN(n14552) );
  INV_X1 U18039 ( .A(n14552), .ZN(n14551) );
  AOI22_X1 U18040 ( .A1(n14551), .A2(n15926), .B1(n14556), .B2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14581) );
  OAI21_X1 U18041 ( .B1(n14554), .B2(n14553), .A(n14552), .ZN(n14555) );
  AOI22_X1 U18042 ( .A1(n20923), .A2(n14579), .B1(
        P1_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n14578), .ZN(n14557) );
  OAI21_X1 U18043 ( .B1(n14581), .B2(n20931), .A(n14557), .ZN(n14558) );
  AOI21_X1 U18044 ( .B1(n20924), .B2(n20688), .A(n14558), .ZN(n14559) );
  OAI21_X1 U18045 ( .B1(n20858), .B2(n14584), .A(n14559), .ZN(P1_U3160) );
  AOI22_X1 U18046 ( .A1(n20892), .A2(n14579), .B1(
        P1_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n14578), .ZN(n14560) );
  OAI21_X1 U18047 ( .B1(n14581), .B2(n20897), .A(n14560), .ZN(n14561) );
  AOI21_X1 U18048 ( .B1(n20893), .B2(n20688), .A(n14561), .ZN(n14562) );
  OAI21_X1 U18049 ( .B1(n20832), .B2(n14584), .A(n14562), .ZN(P1_U3155) );
  AOI22_X1 U18050 ( .A1(n20916), .A2(n14579), .B1(
        P1_INSTQUEUE_REG_15__6__SCAN_IN), .B2(n14578), .ZN(n14563) );
  OAI21_X1 U18051 ( .B1(n14581), .B2(n20921), .A(n14563), .ZN(n14564) );
  AOI21_X1 U18052 ( .B1(n20917), .B2(n20688), .A(n14564), .ZN(n14565) );
  OAI21_X1 U18053 ( .B1(n20852), .B2(n14584), .A(n14565), .ZN(P1_U3159) );
  AOI22_X1 U18054 ( .A1(n20910), .A2(n14579), .B1(
        P1_INSTQUEUE_REG_15__5__SCAN_IN), .B2(n14578), .ZN(n14566) );
  OAI21_X1 U18055 ( .B1(n14581), .B2(n20915), .A(n14566), .ZN(n14567) );
  AOI21_X1 U18056 ( .B1(n20911), .B2(n20688), .A(n14567), .ZN(n14568) );
  OAI21_X1 U18057 ( .B1(n20847), .B2(n14584), .A(n14568), .ZN(P1_U3158) );
  AOI22_X1 U18058 ( .A1(n20904), .A2(n14579), .B1(
        P1_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n14578), .ZN(n14569) );
  OAI21_X1 U18059 ( .B1(n14581), .B2(n20909), .A(n14569), .ZN(n14570) );
  AOI21_X1 U18060 ( .B1(n20905), .B2(n20688), .A(n14570), .ZN(n14571) );
  OAI21_X1 U18061 ( .B1(n20842), .B2(n14584), .A(n14571), .ZN(P1_U3157) );
  AOI22_X1 U18062 ( .A1(n20898), .A2(n14579), .B1(
        P1_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n14578), .ZN(n14572) );
  OAI21_X1 U18063 ( .B1(n14581), .B2(n20903), .A(n14572), .ZN(n14573) );
  AOI21_X1 U18064 ( .B1(n20899), .B2(n20688), .A(n14573), .ZN(n14574) );
  OAI21_X1 U18065 ( .B1(n20837), .B2(n14584), .A(n14574), .ZN(P1_U3156) );
  AOI22_X1 U18066 ( .A1(n20886), .A2(n14579), .B1(
        P1_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n14578), .ZN(n14575) );
  OAI21_X1 U18067 ( .B1(n14581), .B2(n20891), .A(n14575), .ZN(n14576) );
  AOI21_X1 U18068 ( .B1(n20887), .B2(n20688), .A(n14576), .ZN(n14577) );
  OAI21_X1 U18069 ( .B1(n20827), .B2(n14584), .A(n14577), .ZN(P1_U3154) );
  AOI22_X1 U18070 ( .A1(n20874), .A2(n14579), .B1(
        P1_INSTQUEUE_REG_15__0__SCAN_IN), .B2(n14578), .ZN(n14580) );
  OAI21_X1 U18071 ( .B1(n14581), .B2(n20885), .A(n14580), .ZN(n14582) );
  AOI21_X1 U18072 ( .B1(n20875), .B2(n20688), .A(n14582), .ZN(n14583) );
  OAI21_X1 U18073 ( .B1(n20816), .B2(n14584), .A(n14583), .ZN(P1_U3153) );
  INV_X1 U18074 ( .A(n14585), .ZN(n14586) );
  INV_X1 U18075 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16849) );
  NAND2_X1 U18076 ( .A1(n14586), .A2(n16849), .ZN(n14587) );
  INV_X1 U18077 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16840) );
  XNOR2_X1 U18078 ( .A(n9714), .B(n16840), .ZN(n14588) );
  XNOR2_X1 U18079 ( .A(n15194), .B(n14588), .ZN(n16838) );
  AOI22_X1 U18080 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14589) );
  OAI21_X1 U18081 ( .B1(n16769), .B2(n14590), .A(n14589), .ZN(n14591) );
  AOI21_X1 U18082 ( .B1(n21043), .B2(n16764), .A(n14591), .ZN(n14592) );
  OAI21_X1 U18083 ( .B1(n16838), .B2(n20516), .A(n14592), .ZN(P1_U2990) );
  NAND2_X1 U18084 ( .A1(n13958), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n14597) );
  OAI21_X1 U18085 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n14595), .A(
        n14626), .ZN(n16755) );
  AOI22_X1 U18086 ( .A1(n14983), .A2(n16755), .B1(n15245), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14596) );
  AND2_X1 U18087 ( .A1(n14597), .A2(n14596), .ZN(n14598) );
  AOI22_X1 U18088 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14602) );
  AOI22_X1 U18089 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15081), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14601) );
  AOI22_X1 U18090 ( .A1(n15040), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14600) );
  AOI22_X1 U18091 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14599) );
  NAND4_X1 U18092 ( .A1(n14602), .A2(n14601), .A3(n14600), .A4(n14599), .ZN(
        n14608) );
  AOI22_X1 U18093 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14606) );
  AOI22_X1 U18094 ( .A1(n15083), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14605) );
  AOI22_X1 U18095 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14604) );
  AOI22_X1 U18096 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9702), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14603) );
  NAND4_X1 U18097 ( .A1(n14606), .A2(n14605), .A3(n14604), .A4(n14603), .ZN(
        n14607) );
  OR2_X1 U18098 ( .A1(n14608), .A2(n14607), .ZN(n14609) );
  AND2_X1 U18099 ( .A1(n14780), .A2(n14609), .ZN(n14611) );
  INV_X1 U18100 ( .A(n14611), .ZN(n14610) );
  NAND2_X1 U18101 ( .A1(n9770), .A2(n14610), .ZN(n14612) );
  AND2_X1 U18102 ( .A1(n14612), .A2(n14625), .ZN(n16752) );
  INV_X1 U18103 ( .A(n16752), .ZN(n14614) );
  AOI22_X1 U18104 ( .A1(n15612), .A2(n15545), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15610), .ZN(n14613) );
  OAI21_X1 U18105 ( .B1(n14614), .B2(n15614), .A(n14613), .ZN(P1_U2893) );
  INV_X1 U18106 ( .A(n15529), .ZN(n21042) );
  OR2_X1 U18107 ( .A1(n15165), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n14618) );
  INV_X1 U18108 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16750) );
  NAND2_X1 U18109 ( .A1(n15149), .A2(n16750), .ZN(n14616) );
  INV_X1 U18110 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n16724) );
  NAND2_X1 U18111 ( .A1(n15162), .A2(n16724), .ZN(n14615) );
  NAND3_X1 U18112 ( .A1(n14616), .A2(n15129), .A3(n14615), .ZN(n14617) );
  NAND2_X1 U18113 ( .A1(n14618), .A2(n14617), .ZN(n14619) );
  OR2_X1 U18114 ( .A1(n14620), .A2(n14619), .ZN(n14621) );
  NAND2_X1 U18115 ( .A1(n14649), .A2(n14621), .ZN(n16821) );
  OAI22_X1 U18116 ( .A1(n16821), .A2(n16730), .B1(n16724), .B2(n20618), .ZN(
        n14622) );
  AOI21_X1 U18117 ( .B1(n16752), .B2(n21042), .A(n14622), .ZN(n14623) );
  INV_X1 U18118 ( .A(n14623), .ZN(P1_U2861) );
  NAND2_X1 U18119 ( .A1(n14625), .A2(n14624), .ZN(n14641) );
  XOR2_X1 U18120 ( .A(n14645), .B(n14626), .Z(n16741) );
  AOI22_X1 U18121 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14630) );
  AOI22_X1 U18122 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14629) );
  AOI22_X1 U18123 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14628) );
  AOI22_X1 U18124 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n15086), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14627) );
  NAND4_X1 U18125 ( .A1(n14630), .A2(n14629), .A3(n14628), .A4(n14627), .ZN(
        n14636) );
  AOI22_X1 U18126 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n14985), .B1(
        n15082), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14634) );
  AOI22_X1 U18127 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n15076), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14633) );
  AOI22_X1 U18128 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n15081), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14632) );
  AOI22_X1 U18129 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14631) );
  NAND4_X1 U18130 ( .A1(n14634), .A2(n14633), .A3(n14632), .A4(n14631), .ZN(
        n14635) );
  OR2_X1 U18131 ( .A1(n14636), .A2(n14635), .ZN(n14637) );
  AOI22_X1 U18132 ( .A1(n14780), .A2(n14637), .B1(n15245), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14639) );
  NAND2_X1 U18133 ( .A1(n13958), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n14638) );
  OAI211_X1 U18134 ( .C1(n16741), .C2(n15101), .A(n14639), .B(n14638), .ZN(
        n14640) );
  OAI21_X1 U18135 ( .B1(n14641), .B2(n14640), .A(n14767), .ZN(n16740) );
  AOI22_X1 U18136 ( .A1(n15612), .A2(n15541), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15610), .ZN(n14642) );
  OAI21_X1 U18137 ( .B1(n16740), .B2(n15614), .A(n14642), .ZN(P1_U2892) );
  INV_X1 U18138 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21326) );
  INV_X1 U18139 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n16728) );
  NOR2_X1 U18140 ( .A1(n21326), .A2(n16728), .ZN(n15171) );
  OAI21_X1 U18141 ( .B1(n15171), .B2(n20578), .A(n16727), .ZN(n15474) );
  NAND2_X1 U18142 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n14643), .ZN(n16729) );
  OAI21_X1 U18143 ( .B1(n16728), .B2(n16729), .A(n21326), .ZN(n14655) );
  INV_X1 U18144 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14644) );
  OAI22_X1 U18145 ( .A1(n14645), .A2(n20581), .B1(n14644), .B2(n20592), .ZN(
        n14654) );
  NAND2_X1 U18146 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14646) );
  OAI211_X1 U18147 ( .C1(n15287), .C2(P1_EBX_REG_12__SCAN_IN), .A(n15149), .B(
        n14646), .ZN(n14647) );
  OAI21_X1 U18148 ( .B1(n15159), .B2(P1_EBX_REG_12__SCAN_IN), .A(n14647), .ZN(
        n14648) );
  NAND2_X1 U18149 ( .A1(n14649), .A2(n14648), .ZN(n14650) );
  AND2_X1 U18150 ( .A1(n15469), .A2(n14650), .ZN(n15920) );
  INV_X1 U18151 ( .A(n15920), .ZN(n14652) );
  AOI21_X1 U18152 ( .B1(n20604), .B2(n16741), .A(n13116), .ZN(n14651) );
  OAI21_X1 U18153 ( .B1(n14652), .B2(n20580), .A(n14651), .ZN(n14653) );
  AOI211_X1 U18154 ( .C1(n15474), .C2(n14655), .A(n14654), .B(n14653), .ZN(
        n14656) );
  OAI21_X1 U18155 ( .B1(n16740), .B2(n15476), .A(n14656), .ZN(P1_U2828) );
  AOI22_X1 U18156 ( .A1(n15920), .A2(n21040), .B1(n21041), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n14657) );
  OAI21_X1 U18157 ( .B1(n16740), .B2(n15529), .A(n14657), .ZN(P1_U2860) );
  AND2_X1 U18158 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17660) );
  INV_X1 U18159 ( .A(n18929), .ZN(n17969) );
  AND2_X1 U18160 ( .A1(n18929), .A2(n18914), .ZN(n14660) );
  INV_X1 U18161 ( .A(n19321), .ZN(n14659) );
  NOR2_X1 U18162 ( .A1(n17969), .A2(n17911), .ZN(n17920) );
  INV_X1 U18163 ( .A(n17920), .ZN(n17918) );
  NOR2_X2 U18164 ( .A1(n17911), .A2(n18929), .ZN(n17921) );
  INV_X1 U18165 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17627) );
  INV_X1 U18166 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17625) );
  INV_X1 U18167 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17812) );
  INV_X1 U18168 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17890) );
  INV_X1 U18169 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17910) );
  NAND2_X1 U18170 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17912) );
  NOR2_X1 U18171 ( .A1(n17910), .A2(n17912), .ZN(n17902) );
  NAND3_X1 U18172 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17902), .ZN(n17903) );
  NAND2_X1 U18173 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17895), .ZN(n17891) );
  NAND2_X1 U18174 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17685), .ZN(n17679) );
  AOI22_X1 U18175 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14665) );
  AOI22_X1 U18176 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14664) );
  AOI22_X1 U18177 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17820), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14663) );
  AOI22_X1 U18178 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14662) );
  NAND4_X1 U18179 ( .A1(n14665), .A2(n14664), .A3(n14663), .A4(n14662), .ZN(
        n14671) );
  AOI22_X1 U18180 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14669) );
  AOI22_X1 U18181 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14668) );
  AOI22_X1 U18182 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14667) );
  AOI22_X1 U18183 ( .A1(n12093), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14666) );
  NAND4_X1 U18184 ( .A1(n14669), .A2(n14668), .A3(n14667), .A4(n14666), .ZN(
        n14670) );
  NOR2_X1 U18185 ( .A1(n14671), .A2(n14670), .ZN(n17669) );
  AOI22_X1 U18186 ( .A1(n17820), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14675) );
  AOI22_X1 U18187 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14674) );
  AOI22_X1 U18188 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12130), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14673) );
  AOI22_X1 U18189 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17855), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14672) );
  NAND4_X1 U18190 ( .A1(n14675), .A2(n14674), .A3(n14673), .A4(n14672), .ZN(
        n14681) );
  AOI22_X1 U18191 ( .A1(n16555), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14679) );
  AOI22_X1 U18192 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14678) );
  AOI22_X1 U18193 ( .A1(n12175), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17826), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14677) );
  AOI22_X1 U18194 ( .A1(n12093), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14676) );
  NAND4_X1 U18195 ( .A1(n14679), .A2(n14678), .A3(n14677), .A4(n14676), .ZN(
        n14680) );
  NOR2_X1 U18196 ( .A1(n14681), .A2(n14680), .ZN(n17676) );
  AOI22_X1 U18197 ( .A1(n17879), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14685) );
  AOI22_X1 U18198 ( .A1(n17758), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14684) );
  AOI22_X1 U18199 ( .A1(n9698), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17826), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14683) );
  AOI22_X1 U18200 ( .A1(n17844), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14682) );
  NAND4_X1 U18201 ( .A1(n14685), .A2(n14684), .A3(n14683), .A4(n14682), .ZN(
        n14691) );
  AOI22_X1 U18202 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14689) );
  AOI22_X1 U18203 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14688) );
  AOI22_X1 U18204 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17839), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14687) );
  AOI22_X1 U18205 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14686) );
  NAND4_X1 U18206 ( .A1(n14689), .A2(n14688), .A3(n14687), .A4(n14686), .ZN(
        n14690) );
  NOR2_X1 U18207 ( .A1(n14691), .A2(n14690), .ZN(n17687) );
  AOI22_X1 U18208 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17855), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14695) );
  AOI22_X1 U18209 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14694) );
  AOI22_X1 U18210 ( .A1(n12105), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14693) );
  AOI22_X1 U18211 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14692) );
  NAND4_X1 U18212 ( .A1(n14695), .A2(n14694), .A3(n14693), .A4(n14692), .ZN(
        n14701) );
  AOI22_X1 U18213 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14699) );
  AOI22_X1 U18214 ( .A1(n17820), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14698) );
  AOI22_X1 U18215 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14697) );
  AOI22_X1 U18216 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14696) );
  NAND4_X1 U18217 ( .A1(n14699), .A2(n14698), .A3(n14697), .A4(n14696), .ZN(
        n14700) );
  NOR2_X1 U18218 ( .A1(n14701), .A2(n14700), .ZN(n17686) );
  NOR2_X1 U18219 ( .A1(n17687), .A2(n17686), .ZN(n17682) );
  AOI22_X1 U18220 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17860), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14711) );
  AOI22_X1 U18221 ( .A1(n17879), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14710) );
  INV_X1 U18222 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n21147) );
  AOI22_X1 U18223 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14702) );
  OAI21_X1 U18224 ( .B1(n21147), .B2(n17745), .A(n14702), .ZN(n14708) );
  AOI22_X1 U18225 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17839), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n16556), .ZN(n14706) );
  AOI22_X1 U18226 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17826), .B1(
        n12093), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14705) );
  AOI22_X1 U18227 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9697), .ZN(n14704) );
  AOI22_X1 U18228 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12130), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14703) );
  NAND4_X1 U18229 ( .A1(n14706), .A2(n14705), .A3(n14704), .A4(n14703), .ZN(
        n14707) );
  AOI211_X1 U18230 ( .C1(n17763), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n14708), .B(n14707), .ZN(n14709) );
  NAND3_X1 U18231 ( .A1(n14711), .A2(n14710), .A3(n14709), .ZN(n17681) );
  NAND2_X1 U18232 ( .A1(n17682), .A2(n17681), .ZN(n17680) );
  NOR2_X1 U18233 ( .A1(n17676), .A2(n17680), .ZN(n17949) );
  AOI22_X1 U18234 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14721) );
  AOI22_X1 U18235 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17839), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14720) );
  INV_X1 U18236 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n21137) );
  AOI22_X1 U18237 ( .A1(n9698), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14712) );
  OAI21_X1 U18238 ( .B1(n17877), .B2(n21137), .A(n14712), .ZN(n14718) );
  AOI22_X1 U18239 ( .A1(n17873), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14716) );
  AOI22_X1 U18240 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14715) );
  AOI22_X1 U18241 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14714) );
  AOI22_X1 U18242 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14713) );
  NAND4_X1 U18243 ( .A1(n14716), .A2(n14715), .A3(n14714), .A4(n14713), .ZN(
        n14717) );
  AOI211_X1 U18244 ( .C1(n17752), .C2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n14718), .B(n14717), .ZN(n14719) );
  NAND3_X1 U18245 ( .A1(n14721), .A2(n14720), .A3(n14719), .ZN(n17948) );
  NAND2_X1 U18246 ( .A1(n17949), .A2(n17948), .ZN(n17947) );
  NOR2_X1 U18247 ( .A1(n17669), .A2(n17947), .ZN(n17668) );
  INV_X1 U18248 ( .A(n17668), .ZN(n17662) );
  AOI22_X1 U18249 ( .A1(n9698), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14725) );
  AOI22_X1 U18250 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14724) );
  AOI22_X1 U18251 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14723) );
  AOI22_X1 U18252 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14722) );
  NAND4_X1 U18253 ( .A1(n14725), .A2(n14724), .A3(n14723), .A4(n14722), .ZN(
        n14731) );
  AOI22_X1 U18254 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12093), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14729) );
  AOI22_X1 U18255 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14728) );
  AOI22_X1 U18256 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14727) );
  AOI22_X1 U18257 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14726) );
  NAND4_X1 U18258 ( .A1(n14729), .A2(n14728), .A3(n14727), .A4(n14726), .ZN(
        n14730) );
  NOR2_X1 U18259 ( .A1(n14731), .A2(n14730), .ZN(n17661) );
  XOR2_X1 U18260 ( .A(n17662), .B(n17661), .Z(n17939) );
  AOI22_X1 U18261 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17665), .B1(n17921), 
        .B2(n17939), .ZN(n14735) );
  INV_X1 U18262 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14733) );
  INV_X1 U18263 ( .A(n17672), .ZN(n14732) );
  NAND3_X1 U18264 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14733), .A3(n14732), 
        .ZN(n14734) );
  NAND2_X1 U18265 ( .A1(n14735), .A2(n14734), .ZN(P3_U2675) );
  NOR3_X1 U18266 ( .A1(n14739), .A2(n14740), .A3(n21010), .ZN(n14738) );
  NAND2_X1 U18267 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21007) );
  AOI22_X1 U18268 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14736), .B2(n15217), .ZN(
        n21005) );
  NOR2_X1 U18269 ( .A1(n21007), .A2(n21005), .ZN(n14737) );
  OAI21_X1 U18270 ( .B1(n14738), .B2(n14737), .A(n21014), .ZN(n14748) );
  NOR3_X1 U18271 ( .A1(n12761), .A2(n14740), .A3(n14739), .ZN(n14741) );
  AOI21_X1 U18272 ( .B1(n14742), .B2(n9712), .A(n14741), .ZN(n14743) );
  OAI21_X1 U18273 ( .B1(n13840), .B2(n14744), .A(n14743), .ZN(n16617) );
  INV_X1 U18274 ( .A(n14745), .ZN(n14746) );
  NAND2_X1 U18275 ( .A1(n16617), .A2(n14746), .ZN(n14747) );
  OAI211_X1 U18276 ( .C1(n21014), .C2(n9712), .A(n14748), .B(n14747), .ZN(
        P1_U3473) );
  INV_X1 U18277 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14749) );
  XNOR2_X1 U18278 ( .A(n14750), .B(n14749), .ZN(n15772) );
  OR2_X1 U18279 ( .A1(n15772), .A2(n15101), .ZN(n14766) );
  AOI22_X1 U18280 ( .A1(n15082), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15081), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14754) );
  AOI22_X1 U18281 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15071), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14753) );
  AOI22_X1 U18282 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14752) );
  AOI22_X1 U18283 ( .A1(n14930), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14751) );
  NAND4_X1 U18284 ( .A1(n14754), .A2(n14753), .A3(n14752), .A4(n14751), .ZN(
        n14760) );
  AOI22_X1 U18285 ( .A1(n15083), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14758) );
  AOI22_X1 U18286 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14757) );
  AOI22_X1 U18287 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14756) );
  AOI22_X1 U18288 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14755) );
  NAND4_X1 U18289 ( .A1(n14758), .A2(n14757), .A3(n14756), .A4(n14755), .ZN(
        n14759) );
  NOR2_X1 U18290 ( .A1(n14760), .A2(n14759), .ZN(n14763) );
  NAND2_X1 U18291 ( .A1(n13958), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n14762) );
  NAND2_X1 U18292 ( .A1(n15245), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14761) );
  OAI211_X1 U18293 ( .C1(n14797), .C2(n14763), .A(n14762), .B(n14761), .ZN(
        n14764) );
  INV_X1 U18294 ( .A(n14764), .ZN(n14765) );
  XOR2_X1 U18295 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n14768), .Z(
        n16735) );
  AOI22_X1 U18296 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14772) );
  AOI22_X1 U18297 ( .A1(n15082), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14771) );
  AOI22_X1 U18298 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14770) );
  AOI22_X1 U18299 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14769) );
  NAND4_X1 U18300 ( .A1(n14772), .A2(n14771), .A3(n14770), .A4(n14769), .ZN(
        n14778) );
  AOI22_X1 U18301 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14776) );
  AOI22_X1 U18302 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14775) );
  AOI22_X1 U18303 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14929), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14774) );
  AOI22_X1 U18304 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14773) );
  NAND4_X1 U18305 ( .A1(n14776), .A2(n14775), .A3(n14774), .A4(n14773), .ZN(
        n14777) );
  OR2_X1 U18306 ( .A1(n14778), .A2(n14777), .ZN(n14779) );
  AOI22_X1 U18307 ( .A1(n14780), .A2(n14779), .B1(n15245), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U18308 ( .A1(n13958), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n14781) );
  OAI211_X1 U18309 ( .C1(n16735), .C2(n15101), .A(n14782), .B(n14781), .ZN(
        n15521) );
  XNOR2_X1 U18310 ( .A(n14783), .B(n16704), .ZN(n16710) );
  NAND2_X1 U18311 ( .A1(n16710), .A2(n14983), .ZN(n14800) );
  AOI22_X1 U18312 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14787) );
  AOI22_X1 U18313 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14908), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14786) );
  AOI22_X1 U18314 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14785) );
  AOI22_X1 U18315 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14784) );
  NAND4_X1 U18316 ( .A1(n14787), .A2(n14786), .A3(n14785), .A4(n14784), .ZN(
        n14793) );
  AOI22_X1 U18317 ( .A1(n15040), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14791) );
  AOI22_X1 U18318 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14790) );
  AOI22_X1 U18319 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14929), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14789) );
  AOI22_X1 U18320 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14788) );
  NAND4_X1 U18321 ( .A1(n14791), .A2(n14790), .A3(n14789), .A4(n14788), .ZN(
        n14792) );
  NOR2_X1 U18322 ( .A1(n14793), .A2(n14792), .ZN(n14796) );
  NAND2_X1 U18323 ( .A1(n15246), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n14795) );
  NAND2_X1 U18324 ( .A1(n15245), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14794) );
  OAI211_X1 U18325 ( .C1(n14797), .C2(n14796), .A(n14795), .B(n14794), .ZN(
        n14798) );
  INV_X1 U18326 ( .A(n14798), .ZN(n14799) );
  NAND2_X1 U18327 ( .A1(n14800), .A2(n14799), .ZN(n15515) );
  INV_X1 U18328 ( .A(n15514), .ZN(n14818) );
  INV_X1 U18329 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15749) );
  INV_X1 U18330 ( .A(n14801), .ZN(n14802) );
  NAND2_X1 U18331 ( .A1(n15749), .A2(n14802), .ZN(n14803) );
  AND2_X1 U18332 ( .A1(n14803), .A2(n14829), .ZN(n16696) );
  AOI22_X1 U18333 ( .A1(n15082), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15081), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14807) );
  AOI22_X1 U18334 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14806) );
  AOI22_X1 U18335 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14805) );
  AOI22_X1 U18336 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9702), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14804) );
  NAND4_X1 U18337 ( .A1(n14807), .A2(n14806), .A3(n14805), .A4(n14804), .ZN(
        n14813) );
  AOI22_X1 U18338 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14811) );
  AOI22_X1 U18339 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14992), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14810) );
  AOI22_X1 U18340 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14929), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U18341 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14808) );
  NAND4_X1 U18342 ( .A1(n14811), .A2(n14810), .A3(n14809), .A4(n14808), .ZN(
        n14812) );
  OR2_X1 U18343 ( .A1(n14813), .A2(n14812), .ZN(n14815) );
  OAI22_X1 U18344 ( .A1(n13616), .A2(n15593), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15749), .ZN(n14814) );
  AOI21_X1 U18345 ( .B1(n15067), .B2(n14815), .A(n14814), .ZN(n14816) );
  MUX2_X1 U18346 ( .A(n16696), .B(n14816), .S(n15101), .Z(n15591) );
  NAND2_X1 U18347 ( .A1(n14818), .A2(n14817), .ZN(n15504) );
  INV_X1 U18348 ( .A(n15504), .ZN(n14835) );
  AOI22_X1 U18349 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14822) );
  AOI22_X1 U18350 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14908), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14821) );
  AOI22_X1 U18351 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14820) );
  AOI22_X1 U18352 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14819) );
  NAND4_X1 U18353 ( .A1(n14822), .A2(n14821), .A3(n14820), .A4(n14819), .ZN(
        n14828) );
  AOI22_X1 U18354 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14826) );
  AOI22_X1 U18355 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14825) );
  AOI22_X1 U18356 ( .A1(n9707), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14824) );
  AOI22_X1 U18357 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9701), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14823) );
  NAND4_X1 U18358 ( .A1(n14826), .A2(n14825), .A3(n14824), .A4(n14823), .ZN(
        n14827) );
  OAI21_X1 U18359 ( .B1(n14828), .B2(n14827), .A(n15067), .ZN(n14833) );
  XNOR2_X1 U18360 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n14829), .ZN(
        n16685) );
  INV_X1 U18361 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15739) );
  OAI22_X1 U18362 ( .A1(n16685), .A2(n15101), .B1(n14830), .B2(n15739), .ZN(
        n14831) );
  AOI21_X1 U18363 ( .B1(n13958), .B2(P1_EAX_REG_17__SCAN_IN), .A(n14831), .ZN(
        n14832) );
  INV_X1 U18364 ( .A(n15505), .ZN(n14834) );
  INV_X1 U18365 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14849) );
  INV_X1 U18366 ( .A(n14836), .ZN(n14837) );
  NAND2_X1 U18367 ( .A1(n14849), .A2(n14837), .ZN(n14838) );
  NAND2_X1 U18368 ( .A1(n14855), .A2(n14838), .ZN(n15727) );
  INV_X1 U18369 ( .A(n15727), .ZN(n14853) );
  AOI22_X1 U18370 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14842) );
  AOI22_X1 U18371 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14841) );
  AOI22_X1 U18372 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14840) );
  AOI22_X1 U18373 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9702), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14839) );
  NAND4_X1 U18374 ( .A1(n14842), .A2(n14841), .A3(n14840), .A4(n14839), .ZN(
        n14848) );
  AOI22_X1 U18375 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15082), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14846) );
  AOI22_X1 U18376 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14845) );
  AOI22_X1 U18377 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14844) );
  AOI22_X1 U18378 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14929), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14843) );
  NAND4_X1 U18379 ( .A1(n14846), .A2(n14845), .A3(n14844), .A4(n14843), .ZN(
        n14847) );
  OR2_X1 U18380 ( .A1(n14848), .A2(n14847), .ZN(n14851) );
  OAI22_X1 U18381 ( .A1(n13616), .A2(n13062), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14849), .ZN(n14850) );
  AOI21_X1 U18382 ( .B1(n15067), .B2(n14851), .A(n14850), .ZN(n14852) );
  MUX2_X1 U18383 ( .A(n14853), .B(n14852), .S(n15101), .Z(n15455) );
  XNOR2_X1 U18384 ( .A(n14855), .B(n14854), .ZN(n15719) );
  AOI22_X1 U18385 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14859) );
  AOI22_X1 U18386 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14858) );
  AOI22_X1 U18387 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14857) );
  AOI22_X1 U18388 ( .A1(n9708), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14929), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14856) );
  NAND4_X1 U18389 ( .A1(n14859), .A2(n14858), .A3(n14857), .A4(n14856), .ZN(
        n14865) );
  AOI22_X1 U18390 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14863) );
  AOI22_X1 U18391 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14862) );
  AOI22_X1 U18392 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14861) );
  AOI22_X1 U18393 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9701), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14860) );
  NAND4_X1 U18394 ( .A1(n14863), .A2(n14862), .A3(n14861), .A4(n14860), .ZN(
        n14864) );
  NOR2_X1 U18395 ( .A1(n14865), .A2(n14864), .ZN(n14867) );
  AOI22_X1 U18396 ( .A1(n15246), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n14046), .ZN(n14866) );
  OAI21_X1 U18397 ( .B1(n15099), .B2(n14867), .A(n14866), .ZN(n14868) );
  MUX2_X1 U18398 ( .A(n15719), .B(n14868), .S(n15101), .Z(n15440) );
  AOI22_X1 U18399 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14872) );
  AOI22_X1 U18400 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n14985), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14871) );
  AOI22_X1 U18401 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14870) );
  AOI22_X1 U18402 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n15081), .B1(
        n14929), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14869) );
  NAND4_X1 U18403 ( .A1(n14872), .A2(n14871), .A3(n14870), .A4(n14869), .ZN(
        n14878) );
  AOI22_X1 U18404 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14876) );
  AOI22_X1 U18405 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n15040), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14875) );
  AOI22_X1 U18406 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9702), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14874) );
  AOI22_X1 U18407 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14930), .B1(
        n14992), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14873) );
  NAND4_X1 U18408 ( .A1(n14876), .A2(n14875), .A3(n14874), .A4(n14873), .ZN(
        n14877) );
  NOR2_X1 U18409 ( .A1(n14878), .A2(n14877), .ZN(n14882) );
  OAI21_X1 U18410 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20514), .A(
        n14046), .ZN(n14879) );
  INV_X1 U18411 ( .A(n14879), .ZN(n14880) );
  AOI21_X1 U18412 ( .B1(n13958), .B2(P1_EAX_REG_20__SCAN_IN), .A(n14880), .ZN(
        n14881) );
  OAI21_X1 U18413 ( .B1(n15099), .B2(n14882), .A(n14881), .ZN(n14887) );
  INV_X1 U18414 ( .A(n14883), .ZN(n14884) );
  INV_X1 U18415 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15428) );
  NAND2_X1 U18416 ( .A1(n14884), .A2(n15428), .ZN(n14885) );
  NAND2_X1 U18417 ( .A1(n14888), .A2(n14885), .ZN(n15712) );
  OR2_X1 U18418 ( .A1(n15712), .A2(n15101), .ZN(n14886) );
  INV_X1 U18419 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15419) );
  XNOR2_X1 U18420 ( .A(n14888), .B(n15419), .ZN(n15704) );
  AOI22_X1 U18421 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14892) );
  AOI22_X1 U18422 ( .A1(n15082), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14891) );
  AOI22_X1 U18423 ( .A1(n15035), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9701), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14890) );
  AOI22_X1 U18424 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14889) );
  NAND4_X1 U18425 ( .A1(n14892), .A2(n14891), .A3(n14890), .A4(n14889), .ZN(
        n14898) );
  AOI22_X1 U18426 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15086), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14896) );
  AOI22_X1 U18427 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14992), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14895) );
  AOI22_X1 U18428 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14929), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14894) );
  AOI22_X1 U18429 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14893) );
  NAND4_X1 U18430 ( .A1(n14896), .A2(n14895), .A3(n14894), .A4(n14893), .ZN(
        n14897) );
  NOR2_X1 U18431 ( .A1(n14898), .A2(n14897), .ZN(n14900) );
  AOI22_X1 U18432 ( .A1(n15246), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n14046), .ZN(n14899) );
  OAI21_X1 U18433 ( .B1(n15099), .B2(n14900), .A(n14899), .ZN(n14901) );
  MUX2_X1 U18434 ( .A(n15704), .B(n14901), .S(n15101), .Z(n15415) );
  AND2_X2 U18435 ( .A1(n15413), .A2(n15415), .ZN(n15338) );
  NAND2_X1 U18436 ( .A1(n14902), .A2(n15344), .ZN(n14903) );
  NAND2_X1 U18437 ( .A1(n15012), .A2(n14903), .ZN(n15662) );
  AOI22_X1 U18438 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14907) );
  AOI22_X1 U18439 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14906) );
  AOI22_X1 U18440 ( .A1(n14930), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14905) );
  AOI22_X1 U18441 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14904) );
  NAND4_X1 U18442 ( .A1(n14907), .A2(n14906), .A3(n14905), .A4(n14904), .ZN(
        n14914) );
  AOI22_X1 U18443 ( .A1(n15083), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14912) );
  AOI22_X1 U18444 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14908), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14911) );
  AOI22_X1 U18445 ( .A1(n9708), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15081), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14910) );
  AOI22_X1 U18446 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14909) );
  NAND4_X1 U18447 ( .A1(n14912), .A2(n14911), .A3(n14910), .A4(n14909), .ZN(
        n14913) );
  NOR2_X1 U18448 ( .A1(n14914), .A2(n14913), .ZN(n14962) );
  AOI22_X1 U18449 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14918) );
  AOI22_X1 U18450 ( .A1(n14948), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14917) );
  AOI22_X1 U18451 ( .A1(n9710), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14916) );
  AOI22_X1 U18452 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14915) );
  NAND4_X1 U18453 ( .A1(n14918), .A2(n14917), .A3(n14916), .A4(n14915), .ZN(
        n14924) );
  AOI22_X1 U18454 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15071), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14922) );
  AOI22_X1 U18455 ( .A1(n15082), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14921) );
  AOI22_X1 U18456 ( .A1(n15015), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14920) );
  AOI22_X1 U18457 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9694), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14919) );
  NAND4_X1 U18458 ( .A1(n14922), .A2(n14921), .A3(n14920), .A4(n14919), .ZN(
        n14923) );
  NOR2_X1 U18459 ( .A1(n14924), .A2(n14923), .ZN(n14979) );
  AOI22_X1 U18460 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15071), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14928) );
  AOI22_X1 U18461 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13960), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14927) );
  AOI22_X1 U18462 ( .A1(n15083), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14926) );
  AOI22_X1 U18463 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14925) );
  NAND4_X1 U18464 ( .A1(n14928), .A2(n14927), .A3(n14926), .A4(n14925), .ZN(
        n14936) );
  AOI22_X1 U18465 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15040), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14934) );
  AOI22_X1 U18466 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14929), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14933) );
  AOI22_X1 U18467 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14932) );
  AOI22_X1 U18468 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15074), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14931) );
  NAND4_X1 U18469 ( .A1(n14934), .A2(n14933), .A3(n14932), .A4(n14931), .ZN(
        n14935) );
  NOR2_X1 U18470 ( .A1(n14936), .A2(n14935), .ZN(n14980) );
  NOR2_X1 U18471 ( .A1(n14979), .A2(n14980), .ZN(n14975) );
  AOI22_X1 U18472 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15059), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14940) );
  AOI22_X1 U18473 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14939) );
  AOI22_X1 U18474 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14938) );
  AOI22_X1 U18475 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14937) );
  NAND4_X1 U18476 ( .A1(n14940), .A2(n14939), .A3(n14938), .A4(n14937), .ZN(
        n14946) );
  AOI22_X1 U18477 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n15082), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U18478 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14943) );
  AOI22_X1 U18479 ( .A1(n14948), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14942) );
  AOI22_X1 U18480 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14941) );
  NAND4_X1 U18481 ( .A1(n14944), .A2(n14943), .A3(n14942), .A4(n14941), .ZN(
        n14945) );
  OR2_X1 U18482 ( .A1(n14946), .A2(n14945), .ZN(n14974) );
  NAND2_X1 U18483 ( .A1(n14975), .A2(n14974), .ZN(n14963) );
  NOR2_X1 U18484 ( .A1(n14962), .A2(n14963), .ZN(n15014) );
  AOI22_X1 U18485 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14952) );
  AOI22_X1 U18486 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14951) );
  AOI22_X1 U18487 ( .A1(n14948), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14950) );
  AOI22_X1 U18488 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14949) );
  NAND4_X1 U18489 ( .A1(n14952), .A2(n14951), .A3(n14950), .A4(n14949), .ZN(
        n14958) );
  AOI22_X1 U18490 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15059), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14956) );
  AOI22_X1 U18491 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14955) );
  AOI22_X1 U18492 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14954) );
  AOI22_X1 U18493 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14953) );
  NAND4_X1 U18494 ( .A1(n14956), .A2(n14955), .A3(n14954), .A4(n14953), .ZN(
        n14957) );
  OR2_X1 U18495 ( .A1(n14958), .A2(n14957), .ZN(n15013) );
  XNOR2_X1 U18496 ( .A(n15014), .B(n15013), .ZN(n14960) );
  AOI22_X1 U18497 ( .A1(n15246), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n14046), .ZN(n14959) );
  OAI21_X1 U18498 ( .B1(n14960), .B2(n15099), .A(n14959), .ZN(n14961) );
  MUX2_X1 U18499 ( .A(n15662), .B(n14961), .S(n15101), .Z(n15340) );
  XOR2_X1 U18500 ( .A(n14963), .B(n14962), .Z(n14964) );
  NAND2_X1 U18501 ( .A1(n14964), .A2(n15067), .ZN(n14968) );
  AOI21_X1 U18502 ( .B1(n15667), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14965) );
  AOI21_X1 U18503 ( .B1(n13958), .B2(P1_EAX_REG_25__SCAN_IN), .A(n14965), .ZN(
        n14967) );
  XNOR2_X1 U18504 ( .A(n14973), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15669) );
  AND2_X1 U18505 ( .A1(n15669), .A2(n14983), .ZN(n14966) );
  AOI21_X1 U18506 ( .B1(n14968), .B2(n14967), .A(n14966), .ZN(n15357) );
  INV_X1 U18507 ( .A(n15357), .ZN(n15010) );
  INV_X1 U18508 ( .A(n14969), .ZN(n14971) );
  INV_X1 U18509 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14970) );
  NAND2_X1 U18510 ( .A1(n14971), .A2(n14970), .ZN(n14972) );
  NAND2_X1 U18511 ( .A1(n14973), .A2(n14972), .ZN(n15674) );
  XNOR2_X1 U18512 ( .A(n14975), .B(n14974), .ZN(n14977) );
  AOI22_X1 U18513 ( .A1(n15246), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n14046), .ZN(n14976) );
  OAI21_X1 U18514 ( .B1(n14977), .B2(n15099), .A(n14976), .ZN(n14978) );
  MUX2_X1 U18515 ( .A(n15674), .B(n14978), .S(n15101), .Z(n15373) );
  INV_X1 U18516 ( .A(n15373), .ZN(n15009) );
  XOR2_X1 U18517 ( .A(n14980), .B(n14979), .Z(n14982) );
  INV_X1 U18518 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15686) );
  OAI22_X1 U18519 ( .A1(n13616), .A2(n13064), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15686), .ZN(n14981) );
  AOI21_X1 U18520 ( .B1(n14982), .B2(n15067), .A(n14981), .ZN(n14984) );
  XNOR2_X1 U18521 ( .A(n15006), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15684) );
  MUX2_X1 U18522 ( .A(n14984), .B(n15684), .S(n14983), .Z(n15386) );
  AOI22_X1 U18523 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14989) );
  AOI22_X1 U18524 ( .A1(n14985), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15081), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14988) );
  AOI22_X1 U18525 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14987) );
  AOI22_X1 U18526 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14986) );
  NAND4_X1 U18527 ( .A1(n14989), .A2(n14988), .A3(n14987), .A4(n14986), .ZN(
        n14998) );
  AOI22_X1 U18528 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14996) );
  AOI22_X1 U18529 ( .A1(n14991), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14990), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14995) );
  AOI22_X1 U18530 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14994) );
  AOI22_X1 U18531 ( .A1(n14992), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14993) );
  NAND4_X1 U18532 ( .A1(n14996), .A2(n14995), .A3(n14994), .A4(n14993), .ZN(
        n14997) );
  NOR2_X1 U18533 ( .A1(n14998), .A2(n14997), .ZN(n15002) );
  OAI21_X1 U18534 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20514), .A(
        n14046), .ZN(n14999) );
  INV_X1 U18535 ( .A(n14999), .ZN(n15000) );
  AOI21_X1 U18536 ( .B1(n13958), .B2(P1_EAX_REG_22__SCAN_IN), .A(n15000), .ZN(
        n15001) );
  OAI21_X1 U18537 ( .B1(n15099), .B2(n15002), .A(n15001), .ZN(n15008) );
  INV_X1 U18538 ( .A(n15003), .ZN(n15004) );
  INV_X1 U18539 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15405) );
  NAND2_X1 U18540 ( .A1(n15004), .A2(n15405), .ZN(n15005) );
  NAND2_X1 U18541 ( .A1(n15006), .A2(n15005), .ZN(n15694) );
  OR2_X1 U18542 ( .A1(n15694), .A2(n15101), .ZN(n15007) );
  NAND2_X1 U18543 ( .A1(n15008), .A2(n15007), .ZN(n15398) );
  OR2_X1 U18544 ( .A1(n15386), .A2(n15398), .ZN(n15370) );
  NOR2_X1 U18545 ( .A1(n15010), .A2(n15354), .ZN(n15339) );
  XNOR2_X1 U18546 ( .A(n15012), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15654) );
  NAND2_X1 U18547 ( .A1(n15014), .A2(n15013), .ZN(n15033) );
  AOI22_X1 U18548 ( .A1(n15015), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15019) );
  AOI22_X1 U18549 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n9708), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15018) );
  AOI22_X1 U18550 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15017) );
  AOI22_X1 U18551 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15016) );
  NAND4_X1 U18552 ( .A1(n15019), .A2(n15018), .A3(n15017), .A4(n15016), .ZN(
        n15025) );
  AOI22_X1 U18553 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n15086), .B1(
        n15071), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15023) );
  AOI22_X1 U18554 ( .A1(n15035), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14992), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15022) );
  AOI22_X1 U18555 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n15081), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U18556 ( .A1(n15083), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15074), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15020) );
  NAND4_X1 U18557 ( .A1(n15023), .A2(n15022), .A3(n15021), .A4(n15020), .ZN(
        n15024) );
  NOR2_X1 U18558 ( .A1(n15025), .A2(n15024), .ZN(n15034) );
  XOR2_X1 U18559 ( .A(n15033), .B(n15034), .Z(n15027) );
  OAI22_X1 U18560 ( .A1(n13616), .A2(n12930), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15652), .ZN(n15026) );
  AOI21_X1 U18561 ( .B1(n15027), .B2(n15067), .A(n15026), .ZN(n15028) );
  MUX2_X1 U18562 ( .A(n15654), .B(n15028), .S(n15101), .Z(n15325) );
  INV_X1 U18563 ( .A(n15029), .ZN(n15031) );
  INV_X1 U18564 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15030) );
  NAND2_X1 U18565 ( .A1(n15031), .A2(n15030), .ZN(n15032) );
  NAND2_X1 U18566 ( .A1(n15050), .A2(n15032), .ZN(n15637) );
  NOR2_X1 U18567 ( .A1(n15034), .A2(n15033), .ZN(n15052) );
  AOI22_X1 U18568 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15059), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15039) );
  AOI22_X1 U18569 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15038) );
  AOI22_X1 U18570 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15037) );
  AOI22_X1 U18571 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15036) );
  NAND4_X1 U18572 ( .A1(n15039), .A2(n15038), .A3(n15037), .A4(n15036), .ZN(
        n15046) );
  AOI22_X1 U18573 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9707), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15044) );
  AOI22_X1 U18574 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15043) );
  AOI22_X1 U18575 ( .A1(n15081), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14930), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15042) );
  AOI22_X1 U18576 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9702), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15041) );
  NAND4_X1 U18577 ( .A1(n15044), .A2(n15043), .A3(n15042), .A4(n15041), .ZN(
        n15045) );
  OR2_X1 U18578 ( .A1(n15046), .A2(n15045), .ZN(n15051) );
  XNOR2_X1 U18579 ( .A(n15052), .B(n15051), .ZN(n15048) );
  AOI22_X1 U18580 ( .A1(n15246), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n14046), .ZN(n15047) );
  OAI21_X1 U18581 ( .B1(n15048), .B2(n15099), .A(n15047), .ZN(n15049) );
  MUX2_X1 U18582 ( .A(n15637), .B(n15049), .S(n15101), .Z(n15311) );
  XNOR2_X1 U18583 ( .A(n15050), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15631) );
  NAND2_X1 U18584 ( .A1(n15052), .A2(n15051), .ZN(n15094) );
  AOI22_X1 U18585 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15076), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U18586 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13700), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15057) );
  AOI22_X1 U18587 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15053), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U18588 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15075), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15055) );
  NAND4_X1 U18589 ( .A1(n15058), .A2(n15057), .A3(n15056), .A4(n15055), .ZN(
        n15065) );
  AOI22_X1 U18590 ( .A1(n15040), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15081), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15063) );
  AOI22_X1 U18591 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15059), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15062) );
  AOI22_X1 U18592 ( .A1(n15035), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15074), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15061) );
  AOI22_X1 U18593 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15060) );
  NAND4_X1 U18594 ( .A1(n15063), .A2(n15062), .A3(n15061), .A4(n15060), .ZN(
        n15064) );
  NOR2_X1 U18595 ( .A1(n15065), .A2(n15064), .ZN(n15095) );
  XOR2_X1 U18596 ( .A(n15094), .B(n15095), .Z(n15068) );
  OAI22_X1 U18597 ( .A1(n13616), .A2(n12943), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15633), .ZN(n15066) );
  AOI21_X1 U18598 ( .B1(n15068), .B2(n15067), .A(n15066), .ZN(n15069) );
  MUX2_X1 U18599 ( .A(n15631), .B(n15069), .S(n15101), .Z(n15300) );
  XNOR2_X1 U18600 ( .A(n15070), .B(n15187), .ZN(n15621) );
  AOI22_X1 U18601 ( .A1(n15071), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15035), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15080) );
  AOI22_X1 U18602 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13700), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15079) );
  AOI22_X1 U18603 ( .A1(n15074), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15073), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15078) );
  AOI22_X1 U18604 ( .A1(n15076), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9702), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15077) );
  NAND4_X1 U18605 ( .A1(n15080), .A2(n15079), .A3(n15078), .A4(n15077), .ZN(
        n15093) );
  AOI22_X1 U18606 ( .A1(n9708), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15081), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15091) );
  AOI22_X1 U18607 ( .A1(n15084), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15083), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15090) );
  AOI22_X1 U18608 ( .A1(n15086), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15085), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15089) );
  AOI22_X1 U18609 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15087), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15088) );
  NAND4_X1 U18610 ( .A1(n15091), .A2(n15090), .A3(n15089), .A4(n15088), .ZN(
        n15092) );
  NOR2_X1 U18611 ( .A1(n15093), .A2(n15092), .ZN(n15097) );
  NOR2_X1 U18612 ( .A1(n15095), .A2(n15094), .ZN(n15096) );
  XOR2_X1 U18613 ( .A(n15097), .B(n15096), .Z(n15100) );
  AOI22_X1 U18614 ( .A1(n15246), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n14046), .ZN(n15098) );
  OAI21_X1 U18615 ( .B1(n15100), .B2(n15099), .A(n15098), .ZN(n15102) );
  MUX2_X1 U18616 ( .A(n15621), .B(n15102), .S(n15101), .Z(n15104) );
  NAND2_X1 U18617 ( .A1(n15103), .A2(n15104), .ZN(n15249) );
  NOR2_X1 U18618 ( .A1(n15108), .A2(n15105), .ZN(n15106) );
  NAND2_X1 U18619 ( .A1(n15606), .A2(n15106), .ZN(n15594) );
  AOI22_X1 U18620 ( .A1(n15587), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n15610), .ZN(n15112) );
  NOR3_X4 U18621 ( .A1(n15610), .A2(n15533), .A3(n15107), .ZN(n15595) );
  NOR3_X1 U18622 ( .A1(n15610), .A2(n15109), .A3(n15108), .ZN(n15110) );
  AOI22_X1 U18623 ( .A1(n15595), .A2(n15605), .B1(n15600), .B2(DATAI_30_), 
        .ZN(n15111) );
  OAI211_X1 U18624 ( .C1(n15624), .C2(n15614), .A(n15112), .B(n15111), .ZN(
        P1_U2874) );
  INV_X1 U18625 ( .A(n15165), .ZN(n15124) );
  INV_X1 U18626 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15530) );
  NAND2_X1 U18627 ( .A1(n15124), .A2(n15530), .ZN(n15116) );
  INV_X1 U18628 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16813) );
  NAND2_X1 U18629 ( .A1(n15149), .A2(n16813), .ZN(n15114) );
  NAND2_X1 U18630 ( .A1(n15162), .A2(n15530), .ZN(n15113) );
  NAND3_X1 U18631 ( .A1(n15114), .A2(n15129), .A3(n15113), .ZN(n15115) );
  AND2_X1 U18632 ( .A1(n15116), .A2(n15115), .ZN(n15468) );
  MUX2_X1 U18633 ( .A(n15159), .B(n15129), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n15117) );
  OAI21_X1 U18634 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15218), .A(
        n15117), .ZN(n15527) );
  OR2_X1 U18635 ( .A1(n15165), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n15121) );
  INV_X1 U18636 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16805) );
  NAND2_X1 U18637 ( .A1(n15149), .A2(n16805), .ZN(n15119) );
  INV_X1 U18638 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n16707) );
  NAND2_X1 U18639 ( .A1(n15162), .A2(n16707), .ZN(n15118) );
  NAND3_X1 U18640 ( .A1(n15119), .A2(n15129), .A3(n15118), .ZN(n15120) );
  NAND2_X1 U18641 ( .A1(n15121), .A2(n15120), .ZN(n15517) );
  NAND2_X1 U18642 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15122) );
  OAI211_X1 U18643 ( .C1(n15287), .C2(P1_EBX_REG_16__SCAN_IN), .A(n15149), .B(
        n15122), .ZN(n15123) );
  OAI21_X1 U18644 ( .B1(n15159), .B2(P1_EBX_REG_16__SCAN_IN), .A(n15123), .ZN(
        n15883) );
  INV_X1 U18645 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15510) );
  NAND2_X1 U18646 ( .A1(n15124), .A2(n15510), .ZN(n15128) );
  INV_X1 U18647 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16792) );
  NAND2_X1 U18648 ( .A1(n15149), .A2(n16792), .ZN(n15126) );
  NAND2_X1 U18649 ( .A1(n15162), .A2(n15510), .ZN(n15125) );
  NAND3_X1 U18650 ( .A1(n15126), .A2(n15129), .A3(n15125), .ZN(n15127) );
  AND2_X1 U18651 ( .A1(n15128), .A2(n15127), .ZN(n15507) );
  MUX2_X1 U18652 ( .A(n15159), .B(n15129), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n15131) );
  OR2_X1 U18653 ( .A1(n15218), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15130) );
  NAND2_X1 U18654 ( .A1(n15131), .A2(n15130), .ZN(n15458) );
  INV_X1 U18655 ( .A(n15458), .ZN(n15132) );
  INV_X1 U18656 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16786) );
  NAND2_X1 U18657 ( .A1(n15149), .A2(n16786), .ZN(n15133) );
  OAI211_X1 U18658 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n15287), .A(n15133), .B(
        n15129), .ZN(n15135) );
  OR2_X1 U18659 ( .A1(n15165), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n15134) );
  NAND2_X1 U18660 ( .A1(n15135), .A2(n15134), .ZN(n15444) );
  NAND2_X1 U18661 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15136) );
  OAI211_X1 U18662 ( .C1(P1_EBX_REG_20__SCAN_IN), .C2(n15287), .A(n15149), .B(
        n15136), .ZN(n15137) );
  OAI21_X1 U18663 ( .B1(n15159), .B2(P1_EBX_REG_20__SCAN_IN), .A(n15137), .ZN(
        n15430) );
  OR2_X1 U18664 ( .A1(n15165), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n15140) );
  INV_X1 U18665 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15700) );
  NAND2_X1 U18666 ( .A1(n15149), .A2(n15700), .ZN(n15138) );
  OAI211_X1 U18667 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n15287), .A(n15138), .B(
        n15129), .ZN(n15139) );
  AND2_X1 U18668 ( .A1(n15140), .A2(n15139), .ZN(n15416) );
  NAND2_X1 U18669 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15141) );
  OAI211_X1 U18670 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n15287), .A(n15149), .B(
        n15141), .ZN(n15142) );
  OAI21_X1 U18671 ( .B1(n15159), .B2(P1_EBX_REG_22__SCAN_IN), .A(n15142), .ZN(
        n15400) );
  INV_X1 U18672 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15858) );
  NAND2_X1 U18673 ( .A1(n15149), .A2(n15858), .ZN(n15143) );
  OAI211_X1 U18674 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n15287), .A(n15143), .B(
        n15129), .ZN(n15145) );
  OR2_X1 U18675 ( .A1(n15165), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n15144) );
  NAND2_X1 U18676 ( .A1(n15145), .A2(n15144), .ZN(n15387) );
  INV_X1 U18677 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15496) );
  NAND2_X1 U18678 ( .A1(n15146), .A2(n15496), .ZN(n15151) );
  NAND2_X1 U18679 ( .A1(n15147), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15148) );
  OAI211_X1 U18680 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n15287), .A(n15149), .B(
        n15148), .ZN(n15150) );
  AND2_X1 U18681 ( .A1(n15151), .A2(n15150), .ZN(n15375) );
  INV_X1 U18682 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21321) );
  NAND2_X1 U18683 ( .A1(n15149), .A2(n21321), .ZN(n15152) );
  OAI211_X1 U18684 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n15287), .A(n15152), .B(
        n15129), .ZN(n15154) );
  OR2_X1 U18685 ( .A1(n15165), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n15153) );
  NAND2_X1 U18686 ( .A1(n15154), .A2(n15153), .ZN(n15359) );
  MUX2_X1 U18687 ( .A(n15159), .B(n15129), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n15155) );
  OAI21_X1 U18688 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15218), .A(
        n15155), .ZN(n15343) );
  OR2_X1 U18689 ( .A1(n15165), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n15158) );
  INV_X1 U18690 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15648) );
  NAND2_X1 U18691 ( .A1(n15149), .A2(n15648), .ZN(n15156) );
  OAI211_X1 U18692 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n15287), .A(n15156), .B(
        n15129), .ZN(n15157) );
  AND2_X1 U18693 ( .A1(n15158), .A2(n15157), .ZN(n15327) );
  MUX2_X1 U18694 ( .A(n15159), .B(n15129), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n15161) );
  OR2_X1 U18695 ( .A1(n15218), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15160) );
  AND2_X1 U18696 ( .A1(n15161), .A2(n15160), .ZN(n15312) );
  OR2_X1 U18697 ( .A1(n15218), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15164) );
  INV_X1 U18698 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15487) );
  NAND2_X1 U18699 ( .A1(n15162), .A2(n15487), .ZN(n15163) );
  NAND2_X1 U18700 ( .A1(n15164), .A2(n15163), .ZN(n15167) );
  OAI22_X1 U18701 ( .A1(n15167), .A2(n12765), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n15165), .ZN(n15296) );
  NAND2_X1 U18702 ( .A1(n15298), .A2(n12765), .ZN(n15168) );
  INV_X1 U18703 ( .A(n15314), .ZN(n15166) );
  AOI22_X1 U18704 ( .A1(n15168), .A2(n15167), .B1(n15166), .B2(n15129), .ZN(
        n15169) );
  AOI22_X1 U18705 ( .A1(n15218), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15287), .ZN(n15219) );
  XNOR2_X1 U18706 ( .A(n15169), .B(n15219), .ZN(n15796) );
  AOI22_X1 U18707 ( .A1(n15796), .A2(n21040), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n21041), .ZN(n15170) );
  OAI21_X1 U18708 ( .B1(n15624), .B2(n15513), .A(n15170), .ZN(P1_U2842) );
  INV_X1 U18709 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20972) );
  INV_X1 U18710 ( .A(n15171), .ZN(n15467) );
  NOR3_X1 U18711 ( .A1(n15173), .A2(n15172), .A3(n15467), .ZN(n15174) );
  NAND3_X1 U18712 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n15174), .ZN(n16706) );
  NOR2_X1 U18713 ( .A1(n20972), .A2(n16706), .ZN(n15179) );
  NAND2_X1 U18714 ( .A1(n20596), .A2(n15179), .ZN(n16698) );
  NOR2_X1 U18715 ( .A1(n15748), .A2(n16698), .ZN(n16691) );
  NAND2_X1 U18716 ( .A1(n16691), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U18717 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15175) );
  NOR2_X1 U18718 ( .A1(n15459), .A2(n15175), .ZN(n15437) );
  NAND2_X1 U18719 ( .A1(n15437), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15412) );
  AND2_X1 U18720 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15391) );
  NAND2_X1 U18721 ( .A1(n15391), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15178) );
  AND2_X1 U18722 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n15350) );
  AND2_X1 U18723 ( .A1(n15350), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15330) );
  AND2_X1 U18724 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n15176) );
  NAND2_X1 U18725 ( .A1(n15330), .A2(n15176), .ZN(n15177) );
  NOR2_X1 U18726 ( .A1(n15384), .A2(n15177), .ZN(n15307) );
  AOI21_X1 U18727 ( .B1(n15307), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n15190) );
  INV_X1 U18728 ( .A(n15177), .ZN(n15184) );
  INV_X1 U18729 ( .A(n15178), .ZN(n15183) );
  INV_X1 U18730 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15182) );
  INV_X1 U18731 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15181) );
  AND4_X1 U18732 ( .A1(n15180), .A2(P1_REIP_REG_17__SCAN_IN), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(n15179), .ZN(n15460) );
  NAND2_X1 U18733 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15460), .ZN(n15448) );
  NOR3_X1 U18734 ( .A1(n15182), .A2(n15181), .A3(n15448), .ZN(n15403) );
  AND2_X1 U18735 ( .A1(n15183), .A2(n15403), .ZN(n15362) );
  AND2_X1 U18736 ( .A1(n15184), .A2(n15362), .ZN(n15301) );
  AND2_X1 U18737 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n15185) );
  NAND2_X1 U18738 ( .A1(n15301), .A2(n15185), .ZN(n15186) );
  NAND2_X1 U18739 ( .A1(n16694), .A2(n15186), .ZN(n15291) );
  OAI22_X1 U18740 ( .A1(n15187), .A2(n20581), .B1(n20583), .B2(n15621), .ZN(
        n15188) );
  AOI21_X1 U18741 ( .B1(P1_EBX_REG_30__SCAN_IN), .B2(n20602), .A(n15188), .ZN(
        n15189) );
  OAI21_X1 U18742 ( .B1(n15190), .B2(n15291), .A(n15189), .ZN(n15191) );
  AOI21_X1 U18743 ( .B1(n15796), .B2(n20595), .A(n15191), .ZN(n15192) );
  OAI21_X1 U18744 ( .B1(n15624), .B2(n15476), .A(n15192), .ZN(P1_U2810) );
  NAND2_X1 U18745 ( .A1(n9714), .A2(n16840), .ZN(n15195) );
  NAND2_X1 U18746 ( .A1(n15782), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15890) );
  NAND2_X1 U18747 ( .A1(n15193), .A2(n16813), .ZN(n15196) );
  NAND2_X1 U18748 ( .A1(n15890), .A2(n15196), .ZN(n15770) );
  INV_X1 U18749 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15919) );
  NAND2_X1 U18750 ( .A1(n9713), .A2(n15919), .ZN(n15769) );
  NAND2_X1 U18751 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15197) );
  NAND2_X1 U18752 ( .A1(n9713), .A2(n15197), .ZN(n15767) );
  NAND2_X1 U18753 ( .A1(n15769), .A2(n15767), .ZN(n15198) );
  NOR2_X1 U18754 ( .A1(n15770), .A2(n15198), .ZN(n15892) );
  INV_X1 U18755 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21244) );
  NAND2_X1 U18756 ( .A1(n9714), .A2(n21244), .ZN(n15199) );
  OAI21_X1 U18757 ( .B1(n15209), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15756), .ZN(n15200) );
  INV_X1 U18758 ( .A(n15200), .ZN(n15202) );
  XNOR2_X1 U18759 ( .A(n9714), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15746) );
  NAND2_X1 U18760 ( .A1(n9714), .A2(n16805), .ZN(n15754) );
  NAND2_X1 U18761 ( .A1(n15746), .A2(n15754), .ZN(n15744) );
  NAND2_X1 U18762 ( .A1(n15209), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15203) );
  AND2_X1 U18763 ( .A1(n15890), .A2(n15203), .ZN(n15733) );
  INV_X1 U18764 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15781) );
  NAND2_X1 U18765 ( .A1(n16750), .A2(n15781), .ZN(n15732) );
  OAI21_X1 U18766 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15732), .A(
        n15209), .ZN(n15204) );
  NAND2_X1 U18767 ( .A1(n15733), .A2(n15204), .ZN(n15757) );
  NOR2_X1 U18768 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15880) );
  AND2_X1 U18769 ( .A1(n15880), .A2(n16792), .ZN(n15205) );
  NOR2_X1 U18770 ( .A1(n9714), .A2(n15205), .ZN(n15206) );
  NOR2_X1 U18771 ( .A1(n15757), .A2(n15206), .ZN(n15207) );
  XNOR2_X1 U18772 ( .A(n9714), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15723) );
  NAND2_X1 U18773 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16672) );
  INV_X1 U18774 ( .A(n16672), .ZN(n15208) );
  AND2_X2 U18775 ( .A1(n15690), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15213) );
  INV_X1 U18776 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21206) );
  INV_X1 U18777 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15210) );
  NAND2_X1 U18778 ( .A1(n15700), .A2(n15210), .ZN(n15211) );
  INV_X1 U18779 ( .A(n15691), .ZN(n15212) );
  INV_X1 U18780 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15676) );
  NAND3_X1 U18781 ( .A1(n21321), .A2(n15858), .A3(n15676), .ZN(n15639) );
  NOR3_X1 U18782 ( .A1(n15647), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15618) );
  AND2_X1 U18783 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15670) );
  NAND2_X1 U18784 ( .A1(n15670), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15826) );
  AND2_X1 U18785 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15232) );
  OAI21_X1 U18786 ( .B1(n15618), .B2(n9714), .A(n15215), .ZN(n15627) );
  INV_X1 U18787 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21241) );
  NAND2_X1 U18788 ( .A1(n15209), .A2(n21241), .ZN(n15629) );
  NAND2_X1 U18789 ( .A1(n9714), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15628) );
  AOI22_X1 U18790 ( .A1(n15218), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n15287), .ZN(n15220) );
  INV_X1 U18791 ( .A(n15670), .ZN(n15830) );
  INV_X1 U18792 ( .A(n15871), .ZN(n15870) );
  NAND2_X1 U18793 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16793) );
  NOR2_X1 U18794 ( .A1(n16792), .A2(n16793), .ZN(n15873) );
  NAND2_X1 U18795 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15873), .ZN(
        n15238) );
  NOR2_X1 U18796 ( .A1(n21244), .A2(n15238), .ZN(n15226) );
  NAND3_X1 U18797 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16836) );
  NOR3_X1 U18798 ( .A1(n15781), .A2(n16840), .A3(n16836), .ZN(n15911) );
  NAND2_X1 U18799 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15911), .ZN(
        n15916) );
  NOR2_X1 U18800 ( .A1(n15919), .A2(n15916), .ZN(n15235) );
  NAND2_X1 U18801 ( .A1(n15235), .A2(n16823), .ZN(n15862) );
  NOR2_X1 U18802 ( .A1(n16813), .A2(n15862), .ZN(n15900) );
  NOR2_X1 U18803 ( .A1(n15222), .A2(n15221), .ZN(n15910) );
  AND2_X1 U18804 ( .A1(n15235), .A2(n15910), .ZN(n15865) );
  NAND2_X1 U18805 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15865), .ZN(
        n15868) );
  INV_X1 U18806 ( .A(n15226), .ZN(n15223) );
  AOI221_X1 U18807 ( .B1(n15868), .B2(n15224), .C1(n15223), .C2(n15224), .A(
        n20658), .ZN(n15225) );
  OAI221_X1 U18808 ( .B1(n15863), .B2(n15226), .C1(n15863), .C2(n15900), .A(
        n15225), .ZN(n16784) );
  INV_X1 U18809 ( .A(n16784), .ZN(n15227) );
  NAND2_X1 U18810 ( .A1(n15227), .A2(n15208), .ZN(n15229) );
  NAND2_X1 U18811 ( .A1(n15871), .A2(n15228), .ZN(n16824) );
  AND2_X1 U18812 ( .A1(n15229), .A2(n16824), .ZN(n16776) );
  NAND2_X1 U18813 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16775) );
  INV_X1 U18814 ( .A(n16775), .ZN(n15230) );
  NOR2_X1 U18815 ( .A1(n15871), .A2(n15230), .ZN(n15231) );
  NOR2_X1 U18816 ( .A1(n16776), .A2(n15231), .ZN(n15856) );
  OAI21_X1 U18817 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15863), .A(
        n15856), .ZN(n15848) );
  AOI21_X1 U18818 ( .B1(n15830), .B2(n15870), .A(n15848), .ZN(n15841) );
  NAND3_X1 U18819 ( .A1(n15841), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15818) );
  INV_X1 U18820 ( .A(n15232), .ZN(n15240) );
  NAND2_X1 U18821 ( .A1(n15856), .A2(n15871), .ZN(n15817) );
  OAI21_X1 U18822 ( .B1(n15818), .B2(n15240), .A(n15817), .ZN(n15801) );
  OAI211_X1 U18823 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15871), .A(
        n15801), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15791) );
  NAND3_X1 U18824 ( .A1(n15791), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15817), .ZN(n15242) );
  NAND2_X1 U18825 ( .A1(n13116), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n15251) );
  NAND2_X1 U18826 ( .A1(n15234), .A2(n15233), .ZN(n15915) );
  INV_X1 U18827 ( .A(n15235), .ZN(n15236) );
  OAI22_X1 U18828 ( .A1(n15915), .A2(n15236), .B1(n15862), .B2(n15863), .ZN(
        n15869) );
  AND2_X1 U18829 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15237) );
  NAND2_X1 U18830 ( .A1(n15869), .A2(n15237), .ZN(n16806) );
  NOR2_X1 U18831 ( .A1(n16806), .A2(n15238), .ZN(n16787) );
  NAND2_X1 U18832 ( .A1(n16787), .A2(n15208), .ZN(n16783) );
  INV_X1 U18833 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15239) );
  NOR2_X1 U18834 ( .A1(n15821), .A2(n15240), .ZN(n15804) );
  NAND4_X1 U18835 ( .A1(n15804), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n15217), .ZN(n15241) );
  NAND3_X1 U18836 ( .A1(n15242), .A2(n15251), .A3(n15241), .ZN(n15243) );
  AOI21_X1 U18837 ( .B1(n15484), .B2(n16857), .A(n15243), .ZN(n15244) );
  AOI22_X1 U18838 ( .A1(n15246), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n15245), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15247) );
  INV_X1 U18839 ( .A(n15247), .ZN(n15248) );
  NAND2_X1 U18840 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15250) );
  OAI211_X1 U18841 ( .C1(n16769), .C2(n15252), .A(n15251), .B(n15250), .ZN(
        n15253) );
  OAI21_X1 U18842 ( .B1(n15255), .B2(n20516), .A(n15254), .ZN(P1_U2968) );
  INV_X1 U18843 ( .A(n15256), .ZN(n15259) );
  NOR2_X1 U18844 ( .A1(n17039), .A2(n15257), .ZN(n15258) );
  AOI211_X1 U18845 ( .C1(n15260), .C2(n19828), .A(n15259), .B(n15258), .ZN(
        n15263) );
  OAI21_X1 U18846 ( .B1(n19837), .B2(n15261), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15262) );
  OAI211_X1 U18847 ( .C1(n16307), .C2(n15264), .A(n15263), .B(n15262), .ZN(
        P2_U3014) );
  NOR2_X1 U18848 ( .A1(n9693), .A2(n19716), .ZN(n15266) );
  AOI21_X1 U18849 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19716), .A(n15266), .ZN(
        n15267) );
  OAI21_X1 U18850 ( .B1(n15268), .B2(n19713), .A(n15267), .ZN(P2_U2857) );
  NAND2_X1 U18851 ( .A1(n13540), .A2(n20514), .ZN(n15269) );
  AOI211_X1 U18852 ( .C1(n15270), .C2(n15269), .A(n20807), .B(n20663), .ZN(
        n15271) );
  AOI21_X1 U18853 ( .B1(n20663), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15271), .ZN(n15272) );
  OAI21_X1 U18854 ( .B1(n13840), .B2(n15273), .A(n15272), .ZN(P1_U3477) );
  INV_X1 U18855 ( .A(n15274), .ZN(n15276) );
  AND3_X1 U18856 ( .A1(n15276), .A2(n12767), .A3(n15275), .ZN(n15277) );
  OR2_X1 U18857 ( .A1(n16614), .A2(n15277), .ZN(n15280) );
  NAND2_X1 U18858 ( .A1(n16614), .A2(n15278), .ZN(n15279) );
  OAI211_X1 U18859 ( .C1(n15281), .C2(n12766), .A(n15280), .B(n15279), .ZN(
        n16629) );
  OR2_X1 U18860 ( .A1(n16614), .A2(n12779), .ZN(n15285) );
  INV_X1 U18861 ( .A(n15282), .ZN(n15283) );
  NAND2_X1 U18862 ( .A1(n15283), .A2(n12767), .ZN(n15284) );
  NAND2_X1 U18863 ( .A1(n15285), .A2(n15284), .ZN(n20509) );
  NAND3_X1 U18864 ( .A1(n15287), .A2(n15286), .A3(n16666), .ZN(n15288) );
  AND2_X1 U18865 ( .A1(n15288), .A2(n21028), .ZN(n21030) );
  NOR2_X1 U18866 ( .A1(n20509), .A2(n21030), .ZN(n16632) );
  OR2_X1 U18867 ( .A1(n16632), .A2(n20508), .ZN(n20515) );
  MUX2_X1 U18868 ( .A(n16629), .B(P1_MORE_REG_SCAN_IN), .S(n20515), .Z(
        P1_U3484) );
  INV_X1 U18869 ( .A(n15534), .ZN(n15295) );
  INV_X1 U18870 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n15292) );
  NAND4_X1 U18871 ( .A1(n15307), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_30__SCAN_IN), .A4(n15292), .ZN(n15290) );
  AOI22_X1 U18872 ( .A1(n20602), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20593), .ZN(n15289) );
  OAI211_X1 U18873 ( .C1(n15292), .C2(n15291), .A(n15290), .B(n15289), .ZN(
        n15293) );
  OAI21_X1 U18874 ( .B1(n15295), .B2(n15476), .A(n15294), .ZN(P1_U2809) );
  OR2_X1 U18875 ( .A1(n15314), .A2(n15296), .ZN(n15297) );
  NAND2_X1 U18876 ( .A1(n15298), .A2(n15297), .ZN(n15800) );
  NAND2_X1 U18877 ( .A1(n15635), .A2(n20554), .ZN(n15309) );
  INV_X1 U18878 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n15306) );
  INV_X1 U18879 ( .A(n15301), .ZN(n15302) );
  NAND2_X1 U18880 ( .A1(n16694), .A2(n15302), .ZN(n15315) );
  AOI22_X1 U18881 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20593), .B1(
        n20604), .B2(n15631), .ZN(n15304) );
  NAND2_X1 U18882 ( .A1(n20602), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n15303) );
  OAI211_X1 U18883 ( .C1(n15315), .C2(n15306), .A(n15304), .B(n15303), .ZN(
        n15305) );
  AOI21_X1 U18884 ( .B1(n15307), .B2(n15306), .A(n15305), .ZN(n15308) );
  OAI211_X1 U18885 ( .C1(n20580), .C2(n15800), .A(n15309), .B(n15308), .ZN(
        P1_U2811) );
  OAI21_X1 U18886 ( .B1(n15310), .B2(n15311), .A(n15299), .ZN(n15646) );
  NOR2_X1 U18887 ( .A1(n15326), .A2(n15312), .ZN(n15313) );
  OR2_X1 U18888 ( .A1(n15314), .A2(n15313), .ZN(n15488) );
  INV_X1 U18889 ( .A(n15488), .ZN(n15808) );
  INV_X1 U18890 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21319) );
  NAND3_X1 U18891 ( .A1(n15330), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n21319), 
        .ZN(n15321) );
  INV_X1 U18892 ( .A(n15315), .ZN(n15319) );
  INV_X1 U18893 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15489) );
  INV_X1 U18894 ( .A(n15637), .ZN(n15316) );
  AOI22_X1 U18895 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20593), .B1(
        n20604), .B2(n15316), .ZN(n15317) );
  OAI21_X1 U18896 ( .B1(n20592), .B2(n15489), .A(n15317), .ZN(n15318) );
  AOI21_X1 U18897 ( .B1(n15319), .B2(P1_REIP_REG_28__SCAN_IN), .A(n15318), 
        .ZN(n15320) );
  OAI21_X1 U18898 ( .B1(n15384), .B2(n15321), .A(n15320), .ZN(n15322) );
  AOI21_X1 U18899 ( .B1(n15808), .B2(n20595), .A(n15322), .ZN(n15323) );
  OAI21_X1 U18900 ( .B1(n15646), .B2(n15476), .A(n15323), .ZN(P1_U2812) );
  INV_X1 U18901 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15651) );
  NAND2_X1 U18902 ( .A1(n15330), .A2(n15651), .ZN(n15337) );
  AOI21_X1 U18903 ( .B1(n15325), .B2(n15324), .A(n15310), .ZN(n15650) );
  NAND2_X1 U18904 ( .A1(n15650), .A2(n20554), .ZN(n15336) );
  INV_X1 U18905 ( .A(n15326), .ZN(n15329) );
  NAND2_X1 U18906 ( .A1(n15341), .A2(n15327), .ZN(n15328) );
  NAND2_X1 U18907 ( .A1(n15329), .A2(n15328), .ZN(n15490) );
  INV_X1 U18908 ( .A(n15490), .ZN(n15816) );
  NAND2_X1 U18909 ( .A1(n15362), .A2(n15330), .ZN(n15331) );
  NAND2_X1 U18910 ( .A1(n16694), .A2(n15331), .ZN(n15347) );
  AOI22_X1 U18911 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20593), .B1(
        n20604), .B2(n15654), .ZN(n15333) );
  NAND2_X1 U18912 ( .A1(n20602), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n15332) );
  OAI211_X1 U18913 ( .C1(n15347), .C2(n15651), .A(n15333), .B(n15332), .ZN(
        n15334) );
  AOI21_X1 U18914 ( .B1(n15816), .B2(n20595), .A(n15334), .ZN(n15335) );
  OAI211_X1 U18915 ( .C1(n15384), .C2(n15337), .A(n15336), .B(n15335), .ZN(
        P1_U2813) );
  AND2_X1 U18916 ( .A1(n15338), .A2(n15339), .ZN(n15355) );
  OAI21_X1 U18917 ( .B1(n15355), .B2(n15340), .A(n15324), .ZN(n15660) );
  INV_X1 U18918 ( .A(n15341), .ZN(n15342) );
  AOI21_X1 U18919 ( .B1(n15343), .B2(n15361), .A(n15342), .ZN(n15829) );
  INV_X1 U18920 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15349) );
  OAI22_X1 U18921 ( .A1(n15344), .A2(n20581), .B1(n20583), .B2(n15662), .ZN(
        n15345) );
  AOI21_X1 U18922 ( .B1(n20602), .B2(P1_EBX_REG_26__SCAN_IN), .A(n15345), .ZN(
        n15346) );
  OAI21_X1 U18923 ( .B1(n15349), .B2(n15347), .A(n15346), .ZN(n15348) );
  AOI21_X1 U18924 ( .B1(n15829), .B2(n20595), .A(n15348), .ZN(n15353) );
  INV_X1 U18925 ( .A(n15384), .ZN(n15351) );
  NAND3_X1 U18926 ( .A1(n15351), .A2(n15350), .A3(n15349), .ZN(n15352) );
  OAI211_X1 U18927 ( .C1(n15660), .C2(n15476), .A(n15353), .B(n15352), .ZN(
        P1_U2814) );
  XNOR2_X1 U18928 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n15369) );
  INV_X2 U18929 ( .A(n15338), .ZN(n15414) );
  NOR2_X1 U18930 ( .A1(n15414), .A2(n15354), .ZN(n15371) );
  INV_X1 U18931 ( .A(n15355), .ZN(n15356) );
  OAI21_X1 U18932 ( .B1(n15357), .B2(n15371), .A(n15356), .ZN(n15673) );
  INV_X1 U18933 ( .A(n15673), .ZN(n15358) );
  NAND2_X1 U18934 ( .A1(n15358), .A2(n20554), .ZN(n15368) );
  OR2_X1 U18935 ( .A1(n15377), .A2(n15359), .ZN(n15360) );
  NAND2_X1 U18936 ( .A1(n15361), .A2(n15360), .ZN(n15493) );
  INV_X1 U18937 ( .A(n15493), .ZN(n15838) );
  INV_X1 U18938 ( .A(n15362), .ZN(n15363) );
  NAND2_X1 U18939 ( .A1(n16694), .A2(n15363), .ZN(n15392) );
  INV_X1 U18940 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15666) );
  AOI22_X1 U18941 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20593), .B1(
        n20604), .B2(n15669), .ZN(n15365) );
  NAND2_X1 U18942 ( .A1(n20602), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n15364) );
  OAI211_X1 U18943 ( .C1(n15392), .C2(n15666), .A(n15365), .B(n15364), .ZN(
        n15366) );
  AOI21_X1 U18944 ( .B1(n15838), .B2(n20595), .A(n15366), .ZN(n15367) );
  OAI211_X1 U18945 ( .C1(n15384), .C2(n15369), .A(n15368), .B(n15367), .ZN(
        P1_U2815) );
  NOR2_X1 U18946 ( .A1(n15414), .A2(n15370), .ZN(n15385) );
  INV_X1 U18947 ( .A(n15371), .ZN(n15372) );
  INV_X1 U18948 ( .A(n15681), .ZN(n15374) );
  NAND2_X1 U18949 ( .A1(n15374), .A2(n20554), .ZN(n15383) );
  NOR2_X1 U18950 ( .A1(n15389), .A2(n15375), .ZN(n15376) );
  OR2_X1 U18951 ( .A1(n15377), .A2(n15376), .ZN(n15495) );
  INV_X1 U18952 ( .A(n15495), .ZN(n15845) );
  INV_X1 U18953 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20985) );
  INV_X1 U18954 ( .A(n15674), .ZN(n15378) );
  AOI22_X1 U18955 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20593), .B1(
        n20604), .B2(n15378), .ZN(n15380) );
  NAND2_X1 U18956 ( .A1(n20602), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n15379) );
  OAI211_X1 U18957 ( .C1(n15392), .C2(n20985), .A(n15380), .B(n15379), .ZN(
        n15381) );
  AOI21_X1 U18958 ( .B1(n15845), .B2(n20595), .A(n15381), .ZN(n15382) );
  OAI211_X1 U18959 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n15384), .A(n15383), 
        .B(n15382), .ZN(P1_U2816) );
  INV_X1 U18960 ( .A(n15688), .ZN(n15563) );
  NOR2_X1 U18961 ( .A1(n15402), .A2(n15387), .ZN(n15388) );
  OR2_X1 U18962 ( .A1(n15389), .A2(n15388), .ZN(n15497) );
  INV_X1 U18963 ( .A(n15497), .ZN(n15853) );
  INV_X1 U18964 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15498) );
  AOI22_X1 U18965 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20593), .B1(
        n20604), .B2(n15684), .ZN(n15390) );
  OAI21_X1 U18966 ( .B1(n20592), .B2(n15498), .A(n15390), .ZN(n15395) );
  INV_X1 U18967 ( .A(n15412), .ZN(n15425) );
  AOI21_X1 U18968 ( .B1(n15425), .B2(n15391), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n15393) );
  NOR2_X1 U18969 ( .A1(n15393), .A2(n15392), .ZN(n15394) );
  AOI211_X1 U18970 ( .C1(n15853), .C2(n20595), .A(n15395), .B(n15394), .ZN(
        n15396) );
  OAI21_X1 U18971 ( .B1(n15563), .B2(n15476), .A(n15396), .ZN(P1_U2817) );
  XNOR2_X1 U18972 ( .A(P1_REIP_REG_21__SCAN_IN), .B(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15411) );
  NAND2_X1 U18973 ( .A1(n15414), .A2(n15398), .ZN(n15399) );
  INV_X1 U18974 ( .A(n15569), .ZN(n15696) );
  NAND2_X1 U18975 ( .A1(n15696), .A2(n20554), .ZN(n15410) );
  AND2_X1 U18976 ( .A1(n15418), .A2(n15400), .ZN(n15401) );
  NOR2_X1 U18977 ( .A1(n15402), .A2(n15401), .ZN(n16778) );
  INV_X1 U18978 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20982) );
  INV_X1 U18979 ( .A(n15403), .ZN(n15404) );
  NAND2_X1 U18980 ( .A1(n16694), .A2(n15404), .ZN(n15435) );
  OAI22_X1 U18981 ( .A1(n15405), .A2(n20581), .B1(n20583), .B2(n15694), .ZN(
        n15406) );
  AOI21_X1 U18982 ( .B1(n20602), .B2(P1_EBX_REG_22__SCAN_IN), .A(n15406), .ZN(
        n15407) );
  OAI21_X1 U18983 ( .B1(n20982), .B2(n15435), .A(n15407), .ZN(n15408) );
  AOI21_X1 U18984 ( .B1(n16778), .B2(n20595), .A(n15408), .ZN(n15409) );
  OAI211_X1 U18985 ( .C1(n15412), .C2(n15411), .A(n15410), .B(n15409), .ZN(
        P1_U2818) );
  OAI21_X1 U18986 ( .B1(n15413), .B2(n15415), .A(n15414), .ZN(n15702) );
  INV_X1 U18987 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15424) );
  NAND2_X1 U18988 ( .A1(n15432), .A2(n15416), .ZN(n15417) );
  NAND2_X1 U18989 ( .A1(n15418), .A2(n15417), .ZN(n16657) );
  OAI22_X1 U18990 ( .A1(n15419), .A2(n20581), .B1(n20583), .B2(n15704), .ZN(
        n15421) );
  NOR2_X1 U18991 ( .A1(n15435), .A2(n15424), .ZN(n15420) );
  AOI211_X1 U18992 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n20602), .A(n15421), .B(
        n15420), .ZN(n15422) );
  OAI21_X1 U18993 ( .B1(n16657), .B2(n20580), .A(n15422), .ZN(n15423) );
  AOI21_X1 U18994 ( .B1(n15425), .B2(n15424), .A(n15423), .ZN(n15426) );
  OAI21_X1 U18995 ( .B1(n15702), .B2(n15476), .A(n15426), .ZN(P1_U2819) );
  AOI21_X1 U18996 ( .B1(n10329), .B2(n15427), .A(n15413), .ZN(n15714) );
  INV_X1 U18997 ( .A(n15714), .ZN(n15578) );
  OAI22_X1 U18998 ( .A1(n15428), .A2(n20581), .B1(n20583), .B2(n15712), .ZN(
        n15434) );
  NAND2_X1 U18999 ( .A1(n15429), .A2(n15430), .ZN(n15431) );
  NAND2_X1 U19000 ( .A1(n15432), .A2(n15431), .ZN(n16669) );
  NOR2_X1 U19001 ( .A1(n16669), .A2(n20580), .ZN(n15433) );
  AOI211_X1 U19002 ( .C1(P1_EBX_REG_20__SCAN_IN), .C2(n20602), .A(n15434), .B(
        n15433), .ZN(n15439) );
  INV_X1 U19003 ( .A(n15435), .ZN(n15436) );
  OAI21_X1 U19004 ( .B1(n15437), .B2(P1_REIP_REG_20__SCAN_IN), .A(n15436), 
        .ZN(n15438) );
  OAI211_X1 U19005 ( .C1(n15578), .C2(n15476), .A(n15439), .B(n15438), .ZN(
        P1_U2820) );
  INV_X1 U19006 ( .A(n15440), .ZN(n15443) );
  AOI21_X1 U19007 ( .B1(n15443), .B2(n10208), .A(n15442), .ZN(n15721) );
  INV_X1 U19008 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n15725) );
  NOR3_X1 U19009 ( .A1(n15459), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n15725), 
        .ZN(n15452) );
  OR2_X1 U19010 ( .A1(n15456), .A2(n15444), .ZN(n15445) );
  NAND2_X1 U19011 ( .A1(n15429), .A2(n15445), .ZN(n16791) );
  AOI21_X1 U19012 ( .B1(n20593), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n13116), .ZN(n15446) );
  OAI21_X1 U19013 ( .B1(n20583), .B2(n15719), .A(n15446), .ZN(n15447) );
  AOI21_X1 U19014 ( .B1(n20602), .B2(P1_EBX_REG_19__SCAN_IN), .A(n15447), .ZN(
        n15450) );
  NAND3_X1 U19015 ( .A1(n15448), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n16694), 
        .ZN(n15449) );
  OAI211_X1 U19016 ( .C1(n16791), .C2(n20580), .A(n15450), .B(n15449), .ZN(
        n15451) );
  AOI211_X1 U19017 ( .C1(n15721), .C2(n20554), .A(n15452), .B(n15451), .ZN(
        n15453) );
  INV_X1 U19018 ( .A(n15453), .ZN(P1_U2821) );
  AOI21_X1 U19019 ( .B1(n15455), .B2(n15454), .A(n15441), .ZN(n15729) );
  INV_X1 U19020 ( .A(n15729), .ZN(n15586) );
  INV_X1 U19021 ( .A(n15508), .ZN(n15457) );
  AOI21_X1 U19022 ( .B1(n15458), .B2(n15457), .A(n15456), .ZN(n15876) );
  OAI22_X1 U19023 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15459), .B1(n15727), 
        .B2(n20583), .ZN(n15463) );
  INV_X1 U19024 ( .A(n16694), .ZN(n15479) );
  NOR2_X1 U19025 ( .A1(n15479), .A2(n15460), .ZN(n16690) );
  AOI22_X1 U19026 ( .A1(P1_EBX_REG_18__SCAN_IN), .A2(n20602), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n16690), .ZN(n15461) );
  OAI211_X1 U19027 ( .C1(n20581), .C2(n14849), .A(n15461), .B(n16808), .ZN(
        n15462) );
  AOI211_X1 U19028 ( .C1(n15876), .C2(n20595), .A(n15463), .B(n15462), .ZN(
        n15464) );
  OAI21_X1 U19029 ( .B1(n15586), .B2(n15476), .A(n15464), .ZN(P1_U2822) );
  AOI21_X1 U19030 ( .B1(n15466), .B2(n14767), .A(n15465), .ZN(n15776) );
  INV_X1 U19031 ( .A(n15776), .ZN(n15615) );
  NOR2_X1 U19032 ( .A1(n15467), .A2(n16729), .ZN(n16717) );
  INV_X1 U19033 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20970) );
  AND2_X1 U19034 ( .A1(n15469), .A2(n15468), .ZN(n15470) );
  OR2_X1 U19035 ( .A1(n15470), .A2(n15524), .ZN(n16809) );
  AOI21_X1 U19036 ( .B1(n20593), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n13116), .ZN(n15472) );
  AOI22_X1 U19037 ( .A1(n15772), .A2(n20604), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n20602), .ZN(n15471) );
  OAI211_X1 U19038 ( .C1(n20580), .C2(n16809), .A(n15472), .B(n15471), .ZN(
        n15473) );
  AOI221_X1 U19039 ( .B1(n16717), .B2(n20970), .C1(n15474), .C2(
        P1_REIP_REG_13__SCAN_IN), .A(n15473), .ZN(n15475) );
  OAI21_X1 U19040 ( .B1(n15615), .B2(n15476), .A(n15475), .ZN(P1_U2827) );
  NAND2_X1 U19041 ( .A1(n20581), .A2(n20583), .ZN(n15477) );
  INV_X1 U19042 ( .A(n20599), .ZN(n20575) );
  AOI22_X1 U19043 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n15477), .B1(
        n20575), .B2(n15925), .ZN(n15478) );
  OAI21_X1 U19044 ( .B1(n20580), .B2(n20651), .A(n15478), .ZN(n15481) );
  NOR2_X1 U19045 ( .A1(n15479), .A2(n12980), .ZN(n15480) );
  AOI211_X1 U19046 ( .C1(n20602), .C2(P1_EBX_REG_0__SCAN_IN), .A(n15481), .B(
        n15480), .ZN(n15482) );
  OAI21_X1 U19047 ( .B1(n20585), .B2(n15483), .A(n15482), .ZN(P1_U2840) );
  INV_X1 U19048 ( .A(n15484), .ZN(n15486) );
  INV_X1 U19049 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15485) );
  OAI22_X1 U19050 ( .A1(n15486), .A2(n16730), .B1(n15485), .B2(n20618), .ZN(
        P1_U2841) );
  INV_X1 U19051 ( .A(n15635), .ZN(n15540) );
  OAI222_X1 U19052 ( .A1(n15487), .A2(n20618), .B1(n16730), .B2(n15800), .C1(
        n15540), .C2(n15513), .ZN(P1_U2843) );
  OAI222_X1 U19053 ( .A1(n15489), .A2(n20618), .B1(n16730), .B2(n15488), .C1(
        n15646), .C2(n15513), .ZN(P1_U2844) );
  INV_X1 U19054 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15491) );
  INV_X1 U19055 ( .A(n15650), .ZN(n15548) );
  OAI222_X1 U19056 ( .A1(n15491), .A2(n20618), .B1(n16730), .B2(n15490), .C1(
        n15548), .C2(n15513), .ZN(P1_U2845) );
  AOI22_X1 U19057 ( .A1(n15829), .A2(n21040), .B1(n21041), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n15492) );
  OAI21_X1 U19058 ( .B1(n15660), .B2(n15513), .A(n15492), .ZN(P1_U2846) );
  INV_X1 U19059 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15494) );
  OAI222_X1 U19060 ( .A1(n15494), .A2(n20618), .B1(n16730), .B2(n15493), .C1(
        n15673), .C2(n15513), .ZN(P1_U2847) );
  OAI222_X1 U19061 ( .A1(n15496), .A2(n20618), .B1(n16730), .B2(n15495), .C1(
        n15681), .C2(n15513), .ZN(P1_U2848) );
  OAI222_X1 U19062 ( .A1(n15498), .A2(n20618), .B1(n16730), .B2(n15497), .C1(
        n15563), .C2(n15513), .ZN(P1_U2849) );
  INV_X1 U19063 ( .A(n16778), .ZN(n15499) );
  INV_X1 U19064 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n21111) );
  OAI222_X1 U19065 ( .A1(n15499), .A2(n16730), .B1(n21111), .B2(n20618), .C1(
        n15569), .C2(n15513), .ZN(P1_U2850) );
  INV_X1 U19066 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15500) );
  OAI222_X1 U19067 ( .A1(n16657), .A2(n16730), .B1(n15500), .B2(n20618), .C1(
        n15513), .C2(n15702), .ZN(P1_U2851) );
  INV_X1 U19068 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15501) );
  OAI222_X1 U19069 ( .A1(n16669), .A2(n16730), .B1(n15501), .B2(n20618), .C1(
        n15578), .C2(n15513), .ZN(P1_U2852) );
  INV_X1 U19070 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15502) );
  INV_X1 U19071 ( .A(n15721), .ZN(n15582) );
  OAI222_X1 U19072 ( .A1(n16791), .A2(n16730), .B1(n15502), .B2(n20618), .C1(
        n15513), .C2(n15582), .ZN(P1_U2853) );
  AOI22_X1 U19073 ( .A1(n15876), .A2(n21040), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n21041), .ZN(n15503) );
  OAI21_X1 U19074 ( .B1(n15586), .B2(n15529), .A(n15503), .ZN(P1_U2854) );
  NAND2_X1 U19075 ( .A1(n15504), .A2(n15505), .ZN(n15506) );
  AND2_X1 U19076 ( .A1(n15454), .A2(n15506), .ZN(n16689) );
  AND2_X1 U19077 ( .A1(n9717), .A2(n15507), .ZN(n15509) );
  OR2_X1 U19078 ( .A1(n15509), .A2(n15508), .ZN(n16799) );
  OAI22_X1 U19079 ( .A1(n16799), .A2(n16730), .B1(n15510), .B2(n20618), .ZN(
        n15511) );
  INV_X1 U19080 ( .A(n15511), .ZN(n15512) );
  OAI21_X1 U19081 ( .B1(n15743), .B2(n15513), .A(n15512), .ZN(P1_U2855) );
  OR2_X1 U19082 ( .A1(n9731), .A2(n15515), .ZN(n15516) );
  AND2_X1 U19083 ( .A1(n15514), .A2(n15516), .ZN(n16712) );
  OR2_X1 U19084 ( .A1(n15525), .A2(n15517), .ZN(n15518) );
  NAND2_X1 U19085 ( .A1(n9800), .A2(n15518), .ZN(n16801) );
  OAI22_X1 U19086 ( .A1(n16801), .A2(n16730), .B1(n16707), .B2(n20618), .ZN(
        n15519) );
  AOI21_X1 U19087 ( .B1(n16712), .B2(n21042), .A(n15519), .ZN(n15520) );
  INV_X1 U19088 ( .A(n15520), .ZN(P1_U2857) );
  INV_X1 U19089 ( .A(n15521), .ZN(n15523) );
  INV_X1 U19090 ( .A(n15465), .ZN(n15522) );
  AOI21_X1 U19091 ( .B1(n15523), .B2(n15522), .A(n9731), .ZN(n16736) );
  INV_X1 U19092 ( .A(n16736), .ZN(n15609) );
  INV_X1 U19093 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15528) );
  INV_X1 U19094 ( .A(n15524), .ZN(n15526) );
  AOI21_X1 U19095 ( .B1(n15527), .B2(n15526), .A(n15525), .ZN(n16715) );
  INV_X1 U19096 ( .A(n16715), .ZN(n15898) );
  OAI222_X1 U19097 ( .A1(n15609), .A2(n15529), .B1(n20618), .B2(n15528), .C1(
        n15898), .C2(n16730), .ZN(P1_U2858) );
  OAI22_X1 U19098 ( .A1(n16809), .A2(n16730), .B1(n15530), .B2(n20618), .ZN(
        n15531) );
  AOI21_X1 U19099 ( .B1(n15776), .B2(n21042), .A(n15531), .ZN(n15532) );
  INV_X1 U19100 ( .A(n15532), .ZN(P1_U2859) );
  NAND3_X1 U19101 ( .A1(n15534), .A2(n15533), .A3(n15606), .ZN(n15536) );
  AOI22_X1 U19102 ( .A1(n15600), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15610), .ZN(n15535) );
  OAI211_X1 U19103 ( .C1(n15594), .C2(n19903), .A(n15536), .B(n15535), .ZN(
        P1_U2873) );
  OAI22_X1 U19104 ( .A1(n15594), .A2(n17170), .B1(n12943), .B2(n15606), .ZN(
        n15537) );
  INV_X1 U19105 ( .A(n15537), .ZN(n15539) );
  AOI22_X1 U19106 ( .A1(n15595), .A2(n15611), .B1(n15600), .B2(DATAI_29_), 
        .ZN(n15538) );
  OAI211_X1 U19107 ( .C1(n15540), .C2(n15614), .A(n15539), .B(n15538), .ZN(
        P1_U2875) );
  AOI22_X1 U19108 ( .A1(n15587), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n15610), .ZN(n15543) );
  AOI22_X1 U19109 ( .A1(n15595), .A2(n15541), .B1(n15600), .B2(DATAI_28_), 
        .ZN(n15542) );
  OAI211_X1 U19110 ( .C1(n15646), .C2(n15614), .A(n15543), .B(n15542), .ZN(
        P1_U2876) );
  OAI22_X1 U19111 ( .A1(n15594), .A2(n19885), .B1(n12930), .B2(n15606), .ZN(
        n15544) );
  INV_X1 U19112 ( .A(n15544), .ZN(n15547) );
  AOI22_X1 U19113 ( .A1(n15595), .A2(n15545), .B1(n15600), .B2(DATAI_27_), 
        .ZN(n15546) );
  OAI211_X1 U19114 ( .C1(n15548), .C2(n15614), .A(n15547), .B(n15546), .ZN(
        P1_U2877) );
  AOI22_X1 U19115 ( .A1(n15587), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n15610), .ZN(n15551) );
  AOI22_X1 U19116 ( .A1(n15595), .A2(n15549), .B1(n15600), .B2(DATAI_26_), 
        .ZN(n15550) );
  OAI211_X1 U19117 ( .C1(n15660), .C2(n15614), .A(n15551), .B(n15550), .ZN(
        P1_U2878) );
  AOI22_X1 U19118 ( .A1(n15587), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n15610), .ZN(n15554) );
  AOI22_X1 U19119 ( .A1(n15595), .A2(n15552), .B1(n15600), .B2(DATAI_25_), 
        .ZN(n15553) );
  OAI211_X1 U19120 ( .C1(n15673), .C2(n15614), .A(n15554), .B(n15553), .ZN(
        P1_U2879) );
  OAI22_X1 U19121 ( .A1(n15594), .A2(n17178), .B1(n12940), .B2(n15606), .ZN(
        n15555) );
  INV_X1 U19122 ( .A(n15555), .ZN(n15558) );
  AOI22_X1 U19123 ( .A1(n15595), .A2(n15556), .B1(n15600), .B2(DATAI_24_), 
        .ZN(n15557) );
  OAI211_X1 U19124 ( .C1(n15681), .C2(n15614), .A(n15558), .B(n15557), .ZN(
        P1_U2880) );
  OAI22_X1 U19125 ( .A1(n15594), .A2(n17180), .B1(n13064), .B2(n15606), .ZN(
        n15559) );
  INV_X1 U19126 ( .A(n15559), .ZN(n15562) );
  AOI22_X1 U19127 ( .A1(n15595), .A2(n15560), .B1(n15600), .B2(DATAI_23_), 
        .ZN(n15561) );
  OAI211_X1 U19128 ( .C1(n15563), .C2(n15614), .A(n15562), .B(n15561), .ZN(
        P1_U2881) );
  OAI22_X1 U19129 ( .A1(n15594), .A2(n17182), .B1(n15564), .B2(n15606), .ZN(
        n15565) );
  INV_X1 U19130 ( .A(n15565), .ZN(n15568) );
  AOI22_X1 U19131 ( .A1(n15595), .A2(n15566), .B1(n15600), .B2(DATAI_22_), 
        .ZN(n15567) );
  OAI211_X1 U19132 ( .C1(n15569), .C2(n15614), .A(n15568), .B(n15567), .ZN(
        P1_U2882) );
  AOI22_X1 U19133 ( .A1(n15587), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n15610), .ZN(n15572) );
  AOI22_X1 U19134 ( .A1(n15595), .A2(n15570), .B1(n15600), .B2(DATAI_21_), 
        .ZN(n15571) );
  OAI211_X1 U19135 ( .C1(n15702), .C2(n15614), .A(n15572), .B(n15571), .ZN(
        P1_U2883) );
  OAI22_X1 U19136 ( .A1(n15594), .A2(n21269), .B1(n15573), .B2(n15606), .ZN(
        n15574) );
  INV_X1 U19137 ( .A(n15574), .ZN(n15577) );
  AOI22_X1 U19138 ( .A1(n15595), .A2(n15575), .B1(n15600), .B2(DATAI_20_), 
        .ZN(n15576) );
  OAI211_X1 U19139 ( .C1(n15578), .C2(n15614), .A(n15577), .B(n15576), .ZN(
        P1_U2884) );
  AOI22_X1 U19140 ( .A1(n15587), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n15610), .ZN(n15581) );
  AOI22_X1 U19141 ( .A1(n15595), .A2(n15579), .B1(n15600), .B2(DATAI_19_), 
        .ZN(n15580) );
  OAI211_X1 U19142 ( .C1(n15582), .C2(n15614), .A(n15581), .B(n15580), .ZN(
        P1_U2885) );
  AOI22_X1 U19143 ( .A1(n15587), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n15610), .ZN(n15585) );
  AOI22_X1 U19144 ( .A1(n15595), .A2(n15583), .B1(n15600), .B2(DATAI_18_), 
        .ZN(n15584) );
  OAI211_X1 U19145 ( .C1(n15586), .C2(n15614), .A(n15585), .B(n15584), .ZN(
        P1_U2886) );
  AOI22_X1 U19146 ( .A1(n15587), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n15610), .ZN(n15590) );
  AOI22_X1 U19147 ( .A1(n15595), .A2(n15588), .B1(n15600), .B2(DATAI_17_), 
        .ZN(n15589) );
  OAI211_X1 U19148 ( .C1(n15743), .C2(n15614), .A(n15590), .B(n15589), .ZN(
        P1_U2887) );
  NAND2_X1 U19149 ( .A1(n15514), .A2(n15591), .ZN(n15592) );
  AND2_X1 U19150 ( .A1(n15504), .A2(n15592), .ZN(n16733) );
  INV_X1 U19151 ( .A(n16733), .ZN(n15602) );
  OAI22_X1 U19152 ( .A1(n15594), .A2(n21227), .B1(n15593), .B2(n15606), .ZN(
        n15599) );
  INV_X1 U19153 ( .A(n15595), .ZN(n15597) );
  NOR2_X1 U19154 ( .A1(n15597), .A2(n15596), .ZN(n15598) );
  AOI211_X1 U19155 ( .C1(n15600), .C2(DATAI_16_), .A(n15599), .B(n15598), .ZN(
        n15601) );
  OAI21_X1 U19156 ( .B1(n15602), .B2(n15614), .A(n15601), .ZN(P1_U2888) );
  INV_X1 U19157 ( .A(n16712), .ZN(n15604) );
  OAI222_X1 U19158 ( .A1(n15604), .A2(n15614), .B1(n15608), .B2(n15603), .C1(
        n15606), .C2(n20621), .ZN(P1_U2889) );
  INV_X1 U19159 ( .A(n15605), .ZN(n15607) );
  INV_X1 U19160 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21179) );
  OAI222_X1 U19161 ( .A1(n15609), .A2(n15614), .B1(n15608), .B2(n15607), .C1(
        n15606), .C2(n21179), .ZN(P1_U2890) );
  AOI22_X1 U19162 ( .A1(n15612), .A2(n15611), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15610), .ZN(n15613) );
  OAI21_X1 U19163 ( .B1(n15615), .B2(n15614), .A(n15613), .ZN(P1_U2891) );
  INV_X1 U19164 ( .A(n15629), .ZN(n15617) );
  AOI21_X1 U19165 ( .B1(n15618), .B2(n15617), .A(n15616), .ZN(n15619) );
  XOR2_X1 U19166 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n15619), .Z(
        n15798) );
  NAND2_X1 U19167 ( .A1(n13116), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15792) );
  NAND2_X1 U19168 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15620) );
  OAI211_X1 U19169 ( .C1(n16769), .C2(n15621), .A(n15792), .B(n15620), .ZN(
        n15622) );
  INV_X1 U19170 ( .A(n15622), .ZN(n15623) );
  INV_X1 U19171 ( .A(n15625), .ZN(n15626) );
  OAI21_X1 U19172 ( .B1(n15798), .B2(n20516), .A(n15626), .ZN(P1_U2969) );
  NAND2_X1 U19173 ( .A1(n15629), .A2(n15628), .ZN(n15630) );
  XNOR2_X1 U19174 ( .A(n15627), .B(n15630), .ZN(n15806) );
  NAND2_X1 U19175 ( .A1(n16742), .A2(n15631), .ZN(n15632) );
  NAND2_X1 U19176 ( .A1(n13116), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15799) );
  OAI211_X1 U19177 ( .C1(n16774), .C2(n15633), .A(n15632), .B(n15799), .ZN(
        n15634) );
  AOI21_X1 U19178 ( .B1(n15635), .B2(n16764), .A(n15634), .ZN(n15636) );
  OAI21_X1 U19179 ( .B1(n20516), .B2(n15806), .A(n15636), .ZN(P1_U2970) );
  NOR2_X1 U19180 ( .A1(n16808), .A2(n21319), .ZN(n15807) );
  NOR2_X1 U19181 ( .A1(n16769), .A2(n15637), .ZN(n15638) );
  AOI211_X1 U19182 ( .C1(n16759), .C2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15807), .B(n15638), .ZN(n15645) );
  NAND3_X1 U19183 ( .A1(n9714), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15642) );
  OR4_X1 U19184 ( .A1(n9714), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(n15639), .ZN(n15641) );
  NAND2_X1 U19185 ( .A1(n9714), .A2(n15826), .ZN(n15657) );
  NAND2_X1 U19186 ( .A1(n15683), .A2(n15657), .ZN(n15640) );
  MUX2_X1 U19187 ( .A(n15642), .B(n15641), .S(n15640), .Z(n15643) );
  XNOR2_X1 U19188 ( .A(n15643), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15813) );
  NAND2_X1 U19189 ( .A1(n15813), .A2(n16772), .ZN(n15644) );
  OAI211_X1 U19190 ( .C1(n15646), .C2(n16770), .A(n15645), .B(n15644), .ZN(
        P1_U2971) );
  MUX2_X1 U19191 ( .A(n9773), .B(n15647), .S(n15209), .Z(n15649) );
  XNOR2_X1 U19192 ( .A(n15649), .B(n15648), .ZN(n15824) );
  NAND2_X1 U19193 ( .A1(n15650), .A2(n16764), .ZN(n15656) );
  NOR2_X1 U19194 ( .A1(n16808), .A2(n15651), .ZN(n15815) );
  NOR2_X1 U19195 ( .A1(n16774), .A2(n15652), .ZN(n15653) );
  AOI211_X1 U19196 ( .C1(n16742), .C2(n15654), .A(n15815), .B(n15653), .ZN(
        n15655) );
  OAI211_X1 U19197 ( .C1(n15824), .C2(n20516), .A(n15656), .B(n15655), .ZN(
        P1_U2972) );
  OAI211_X1 U19198 ( .C1(n15658), .C2(n9714), .A(n9943), .B(n15657), .ZN(
        n15659) );
  XOR2_X1 U19199 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15659), .Z(
        n15834) );
  INV_X1 U19200 ( .A(n15660), .ZN(n15664) );
  NAND2_X1 U19201 ( .A1(n13116), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15825) );
  NAND2_X1 U19202 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15661) );
  OAI211_X1 U19203 ( .C1(n16769), .C2(n15662), .A(n15825), .B(n15661), .ZN(
        n15663) );
  AOI21_X1 U19204 ( .B1(n15664), .B2(n16764), .A(n15663), .ZN(n15665) );
  OAI21_X1 U19205 ( .B1(n20516), .B2(n15834), .A(n15665), .ZN(P1_U2973) );
  NOR2_X1 U19206 ( .A1(n16808), .A2(n15666), .ZN(n15837) );
  NOR2_X1 U19207 ( .A1(n16774), .A2(n15667), .ZN(n15668) );
  AOI211_X1 U19208 ( .C1(n16742), .C2(n15669), .A(n15837), .B(n15668), .ZN(
        n15672) );
  NAND2_X1 U19209 ( .A1(n15835), .A2(n16772), .ZN(n15671) );
  OAI211_X1 U19210 ( .C1(n15673), .C2(n16770), .A(n15672), .B(n15671), .ZN(
        P1_U2974) );
  NOR2_X1 U19211 ( .A1(n16808), .A2(n20985), .ZN(n15844) );
  NOR2_X1 U19212 ( .A1(n16769), .A2(n15674), .ZN(n15675) );
  AOI211_X1 U19213 ( .C1(n16759), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15844), .B(n15675), .ZN(n15680) );
  AOI21_X1 U19214 ( .B1(n15858), .B2(n9714), .A(n9780), .ZN(n15678) );
  XNOR2_X1 U19215 ( .A(n9714), .B(n15676), .ZN(n15677) );
  XNOR2_X1 U19216 ( .A(n15678), .B(n15677), .ZN(n15842) );
  NAND2_X1 U19217 ( .A1(n15842), .A2(n16772), .ZN(n15679) );
  OAI211_X1 U19218 ( .C1(n15681), .C2(n16770), .A(n15680), .B(n15679), .ZN(
        P1_U2975) );
  XNOR2_X1 U19219 ( .A(n9714), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15682) );
  XNOR2_X1 U19220 ( .A(n15683), .B(n15682), .ZN(n15861) );
  NAND2_X1 U19221 ( .A1(n16742), .A2(n15684), .ZN(n15685) );
  NAND2_X1 U19222 ( .A1(n13116), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15854) );
  OAI211_X1 U19223 ( .C1(n16774), .C2(n15686), .A(n15685), .B(n15854), .ZN(
        n15687) );
  AOI21_X1 U19224 ( .B1(n15688), .B2(n16764), .A(n15687), .ZN(n15689) );
  OAI21_X1 U19225 ( .B1(n20516), .B2(n15861), .A(n15689), .ZN(P1_U2976) );
  OAI21_X1 U19226 ( .B1(n15691), .B2(n9714), .A(n15690), .ZN(n15692) );
  XOR2_X1 U19227 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15692), .Z(
        n16777) );
  AOI22_X1 U19228 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15693) );
  OAI21_X1 U19229 ( .B1(n15694), .B2(n16769), .A(n15693), .ZN(n15695) );
  AOI21_X1 U19230 ( .B1(n15696), .B2(n16764), .A(n15695), .ZN(n15697) );
  OAI21_X1 U19231 ( .B1(n20516), .B2(n16777), .A(n15697), .ZN(P1_U2977) );
  OR2_X1 U19232 ( .A1(n15698), .A2(n9714), .ZN(n15709) );
  OR3_X1 U19233 ( .A1(n15699), .A2(n15209), .A3(n16786), .ZN(n15708) );
  MUX2_X1 U19234 ( .A(n15709), .B(n15708), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n15701) );
  XNOR2_X1 U19235 ( .A(n15701), .B(n15700), .ZN(n16651) );
  INV_X1 U19236 ( .A(n15702), .ZN(n15706) );
  NAND2_X1 U19237 ( .A1(n13116), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16652) );
  NAND2_X1 U19238 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15703) );
  OAI211_X1 U19239 ( .C1(n16769), .C2(n15704), .A(n16652), .B(n15703), .ZN(
        n15705) );
  AOI21_X1 U19240 ( .B1(n15706), .B2(n16764), .A(n15705), .ZN(n15707) );
  OAI21_X1 U19241 ( .B1(n16651), .B2(n20516), .A(n15707), .ZN(P1_U2978) );
  NAND2_X1 U19242 ( .A1(n15709), .A2(n15708), .ZN(n15710) );
  XNOR2_X1 U19243 ( .A(n15710), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16668) );
  AOI22_X1 U19244 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15711) );
  OAI21_X1 U19245 ( .B1(n15712), .B2(n16769), .A(n15711), .ZN(n15713) );
  AOI21_X1 U19246 ( .B1(n15714), .B2(n16764), .A(n15713), .ZN(n15715) );
  OAI21_X1 U19247 ( .B1(n16668), .B2(n20516), .A(n15715), .ZN(P1_U2979) );
  OAI21_X1 U19248 ( .B1(n9714), .B2(n21206), .A(n15699), .ZN(n15717) );
  XNOR2_X1 U19249 ( .A(n9714), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15716) );
  XNOR2_X1 U19250 ( .A(n15717), .B(n15716), .ZN(n16785) );
  AOI22_X1 U19251 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15718) );
  OAI21_X1 U19252 ( .B1(n15719), .B2(n16769), .A(n15718), .ZN(n15720) );
  AOI21_X1 U19253 ( .B1(n15721), .B2(n16764), .A(n15720), .ZN(n15722) );
  OAI21_X1 U19254 ( .B1(n16785), .B2(n20516), .A(n15722), .ZN(P1_U2980) );
  OAI21_X1 U19255 ( .B1(n15724), .B2(n15723), .A(n15699), .ZN(n15879) );
  NOR2_X1 U19256 ( .A1(n16808), .A2(n15725), .ZN(n15875) );
  AOI21_X1 U19257 ( .B1(n16759), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15875), .ZN(n15726) );
  OAI21_X1 U19258 ( .B1(n15727), .B2(n16769), .A(n15726), .ZN(n15728) );
  AOI21_X1 U19259 ( .B1(n15729), .B2(n16764), .A(n15728), .ZN(n15730) );
  OAI21_X1 U19260 ( .B1(n20516), .B2(n15879), .A(n15730), .ZN(P1_U2981) );
  NOR2_X1 U19261 ( .A1(n9714), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15736) );
  NAND2_X1 U19262 ( .A1(n15209), .A2(n15732), .ZN(n15765) );
  NAND2_X1 U19263 ( .A1(n15209), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15768) );
  NAND3_X1 U19264 ( .A1(n15731), .A2(n15765), .A3(n15768), .ZN(n15893) );
  NOR2_X1 U19265 ( .A1(n9714), .A2(n16805), .ZN(n15753) );
  INV_X1 U19266 ( .A(n15733), .ZN(n15734) );
  AOI211_X1 U19267 ( .C1(n15893), .C2(n15756), .A(n15753), .B(n15734), .ZN(
        n15745) );
  NOR2_X1 U19268 ( .A1(n15745), .A2(n15744), .ZN(n15735) );
  MUX2_X1 U19269 ( .A(n15736), .B(n9714), .S(n15735), .Z(n15737) );
  XNOR2_X1 U19270 ( .A(n15737), .B(n16792), .ZN(n16796) );
  NAND2_X1 U19271 ( .A1(n16796), .A2(n16772), .ZN(n15742) );
  INV_X1 U19272 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15738) );
  OAI22_X1 U19273 ( .A1(n16774), .A2(n15739), .B1(n16808), .B2(n15738), .ZN(
        n15740) );
  AOI21_X1 U19274 ( .B1(n16742), .B2(n16685), .A(n15740), .ZN(n15741) );
  OAI211_X1 U19275 ( .C1(n16770), .C2(n15743), .A(n15742), .B(n15741), .ZN(
        P1_U2982) );
  NOR2_X1 U19276 ( .A1(n15745), .A2(n15880), .ZN(n15747) );
  OAI22_X1 U19277 ( .A1(n15747), .A2(n15746), .B1(n15745), .B2(n15744), .ZN(
        n15889) );
  INV_X1 U19278 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15748) );
  NOR2_X1 U19279 ( .A1(n16808), .A2(n15748), .ZN(n15885) );
  NOR2_X1 U19280 ( .A1(n16774), .A2(n15749), .ZN(n15750) );
  AOI211_X1 U19281 ( .C1(n16742), .C2(n16696), .A(n15885), .B(n15750), .ZN(
        n15752) );
  NAND2_X1 U19282 ( .A1(n16733), .A2(n16764), .ZN(n15751) );
  OAI211_X1 U19283 ( .C1(n15889), .C2(n20516), .A(n15752), .B(n15751), .ZN(
        P1_U2983) );
  INV_X1 U19284 ( .A(n15753), .ZN(n15755) );
  NAND2_X1 U19285 ( .A1(n15755), .A2(n15754), .ZN(n15761) );
  INV_X1 U19286 ( .A(n15756), .ZN(n15759) );
  INV_X1 U19287 ( .A(n15757), .ZN(n15758) );
  OAI21_X1 U19288 ( .B1(n15731), .B2(n15759), .A(n15758), .ZN(n15760) );
  XOR2_X1 U19289 ( .A(n15761), .B(n15760), .Z(n16800) );
  AOI22_X1 U19290 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15762) );
  OAI21_X1 U19291 ( .B1(n16710), .B2(n16769), .A(n15762), .ZN(n15763) );
  AOI21_X1 U19292 ( .B1(n16712), .B2(n16764), .A(n15763), .ZN(n15764) );
  OAI21_X1 U19293 ( .B1(n16800), .B2(n20516), .A(n15764), .ZN(P1_U2984) );
  INV_X1 U19294 ( .A(n15731), .ZN(n16747) );
  INV_X1 U19295 ( .A(n15765), .ZN(n15766) );
  AOI21_X1 U19296 ( .B1(n16747), .B2(n15767), .A(n15766), .ZN(n15907) );
  AND2_X1 U19297 ( .A1(n15768), .A2(n15769), .ZN(n15906) );
  NAND2_X1 U19298 ( .A1(n15907), .A2(n15906), .ZN(n15905) );
  NAND2_X1 U19299 ( .A1(n15905), .A2(n15769), .ZN(n15771) );
  XNOR2_X1 U19300 ( .A(n15771), .B(n15770), .ZN(n16807) );
  INV_X1 U19301 ( .A(n15772), .ZN(n15774) );
  AOI22_X1 U19302 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n15773) );
  OAI21_X1 U19303 ( .B1(n15774), .B2(n16769), .A(n15773), .ZN(n15775) );
  AOI21_X1 U19304 ( .B1(n15776), .B2(n16764), .A(n15775), .ZN(n15777) );
  OAI21_X1 U19305 ( .B1(n16807), .B2(n20516), .A(n15777), .ZN(P1_U2986) );
  NAND2_X1 U19306 ( .A1(n15778), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15780) );
  XNOR2_X1 U19307 ( .A(n15731), .B(n15781), .ZN(n15779) );
  MUX2_X1 U19308 ( .A(n15780), .B(n15779), .S(n15193), .Z(n15784) );
  INV_X1 U19309 ( .A(n15778), .ZN(n15783) );
  NAND3_X1 U19310 ( .A1(n15783), .A2(n15209), .A3(n15781), .ZN(n16748) );
  NAND2_X1 U19311 ( .A1(n15784), .A2(n16748), .ZN(n16829) );
  NAND2_X1 U19312 ( .A1(n16829), .A2(n16772), .ZN(n15789) );
  OAI22_X1 U19313 ( .A1(n16774), .A2(n15785), .B1(n16808), .B2(n14388), .ZN(
        n15786) );
  AOI21_X1 U19314 ( .B1(n16742), .B2(n15787), .A(n15786), .ZN(n15788) );
  OAI211_X1 U19315 ( .C1(n15790), .C2(n16770), .A(n15789), .B(n15788), .ZN(
        P1_U2989) );
  INV_X1 U19316 ( .A(n15791), .ZN(n15794) );
  AOI21_X1 U19317 ( .B1(n15804), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15793) );
  OAI21_X1 U19318 ( .B1(n15794), .B2(n15793), .A(n15792), .ZN(n15795) );
  AOI21_X1 U19319 ( .B1(n16857), .B2(n15796), .A(n15795), .ZN(n15797) );
  OAI21_X1 U19320 ( .B1(n15798), .B2(n20653), .A(n15797), .ZN(P1_U3001) );
  OAI21_X1 U19321 ( .B1(n15800), .B2(n20652), .A(n15799), .ZN(n15803) );
  NOR2_X1 U19322 ( .A1(n15801), .A2(n21241), .ZN(n15802) );
  AOI211_X1 U19323 ( .C1(n15804), .C2(n21241), .A(n15803), .B(n15802), .ZN(
        n15805) );
  OAI21_X1 U19324 ( .B1(n15806), .B2(n20653), .A(n15805), .ZN(P1_U3002) );
  XNOR2_X1 U19325 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15811) );
  AOI21_X1 U19326 ( .B1(n15808), .B2(n16857), .A(n15807), .ZN(n15810) );
  NAND3_X1 U19327 ( .A1(n15818), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15817), .ZN(n15809) );
  OAI211_X1 U19328 ( .C1(n15821), .C2(n15811), .A(n15810), .B(n15809), .ZN(
        n15812) );
  AOI21_X1 U19329 ( .B1(n15813), .B2(n16861), .A(n15812), .ZN(n15814) );
  INV_X1 U19330 ( .A(n15814), .ZN(P1_U3003) );
  AOI21_X1 U19331 ( .B1(n15816), .B2(n16857), .A(n15815), .ZN(n15820) );
  NAND3_X1 U19332 ( .A1(n15818), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15817), .ZN(n15819) );
  OAI211_X1 U19333 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15821), .A(
        n15820), .B(n15819), .ZN(n15822) );
  INV_X1 U19334 ( .A(n15822), .ZN(n15823) );
  OAI21_X1 U19335 ( .B1(n15824), .B2(n20653), .A(n15823), .ZN(P1_U3004) );
  INV_X1 U19336 ( .A(n15825), .ZN(n15828) );
  NOR3_X1 U19337 ( .A1(n15852), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15826), .ZN(n15827) );
  AOI211_X1 U19338 ( .C1(n15829), .C2(n16857), .A(n15828), .B(n15827), .ZN(
        n15833) );
  INV_X1 U19339 ( .A(n15841), .ZN(n15831) );
  NOR3_X1 U19340 ( .A1(n15852), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15830), .ZN(n15836) );
  OAI21_X1 U19341 ( .B1(n15831), .B2(n15836), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15832) );
  OAI211_X1 U19342 ( .C1(n15834), .C2(n20653), .A(n15833), .B(n15832), .ZN(
        P1_U3005) );
  NAND2_X1 U19343 ( .A1(n15835), .A2(n16861), .ZN(n15840) );
  AOI211_X1 U19344 ( .C1(n16857), .C2(n15838), .A(n15837), .B(n15836), .ZN(
        n15839) );
  OAI211_X1 U19345 ( .C1(n15841), .C2(n21321), .A(n15840), .B(n15839), .ZN(
        P1_U3006) );
  INV_X1 U19346 ( .A(n15842), .ZN(n15851) );
  NOR3_X1 U19347 ( .A1(n15852), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15858), .ZN(n15843) );
  AOI211_X1 U19348 ( .C1(n16857), .C2(n15845), .A(n15844), .B(n15843), .ZN(
        n15850) );
  NOR2_X1 U19349 ( .A1(n15846), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15847) );
  OAI21_X1 U19350 ( .B1(n15848), .B2(n15847), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15849) );
  OAI211_X1 U19351 ( .C1(n15851), .C2(n20653), .A(n15850), .B(n15849), .ZN(
        P1_U3007) );
  INV_X1 U19352 ( .A(n15852), .ZN(n15859) );
  NAND2_X1 U19353 ( .A1(n15853), .A2(n16857), .ZN(n15855) );
  OAI211_X1 U19354 ( .C1(n15856), .C2(n15858), .A(n15855), .B(n15854), .ZN(
        n15857) );
  AOI21_X1 U19355 ( .B1(n15859), .B2(n15858), .A(n15857), .ZN(n15860) );
  OAI21_X1 U19356 ( .B1(n15861), .B2(n20653), .A(n15860), .ZN(P1_U3008) );
  INV_X1 U19357 ( .A(n20656), .ZN(n15866) );
  INV_X1 U19358 ( .A(n15862), .ZN(n15864) );
  OAI22_X1 U19359 ( .A1(n15866), .A2(n15865), .B1(n15864), .B2(n15863), .ZN(
        n15867) );
  AOI211_X1 U19360 ( .C1(n20657), .C2(n15868), .A(n20658), .B(n15867), .ZN(
        n16814) );
  NAND2_X1 U19361 ( .A1(n16813), .A2(n15869), .ZN(n16811) );
  NAND2_X1 U19362 ( .A1(n16814), .A2(n16811), .ZN(n15902) );
  AOI21_X1 U19363 ( .B1(n21244), .B2(n15870), .A(n15902), .ZN(n16804) );
  OAI21_X1 U19364 ( .B1(n15871), .B2(n15873), .A(n16804), .ZN(n16795) );
  NOR2_X1 U19365 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16806), .ZN(
        n15872) );
  AND2_X1 U19366 ( .A1(n15873), .A2(n15872), .ZN(n15874) );
  AOI211_X1 U19367 ( .C1(n16795), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15875), .B(n15874), .ZN(n15878) );
  NAND2_X1 U19368 ( .A1(n15876), .A2(n16857), .ZN(n15877) );
  OAI211_X1 U19369 ( .C1(n15879), .C2(n20653), .A(n15878), .B(n15877), .ZN(
        P1_U3013) );
  INV_X1 U19370 ( .A(n16804), .ZN(n15882) );
  NOR2_X1 U19371 ( .A1(n15880), .A2(n16806), .ZN(n15881) );
  AOI22_X1 U19372 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15882), .B1(
        n15881), .B2(n16793), .ZN(n15888) );
  NAND2_X1 U19373 ( .A1(n9800), .A2(n15883), .ZN(n15884) );
  NAND2_X1 U19374 ( .A1(n9717), .A2(n15884), .ZN(n16731) );
  INV_X1 U19375 ( .A(n16731), .ZN(n15886) );
  AOI21_X1 U19376 ( .B1(n15886), .B2(n16857), .A(n15885), .ZN(n15887) );
  OAI211_X1 U19377 ( .C1(n15889), .C2(n20653), .A(n15888), .B(n15887), .ZN(
        P1_U3015) );
  INV_X1 U19378 ( .A(n15890), .ZN(n15891) );
  AOI21_X1 U19379 ( .B1(n15893), .B2(n15892), .A(n15891), .ZN(n15895) );
  XNOR2_X1 U19380 ( .A(n15193), .B(n21244), .ZN(n15894) );
  XNOR2_X1 U19381 ( .A(n15895), .B(n15894), .ZN(n16739) );
  NOR2_X1 U19382 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15896), .ZN(
        n15901) );
  INV_X1 U19383 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15897) );
  OAI22_X1 U19384 ( .A1(n15898), .A2(n20652), .B1(n16808), .B2(n15897), .ZN(
        n15899) );
  AOI21_X1 U19385 ( .B1(n15901), .B2(n15900), .A(n15899), .ZN(n15904) );
  NAND2_X1 U19386 ( .A1(n15902), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15903) );
  OAI211_X1 U19387 ( .C1(n16739), .C2(n20653), .A(n15904), .B(n15903), .ZN(
        P1_U3017) );
  OAI21_X1 U19388 ( .B1(n15907), .B2(n15906), .A(n15905), .ZN(n15908) );
  INV_X1 U19389 ( .A(n15908), .ZN(n16746) );
  NAND2_X1 U19390 ( .A1(n15911), .A2(n16750), .ZN(n16815) );
  AOI21_X1 U19391 ( .B1(n15911), .B2(n15910), .A(n15909), .ZN(n15913) );
  AOI211_X1 U19392 ( .C1(n15914), .C2(n15916), .A(n15913), .B(n15912), .ZN(
        n16816) );
  OAI21_X1 U19393 ( .B1(n15915), .B2(n16815), .A(n16816), .ZN(n15918) );
  OAI21_X1 U19394 ( .B1(n15916), .B2(n16859), .A(n15919), .ZN(n15917) );
  OAI21_X1 U19395 ( .B1(n15919), .B2(n15918), .A(n15917), .ZN(n15922) );
  AOI22_X1 U19396 ( .A1(n15920), .A2(n16857), .B1(n13116), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15921) );
  OAI211_X1 U19397 ( .C1(n16746), .C2(n20653), .A(n15922), .B(n15921), .ZN(
        P1_U3019) );
  NAND2_X1 U19398 ( .A1(n15923), .A2(n21290), .ZN(n16643) );
  AOI22_X1 U19399 ( .A1(n15927), .A2(n15926), .B1(n15925), .B2(n15924), .ZN(
        n15928) );
  NAND2_X1 U19400 ( .A1(n16643), .A2(n15928), .ZN(n15929) );
  MUX2_X1 U19401 ( .A(n15929), .B(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(
        n20663), .Z(P1_U3478) );
  NAND2_X1 U19402 ( .A1(n15930), .A2(n15931), .ZN(n15932) );
  AND2_X1 U19403 ( .A1(n16033), .A2(n15932), .ZN(n16330) );
  INV_X1 U19404 ( .A(n16330), .ZN(n15947) );
  AOI211_X1 U19405 ( .C1(n15935), .C2(n15934), .A(n19704), .B(n15933), .ZN(
        n15936) );
  INV_X1 U19406 ( .A(n15936), .ZN(n15946) );
  OR2_X1 U19407 ( .A1(n15939), .A2(n15938), .ZN(n15940) );
  NAND2_X1 U19408 ( .A1(n15937), .A2(n15940), .ZN(n16326) );
  AOI22_X1 U19409 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19697), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19672), .ZN(n15942) );
  NAND2_X1 U19410 ( .A1(n19678), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15941) );
  OAI211_X1 U19411 ( .C1(n16326), .C2(n19703), .A(n15942), .B(n15941), .ZN(
        n15943) );
  AOI21_X1 U19412 ( .B1(n15944), .B2(n19679), .A(n15943), .ZN(n15945) );
  OAI211_X1 U19413 ( .C1(n15947), .C2(n19687), .A(n15946), .B(n15945), .ZN(
        P2_U2829) );
  INV_X1 U19414 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15948) );
  XNOR2_X1 U19415 ( .A(n15949), .B(n15948), .ZN(n15960) );
  AOI21_X1 U19416 ( .B1(n15950), .B2(n16057), .A(n16049), .ZN(n15951) );
  INV_X1 U19417 ( .A(n15951), .ZN(n16960) );
  AOI21_X1 U19418 ( .B1(n15952), .B2(n9725), .A(n10235), .ZN(n16974) );
  INV_X1 U19419 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n15954) );
  AOI22_X1 U19420 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19678), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19672), .ZN(n15953) );
  OAI21_X1 U19421 ( .B1(n19676), .B2(n15954), .A(n15953), .ZN(n15955) );
  AOI21_X1 U19422 ( .B1(n16974), .B2(n19671), .A(n15955), .ZN(n15956) );
  OAI21_X1 U19423 ( .B1(n16960), .B2(n19687), .A(n15956), .ZN(n15959) );
  AOI211_X1 U19424 ( .C1(n15957), .C2(n16201), .A(n19704), .B(n10137), .ZN(
        n15958) );
  AOI211_X1 U19425 ( .C1(n19679), .C2(n15960), .A(n15959), .B(n15958), .ZN(
        n15961) );
  INV_X1 U19426 ( .A(n15961), .ZN(P2_U2831) );
  AOI211_X1 U19427 ( .C1(n9783), .C2(n15973), .A(n15962), .B(n19704), .ZN(
        n15964) );
  INV_X1 U19428 ( .A(n19678), .ZN(n19694) );
  INV_X1 U19429 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20429) );
  OAI22_X1 U19430 ( .A1(n19694), .A2(n11106), .B1(n20429), .B2(n19676), .ZN(
        n15963) );
  AOI211_X1 U19431 ( .C1(n19672), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15964), .B(n15963), .ZN(n15971) );
  NOR2_X1 U19432 ( .A1(n15979), .A2(n15965), .ZN(n15966) );
  OR2_X1 U19433 ( .A1(n16064), .A2(n15966), .ZN(n16961) );
  AND2_X1 U19434 ( .A1(n15983), .A2(n15967), .ZN(n15968) );
  OR2_X1 U19435 ( .A1(n15968), .A2(n16118), .ZN(n16386) );
  OAI22_X1 U19436 ( .A1(n16961), .A2(n19687), .B1(n16386), .B2(n19703), .ZN(
        n15969) );
  INV_X1 U19437 ( .A(n15969), .ZN(n15970) );
  OAI211_X1 U19438 ( .C1(n15972), .C2(n19692), .A(n15971), .B(n15970), .ZN(
        P2_U2834) );
  AOI22_X1 U19439 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19678), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19697), .ZN(n15976) );
  OAI211_X1 U19440 ( .C1(n15974), .C2(n16253), .A(n19684), .B(n15973), .ZN(
        n15975) );
  OAI211_X1 U19441 ( .C1(n19710), .C2(n16253), .A(n15976), .B(n15975), .ZN(
        n15977) );
  AOI21_X1 U19442 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19672), .A(
        n15977), .ZN(n15985) );
  AND2_X1 U19443 ( .A1(n15994), .A2(n15978), .ZN(n15980) );
  OR2_X1 U19444 ( .A1(n15980), .A2(n15979), .ZN(n16399) );
  INV_X1 U19445 ( .A(n16399), .ZN(n16258) );
  NAND2_X1 U19446 ( .A1(n15997), .A2(n15981), .ZN(n15982) );
  NAND2_X1 U19447 ( .A1(n15983), .A2(n15982), .ZN(n16398) );
  INV_X1 U19448 ( .A(n16398), .ZN(n16142) );
  AOI22_X1 U19449 ( .A1(n16258), .A2(n19698), .B1(n16142), .B2(n19671), .ZN(
        n15984) );
  OAI211_X1 U19450 ( .C1(n15986), .C2(n19692), .A(n15985), .B(n15984), .ZN(
        P2_U2835) );
  INV_X1 U19451 ( .A(n15987), .ZN(n16005) );
  NAND2_X1 U19452 ( .A1(n16007), .A2(n15988), .ZN(n15989) );
  XNOR2_X1 U19453 ( .A(n16268), .B(n15989), .ZN(n15990) );
  NAND2_X1 U19454 ( .A1(n15990), .A2(n19684), .ZN(n16004) );
  NAND2_X1 U19455 ( .A1(n15991), .A2(n15992), .ZN(n15993) );
  NAND2_X1 U19456 ( .A1(n15994), .A2(n15993), .ZN(n16965) );
  INV_X1 U19457 ( .A(n16965), .ZN(n16002) );
  OR2_X1 U19458 ( .A1(n9792), .A2(n15995), .ZN(n15996) );
  NAND2_X1 U19459 ( .A1(n15997), .A2(n15996), .ZN(n16404) );
  INV_X1 U19460 ( .A(n16404), .ZN(n16150) );
  OAI21_X1 U19461 ( .B1(n20425), .B2(n19676), .A(n19856), .ZN(n15999) );
  NOR2_X1 U19462 ( .A1(n10144), .A2(n19690), .ZN(n15998) );
  AOI211_X1 U19463 ( .C1(n16150), .C2(n19671), .A(n15999), .B(n15998), .ZN(
        n16000) );
  OAI21_X1 U19464 ( .B1(n16969), .B2(n19694), .A(n16000), .ZN(n16001) );
  AOI21_X1 U19465 ( .B1(n16002), .B2(n19698), .A(n16001), .ZN(n16003) );
  OAI211_X1 U19466 ( .C1(n16005), .C2(n19692), .A(n16004), .B(n16003), .ZN(
        P2_U2836) );
  NAND2_X1 U19467 ( .A1(n16007), .A2(n16006), .ZN(n16008) );
  XNOR2_X1 U19468 ( .A(n16283), .B(n16008), .ZN(n16009) );
  NAND2_X1 U19469 ( .A1(n16009), .A2(n19684), .ZN(n16019) );
  AND2_X1 U19470 ( .A1(n16011), .A2(n16010), .ZN(n16012) );
  INV_X1 U19471 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20420) );
  OAI21_X1 U19472 ( .B1(n20420), .B2(n19676), .A(n19856), .ZN(n16014) );
  NOR2_X1 U19473 ( .A1(n16285), .A2(n19690), .ZN(n16013) );
  AOI211_X1 U19474 ( .C1(n19671), .C2(n16015), .A(n16014), .B(n16013), .ZN(
        n16016) );
  OAI21_X1 U19475 ( .B1(n19694), .B2(n10876), .A(n16016), .ZN(n16017) );
  AOI21_X1 U19476 ( .B1(n10320), .B2(n19698), .A(n16017), .ZN(n16018) );
  OAI211_X1 U19477 ( .C1(n19692), .C2(n16020), .A(n16019), .B(n16018), .ZN(
        P2_U2838) );
  XNOR2_X1 U19478 ( .A(n16022), .B(n16021), .ZN(n16082) );
  NOR2_X1 U19479 ( .A1(n16894), .A2(n19716), .ZN(n16023) );
  AOI21_X1 U19480 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n19716), .A(n16023), .ZN(
        n16024) );
  OAI21_X1 U19481 ( .B1(n16082), .B2(n19713), .A(n16024), .ZN(P2_U2858) );
  INV_X1 U19482 ( .A(n16025), .ZN(n16026) );
  NOR2_X1 U19483 ( .A1(n16027), .A2(n16026), .ZN(n16029) );
  XNOR2_X1 U19484 ( .A(n16029), .B(n16028), .ZN(n16088) );
  NAND2_X1 U19485 ( .A1(n19716), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16031) );
  NAND2_X1 U19486 ( .A1(n16907), .A2(n19712), .ZN(n16030) );
  OAI211_X1 U19487 ( .C1(n16088), .C2(n19713), .A(n16031), .B(n16030), .ZN(
        P2_U2859) );
  NAND2_X1 U19488 ( .A1(n16033), .A2(n16032), .ZN(n16034) );
  NAND2_X1 U19489 ( .A1(n16035), .A2(n16034), .ZN(n16918) );
  AOI21_X1 U19490 ( .B1(n16038), .B2(n16037), .A(n16036), .ZN(n16089) );
  NAND2_X1 U19491 ( .A1(n16089), .A2(n16970), .ZN(n16040) );
  NAND2_X1 U19492 ( .A1(n19716), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16039) );
  OAI211_X1 U19493 ( .C1(n16918), .C2(n19716), .A(n16040), .B(n16039), .ZN(
        P2_U2860) );
  XNOR2_X1 U19494 ( .A(n16042), .B(n16041), .ZN(n16101) );
  NAND2_X1 U19495 ( .A1(n19716), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16044) );
  NAND2_X1 U19496 ( .A1(n16330), .A2(n19712), .ZN(n16043) );
  OAI211_X1 U19497 ( .C1(n16101), .C2(n19713), .A(n16044), .B(n16043), .ZN(
        P2_U2861) );
  OAI21_X1 U19498 ( .B1(n16047), .B2(n16046), .A(n16045), .ZN(n16108) );
  OR2_X1 U19499 ( .A1(n16049), .A2(n16048), .ZN(n16050) );
  NAND2_X1 U19500 ( .A1(n15930), .A2(n16050), .ZN(n16334) );
  MUX2_X1 U19501 ( .A(n10941), .B(n16334), .S(n19712), .Z(n16051) );
  OAI21_X1 U19502 ( .B1(n16108), .B2(n19713), .A(n16051), .ZN(P2_U2862) );
  OAI21_X1 U19503 ( .B1(n16054), .B2(n16053), .A(n16052), .ZN(n16116) );
  NAND2_X1 U19504 ( .A1(n19716), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16059) );
  NAND2_X1 U19505 ( .A1(n16062), .A2(n16055), .ZN(n16056) );
  AND2_X1 U19506 ( .A1(n16057), .A2(n16056), .ZN(n16942) );
  NAND2_X1 U19507 ( .A1(n16942), .A2(n19712), .ZN(n16058) );
  OAI211_X1 U19508 ( .C1(n16116), .C2(n19713), .A(n16059), .B(n16058), .ZN(
        P2_U2864) );
  INV_X1 U19509 ( .A(n16060), .ZN(n16130) );
  OAI21_X1 U19510 ( .B1(n16060), .B2(n10316), .A(n16061), .ZN(n16126) );
  OAI21_X1 U19511 ( .B1(n16064), .B2(n16063), .A(n16062), .ZN(n16219) );
  NOR2_X1 U19512 ( .A1(n16219), .A2(n19716), .ZN(n16065) );
  AOI21_X1 U19513 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n19716), .A(n16065), .ZN(
        n16066) );
  OAI21_X1 U19514 ( .B1(n16126), .B2(n19713), .A(n16066), .ZN(P2_U2865) );
  OAI21_X1 U19515 ( .B1(n16067), .B2(n16069), .A(n16128), .ZN(n16144) );
  MUX2_X1 U19516 ( .A(n16399), .B(n10885), .S(n19716), .Z(n16070) );
  OAI21_X1 U19517 ( .B1(n16144), .B2(n19713), .A(n16070), .ZN(P2_U2867) );
  OAI21_X1 U19518 ( .B1(n14329), .B2(n16072), .A(n16071), .ZN(n16162) );
  OAI21_X1 U19519 ( .B1(n16074), .B2(n16073), .A(n15991), .ZN(n19592) );
  NOR2_X1 U19520 ( .A1(n19592), .A2(n19716), .ZN(n16075) );
  AOI21_X1 U19521 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n19716), .A(n16075), .ZN(
        n16076) );
  OAI21_X1 U19522 ( .B1(n16162), .B2(n19713), .A(n16076), .ZN(P2_U2869) );
  OAI22_X1 U19523 ( .A1(n16155), .A2(n19727), .B1(n19744), .B2(n16077), .ZN(
        n16078) );
  AOI21_X1 U19524 ( .B1(n19717), .B2(BUF2_REG_29__SCAN_IN), .A(n16078), .ZN(
        n16079) );
  OAI21_X1 U19525 ( .B1(n16156), .B2(n17170), .A(n16079), .ZN(n16080) );
  AOI21_X1 U19526 ( .B1(n16895), .B2(n19772), .A(n16080), .ZN(n16081) );
  OAI21_X1 U19527 ( .B1(n16082), .B2(n19754), .A(n16081), .ZN(P2_U2890) );
  AOI22_X1 U19528 ( .A1(n16973), .A2(n19730), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n19771), .ZN(n16084) );
  AOI22_X1 U19529 ( .A1(n19717), .A2(BUF2_REG_28__SCAN_IN), .B1(n19719), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n16083) );
  OAI211_X1 U19530 ( .C1(n16905), .C2(n16085), .A(n16084), .B(n16083), .ZN(
        n16086) );
  INV_X1 U19531 ( .A(n16086), .ZN(n16087) );
  OAI21_X1 U19532 ( .B1(n16088), .B2(n19754), .A(n16087), .ZN(P2_U2891) );
  INV_X1 U19533 ( .A(n16089), .ZN(n16095) );
  NAND2_X1 U19534 ( .A1(n15937), .A2(n16090), .ZN(n16091) );
  AND2_X1 U19535 ( .A1(n9772), .A2(n16091), .ZN(n16311) );
  OAI22_X1 U19536 ( .A1(n16155), .A2(n19733), .B1(n19744), .B2(n21132), .ZN(
        n16092) );
  AOI21_X1 U19537 ( .B1(n16311), .B2(n19772), .A(n16092), .ZN(n16094) );
  AOI22_X1 U19538 ( .A1(n19717), .A2(BUF2_REG_27__SCAN_IN), .B1(n19719), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16093) );
  OAI211_X1 U19539 ( .C1(n16095), .C2(n19754), .A(n16094), .B(n16093), .ZN(
        P2_U2892) );
  INV_X1 U19540 ( .A(n16326), .ZN(n16098) );
  OAI22_X1 U19541 ( .A1(n16155), .A2(n19735), .B1(n19744), .B2(n16096), .ZN(
        n16097) );
  AOI21_X1 U19542 ( .B1(n16098), .B2(n19772), .A(n16097), .ZN(n16100) );
  AOI22_X1 U19543 ( .A1(n19717), .A2(BUF2_REG_26__SCAN_IN), .B1(n19719), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n16099) );
  OAI211_X1 U19544 ( .C1(n16101), .C2(n19754), .A(n16100), .B(n16099), .ZN(
        P2_U2893) );
  XNOR2_X1 U19545 ( .A(n16103), .B(n16102), .ZN(n16338) );
  INV_X1 U19546 ( .A(n16338), .ZN(n16931) );
  OAI22_X1 U19547 ( .A1(n16155), .A2(n19737), .B1(n19744), .B2(n16104), .ZN(
        n16105) );
  AOI21_X1 U19548 ( .B1(n16931), .B2(n19772), .A(n16105), .ZN(n16107) );
  AOI22_X1 U19549 ( .A1(n19717), .A2(BUF2_REG_25__SCAN_IN), .B1(n19719), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n16106) );
  OAI211_X1 U19550 ( .C1(n16108), .C2(n19754), .A(n16107), .B(n16106), .ZN(
        P2_U2894) );
  OR2_X1 U19551 ( .A1(n16120), .A2(n16109), .ZN(n16110) );
  NAND2_X1 U19552 ( .A1(n9725), .A2(n16110), .ZN(n16357) );
  INV_X1 U19553 ( .A(n16357), .ZN(n16941) );
  OAI22_X1 U19554 ( .A1(n16155), .A2(n19908), .B1(n19744), .B2(n16111), .ZN(
        n16114) );
  INV_X1 U19555 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16112) );
  OAI22_X1 U19556 ( .A1(n16158), .A2(n16112), .B1(n16156), .B2(n17180), .ZN(
        n16113) );
  AOI211_X1 U19557 ( .C1(n19772), .C2(n16941), .A(n16114), .B(n16113), .ZN(
        n16115) );
  OAI21_X1 U19558 ( .B1(n16116), .B2(n19754), .A(n16115), .ZN(P2_U2896) );
  NOR2_X1 U19559 ( .A1(n16118), .A2(n16117), .ZN(n16119) );
  OR2_X1 U19560 ( .A1(n16120), .A2(n16119), .ZN(n16372) );
  INV_X1 U19561 ( .A(n16372), .ZN(n16602) );
  OAI22_X1 U19562 ( .A1(n16155), .A2(n19897), .B1(n19744), .B2(n16121), .ZN(
        n16124) );
  INV_X1 U19563 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16122) );
  OAI22_X1 U19564 ( .A1(n16158), .A2(n16122), .B1(n16156), .B2(n17182), .ZN(
        n16123) );
  AOI211_X1 U19565 ( .C1(n19772), .C2(n16602), .A(n16124), .B(n16123), .ZN(
        n16125) );
  OAI21_X1 U19566 ( .B1(n16126), .B2(n19754), .A(n16125), .ZN(P2_U2897) );
  NAND2_X1 U19567 ( .A1(n16128), .A2(n16127), .ZN(n16129) );
  AND2_X1 U19568 ( .A1(n16130), .A2(n16129), .ZN(n16963) );
  INV_X1 U19569 ( .A(n16963), .ZN(n16138) );
  INV_X1 U19570 ( .A(n16386), .ZN(n16136) );
  OAI22_X1 U19571 ( .A1(n16155), .A2(n16132), .B1(n19744), .B2(n16131), .ZN(
        n16135) );
  INV_X1 U19572 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16133) );
  OAI22_X1 U19573 ( .A1(n16158), .A2(n16133), .B1(n16156), .B2(n17184), .ZN(
        n16134) );
  AOI211_X1 U19574 ( .C1(n19772), .C2(n16136), .A(n16135), .B(n16134), .ZN(
        n16137) );
  OAI21_X1 U19575 ( .B1(n16138), .B2(n19754), .A(n16137), .ZN(P2_U2898) );
  OAI22_X1 U19576 ( .A1(n16155), .A2(n19891), .B1(n19744), .B2(n12654), .ZN(
        n16141) );
  INV_X1 U19577 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16139) );
  OAI22_X1 U19578 ( .A1(n16158), .A2(n16139), .B1(n16156), .B2(n21269), .ZN(
        n16140) );
  AOI211_X1 U19579 ( .C1(n19772), .C2(n16142), .A(n16141), .B(n16140), .ZN(
        n16143) );
  OAI21_X1 U19580 ( .B1(n16144), .B2(n19754), .A(n16143), .ZN(P2_U2899) );
  AND2_X1 U19581 ( .A1(n16071), .A2(n16145), .ZN(n16146) );
  OR2_X1 U19582 ( .A1(n16146), .A2(n16067), .ZN(n16966) );
  OAI22_X1 U19583 ( .A1(n16155), .A2(n19886), .B1(n19744), .B2(n12662), .ZN(
        n16149) );
  INV_X1 U19584 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16147) );
  OAI22_X1 U19585 ( .A1(n16158), .A2(n16147), .B1(n16156), .B2(n17187), .ZN(
        n16148) );
  AOI211_X1 U19586 ( .C1(n19772), .C2(n16150), .A(n16149), .B(n16148), .ZN(
        n16151) );
  OAI21_X1 U19587 ( .B1(n16966), .B2(n19754), .A(n16151), .ZN(P2_U2900) );
  AND2_X1 U19588 ( .A1(n16153), .A2(n16152), .ZN(n16154) );
  NOR2_X1 U19589 ( .A1(n9792), .A2(n16154), .ZN(n19593) );
  OAI22_X1 U19590 ( .A1(n16155), .A2(n19881), .B1(n19744), .B2(n21238), .ZN(
        n16160) );
  INV_X1 U19591 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n16157) );
  OAI22_X1 U19592 ( .A1(n16158), .A2(n16157), .B1(n16156), .B2(n17189), .ZN(
        n16159) );
  AOI211_X1 U19593 ( .C1(n19772), .C2(n19593), .A(n16160), .B(n16159), .ZN(
        n16161) );
  OAI21_X1 U19594 ( .B1(n16162), .B2(n19754), .A(n16161), .ZN(P2_U2901) );
  NOR2_X1 U19595 ( .A1(n16164), .A2(n19840), .ZN(n16168) );
  OAI21_X1 U19596 ( .B1(n17046), .B2(n16166), .A(n16165), .ZN(n16167) );
  AOI211_X1 U19597 ( .C1(n16907), .C2(n19848), .A(n16168), .B(n16167), .ZN(
        n16169) );
  XNOR2_X1 U19598 ( .A(n16171), .B(n16312), .ZN(n16321) );
  AOI21_X1 U19599 ( .B1(n16312), .B2(n16172), .A(n9751), .ZN(n16318) );
  NAND2_X1 U19600 ( .A1(n19825), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n16314) );
  OAI21_X1 U19601 ( .B1(n17046), .B2(n16173), .A(n16314), .ZN(n16174) );
  AOI21_X1 U19602 ( .B1(n16922), .B2(n17038), .A(n16174), .ZN(n16175) );
  OAI21_X1 U19603 ( .B1(n16918), .B2(n16307), .A(n16175), .ZN(n16176) );
  AOI21_X1 U19604 ( .B1(n16318), .B2(n11531), .A(n16176), .ZN(n16177) );
  OAI21_X1 U19605 ( .B1(n16321), .B2(n19845), .A(n16177), .ZN(P2_U2987) );
  OAI21_X1 U19606 ( .B1(n16178), .B2(n16186), .A(n16184), .ZN(n16179) );
  XOR2_X1 U19607 ( .A(n16180), .B(n16179), .Z(n16322) );
  NAND2_X1 U19608 ( .A1(n19825), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16325) );
  NAND2_X1 U19609 ( .A1(n19837), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16181) );
  OAI211_X1 U19610 ( .C1(n16182), .C2(n19840), .A(n16325), .B(n16181), .ZN(
        n16183) );
  INV_X1 U19611 ( .A(n16184), .ZN(n16185) );
  NOR2_X1 U19612 ( .A1(n16186), .A2(n16185), .ZN(n16187) );
  XNOR2_X1 U19613 ( .A(n16178), .B(n16187), .ZN(n16346) );
  NAND2_X1 U19614 ( .A1(n19825), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16337) );
  OAI21_X1 U19615 ( .B1(n17046), .B2(n16188), .A(n16337), .ZN(n16190) );
  NOR2_X1 U19616 ( .A1(n16334), .A2(n16307), .ZN(n16189) );
  AOI211_X1 U19617 ( .C1(n17038), .C2(n16935), .A(n16190), .B(n16189), .ZN(
        n16192) );
  NAND2_X1 U19618 ( .A1(n16194), .A2(n16339), .ZN(n16343) );
  NAND3_X1 U19619 ( .A1(n9769), .A2(n11531), .A3(n16343), .ZN(n16191) );
  OAI211_X1 U19620 ( .C1(n16346), .C2(n19845), .A(n16192), .B(n16191), .ZN(
        P2_U2989) );
  OAI21_X1 U19621 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16193), .A(
        n16194), .ZN(n16355) );
  XNOR2_X1 U19622 ( .A(n16196), .B(n16195), .ZN(n16197) );
  XNOR2_X1 U19623 ( .A(n16198), .B(n16197), .ZN(n16353) );
  AND2_X1 U19624 ( .A1(n19825), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16349) );
  NOR2_X1 U19625 ( .A1(n17046), .A2(n16199), .ZN(n16200) );
  AOI211_X1 U19626 ( .C1(n16201), .C2(n17038), .A(n16349), .B(n16200), .ZN(
        n16202) );
  OAI21_X1 U19627 ( .B1(n16960), .B2(n16307), .A(n16202), .ZN(n16203) );
  AOI21_X1 U19628 ( .B1(n16353), .B2(n19828), .A(n16203), .ZN(n16204) );
  OAI21_X1 U19629 ( .B1(n17039), .B2(n16355), .A(n16204), .ZN(P2_U2990) );
  INV_X1 U19630 ( .A(n16205), .ZN(n16207) );
  INV_X1 U19631 ( .A(n16193), .ZN(n16206) );
  OAI21_X1 U19632 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16207), .A(
        n16206), .ZN(n16368) );
  XOR2_X1 U19633 ( .A(n16209), .B(n16208), .Z(n16366) );
  NAND2_X1 U19634 ( .A1(n16366), .A2(n19828), .ZN(n16214) );
  NAND2_X1 U19635 ( .A1(n16945), .A2(n17038), .ZN(n16210) );
  NAND2_X1 U19636 ( .A1(n19825), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16356) );
  OAI211_X1 U19637 ( .C1(n17046), .C2(n16211), .A(n16210), .B(n16356), .ZN(
        n16212) );
  AOI21_X1 U19638 ( .B1(n16942), .B2(n19848), .A(n16212), .ZN(n16213) );
  OAI211_X1 U19639 ( .C1(n16368), .C2(n17039), .A(n16214), .B(n16213), .ZN(
        P2_U2991) );
  NAND2_X1 U19640 ( .A1(n10252), .A2(n16216), .ZN(n16217) );
  XNOR2_X1 U19641 ( .A(n16218), .B(n16217), .ZN(n16382) );
  INV_X1 U19642 ( .A(n16219), .ZN(n16603) );
  NOR2_X1 U19643 ( .A1(n19856), .A2(n16220), .ZN(n16369) );
  AOI21_X1 U19644 ( .B1(n19837), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16369), .ZN(n16221) );
  OAI21_X1 U19645 ( .B1(n16222), .B2(n19840), .A(n16221), .ZN(n16223) );
  AOI21_X1 U19646 ( .B1(n16603), .B2(n19848), .A(n16223), .ZN(n16226) );
  NAND2_X1 U19647 ( .A1(n16224), .A2(n16375), .ZN(n16379) );
  NAND3_X1 U19648 ( .A1(n16205), .A2(n11531), .A3(n16379), .ZN(n16225) );
  OAI211_X1 U19649 ( .C1(n16382), .C2(n19845), .A(n16226), .B(n16225), .ZN(
        P2_U2992) );
  OAI21_X1 U19650 ( .B1(n16227), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16224), .ZN(n16392) );
  INV_X1 U19651 ( .A(n16989), .ZN(n16229) );
  INV_X1 U19652 ( .A(n16987), .ZN(n16228) );
  INV_X1 U19653 ( .A(n16979), .ZN(n16230) );
  INV_X1 U19654 ( .A(n16301), .ZN(n16231) );
  INV_X1 U19655 ( .A(n16232), .ZN(n16290) );
  INV_X1 U19656 ( .A(n16233), .ZN(n16234) );
  NAND2_X1 U19657 ( .A1(n16236), .A2(n16235), .ZN(n16281) );
  INV_X1 U19658 ( .A(n16260), .ZN(n16272) );
  INV_X1 U19659 ( .A(n16238), .ZN(n16248) );
  NAND2_X1 U19660 ( .A1(n16249), .A2(n16248), .ZN(n16239) );
  OAI21_X1 U19661 ( .B1(n16250), .B2(n16239), .A(n16247), .ZN(n16242) );
  NAND2_X1 U19662 ( .A1(n9801), .A2(n16240), .ZN(n16241) );
  XNOR2_X1 U19663 ( .A(n16242), .B(n16241), .ZN(n16383) );
  NAND2_X1 U19664 ( .A1(n16383), .A2(n19828), .ZN(n16246) );
  NAND2_X1 U19665 ( .A1(n19825), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16385) );
  OAI21_X1 U19666 ( .B1(n17046), .B2(n10145), .A(n16385), .ZN(n16244) );
  NOR2_X1 U19667 ( .A1(n16961), .A2(n16307), .ZN(n16243) );
  AOI211_X1 U19668 ( .C1(n17038), .C2(n9783), .A(n16244), .B(n16243), .ZN(
        n16245) );
  OAI211_X1 U19669 ( .C1(n17039), .C2(n16392), .A(n16246), .B(n16245), .ZN(
        P2_U2993) );
  NAND2_X1 U19670 ( .A1(n16248), .A2(n16247), .ZN(n16251) );
  INV_X1 U19671 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20427) );
  NOR2_X1 U19672 ( .A1(n19856), .A2(n20427), .ZN(n16394) );
  AOI21_X1 U19673 ( .B1(n19837), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16394), .ZN(n16252) );
  OAI21_X1 U19674 ( .B1(n16253), .B2(n19840), .A(n16252), .ZN(n16257) );
  NOR2_X1 U19675 ( .A1(n16254), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16255) );
  OR2_X1 U19676 ( .A1(n16227), .A2(n16255), .ZN(n16403) );
  NOR2_X1 U19677 ( .A1(n16403), .A2(n17039), .ZN(n16256) );
  AOI211_X1 U19678 ( .C1(n19848), .C2(n16258), .A(n16257), .B(n16256), .ZN(
        n16259) );
  OAI21_X1 U19679 ( .B1(n16393), .B2(n19845), .A(n16259), .ZN(P2_U2994) );
  INV_X1 U19680 ( .A(n16275), .ZN(n16261) );
  OAI21_X1 U19681 ( .B1(n16261), .B2(n16273), .A(n16260), .ZN(n16265) );
  NOR2_X1 U19682 ( .A1(n16263), .A2(n16262), .ZN(n16264) );
  XNOR2_X1 U19683 ( .A(n16265), .B(n16264), .ZN(n16414) );
  AOI21_X1 U19684 ( .B1(n10313), .B2(n10314), .A(n16254), .ZN(n16411) );
  NAND2_X1 U19685 ( .A1(n19825), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16407) );
  OAI21_X1 U19686 ( .B1(n17046), .B2(n10144), .A(n16407), .ZN(n16267) );
  AOI21_X1 U19687 ( .B1(n16268), .B2(n17038), .A(n16267), .ZN(n16269) );
  OAI21_X1 U19688 ( .B1(n16965), .B2(n16307), .A(n16269), .ZN(n16270) );
  AOI21_X1 U19689 ( .B1(n16411), .B2(n11531), .A(n16270), .ZN(n16271) );
  OAI21_X1 U19690 ( .B1(n16414), .B2(n19845), .A(n16271), .ZN(P2_U2995) );
  NOR2_X1 U19691 ( .A1(n16273), .A2(n16272), .ZN(n16274) );
  XNOR2_X1 U19692 ( .A(n16275), .B(n16274), .ZN(n16426) );
  AOI21_X1 U19693 ( .B1(n16420), .B2(n16276), .A(n16266), .ZN(n16424) );
  NOR2_X1 U19694 ( .A1(n19592), .A2(n16307), .ZN(n16279) );
  NAND2_X1 U19695 ( .A1(n19825), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n16417) );
  NAND2_X1 U19696 ( .A1(n19837), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16277) );
  OAI211_X1 U19697 ( .C1(n19587), .C2(n19840), .A(n16417), .B(n16277), .ZN(
        n16278) );
  AOI211_X1 U19698 ( .C1(n16424), .C2(n11531), .A(n16279), .B(n16278), .ZN(
        n16280) );
  OAI21_X1 U19699 ( .B1(n16426), .B2(n19845), .A(n16280), .ZN(P2_U2996) );
  XNOR2_X1 U19700 ( .A(n16282), .B(n16281), .ZN(n16443) );
  NAND2_X1 U19701 ( .A1(n16283), .A2(n17038), .ZN(n16284) );
  NAND2_X1 U19702 ( .A1(n19825), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16428) );
  OAI211_X1 U19703 ( .C1(n17046), .C2(n16285), .A(n16284), .B(n16428), .ZN(
        n16288) );
  INV_X1 U19704 ( .A(n16276), .ZN(n16286) );
  AOI211_X1 U19705 ( .C1(n16441), .C2(n9761), .A(n17039), .B(n16286), .ZN(
        n16287) );
  AOI211_X1 U19706 ( .C1(n19848), .C2(n10320), .A(n16288), .B(n16287), .ZN(
        n16289) );
  OAI21_X1 U19707 ( .B1(n16443), .B2(n19845), .A(n16289), .ZN(P2_U2997) );
  XNOR2_X1 U19708 ( .A(n16291), .B(n16290), .ZN(n16452) );
  INV_X1 U19709 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n21255) );
  NOR2_X1 U19710 ( .A1(n21255), .A2(n19838), .ZN(n16294) );
  INV_X1 U19711 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16292) );
  OAI22_X1 U19712 ( .A1(n17046), .A2(n16292), .B1(n19840), .B2(n19599), .ZN(
        n16293) );
  AOI211_X1 U19713 ( .C1(n19848), .C2(n19605), .A(n16294), .B(n16293), .ZN(
        n16299) );
  OAI21_X1 U19714 ( .B1(n16296), .B2(n16459), .A(n16444), .ZN(n16297) );
  NAND3_X1 U19715 ( .A1(n9761), .A2(n11531), .A3(n16297), .ZN(n16298) );
  OAI211_X1 U19716 ( .C1(n16452), .C2(n19845), .A(n16299), .B(n16298), .ZN(
        P2_U2998) );
  NAND2_X1 U19717 ( .A1(n16301), .A2(n16300), .ZN(n16302) );
  XNOR2_X1 U19718 ( .A(n16303), .B(n16302), .ZN(n16465) );
  XNOR2_X1 U19719 ( .A(n16296), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16463) );
  OAI22_X1 U19720 ( .A1(n17046), .A2(n16305), .B1(n19840), .B2(n16304), .ZN(
        n16309) );
  INV_X1 U19721 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n16306) );
  OAI22_X1 U19722 ( .A1(n16454), .A2(n16307), .B1(n16306), .B2(n19856), .ZN(
        n16308) );
  AOI211_X1 U19723 ( .C1(n16463), .C2(n11531), .A(n16309), .B(n16308), .ZN(
        n16310) );
  OAI21_X1 U19724 ( .B1(n16465), .B2(n19845), .A(n16310), .ZN(P2_U2999) );
  INV_X1 U19725 ( .A(n16311), .ZN(n16917) );
  NAND3_X1 U19726 ( .A1(n16323), .A2(n16312), .A3(n16335), .ZN(n16313) );
  OAI211_X1 U19727 ( .C1(n16917), .C2(n17070), .A(n16314), .B(n16313), .ZN(
        n16316) );
  NOR2_X1 U19728 ( .A1(n16918), .A2(n19870), .ZN(n16315) );
  AOI211_X1 U19729 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n16317), .A(
        n16316), .B(n16315), .ZN(n16320) );
  NAND2_X1 U19730 ( .A1(n16318), .A2(n11551), .ZN(n16319) );
  OAI211_X1 U19731 ( .C1(n16321), .C2(n16500), .A(n16320), .B(n16319), .ZN(
        P2_U3019) );
  OAI211_X1 U19732 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n9998), .B(n16335), .ZN(n16324) );
  OAI211_X1 U19733 ( .C1(n16326), .C2(n17070), .A(n16325), .B(n16324), .ZN(
        n16329) );
  NOR2_X1 U19734 ( .A1(n16340), .A2(n16327), .ZN(n16328) );
  AOI211_X1 U19735 ( .C1(n16330), .C2(n17086), .A(n16329), .B(n16328), .ZN(
        n16331) );
  OAI211_X1 U19736 ( .C1(n16333), .C2(n19859), .A(n16332), .B(n16331), .ZN(
        P2_U3020) );
  INV_X1 U19737 ( .A(n16334), .ZN(n16932) );
  NAND2_X1 U19738 ( .A1(n16339), .A2(n16335), .ZN(n16336) );
  OAI211_X1 U19739 ( .C1(n17070), .C2(n16338), .A(n16337), .B(n16336), .ZN(
        n16342) );
  NOR2_X1 U19740 ( .A1(n16340), .A2(n16339), .ZN(n16341) );
  AOI211_X1 U19741 ( .C1(n16932), .C2(n17086), .A(n16342), .B(n16341), .ZN(
        n16345) );
  NAND3_X1 U19742 ( .A1(n9769), .A2(n11551), .A3(n16343), .ZN(n16344) );
  OAI211_X1 U19743 ( .C1(n16346), .C2(n16500), .A(n16345), .B(n16344), .ZN(
        P2_U3021) );
  OAI21_X1 U19744 ( .B1(n16348), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16347), .ZN(n16351) );
  AOI21_X1 U19745 ( .B1(n16974), .B2(n19854), .A(n16349), .ZN(n16350) );
  OAI211_X1 U19746 ( .C1(n19870), .C2(n16960), .A(n16351), .B(n16350), .ZN(
        n16352) );
  AOI21_X1 U19747 ( .B1(n16353), .B2(n19866), .A(n16352), .ZN(n16354) );
  OAI21_X1 U19748 ( .B1(n19859), .B2(n16355), .A(n16354), .ZN(P2_U3022) );
  INV_X1 U19749 ( .A(n16376), .ZN(n16389) );
  AOI21_X1 U19750 ( .B1(n16360), .B2(n16374), .A(n16389), .ZN(n16364) );
  OAI21_X1 U19751 ( .B1(n17070), .B2(n16357), .A(n16356), .ZN(n16358) );
  AOI21_X1 U19752 ( .B1(n16942), .B2(n17086), .A(n16358), .ZN(n16362) );
  INV_X1 U19753 ( .A(n16359), .ZN(n16370) );
  NAND3_X1 U19754 ( .A1(n16360), .A2(n16370), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16361) );
  OAI211_X1 U19755 ( .C1(n16364), .C2(n16363), .A(n16362), .B(n16361), .ZN(
        n16365) );
  AOI21_X1 U19756 ( .B1(n16366), .B2(n19866), .A(n16365), .ZN(n16367) );
  OAI21_X1 U19757 ( .B1(n19859), .B2(n16368), .A(n16367), .ZN(P2_U3023) );
  AOI21_X1 U19758 ( .B1(n16370), .B2(n16375), .A(n16369), .ZN(n16371) );
  OAI21_X1 U19759 ( .B1(n17070), .B2(n16372), .A(n16371), .ZN(n16378) );
  NAND2_X1 U19760 ( .A1(n16374), .A2(n16373), .ZN(n16384) );
  AOI21_X1 U19761 ( .B1(n16376), .B2(n16384), .A(n16375), .ZN(n16377) );
  AOI211_X1 U19762 ( .C1(n16603), .C2(n17086), .A(n16378), .B(n16377), .ZN(
        n16381) );
  NAND3_X1 U19763 ( .A1(n16205), .A2(n11551), .A3(n16379), .ZN(n16380) );
  OAI211_X1 U19764 ( .C1(n16382), .C2(n16500), .A(n16381), .B(n16380), .ZN(
        P2_U3024) );
  NAND2_X1 U19765 ( .A1(n16383), .A2(n19866), .ZN(n16391) );
  OAI211_X1 U19766 ( .C1(n17070), .C2(n16386), .A(n16385), .B(n16384), .ZN(
        n16388) );
  NOR2_X1 U19767 ( .A1(n16961), .A2(n19870), .ZN(n16387) );
  AOI211_X1 U19768 ( .C1(n16389), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16388), .B(n16387), .ZN(n16390) );
  OAI211_X1 U19769 ( .C1(n16392), .C2(n19859), .A(n16391), .B(n16390), .ZN(
        P2_U3025) );
  INV_X1 U19770 ( .A(n16394), .ZN(n16397) );
  OAI211_X1 U19771 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16405), .B(n16395), .ZN(
        n16396) );
  OAI211_X1 U19772 ( .C1(n17070), .C2(n16398), .A(n16397), .B(n16396), .ZN(
        n16401) );
  NOR2_X1 U19773 ( .A1(n16399), .A2(n19870), .ZN(n16400) );
  AOI211_X1 U19774 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n16410), .A(
        n16401), .B(n16400), .ZN(n16402) );
  NOR2_X1 U19775 ( .A1(n17070), .A2(n16404), .ZN(n16409) );
  NAND2_X1 U19776 ( .A1(n16405), .A2(n10313), .ZN(n16406) );
  OAI211_X1 U19777 ( .C1(n16965), .C2(n19870), .A(n16407), .B(n16406), .ZN(
        n16408) );
  AOI211_X1 U19778 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16410), .A(
        n16409), .B(n16408), .ZN(n16413) );
  NAND2_X1 U19779 ( .A1(n16411), .A2(n11551), .ZN(n16412) );
  OAI211_X1 U19780 ( .C1(n16414), .C2(n16500), .A(n16413), .B(n16412), .ZN(
        P2_U3027) );
  NAND2_X1 U19781 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16415), .ZN(
        n17052) );
  INV_X1 U19782 ( .A(n17052), .ZN(n17057) );
  NAND2_X1 U19783 ( .A1(n17057), .A2(n11481), .ZN(n16453) );
  NOR3_X1 U19784 ( .A1(n16453), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16416), .ZN(n16423) );
  OAI21_X1 U19785 ( .B1(n19592), .B2(n19870), .A(n16417), .ZN(n16418) );
  AOI21_X1 U19786 ( .B1(n19854), .B2(n19593), .A(n16418), .ZN(n16419) );
  OAI21_X1 U19787 ( .B1(n16421), .B2(n16420), .A(n16419), .ZN(n16422) );
  AOI211_X1 U19788 ( .C1(n16424), .C2(n11551), .A(n16423), .B(n16422), .ZN(
        n16425) );
  OAI21_X1 U19789 ( .B1(n16426), .B2(n16500), .A(n16425), .ZN(P2_U3028) );
  OAI22_X1 U19790 ( .A1(n9761), .A2(n19859), .B1(n16427), .B2(n16453), .ZN(
        n16440) );
  NAND2_X1 U19791 ( .A1(n10320), .A2(n17086), .ZN(n16429) );
  OAI211_X1 U19792 ( .C1(n17070), .C2(n16430), .A(n16429), .B(n16428), .ZN(
        n16439) );
  INV_X1 U19793 ( .A(n16431), .ZN(n19853) );
  OAI21_X1 U19794 ( .B1(n11551), .B2(n19853), .A(n9761), .ZN(n16435) );
  OR2_X1 U19795 ( .A1(n16432), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16433) );
  NAND2_X1 U19796 ( .A1(n16508), .A2(n16433), .ZN(n17053) );
  AOI21_X1 U19797 ( .B1(n16434), .B2(n17054), .A(n17053), .ZN(n16460) );
  OAI211_X1 U19798 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16436), .A(
        n16435), .B(n16460), .ZN(n16450) );
  AOI21_X1 U19799 ( .B1(n16444), .B2(n17054), .A(n16450), .ZN(n16437) );
  NOR2_X1 U19800 ( .A1(n16437), .A2(n16441), .ZN(n16438) );
  OAI21_X1 U19801 ( .B1(n16443), .B2(n16500), .A(n16442), .ZN(P2_U3029) );
  OAI21_X1 U19802 ( .B1(n16296), .B2(n19859), .A(n16453), .ZN(n16445) );
  NAND3_X1 U19803 ( .A1(n16445), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16444), .ZN(n16447) );
  AOI22_X1 U19804 ( .A1(n19605), .A2(n17086), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19825), .ZN(n16446) );
  OAI211_X1 U19805 ( .C1(n17070), .C2(n16448), .A(n16447), .B(n16446), .ZN(
        n16449) );
  AOI21_X1 U19806 ( .B1(n16450), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16449), .ZN(n16451) );
  OAI21_X1 U19807 ( .B1(n16452), .B2(n16500), .A(n16451), .ZN(P2_U3030) );
  NOR2_X1 U19808 ( .A1(n16453), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16462) );
  INV_X1 U19809 ( .A(n16454), .ZN(n16457) );
  NOR2_X1 U19810 ( .A1(n16306), .A2(n19856), .ZN(n16456) );
  NOR2_X1 U19811 ( .A1(n17070), .A2(n19723), .ZN(n16455) );
  AOI211_X1 U19812 ( .C1(n16457), .C2(n17086), .A(n16456), .B(n16455), .ZN(
        n16458) );
  OAI21_X1 U19813 ( .B1(n16460), .B2(n16459), .A(n16458), .ZN(n16461) );
  AOI211_X1 U19814 ( .C1(n16463), .C2(n11551), .A(n16462), .B(n16461), .ZN(
        n16464) );
  OAI21_X1 U19815 ( .B1(n16465), .B2(n16500), .A(n16464), .ZN(P2_U3031) );
  NOR2_X1 U19816 ( .A1(n16466), .A2(n16492), .ZN(n17009) );
  INV_X1 U19817 ( .A(n17058), .ZN(n17055) );
  OAI21_X1 U19818 ( .B1(n17009), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16998), .ZN(n17002) );
  OR2_X1 U19819 ( .A1(n16468), .A2(n16467), .ZN(n16471) );
  NOR2_X1 U19820 ( .A1(n16469), .A2(n9824), .ZN(n16470) );
  XNOR2_X1 U19821 ( .A(n16471), .B(n16470), .ZN(n17001) );
  INV_X1 U19822 ( .A(n17001), .ZN(n16481) );
  AOI211_X1 U19823 ( .C1(n16492), .C2(n16478), .A(n17058), .B(n17052), .ZN(
        n16480) );
  INV_X1 U19824 ( .A(n17053), .ZN(n16493) );
  INV_X1 U19825 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20412) );
  NOR2_X1 U19826 ( .A1(n20412), .A2(n19856), .ZN(n16476) );
  OR2_X1 U19827 ( .A1(n16473), .A2(n16472), .ZN(n16474) );
  NAND2_X1 U19828 ( .A1(n16474), .A2(n17079), .ZN(n19734) );
  NOR2_X1 U19829 ( .A1(n17070), .A2(n19734), .ZN(n16475) );
  AOI211_X1 U19830 ( .C1(n19637), .C2(n17086), .A(n16476), .B(n16475), .ZN(
        n16477) );
  OAI21_X1 U19831 ( .B1(n16493), .B2(n16478), .A(n16477), .ZN(n16479) );
  AOI211_X1 U19832 ( .C1(n16481), .C2(n19866), .A(n16480), .B(n16479), .ZN(
        n16482) );
  OAI21_X1 U19833 ( .B1(n19859), .B2(n17002), .A(n16482), .ZN(P2_U3035) );
  NAND2_X1 U19834 ( .A1(n16483), .A2(n16504), .ZN(n16488) );
  INV_X1 U19835 ( .A(n16484), .ZN(n16486) );
  NAND2_X1 U19836 ( .A1(n16486), .A2(n16485), .ZN(n16487) );
  XNOR2_X1 U19837 ( .A(n16488), .B(n16487), .ZN(n17010) );
  INV_X1 U19838 ( .A(n17010), .ZN(n16501) );
  INV_X1 U19839 ( .A(n17009), .ZN(n16489) );
  NAND2_X1 U19840 ( .A1(n16466), .A2(n16492), .ZN(n17007) );
  NAND3_X1 U19841 ( .A1(n16489), .A2(n11551), .A3(n17007), .ZN(n16499) );
  INV_X1 U19842 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20411) );
  NOR2_X1 U19843 ( .A1(n20411), .A2(n19856), .ZN(n16490) );
  AOI21_X1 U19844 ( .B1(n17086), .B2(n19646), .A(n16490), .ZN(n16491) );
  OAI21_X1 U19845 ( .B1(n16493), .B2(n16492), .A(n16491), .ZN(n16497) );
  XNOR2_X1 U19846 ( .A(n16495), .B(n16494), .ZN(n19736) );
  NOR2_X1 U19847 ( .A1(n19736), .A2(n17070), .ZN(n16496) );
  AOI211_X1 U19848 ( .C1(n16492), .C2(n17057), .A(n16497), .B(n16496), .ZN(
        n16498) );
  OAI211_X1 U19849 ( .C1(n16501), .C2(n16500), .A(n16499), .B(n16498), .ZN(
        P2_U3036) );
  OAI21_X1 U19850 ( .B1(n16502), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16466), .ZN(n17017) );
  INV_X1 U19851 ( .A(n16504), .ZN(n16505) );
  OR2_X1 U19852 ( .A1(n16506), .A2(n16505), .ZN(n16507) );
  XNOR2_X1 U19853 ( .A(n16503), .B(n16507), .ZN(n17016) );
  INV_X1 U19854 ( .A(n17016), .ZN(n16518) );
  INV_X1 U19855 ( .A(n16508), .ZN(n16515) );
  INV_X1 U19856 ( .A(n17019), .ZN(n16513) );
  NOR2_X1 U19857 ( .A1(n20409), .A2(n19856), .ZN(n16511) );
  NOR2_X1 U19858 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16509), .ZN(
        n16510) );
  NOR2_X1 U19859 ( .A1(n16511), .A2(n16510), .ZN(n16512) );
  OAI21_X1 U19860 ( .B1(n19870), .B2(n16513), .A(n16512), .ZN(n16514) );
  AOI21_X1 U19861 ( .B1(n16515), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16514), .ZN(n16516) );
  OAI21_X1 U19862 ( .B1(n19738), .B2(n17070), .A(n16516), .ZN(n16517) );
  AOI21_X1 U19863 ( .B1(n16518), .B2(n19866), .A(n16517), .ZN(n16519) );
  OAI21_X1 U19864 ( .B1(n17017), .B2(n19859), .A(n16519), .ZN(P2_U3037) );
  NOR2_X1 U19865 ( .A1(n16520), .A2(n21108), .ZN(n16521) );
  AOI211_X1 U19866 ( .C1(n11551), .C2(n16523), .A(n16522), .B(n16521), .ZN(
        n16528) );
  AOI22_X1 U19867 ( .A1(n19866), .A2(n16524), .B1(n19854), .B2(n20474), .ZN(
        n16527) );
  NAND2_X1 U19868 ( .A1(n17086), .A2(n9706), .ZN(n16526) );
  OAI211_X1 U19869 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n17054), .B(n19852), .ZN(n16525) );
  NAND4_X1 U19870 ( .A1(n16528), .A2(n16527), .A3(n16526), .A4(n16525), .ZN(
        P2_U3045) );
  AOI22_X1 U19871 ( .A1(n19656), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n16529), .B2(n14277), .ZN(n16538) );
  NAND2_X1 U19872 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n16538), .ZN(n16532) );
  NAND2_X1 U19873 ( .A1(n16530), .A2(n16547), .ZN(n16531) );
  OAI211_X1 U19874 ( .C1(n16533), .C2(n16552), .A(n16532), .B(n16531), .ZN(
        n16534) );
  MUX2_X1 U19875 ( .A(n16534), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n16553), .Z(P2_U3601) );
  OAI21_X1 U19876 ( .B1(n16537), .B2(n16536), .A(n16535), .ZN(n19705) );
  OAI21_X1 U19877 ( .B1(n14277), .B2(n21108), .A(n19705), .ZN(n16545) );
  NOR2_X1 U19878 ( .A1(n16538), .A2(n11007), .ZN(n16546) );
  INV_X1 U19879 ( .A(n16546), .ZN(n16539) );
  OAI22_X1 U19880 ( .A1(n16540), .A2(n20455), .B1(n16545), .B2(n16539), .ZN(
        n16541) );
  AOI21_X1 U19881 ( .B1(n20478), .B2(n16542), .A(n16541), .ZN(n16544) );
  NAND2_X1 U19882 ( .A1(n16553), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16543) );
  OAI21_X1 U19883 ( .B1(n16553), .B2(n16544), .A(n16543), .ZN(P2_U3600) );
  AOI22_X1 U19884 ( .A1(n16548), .A2(n16547), .B1(n16546), .B2(n16545), .ZN(
        n16549) );
  OAI21_X1 U19885 ( .B1(n20466), .B2(n16552), .A(n16549), .ZN(n16550) );
  MUX2_X1 U19886 ( .A(n16550), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n16553), .Z(P2_U3599) );
  OAI22_X1 U19887 ( .A1(n19749), .A2(n16552), .B1(n20455), .B2(n16551), .ZN(
        n16554) );
  MUX2_X1 U19888 ( .A(n16554), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16553), .Z(P2_U3596) );
  NAND2_X1 U19889 ( .A1(n17916), .A2(n17808), .ZN(n17811) );
  AOI22_X1 U19890 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17855), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16567) );
  AOI22_X1 U19891 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16566) );
  AOI22_X1 U19892 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16557) );
  OAI21_X1 U19893 ( .B1(n16558), .B2(n21193), .A(n16557), .ZN(n16564) );
  AOI22_X1 U19894 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16562) );
  AOI22_X1 U19895 ( .A1(n17857), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16561) );
  AOI22_X1 U19896 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16560) );
  AOI22_X1 U19897 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16559) );
  NAND4_X1 U19898 ( .A1(n16562), .A2(n16561), .A3(n16560), .A4(n16559), .ZN(
        n16563) );
  AOI211_X1 U19899 ( .C1(n17880), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n16564), .B(n16563), .ZN(n16565) );
  NAND3_X1 U19900 ( .A1(n16567), .A2(n16566), .A3(n16565), .ZN(n18015) );
  NAND2_X1 U19901 ( .A1(n17921), .A2(n18015), .ZN(n16568) );
  OAI221_X1 U19902 ( .B1(n17811), .B2(n17454), .C1(n17811), .C2(n9784), .A(
        n16568), .ZN(P3_U2690) );
  NOR2_X1 U19903 ( .A1(n19492), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18934) );
  NOR3_X1 U19904 ( .A1(n19503), .A2(n17110), .A3(n19393), .ZN(n16570) );
  AOI211_X1 U19905 ( .C1(n16586), .C2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n17826), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16569) );
  INV_X1 U19906 ( .A(n16569), .ZN(n18880) );
  NAND2_X1 U19907 ( .A1(n19330), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19382) );
  OAI221_X1 U19908 ( .B1(n19393), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n19503), .A(n19382), .ZN(n18891) );
  INV_X1 U19909 ( .A(n19001), .ZN(n19230) );
  INV_X1 U19910 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18881) );
  INV_X1 U19911 ( .A(n16570), .ZN(n19490) );
  NOR2_X1 U19912 ( .A1(n18881), .A2(n19490), .ZN(n16585) );
  AOI211_X1 U19913 ( .C1(n16570), .C2(n18880), .A(n19230), .B(n16585), .ZN(
        n16571) );
  NOR2_X1 U19914 ( .A1(n18934), .A2(n16571), .ZN(n16573) );
  NAND3_X1 U19915 ( .A1(n19393), .A2(n19492), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19227) );
  INV_X1 U19916 ( .A(n16571), .ZN(n18886) );
  NAND2_X1 U19917 ( .A1(n19393), .A2(n19492), .ZN(n17253) );
  AND2_X1 U19918 ( .A1(n19497), .A2(n17253), .ZN(n19534) );
  NOR2_X1 U19919 ( .A1(n19503), .A2(n19538), .ZN(n18452) );
  NAND2_X1 U19920 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18887) );
  OAI21_X1 U19921 ( .B1(n19534), .B2(n18452), .A(n18887), .ZN(n16576) );
  NAND3_X1 U19922 ( .A1(n19366), .A2(n18886), .A3(n16576), .ZN(n16572) );
  OAI221_X1 U19923 ( .B1(n19366), .B2(n16573), .C1(n19366), .C2(n19227), .A(
        n16572), .ZN(P3_U2864) );
  NAND2_X1 U19924 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19047) );
  NOR2_X1 U19925 ( .A1(n19534), .A2(n18452), .ZN(n16575) );
  INV_X1 U19926 ( .A(n16573), .ZN(n16574) );
  AOI221_X1 U19927 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19047), .C1(n16575), 
        .C2(n19047), .A(n16574), .ZN(n18885) );
  INV_X1 U19928 ( .A(n19227), .ZN(n16577) );
  OAI221_X1 U19929 ( .B1(n16577), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n16577), .C2(n16576), .A(n18886), .ZN(n18883) );
  AOI22_X1 U19930 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18885), .B1(
        n18883), .B2(n19371), .ZN(P3_U2865) );
  NAND2_X1 U19931 ( .A1(n19324), .A2(n19540), .ZN(n16584) );
  INV_X1 U19932 ( .A(n19537), .ZN(n16578) );
  NAND2_X1 U19933 ( .A1(n16579), .A2(n16578), .ZN(n18072) );
  NOR2_X1 U19934 ( .A1(n16581), .A2(n16580), .ZN(n16583) );
  OAI211_X1 U19935 ( .C1(n16584), .C2(n18072), .A(n16583), .B(n16679), .ZN(
        n19357) );
  NOR2_X1 U19936 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19492), .ZN(n18892) );
  AOI211_X1 U19937 ( .C1(n19535), .C2(n19357), .A(n18892), .B(n16585), .ZN(
        n19523) );
  INV_X1 U19938 ( .A(n19523), .ZN(n19520) );
  INV_X1 U19939 ( .A(n19497), .ZN(n19518) );
  AOI21_X1 U19940 ( .B1(n16586), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16588) );
  INV_X1 U19941 ( .A(n19349), .ZN(n16587) );
  NOR2_X1 U19942 ( .A1(n16588), .A2(n16587), .ZN(n19381) );
  NAND3_X1 U19943 ( .A1(n19520), .A2(n19518), .A3(n19381), .ZN(n16589) );
  OAI21_X1 U19944 ( .B1(n19520), .B2(n19330), .A(n16589), .ZN(P3_U3284) );
  INV_X1 U19945 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17141) );
  NAND2_X1 U19946 ( .A1(n17116), .A2(n18868), .ZN(n18792) );
  NOR2_X1 U19947 ( .A1(n17142), .A2(n17141), .ZN(n17133) );
  INV_X1 U19948 ( .A(n18572), .ZN(n16598) );
  NAND2_X1 U19949 ( .A1(n17133), .A2(n16598), .ZN(n17134) );
  NOR2_X1 U19950 ( .A1(n18601), .A2(n18871), .ZN(n18864) );
  AOI21_X1 U19951 ( .B1(n18570), .B2(n17133), .A(n18878), .ZN(n16590) );
  AOI21_X1 U19952 ( .B1(n18725), .B2(n17134), .A(n16590), .ZN(n16661) );
  INV_X1 U19953 ( .A(n18783), .ZN(n18690) );
  OAI221_X1 U19954 ( .B1(n16592), .B2(n18690), .C1(n16592), .C2(n16591), .A(
        n18833), .ZN(n16601) );
  INV_X1 U19955 ( .A(n16593), .ZN(n16594) );
  OAI21_X1 U19956 ( .B1(n16595), .B2(n16658), .A(n16594), .ZN(n16596) );
  NOR2_X1 U19957 ( .A1(n17141), .A2(n16596), .ZN(n17120) );
  AOI21_X1 U19958 ( .B1(n17141), .B2(n16596), .A(n17120), .ZN(n17145) );
  NOR2_X1 U19959 ( .A1(n18833), .A2(n19475), .ZN(n17138) );
  NAND3_X1 U19960 ( .A1(n18854), .A2(n17125), .A3(n18586), .ZN(n17154) );
  OAI21_X1 U19961 ( .B1(n18878), .B2(n18195), .A(n17154), .ZN(n16597) );
  AOI21_X1 U19962 ( .B1(n16598), .B2(n18725), .A(n16597), .ZN(n16664) );
  NOR3_X1 U19963 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16664), .A3(
        n17142), .ZN(n16599) );
  AOI211_X1 U19964 ( .C1(n18788), .C2(n17145), .A(n17138), .B(n16599), .ZN(
        n16600) );
  OAI221_X1 U19965 ( .B1(n17141), .B2(n16661), .C1(n17141), .C2(n16601), .A(
        n16600), .ZN(P3_U2833) );
  AOI22_X1 U19966 ( .A1(n16603), .A2(n19698), .B1(n16602), .B2(n19671), .ZN(
        n16613) );
  AOI211_X1 U19967 ( .C1(n16606), .C2(n16605), .A(n16604), .B(n19704), .ZN(
        n16611) );
  INV_X1 U19968 ( .A(n16607), .ZN(n16609) );
  AOI22_X1 U19969 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19697), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19672), .ZN(n16608) );
  OAI21_X1 U19970 ( .B1(n16609), .B2(n19692), .A(n16608), .ZN(n16610) );
  AOI211_X1 U19971 ( .C1(P2_EBX_REG_22__SCAN_IN), .C2(n19678), .A(n16611), .B(
        n16610), .ZN(n16612) );
  NAND2_X1 U19972 ( .A1(n16613), .A2(n16612), .ZN(P2_U2833) );
  INV_X1 U19973 ( .A(n16614), .ZN(n16615) );
  NOR2_X1 U19974 ( .A1(n16615), .A2(n16642), .ZN(n16650) );
  INV_X1 U19975 ( .A(n16623), .ZN(n16625) );
  NAND2_X1 U19976 ( .A1(n16617), .A2(n16616), .ZN(n16619) );
  NAND2_X1 U19977 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16619), .ZN(
        n16621) );
  OAI211_X1 U19978 ( .C1(n16619), .C2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16618), .ZN(n16620) );
  OAI211_X1 U19979 ( .C1(n16623), .C2(n16622), .A(n16621), .B(n16620), .ZN(
        n16624) );
  OAI21_X1 U19980 ( .B1(n16625), .B2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16624), .ZN(n16626) );
  AOI222_X1 U19981 ( .A1(n16627), .A2(n16626), .B1(n16627), .B2(n20737), .C1(
        n16626), .C2(n20737), .ZN(n16635) );
  INV_X1 U19982 ( .A(n16628), .ZN(n16630) );
  NOR3_X1 U19983 ( .A1(n16631), .A2(n16630), .A3(n16629), .ZN(n16634) );
  OAI21_X1 U19984 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n16632), .ZN(n16633) );
  OAI211_X1 U19985 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n16635), .A(
        n16634), .B(n16633), .ZN(n16645) );
  INV_X1 U19986 ( .A(n16645), .ZN(n16641) );
  NOR2_X1 U19987 ( .A1(n16636), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21032) );
  OR2_X1 U19988 ( .A1(n16637), .A2(n21028), .ZN(n16638) );
  AOI22_X1 U19989 ( .A1(n16640), .A2(n21032), .B1(n16639), .B2(n16638), .ZN(
        n16877) );
  OAI221_X1 U19990 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n16641), 
        .A(n16877), .ZN(n16884) );
  NAND2_X1 U19991 ( .A1(n16884), .A2(n9922), .ZN(n16649) );
  OAI211_X1 U19992 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21028), .A(n16643), 
        .B(n16642), .ZN(n16644) );
  AOI21_X1 U19993 ( .B1(n16646), .B2(n16645), .A(n16644), .ZN(n16647) );
  AND2_X1 U19994 ( .A1(n16884), .A2(n16647), .ZN(n16648) );
  OAI22_X1 U19995 ( .A1(n16650), .A2(n16649), .B1(n16648), .B2(n9922), .ZN(
        P1_U3161) );
  INV_X1 U19996 ( .A(n16651), .ZN(n16655) );
  NAND2_X1 U19997 ( .A1(n16776), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16653) );
  OAI211_X1 U19998 ( .C1(n16783), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16653), .B(n16652), .ZN(n16654) );
  AOI21_X1 U19999 ( .B1(n16655), .B2(n16861), .A(n16654), .ZN(n16656) );
  OAI21_X1 U20000 ( .B1(n20652), .B2(n16657), .A(n16656), .ZN(P1_U3010) );
  INV_X1 U20001 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17117) );
  NAND2_X1 U20002 ( .A1(n17133), .A2(n17117), .ZN(n17137) );
  AOI21_X1 U20003 ( .B1(n16658), .B2(n17141), .A(n18463), .ZN(n17121) );
  OAI211_X1 U20004 ( .C1(n18783), .C2(n17133), .A(n18854), .B(n16659), .ZN(
        n16660) );
  NAND2_X1 U20005 ( .A1(n18833), .A2(n16660), .ZN(n17156) );
  AOI21_X1 U20006 ( .B1(n16661), .B2(n17156), .A(n17117), .ZN(n16662) );
  AOI21_X1 U20007 ( .B1(n18788), .B2(n17132), .A(n16662), .ZN(n16663) );
  NAND2_X1 U20008 ( .A1(n18869), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17127) );
  OAI211_X1 U20009 ( .C1(n16664), .C2(n17137), .A(n16663), .B(n17127), .ZN(
        P3_U2832) );
  INV_X1 U20010 ( .A(HOLD), .ZN(n20938) );
  NOR2_X1 U20011 ( .A1(n20951), .A2(n20938), .ZN(n20940) );
  AOI22_X1 U20012 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n16667) );
  NAND2_X1 U20013 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20943), .ZN(n16665) );
  OAI211_X1 U20014 ( .C1(n20940), .C2(n16667), .A(n16666), .B(n16665), .ZN(
        P1_U3195) );
  AOI22_X1 U20015 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16784), .B1(
        n13116), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n16675) );
  INV_X1 U20016 ( .A(n16668), .ZN(n16671) );
  INV_X1 U20017 ( .A(n16669), .ZN(n16670) );
  AOI22_X1 U20018 ( .A1(n16671), .A2(n16861), .B1(n16857), .B2(n16670), .ZN(
        n16674) );
  OAI211_X1 U20019 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16787), .B(n16672), .ZN(
        n16673) );
  NAND3_X1 U20020 ( .A1(n16675), .A2(n16674), .A3(n16673), .ZN(P1_U3011) );
  NOR3_X1 U20021 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16677) );
  NOR2_X1 U20022 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16676) );
  NOR4_X1 U20023 ( .A1(n16677), .A2(n16676), .A3(n17093), .A4(n17094), .ZN(
        P2_U3178) );
  INV_X1 U20024 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n19564) );
  OAI221_X1 U20025 ( .B1(n19564), .B2(n16678), .C1(n20502), .C2(n16678), .A(
        n20074), .ZN(n20491) );
  NOR2_X1 U20026 ( .A1(n21126), .A2(n20491), .ZN(P2_U3047) );
  NAND2_X1 U20027 ( .A1(n18929), .A2(n9913), .ZN(n18064) );
  INV_X1 U20028 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18150) );
  AOI22_X1 U20029 ( .A1(n18068), .A2(BUF2_REG_0__SCAN_IN), .B1(n18067), .B2(
        n16683), .ZN(n16684) );
  OAI221_X1 U20030 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n18064), .C1(n18150), 
        .C2(n9913), .A(n16684), .ZN(P3_U2735) );
  AOI22_X1 U20031 ( .A1(n16685), .A2(n20604), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n20602), .ZN(n16687) );
  NAND2_X1 U20032 ( .A1(n20593), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16686) );
  NAND3_X1 U20033 ( .A1(n16687), .A2(n16808), .A3(n16686), .ZN(n16688) );
  AOI21_X1 U20034 ( .B1(n16689), .B2(n20554), .A(n16688), .ZN(n16693) );
  OAI21_X1 U20035 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n16691), .A(n16690), 
        .ZN(n16692) );
  OAI211_X1 U20036 ( .C1(n16799), .C2(n20580), .A(n16693), .B(n16692), .ZN(
        P1_U2823) );
  OAI21_X1 U20037 ( .B1(n16706), .B2(n20565), .A(n16694), .ZN(n16695) );
  INV_X1 U20038 ( .A(n16695), .ZN(n16716) );
  AOI21_X1 U20039 ( .B1(n20596), .B2(n20972), .A(n16716), .ZN(n16703) );
  AOI22_X1 U20040 ( .A1(n16696), .A2(n20604), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n20602), .ZN(n16697) );
  OAI21_X1 U20041 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n16698), .A(n16697), 
        .ZN(n16699) );
  AOI211_X1 U20042 ( .C1(n20593), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n13116), .B(n16699), .ZN(n16702) );
  NOR2_X1 U20043 ( .A1(n16731), .A2(n20580), .ZN(n16700) );
  AOI21_X1 U20044 ( .B1(n16733), .B2(n20554), .A(n16700), .ZN(n16701) );
  OAI211_X1 U20045 ( .C1(n16703), .C2(n15748), .A(n16702), .B(n16701), .ZN(
        P1_U2824) );
  OAI21_X1 U20046 ( .B1(n20581), .B2(n16704), .A(n16808), .ZN(n16709) );
  NAND2_X1 U20047 ( .A1(n20596), .A2(n20972), .ZN(n16705) );
  OAI22_X1 U20048 ( .A1(n16707), .A2(n20592), .B1(n16706), .B2(n16705), .ZN(
        n16708) );
  AOI211_X1 U20049 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n16716), .A(n16709), 
        .B(n16708), .ZN(n16714) );
  INV_X1 U20050 ( .A(n16710), .ZN(n16711) );
  AOI22_X1 U20051 ( .A1(n16712), .A2(n20554), .B1(n20604), .B2(n16711), .ZN(
        n16713) );
  OAI211_X1 U20052 ( .C1(n20580), .C2(n16801), .A(n16714), .B(n16713), .ZN(
        P1_U2825) );
  AOI22_X1 U20053 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20593), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(n20602), .ZN(n16721) );
  AOI21_X1 U20054 ( .B1(n16715), .B2(n20595), .A(n13116), .ZN(n16720) );
  AOI22_X1 U20055 ( .A1(n16736), .A2(n20554), .B1(n20604), .B2(n16735), .ZN(
        n16719) );
  OAI221_X1 U20056 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(P1_REIP_REG_13__SCAN_IN), .C1(P1_REIP_REG_14__SCAN_IN), .C2(n16717), .A(n16716), .ZN(n16718) );
  NAND4_X1 U20057 ( .A1(n16721), .A2(n16720), .A3(n16719), .A4(n16718), .ZN(
        P1_U2826) );
  OAI22_X1 U20058 ( .A1(n16755), .A2(n20583), .B1(n20580), .B2(n16821), .ZN(
        n16722) );
  AOI211_X1 U20059 ( .C1(n20593), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n13116), .B(n16722), .ZN(n16723) );
  OAI21_X1 U20060 ( .B1(n16724), .B2(n20592), .A(n16723), .ZN(n16725) );
  AOI21_X1 U20061 ( .B1(n16752), .B2(n20554), .A(n16725), .ZN(n16726) );
  OAI221_X1 U20062 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16729), .C1(n16728), 
        .C2(n16727), .A(n16726), .ZN(P1_U2829) );
  INV_X1 U20063 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21109) );
  NOR2_X1 U20064 ( .A1(n16731), .A2(n16730), .ZN(n16732) );
  AOI21_X1 U20065 ( .B1(n16733), .B2(n21042), .A(n16732), .ZN(n16734) );
  OAI21_X1 U20066 ( .B1(n20618), .B2(n21109), .A(n16734), .ZN(P1_U2856) );
  AOI22_X1 U20067 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16738) );
  AOI22_X1 U20068 ( .A1(n16736), .A2(n16764), .B1(n16742), .B2(n16735), .ZN(
        n16737) );
  OAI211_X1 U20069 ( .C1(n16739), .C2(n20516), .A(n16738), .B(n16737), .ZN(
        P1_U2985) );
  AOI22_X1 U20070 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16745) );
  INV_X1 U20071 ( .A(n16740), .ZN(n16743) );
  AOI22_X1 U20072 ( .A1(n16743), .A2(n16764), .B1(n16742), .B2(n16741), .ZN(
        n16744) );
  OAI211_X1 U20073 ( .C1(n16746), .C2(n20516), .A(n16745), .B(n16744), .ZN(
        P1_U2987) );
  AOI22_X1 U20074 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16754) );
  NAND3_X1 U20075 ( .A1(n16747), .A2(n9714), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16749) );
  NAND2_X1 U20076 ( .A1(n16749), .A2(n16748), .ZN(n16751) );
  XNOR2_X1 U20077 ( .A(n16751), .B(n16750), .ZN(n16818) );
  AOI22_X1 U20078 ( .A1(n16818), .A2(n16772), .B1(n16764), .B2(n16752), .ZN(
        n16753) );
  OAI211_X1 U20079 ( .C1(n16769), .C2(n16755), .A(n16754), .B(n16753), .ZN(
        P1_U2988) );
  AOI22_X1 U20080 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16758) );
  AOI22_X1 U20081 ( .A1(n16756), .A2(n16772), .B1(n16764), .B2(n20547), .ZN(
        n16757) );
  OAI211_X1 U20082 ( .C1(n16769), .C2(n20545), .A(n16758), .B(n16757), .ZN(
        P1_U2992) );
  AOI22_X1 U20083 ( .A1(n16759), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n13116), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16766) );
  NAND2_X1 U20084 ( .A1(n16762), .A2(n16761), .ZN(n16763) );
  XNOR2_X1 U20085 ( .A(n16760), .B(n16763), .ZN(n16862) );
  AOI22_X1 U20086 ( .A1(n16862), .A2(n16772), .B1(n16764), .B2(n20611), .ZN(
        n16765) );
  OAI211_X1 U20087 ( .C1(n16769), .C2(n20551), .A(n16766), .B(n16765), .ZN(
        P1_U2993) );
  XOR2_X1 U20088 ( .A(n16767), .B(n16768), .Z(n16866) );
  OAI22_X1 U20089 ( .A1(n20568), .A2(n16770), .B1(n20572), .B2(n16769), .ZN(
        n16771) );
  AOI21_X1 U20090 ( .B1(n16866), .B2(n16772), .A(n16771), .ZN(n16773) );
  NAND2_X1 U20091 ( .A1(n13116), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16873) );
  OAI211_X1 U20092 ( .C1(n20559), .C2(n16774), .A(n16773), .B(n16873), .ZN(
        P1_U2994) );
  OAI21_X1 U20093 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16775), .ZN(n16782) );
  AOI22_X1 U20094 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16776), .B1(
        n13116), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16781) );
  INV_X1 U20095 ( .A(n16777), .ZN(n16779) );
  AOI22_X1 U20096 ( .A1(n16779), .A2(n16861), .B1(n16857), .B2(n16778), .ZN(
        n16780) );
  OAI211_X1 U20097 ( .C1(n16783), .C2(n16782), .A(n16781), .B(n16780), .ZN(
        P1_U3009) );
  AOI22_X1 U20098 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16784), .B1(
        n13116), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16790) );
  INV_X1 U20099 ( .A(n16785), .ZN(n16788) );
  AOI22_X1 U20100 ( .A1(n16788), .A2(n16861), .B1(n16787), .B2(n16786), .ZN(
        n16789) );
  OAI211_X1 U20101 ( .C1(n20652), .C2(n16791), .A(n16790), .B(n16789), .ZN(
        P1_U3012) );
  OAI21_X1 U20102 ( .B1(n16806), .B2(n16793), .A(n16792), .ZN(n16794) );
  AOI22_X1 U20103 ( .A1(n16796), .A2(n16861), .B1(n16795), .B2(n16794), .ZN(
        n16798) );
  NAND2_X1 U20104 ( .A1(n13116), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16797) );
  OAI211_X1 U20105 ( .C1(n20652), .C2(n16799), .A(n16798), .B(n16797), .ZN(
        P1_U3014) );
  OAI222_X1 U20106 ( .A1(n16801), .A2(n20652), .B1(n16808), .B2(n20972), .C1(
        n20653), .C2(n16800), .ZN(n16802) );
  INV_X1 U20107 ( .A(n16802), .ZN(n16803) );
  OAI221_X1 U20108 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16806), 
        .C1(n16805), .C2(n16804), .A(n16803), .ZN(P1_U3016) );
  OAI222_X1 U20109 ( .A1(n16809), .A2(n20652), .B1(n16808), .B2(n20970), .C1(
        n20653), .C2(n16807), .ZN(n16810) );
  INV_X1 U20110 ( .A(n16810), .ZN(n16812) );
  OAI211_X1 U20111 ( .C1(n16814), .C2(n16813), .A(n16812), .B(n16811), .ZN(
        P1_U3018) );
  OAI22_X1 U20112 ( .A1(n16816), .A2(n16750), .B1(n16859), .B2(n16815), .ZN(
        n16817) );
  AOI21_X1 U20113 ( .B1(n16818), .B2(n16861), .A(n16817), .ZN(n16820) );
  NAND2_X1 U20114 ( .A1(n13116), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n16819) );
  OAI211_X1 U20115 ( .C1(n20652), .C2(n16821), .A(n16820), .B(n16819), .ZN(
        P1_U3020) );
  NAND2_X1 U20116 ( .A1(n16823), .A2(n16822), .ZN(n16825) );
  OAI21_X1 U20117 ( .B1(n16836), .B2(n16825), .A(n16824), .ZN(n16837) );
  AOI22_X1 U20118 ( .A1(n13116), .A2(P1_REIP_REG_10__SCAN_IN), .B1(n16857), 
        .B2(n16826), .ZN(n16831) );
  NAND2_X1 U20119 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16828) );
  AOI211_X1 U20120 ( .C1(n15781), .C2(n16840), .A(n16836), .B(n16859), .ZN(
        n16827) );
  AOI22_X1 U20121 ( .A1(n16829), .A2(n16861), .B1(n16828), .B2(n16827), .ZN(
        n16830) );
  OAI211_X1 U20122 ( .C1(n15781), .C2(n16837), .A(n16831), .B(n16830), .ZN(
        P1_U3021) );
  NAND2_X1 U20123 ( .A1(n16833), .A2(n16832), .ZN(n16834) );
  AND2_X1 U20124 ( .A1(n16835), .A2(n16834), .ZN(n21039) );
  INV_X1 U20125 ( .A(n21039), .ZN(n16844) );
  NOR2_X1 U20126 ( .A1(n16836), .A2(n16859), .ZN(n16841) );
  OAI22_X1 U20127 ( .A1(n16838), .A2(n20653), .B1(n16837), .B2(n16840), .ZN(
        n16839) );
  AOI21_X1 U20128 ( .B1(n16841), .B2(n16840), .A(n16839), .ZN(n16843) );
  NAND2_X1 U20129 ( .A1(n13116), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n16842) );
  OAI211_X1 U20130 ( .C1(n20652), .C2(n16844), .A(n16843), .B(n16842), .ZN(
        P1_U3022) );
  AOI22_X1 U20131 ( .A1(n13116), .A2(P1_REIP_REG_8__SCAN_IN), .B1(n16857), 
        .B2(n16845), .ZN(n16852) );
  AOI22_X1 U20132 ( .A1(n16847), .A2(n16861), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16846), .ZN(n16851) );
  OAI221_X1 U20133 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16849), .C2(n14523), .A(
        n16848), .ZN(n16850) );
  NAND3_X1 U20134 ( .A1(n16852), .A2(n16851), .A3(n16850), .ZN(P1_U3023) );
  NOR2_X1 U20135 ( .A1(n16854), .A2(n16853), .ZN(n16855) );
  AOI22_X1 U20136 ( .A1(n13116), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n16857), 
        .B2(n9813), .ZN(n16864) );
  INV_X1 U20137 ( .A(n16859), .ZN(n16860) );
  AOI22_X1 U20138 ( .A1(n16862), .A2(n16861), .B1(n16860), .B2(n21163), .ZN(
        n16863) );
  OAI211_X1 U20139 ( .C1(n16865), .C2(n21163), .A(n16864), .B(n16863), .ZN(
        P1_U3025) );
  INV_X1 U20140 ( .A(n16866), .ZN(n16869) );
  OAI22_X1 U20141 ( .A1(n16869), .A2(n20653), .B1(n16868), .B2(n16867), .ZN(
        n16870) );
  AOI21_X1 U20142 ( .B1(n16872), .B2(n16871), .A(n16870), .ZN(n16874) );
  OAI211_X1 U20143 ( .C1(n20652), .C2(n20560), .A(n16874), .B(n16873), .ZN(
        P1_U3026) );
  AOI21_X1 U20144 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16884), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16882) );
  NAND4_X1 U20145 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n14046), .A4(n21028), .ZN(n16875) );
  AND2_X1 U20146 ( .A1(n16876), .A2(n16875), .ZN(n20934) );
  AOI21_X1 U20147 ( .B1(n20934), .B2(n16878), .A(n16877), .ZN(n16881) );
  AOI21_X1 U20148 ( .B1(n12826), .B2(n21028), .A(n16879), .ZN(n16880) );
  NOR3_X1 U20149 ( .A1(n16882), .A2(n16881), .A3(n16880), .ZN(P1_U3162) );
  OAI221_X1 U20150 ( .B1(n12826), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n12826), 
        .C2(n16884), .A(n16883), .ZN(P1_U3466) );
  INV_X1 U20151 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n16888) );
  INV_X1 U20152 ( .A(n16885), .ZN(n16887) );
  OAI222_X1 U20153 ( .A1(n19676), .A2(n16888), .B1(n19692), .B2(n16887), .C1(
        n16886), .C2(n16952), .ZN(n16889) );
  AOI21_X1 U20154 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19672), .A(
        n16889), .ZN(n16892) );
  OAI211_X1 U20155 ( .C1(n16953), .C2(n19687), .A(n16892), .B(n16891), .ZN(
        P2_U2824) );
  AOI22_X1 U20156 ( .A1(n16893), .A2(n19679), .B1(P2_REIP_REG_29__SCAN_IN), 
        .B2(n19697), .ZN(n16904) );
  AOI22_X1 U20157 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19678), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19672), .ZN(n16903) );
  INV_X1 U20158 ( .A(n16894), .ZN(n16896) );
  AOI22_X1 U20159 ( .A1(n16896), .A2(n19698), .B1(n19671), .B2(n16895), .ZN(
        n16902) );
  AOI21_X1 U20160 ( .B1(n16899), .B2(n16898), .A(n16897), .ZN(n16900) );
  NAND2_X1 U20161 ( .A1(n19684), .A2(n16900), .ZN(n16901) );
  NAND4_X1 U20162 ( .A1(n16904), .A2(n16903), .A3(n16902), .A4(n16901), .ZN(
        P2_U2826) );
  INV_X1 U20163 ( .A(n16905), .ZN(n16906) );
  AOI22_X1 U20164 ( .A1(n16907), .A2(n19698), .B1(n16906), .B2(n19671), .ZN(
        n16916) );
  AOI211_X1 U20165 ( .C1(n16910), .C2(n16909), .A(n16908), .B(n19704), .ZN(
        n16914) );
  AOI22_X1 U20166 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n19697), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19672), .ZN(n16911) );
  OAI21_X1 U20167 ( .B1(n16912), .B2(n19692), .A(n16911), .ZN(n16913) );
  AOI211_X1 U20168 ( .C1(P2_EBX_REG_28__SCAN_IN), .C2(n19678), .A(n16914), .B(
        n16913), .ZN(n16915) );
  NAND2_X1 U20169 ( .A1(n16916), .A2(n16915), .ZN(P2_U2827) );
  OAI22_X1 U20170 ( .A1(n16918), .A2(n19687), .B1(n16917), .B2(n19703), .ZN(
        n16919) );
  INV_X1 U20171 ( .A(n16919), .ZN(n16928) );
  AOI211_X1 U20172 ( .C1(n16922), .C2(n16921), .A(n16920), .B(n19704), .ZN(
        n16926) );
  AOI22_X1 U20173 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19672), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19697), .ZN(n16923) );
  OAI21_X1 U20174 ( .B1(n16924), .B2(n19692), .A(n16923), .ZN(n16925) );
  AOI211_X1 U20175 ( .C1(P2_EBX_REG_27__SCAN_IN), .C2(n19678), .A(n16926), .B(
        n16925), .ZN(n16927) );
  NAND2_X1 U20176 ( .A1(n16928), .A2(n16927), .ZN(P2_U2828) );
  INV_X1 U20177 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n21294) );
  OAI22_X1 U20178 ( .A1(n16929), .A2(n19692), .B1(n21294), .B2(n19676), .ZN(
        n16930) );
  INV_X1 U20179 ( .A(n16930), .ZN(n16940) );
  AOI22_X1 U20180 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19678), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19672), .ZN(n16939) );
  AOI22_X1 U20181 ( .A1(n16932), .A2(n19698), .B1(n19671), .B2(n16931), .ZN(
        n16938) );
  AOI21_X1 U20182 ( .B1(n16935), .B2(n16934), .A(n16933), .ZN(n16936) );
  NAND2_X1 U20183 ( .A1(n19684), .A2(n16936), .ZN(n16937) );
  NAND4_X1 U20184 ( .A1(n16940), .A2(n16939), .A3(n16938), .A4(n16937), .ZN(
        P2_U2830) );
  AOI22_X1 U20185 ( .A1(n16942), .A2(n19698), .B1(n16941), .B2(n19671), .ZN(
        n16951) );
  AOI211_X1 U20186 ( .C1(n16945), .C2(n16944), .A(n16943), .B(n19704), .ZN(
        n16949) );
  AOI22_X1 U20187 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19672), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19697), .ZN(n16946) );
  OAI21_X1 U20188 ( .B1(n16947), .B2(n19692), .A(n16946), .ZN(n16948) );
  AOI211_X1 U20189 ( .C1(P2_EBX_REG_23__SCAN_IN), .C2(n19678), .A(n16949), .B(
        n16948), .ZN(n16950) );
  NAND2_X1 U20190 ( .A1(n16951), .A2(n16950), .ZN(P2_U2832) );
  AOI22_X1 U20191 ( .A1(n19712), .A2(n16953), .B1(n16952), .B2(n19716), .ZN(
        P2_U2856) );
  NOR2_X1 U20192 ( .A1(n16955), .A2(n14265), .ZN(n16956) );
  XNOR2_X1 U20193 ( .A(n16957), .B(n16956), .ZN(n16958) );
  XNOR2_X1 U20194 ( .A(n16954), .B(n16958), .ZN(n16975) );
  AOI22_X1 U20195 ( .A1(n16975), .A2(n16970), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n19716), .ZN(n16959) );
  OAI21_X1 U20196 ( .B1(n19716), .B2(n16960), .A(n16959), .ZN(P2_U2863) );
  NOR2_X1 U20197 ( .A1(n16961), .A2(n19716), .ZN(n16962) );
  AOI21_X1 U20198 ( .B1(n16963), .B2(n16970), .A(n16962), .ZN(n16964) );
  OAI21_X1 U20199 ( .B1(n19712), .B2(n11106), .A(n16964), .ZN(P2_U2866) );
  OAI22_X1 U20200 ( .A1(n16966), .A2(n19713), .B1(n19716), .B2(n16965), .ZN(
        n16967) );
  INV_X1 U20201 ( .A(n16967), .ZN(n16968) );
  OAI21_X1 U20202 ( .B1(n19712), .B2(n16969), .A(n16968), .ZN(P2_U2868) );
  AOI22_X1 U20203 ( .A1(n16971), .A2(n16970), .B1(n19712), .B2(n10320), .ZN(
        n16972) );
  OAI21_X1 U20204 ( .B1(n19712), .B2(n10876), .A(n16972), .ZN(P2_U2870) );
  AOI22_X1 U20205 ( .A1(n16973), .A2(n19740), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19771), .ZN(n16978) );
  AOI22_X1 U20206 ( .A1(n19719), .A2(BUF1_REG_24__SCAN_IN), .B1(n19717), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U20207 ( .A1(n16975), .A2(n19773), .B1(n19772), .B2(n16974), .ZN(
        n16976) );
  NAND3_X1 U20208 ( .A1(n16978), .A2(n16977), .A3(n16976), .ZN(P2_U2895) );
  AOI22_X1 U20209 ( .A1(n19837), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19825), .ZN(n16984) );
  NAND2_X1 U20210 ( .A1(n16980), .A2(n16979), .ZN(n16981) );
  XNOR2_X1 U20211 ( .A(n9732), .B(n16981), .ZN(n17064) );
  INV_X1 U20212 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17090) );
  AOI21_X1 U20213 ( .B1(n16997), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16982) );
  NOR2_X1 U20214 ( .A1(n16982), .A2(n10311), .ZN(n17063) );
  AOI222_X1 U20215 ( .A1(n17064), .A2(n19828), .B1(n11531), .B2(n17063), .C1(
        n19848), .C2(n17062), .ZN(n16983) );
  OAI211_X1 U20216 ( .C1(n19840), .C2(n19613), .A(n16984), .B(n16983), .ZN(
        P2_U3000) );
  AOI22_X1 U20217 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19825), .B1(n17038), 
        .B2(n16985), .ZN(n16991) );
  NAND2_X1 U20218 ( .A1(n16987), .A2(n16986), .ZN(n16988) );
  XNOR2_X1 U20219 ( .A(n16989), .B(n16988), .ZN(n17074) );
  OAI211_X1 U20220 ( .C1(n17046), .C2(n16992), .A(n16991), .B(n16990), .ZN(
        P2_U3001) );
  AOI22_X1 U20221 ( .A1(n19837), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19825), .ZN(n17000) );
  NOR2_X1 U20222 ( .A1(n16994), .A2(n10076), .ZN(n16995) );
  XNOR2_X1 U20223 ( .A(n16996), .B(n16995), .ZN(n17087) );
  AOI21_X1 U20224 ( .B1(n17090), .B2(n16998), .A(n16997), .ZN(n17084) );
  AOI222_X1 U20225 ( .A1(n17087), .A2(n19828), .B1(n19848), .B2(n17085), .C1(
        n11531), .C2(n17084), .ZN(n16999) );
  OAI211_X1 U20226 ( .C1(n19840), .C2(n19622), .A(n17000), .B(n16999), .ZN(
        P2_U3002) );
  AOI22_X1 U20227 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19825), .B1(n17038), 
        .B2(n19634), .ZN(n17005) );
  OAI22_X1 U20228 ( .A1(n17002), .A2(n17039), .B1(n17001), .B2(n19845), .ZN(
        n17003) );
  AOI21_X1 U20229 ( .B1(n19848), .B2(n19637), .A(n17003), .ZN(n17004) );
  OAI211_X1 U20230 ( .C1(n17046), .C2(n17006), .A(n17005), .B(n17004), .ZN(
        P2_U3003) );
  AOI22_X1 U20231 ( .A1(n19837), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19825), .ZN(n17014) );
  NAND2_X1 U20232 ( .A1(n17007), .A2(n11531), .ZN(n17008) );
  OR2_X1 U20233 ( .A1(n17009), .A2(n17008), .ZN(n17012) );
  AOI22_X1 U20234 ( .A1(n17010), .A2(n19828), .B1(n19848), .B2(n19646), .ZN(
        n17011) );
  AND2_X1 U20235 ( .A1(n17012), .A2(n17011), .ZN(n17013) );
  OAI211_X1 U20236 ( .C1(n19840), .C2(n19645), .A(n17014), .B(n17013), .ZN(
        P2_U3004) );
  AOI22_X1 U20237 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19825), .B1(n17038), 
        .B2(n17015), .ZN(n17021) );
  OAI22_X1 U20238 ( .A1(n17017), .A2(n17039), .B1(n19845), .B2(n17016), .ZN(
        n17018) );
  AOI21_X1 U20239 ( .B1(n19848), .B2(n17019), .A(n17018), .ZN(n17020) );
  OAI211_X1 U20240 ( .C1(n17046), .C2(n17022), .A(n17021), .B(n17020), .ZN(
        P2_U3005) );
  AOI22_X1 U20241 ( .A1(n19837), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19825), .ZN(n17028) );
  INV_X1 U20242 ( .A(n17023), .ZN(n17026) );
  AOI222_X1 U20243 ( .A1(n17026), .A2(n11531), .B1(n19848), .B2(n17025), .C1(
        n19828), .C2(n17024), .ZN(n17027) );
  OAI211_X1 U20244 ( .C1(n19840), .C2(n19657), .A(n17028), .B(n17027), .ZN(
        P2_U3006) );
  AOI22_X1 U20245 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19825), .B1(n17038), 
        .B2(n17029), .ZN(n17035) );
  OAI22_X1 U20246 ( .A1(n17031), .A2(n19845), .B1(n17039), .B2(n17030), .ZN(
        n17032) );
  AOI21_X1 U20247 ( .B1(n19848), .B2(n17033), .A(n17032), .ZN(n17034) );
  OAI211_X1 U20248 ( .C1(n17046), .C2(n17036), .A(n17035), .B(n17034), .ZN(
        P2_U3009) );
  AOI22_X1 U20249 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19825), .B1(n17038), 
        .B2(n17037), .ZN(n17045) );
  NOR2_X1 U20250 ( .A1(n17042), .A2(n19845), .ZN(n17043) );
  OAI211_X1 U20251 ( .C1(n17047), .C2(n17046), .A(n17045), .B(n17044), .ZN(
        P2_U3011) );
  NAND2_X1 U20252 ( .A1(n17057), .A2(n17048), .ZN(n17067) );
  AOI21_X1 U20253 ( .B1(n17051), .B2(n17050), .A(n17049), .ZN(n19724) );
  NOR3_X1 U20254 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17055), .A3(
        n17052), .ZN(n17083) );
  AOI21_X1 U20255 ( .B1(n17055), .B2(n17054), .A(n17053), .ZN(n17091) );
  INV_X1 U20256 ( .A(n17091), .ZN(n17056) );
  NOR2_X1 U20257 ( .A1(n17083), .A2(n17056), .ZN(n17069) );
  NAND3_X1 U20258 ( .A1(n17058), .A2(n17057), .A3(n17068), .ZN(n17077) );
  AOI21_X1 U20259 ( .B1(n17069), .B2(n17077), .A(n17059), .ZN(n17061) );
  INV_X1 U20260 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20417) );
  NOR2_X1 U20261 ( .A1(n19838), .A2(n20417), .ZN(n17060) );
  AOI211_X1 U20262 ( .C1(n19724), .C2(n19854), .A(n17061), .B(n17060), .ZN(
        n17066) );
  AOI222_X1 U20263 ( .A1(n17064), .A2(n19866), .B1(n11551), .B2(n17063), .C1(
        n17086), .C2(n17062), .ZN(n17065) );
  OAI211_X1 U20264 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17067), .A(
        n17066), .B(n17065), .ZN(P2_U3032) );
  OAI22_X1 U20265 ( .A1(n19728), .A2(n17070), .B1(n17069), .B2(n17068), .ZN(
        n17071) );
  AOI21_X1 U20266 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(n19825), .A(n17071), 
        .ZN(n17076) );
  AOI222_X1 U20267 ( .A1(n17074), .A2(n19866), .B1(n17073), .B2(n11551), .C1(
        n17086), .C2(n17072), .ZN(n17075) );
  OAI211_X1 U20268 ( .C1(n17090), .C2(n17077), .A(n17076), .B(n17075), .ZN(
        P2_U3033) );
  INV_X1 U20269 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20414) );
  AOI21_X1 U20270 ( .B1(n17080), .B2(n17079), .A(n17078), .ZN(n19729) );
  NAND2_X1 U20271 ( .A1(n19854), .A2(n19729), .ZN(n17081) );
  OAI21_X1 U20272 ( .B1(n20414), .B2(n19856), .A(n17081), .ZN(n17082) );
  NOR2_X1 U20273 ( .A1(n17083), .A2(n17082), .ZN(n17089) );
  AOI222_X1 U20274 ( .A1(n17087), .A2(n19866), .B1(n17086), .B2(n17085), .C1(
        n11551), .C2(n17084), .ZN(n17088) );
  OAI211_X1 U20275 ( .C1(n17091), .C2(n17090), .A(n17089), .B(n17088), .ZN(
        P2_U3034) );
  AOI211_X1 U20276 ( .C1(n20502), .C2(n17094), .A(n17093), .B(n17092), .ZN(
        n17105) );
  INV_X1 U20277 ( .A(n17095), .ZN(n17098) );
  INV_X1 U20278 ( .A(n17096), .ZN(n17097) );
  OAI21_X1 U20279 ( .B1(n17099), .B2(n17098), .A(n17097), .ZN(n17103) );
  NAND3_X1 U20280 ( .A1(n17101), .A2(n17100), .A3(n20385), .ZN(n17102) );
  NAND2_X1 U20281 ( .A1(n17103), .A2(n17102), .ZN(n17104) );
  OAI211_X1 U20282 ( .C1(n17106), .C2(n19561), .A(n17105), .B(n17104), .ZN(
        P2_U3176) );
  INV_X1 U20283 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19505) );
  NAND3_X1 U20284 ( .A1(n18570), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n17133), .ZN(n17107) );
  XNOR2_X1 U20285 ( .A(n19505), .B(n17107), .ZN(n17164) );
  INV_X1 U20286 ( .A(n17108), .ZN(n19325) );
  NOR2_X2 U20287 ( .A1(n18125), .A2(n17260), .ZN(n18547) );
  INV_X1 U20288 ( .A(n18452), .ZN(n18509) );
  NAND2_X2 U20289 ( .A1(n18554), .A2(n18509), .ZN(n18549) );
  INV_X1 U20290 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19477) );
  NOR2_X1 U20291 ( .A1(n19477), .A2(n18833), .ZN(n17158) );
  NAND2_X1 U20292 ( .A1(n17110), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18555) );
  NOR2_X2 U20293 ( .A1(n19001), .A2(n19227), .ZN(n19265) );
  OR2_X1 U20294 ( .A1(n17111), .A2(n18388), .ZN(n17129) );
  XNOR2_X1 U20295 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17114) );
  INV_X1 U20296 ( .A(n18296), .ZN(n18256) );
  NOR2_X1 U20297 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18256), .ZN(
        n17140) );
  INV_X1 U20298 ( .A(n18555), .ZN(n18384) );
  AOI22_X1 U20299 ( .A1(n18384), .A2(n17112), .B1(n19265), .B2(n17111), .ZN(
        n17113) );
  NAND2_X1 U20300 ( .A1(n17113), .A2(n18554), .ZN(n17148) );
  NOR2_X1 U20301 ( .A1(n17140), .A2(n17148), .ZN(n17128) );
  OAI22_X1 U20302 ( .A1(n17129), .A2(n17114), .B1(n17128), .B2(n17276), .ZN(
        n17115) );
  AOI211_X1 U20303 ( .C1(n18401), .C2(n17547), .A(n17158), .B(n17115), .ZN(
        n17124) );
  NAND2_X1 U20304 ( .A1(n17116), .A2(n18502), .ZN(n18467) );
  NAND3_X1 U20305 ( .A1(n17133), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n19505), .ZN(n17155) );
  OAI21_X1 U20306 ( .B1(n17117), .B2(n17134), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17118) );
  OAI21_X1 U20307 ( .B1(n17155), .B2(n18572), .A(n17118), .ZN(n17160) );
  AOI22_X1 U20308 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18382), .B1(
        n18463), .B2(n19505), .ZN(n17122) );
  NOR2_X1 U20309 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19505), .ZN(
        n17161) );
  OAI211_X1 U20310 ( .C1(n17164), .C2(n18560), .A(n17124), .B(n17123), .ZN(
        P3_U2799) );
  OAI22_X1 U20311 ( .A1(n18560), .A2(n18731), .B1(n18467), .B2(n18729), .ZN(
        n18395) );
  NAND2_X1 U20312 ( .A1(n18395), .A2(n18345), .ZN(n18356) );
  NAND2_X1 U20313 ( .A1(n17125), .A2(n18340), .ZN(n18206) );
  OAI21_X1 U20314 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n12371), .A(
        n17126), .ZN(n17285) );
  NOR2_X1 U20315 ( .A1(n18393), .A2(n17285), .ZN(n17131) );
  INV_X1 U20316 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17288) );
  OAI221_X1 U20317 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17129), .C1(
        n17288), .C2(n17128), .A(n17127), .ZN(n17130) );
  AOI21_X1 U20318 ( .B1(n18570), .B2(n17133), .A(n18560), .ZN(n17146) );
  AND2_X1 U20319 ( .A1(n17134), .A2(n18396), .ZN(n17144) );
  OAI21_X1 U20320 ( .B1(n17146), .B2(n17144), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17135) );
  OAI211_X1 U20321 ( .C1(n18206), .C2(n17137), .A(n17136), .B(n17135), .ZN(
        P3_U2800) );
  AOI221_X1 U20322 ( .B1(n17140), .B2(n17139), .C1(n18401), .C2(n17139), .A(
        n17138), .ZN(n17153) );
  OAI21_X1 U20323 ( .B1(n17142), .B2(n18572), .A(n17141), .ZN(n17143) );
  AOI22_X1 U20324 ( .A1(n18464), .A2(n17145), .B1(n17144), .B2(n17143), .ZN(
        n17152) );
  OAI21_X1 U20325 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17147), .A(
        n17146), .ZN(n17151) );
  OAI221_X1 U20326 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19265), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n17149), .A(n17148), .ZN(
        n17150) );
  NAND4_X1 U20327 ( .A1(n17153), .A2(n17152), .A3(n17151), .A4(n17150), .ZN(
        P3_U2801) );
  OAI22_X1 U20328 ( .A1(n19505), .A2(n17156), .B1(n17155), .B2(n17154), .ZN(
        n17157) );
  AOI211_X1 U20329 ( .C1(n17159), .C2(n18788), .A(n17158), .B(n17157), .ZN(
        n17163) );
  NOR2_X1 U20330 ( .A1(n18783), .A2(n18871), .ZN(n18858) );
  OAI221_X1 U20331 ( .B1(n18725), .B2(n17161), .C1(n18725), .C2(n18858), .A(
        n17160), .ZN(n17162) );
  OAI211_X1 U20332 ( .C1(n17164), .C2(n18878), .A(n17163), .B(n17162), .ZN(
        P3_U2831) );
  NOR3_X1 U20333 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n17166) );
  NOR4_X1 U20334 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17165) );
  NAND4_X1 U20335 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17166), .A3(n17165), .A4(
        U215), .ZN(U213) );
  INV_X1 U20336 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19781) );
  NOR2_X1 U20337 ( .A1(n17212), .A2(n17167), .ZN(n17214) );
  INV_X1 U20338 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17246) );
  OAI222_X1 U20339 ( .A1(U212), .A2(n19781), .B1(n17209), .B2(n19903), .C1(
        U214), .C2(n17246), .ZN(U216) );
  AOI222_X1 U20340 ( .A1(n17207), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17214), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n17212), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n17168) );
  INV_X1 U20341 ( .A(n17168), .ZN(U217) );
  AOI22_X1 U20342 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17207), .ZN(n17169) );
  OAI21_X1 U20343 ( .B1(n17170), .B2(n17209), .A(n17169), .ZN(U218) );
  AOI22_X1 U20344 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17207), .ZN(n17171) );
  OAI21_X1 U20345 ( .B1(n19889), .B2(n17209), .A(n17171), .ZN(U219) );
  AOI22_X1 U20346 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17207), .ZN(n17172) );
  OAI21_X1 U20347 ( .B1(n19885), .B2(n17209), .A(n17172), .ZN(U220) );
  AOI22_X1 U20348 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17207), .ZN(n17173) );
  OAI21_X1 U20349 ( .B1(n17174), .B2(n17209), .A(n17173), .ZN(U221) );
  AOI22_X1 U20350 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17207), .ZN(n17175) );
  OAI21_X1 U20351 ( .B1(n17176), .B2(n17209), .A(n17175), .ZN(U222) );
  AOI22_X1 U20352 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17207), .ZN(n17177) );
  OAI21_X1 U20353 ( .B1(n17178), .B2(n17209), .A(n17177), .ZN(U223) );
  AOI22_X1 U20354 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17207), .ZN(n17179) );
  OAI21_X1 U20355 ( .B1(n17180), .B2(n17209), .A(n17179), .ZN(U224) );
  AOI22_X1 U20356 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17207), .ZN(n17181) );
  OAI21_X1 U20357 ( .B1(n17182), .B2(n17209), .A(n17181), .ZN(U225) );
  AOI22_X1 U20358 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17207), .ZN(n17183) );
  OAI21_X1 U20359 ( .B1(n17184), .B2(n17209), .A(n17183), .ZN(U226) );
  AOI22_X1 U20360 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17207), .ZN(n17185) );
  OAI21_X1 U20361 ( .B1(n21269), .B2(n17209), .A(n17185), .ZN(U227) );
  AOI22_X1 U20362 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17207), .ZN(n17186) );
  OAI21_X1 U20363 ( .B1(n17187), .B2(n17209), .A(n17186), .ZN(U228) );
  AOI22_X1 U20364 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17207), .ZN(n17188) );
  OAI21_X1 U20365 ( .B1(n17189), .B2(n17209), .A(n17188), .ZN(U229) );
  AOI22_X1 U20366 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17207), .ZN(n17190) );
  OAI21_X1 U20367 ( .B1(n17191), .B2(n17209), .A(n17190), .ZN(U230) );
  AOI22_X1 U20368 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17207), .ZN(n17192) );
  OAI21_X1 U20369 ( .B1(n21227), .B2(n17209), .A(n17192), .ZN(U231) );
  INV_X1 U20370 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n21246) );
  AOI22_X1 U20371 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n17214), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n17212), .ZN(n17193) );
  OAI21_X1 U20372 ( .B1(n21246), .B2(U212), .A(n17193), .ZN(U232) );
  INV_X1 U20373 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U20374 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n17214), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n17212), .ZN(n17194) );
  OAI21_X1 U20375 ( .B1(n17195), .B2(U212), .A(n17194), .ZN(U233) );
  AOI222_X1 U20376 ( .A1(n17207), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n17214), 
        .B2(BUF1_REG_13__SCAN_IN), .C1(n17212), .C2(P1_DATAO_REG_13__SCAN_IN), 
        .ZN(n17196) );
  INV_X1 U20377 ( .A(n17196), .ZN(U234) );
  AOI22_X1 U20378 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17207), .ZN(n17197) );
  OAI21_X1 U20379 ( .B1(n17198), .B2(n17209), .A(n17197), .ZN(U235) );
  INV_X1 U20380 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20381 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n17214), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n17212), .ZN(n17199) );
  OAI21_X1 U20382 ( .B1(n17227), .B2(U212), .A(n17199), .ZN(U236) );
  INV_X1 U20383 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n21266) );
  AOI22_X1 U20384 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17207), .ZN(n17200) );
  OAI21_X1 U20385 ( .B1(n21266), .B2(n17209), .A(n17200), .ZN(U237) );
  INV_X1 U20386 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20387 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n17214), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n17212), .ZN(n17201) );
  OAI21_X1 U20388 ( .B1(n17202), .B2(U212), .A(n17201), .ZN(U238) );
  AOI22_X1 U20389 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17207), .ZN(n17203) );
  OAI21_X1 U20390 ( .B1(n17204), .B2(n17209), .A(n17203), .ZN(U239) );
  INV_X1 U20391 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20392 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17214), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17212), .ZN(n17205) );
  OAI21_X1 U20393 ( .B1(n17223), .B2(U212), .A(n17205), .ZN(U240) );
  INV_X1 U20394 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17222) );
  INV_X1 U20395 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n21113) );
  INV_X1 U20396 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n21196) );
  OAI222_X1 U20397 ( .A1(U212), .A2(n17222), .B1(n17209), .B2(n21113), .C1(
        U214), .C2(n21196), .ZN(U241) );
  AOI22_X1 U20398 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17207), .ZN(n17206) );
  OAI21_X1 U20399 ( .B1(n21094), .B2(n17209), .A(n17206), .ZN(U242) );
  INV_X1 U20400 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n21063) );
  AOI22_X1 U20401 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17212), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17207), .ZN(n17208) );
  OAI21_X1 U20402 ( .B1(n21063), .B2(n17209), .A(n17208), .ZN(U243) );
  INV_X1 U20403 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17219) );
  AOI22_X1 U20404 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n17214), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17212), .ZN(n17210) );
  OAI21_X1 U20405 ( .B1(n17219), .B2(U212), .A(n17210), .ZN(U244) );
  INV_X1 U20406 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20407 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n17214), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n17212), .ZN(n17211) );
  OAI21_X1 U20408 ( .B1(n17218), .B2(U212), .A(n17211), .ZN(U245) );
  INV_X1 U20409 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20410 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n17214), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n17212), .ZN(n17213) );
  OAI21_X1 U20411 ( .B1(n17217), .B2(U212), .A(n17213), .ZN(U246) );
  INV_X1 U20412 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20413 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n17214), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n17212), .ZN(n17215) );
  OAI21_X1 U20414 ( .B1(n17216), .B2(U212), .A(n17215), .ZN(U247) );
  INV_X1 U20415 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18890) );
  AOI22_X1 U20416 ( .A1(n17245), .A2(n17216), .B1(n18890), .B2(U215), .ZN(U251) );
  INV_X1 U20417 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18899) );
  AOI22_X1 U20418 ( .A1(n17245), .A2(n17217), .B1(n18899), .B2(U215), .ZN(U252) );
  INV_X1 U20419 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18903) );
  AOI22_X1 U20420 ( .A1(n17245), .A2(n17218), .B1(n18903), .B2(U215), .ZN(U253) );
  INV_X1 U20421 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18908) );
  AOI22_X1 U20422 ( .A1(n17245), .A2(n17219), .B1(n18908), .B2(U215), .ZN(U254) );
  OAI22_X1 U20423 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17245), .ZN(n17220) );
  INV_X1 U20424 ( .A(n17220), .ZN(U255) );
  OAI22_X1 U20425 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n17245), .ZN(n17221) );
  INV_X1 U20426 ( .A(n17221), .ZN(U256) );
  INV_X1 U20427 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18921) );
  AOI22_X1 U20428 ( .A1(n17245), .A2(n17222), .B1(n18921), .B2(U215), .ZN(U257) );
  INV_X1 U20429 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18926) );
  AOI22_X1 U20430 ( .A1(n17239), .A2(n17223), .B1(n18926), .B2(U215), .ZN(U258) );
  OAI22_X1 U20431 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17245), .ZN(n17224) );
  INV_X1 U20432 ( .A(n17224), .ZN(U259) );
  OAI22_X1 U20433 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n17245), .ZN(n17225) );
  INV_X1 U20434 ( .A(n17225), .ZN(U260) );
  OAI22_X1 U20435 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17245), .ZN(n17226) );
  INV_X1 U20436 ( .A(n17226), .ZN(U261) );
  INV_X1 U20437 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n18168) );
  AOI22_X1 U20438 ( .A1(n17245), .A2(n17227), .B1(n18168), .B2(U215), .ZN(U262) );
  OAI22_X1 U20439 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n17245), .ZN(n17228) );
  INV_X1 U20440 ( .A(n17228), .ZN(U263) );
  INV_X1 U20441 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n19790) );
  INV_X1 U20442 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n21221) );
  AOI22_X1 U20443 ( .A1(n17239), .A2(n19790), .B1(n21221), .B2(U215), .ZN(U264) );
  OAI22_X1 U20444 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17245), .ZN(n17229) );
  INV_X1 U20445 ( .A(n17229), .ZN(U265) );
  INV_X1 U20446 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n18179) );
  AOI22_X1 U20447 ( .A1(n17239), .A2(n21246), .B1(n18179), .B2(U215), .ZN(U266) );
  OAI22_X1 U20448 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17245), .ZN(n17230) );
  INV_X1 U20449 ( .A(n17230), .ZN(U267) );
  OAI22_X1 U20450 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17245), .ZN(n17231) );
  INV_X1 U20451 ( .A(n17231), .ZN(U268) );
  OAI22_X1 U20452 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17239), .ZN(n17232) );
  INV_X1 U20453 ( .A(n17232), .ZN(U269) );
  OAI22_X1 U20454 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17239), .ZN(n17233) );
  INV_X1 U20455 ( .A(n17233), .ZN(U270) );
  OAI22_X1 U20456 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17239), .ZN(n17234) );
  INV_X1 U20457 ( .A(n17234), .ZN(U271) );
  OAI22_X1 U20458 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17239), .ZN(n17235) );
  INV_X1 U20459 ( .A(n17235), .ZN(U272) );
  OAI22_X1 U20460 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17239), .ZN(n17236) );
  INV_X1 U20461 ( .A(n17236), .ZN(U273) );
  OAI22_X1 U20462 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17239), .ZN(n17237) );
  INV_X1 U20463 ( .A(n17237), .ZN(U274) );
  OAI22_X1 U20464 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17245), .ZN(n17238) );
  INV_X1 U20465 ( .A(n17238), .ZN(U275) );
  OAI22_X1 U20466 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17239), .ZN(n17240) );
  INV_X1 U20467 ( .A(n17240), .ZN(U276) );
  OAI22_X1 U20468 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17245), .ZN(n17241) );
  INV_X1 U20469 ( .A(n17241), .ZN(U277) );
  OAI22_X1 U20470 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17245), .ZN(n17242) );
  INV_X1 U20471 ( .A(n17242), .ZN(U278) );
  OAI22_X1 U20472 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17245), .ZN(n17243) );
  INV_X1 U20473 ( .A(n17243), .ZN(U279) );
  OAI22_X1 U20474 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17245), .ZN(n17244) );
  INV_X1 U20475 ( .A(n17244), .ZN(U280) );
  INV_X1 U20476 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19785) );
  INV_X1 U20477 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U20478 ( .A1(n17245), .A2(n19785), .B1(n19894), .B2(U215), .ZN(U281) );
  INV_X1 U20479 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19901) );
  AOI22_X1 U20480 ( .A1(n17245), .A2(n19781), .B1(n19901), .B2(U215), .ZN(U282) );
  INV_X1 U20481 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18073) );
  AOI222_X1 U20482 ( .A1(n17246), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19781), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n18073), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17247) );
  INV_X1 U20483 ( .A(n17249), .ZN(n17248) );
  INV_X1 U20484 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19440) );
  INV_X1 U20485 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n21224) );
  AOI22_X1 U20486 ( .A1(n17248), .A2(n19440), .B1(n21224), .B2(n17249), .ZN(
        U347) );
  INV_X1 U20487 ( .A(n17249), .ZN(n17250) );
  INV_X1 U20488 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19438) );
  INV_X1 U20489 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20410) );
  AOI22_X1 U20490 ( .A1(n17250), .A2(n19438), .B1(n20410), .B2(n17249), .ZN(
        U348) );
  INV_X1 U20491 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19436) );
  INV_X1 U20492 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20408) );
  AOI22_X1 U20493 ( .A1(n17248), .A2(n19436), .B1(n20408), .B2(n17249), .ZN(
        U349) );
  INV_X1 U20494 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19435) );
  INV_X1 U20495 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20406) );
  AOI22_X1 U20496 ( .A1(n17248), .A2(n19435), .B1(n20406), .B2(n17249), .ZN(
        U350) );
  INV_X1 U20497 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19433) );
  INV_X1 U20498 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20404) );
  AOI22_X1 U20499 ( .A1(n17248), .A2(n19433), .B1(n20404), .B2(n17249), .ZN(
        U351) );
  INV_X1 U20500 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19430) );
  INV_X1 U20501 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20402) );
  AOI22_X1 U20502 ( .A1(n17248), .A2(n19430), .B1(n20402), .B2(n17249), .ZN(
        U352) );
  INV_X1 U20503 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19429) );
  INV_X1 U20504 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20401) );
  AOI22_X1 U20505 ( .A1(n17250), .A2(n19429), .B1(n20401), .B2(n17249), .ZN(
        U353) );
  INV_X1 U20506 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19427) );
  AOI22_X1 U20507 ( .A1(n17248), .A2(n19427), .B1(n20399), .B2(n17249), .ZN(
        U354) );
  INV_X1 U20508 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19478) );
  INV_X1 U20509 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20446) );
  AOI22_X1 U20510 ( .A1(n17248), .A2(n19478), .B1(n20446), .B2(n17249), .ZN(
        U355) );
  INV_X1 U20511 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19476) );
  INV_X1 U20512 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20443) );
  AOI22_X1 U20513 ( .A1(n17248), .A2(n19476), .B1(n20443), .B2(n17249), .ZN(
        U356) );
  INV_X1 U20514 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19473) );
  INV_X1 U20515 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20441) );
  AOI22_X1 U20516 ( .A1(n17248), .A2(n19473), .B1(n20441), .B2(n17249), .ZN(
        U357) );
  INV_X1 U20517 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19470) );
  INV_X1 U20518 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20438) );
  AOI22_X1 U20519 ( .A1(n17248), .A2(n19470), .B1(n20438), .B2(n17249), .ZN(
        U358) );
  INV_X1 U20520 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19467) );
  INV_X1 U20521 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20437) );
  AOI22_X1 U20522 ( .A1(n17248), .A2(n19467), .B1(n20437), .B2(n17249), .ZN(
        U359) );
  INV_X1 U20523 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19466) );
  INV_X1 U20524 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20435) );
  AOI22_X1 U20525 ( .A1(n17248), .A2(n19466), .B1(n20435), .B2(n17249), .ZN(
        U360) );
  INV_X1 U20526 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19464) );
  INV_X1 U20527 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20434) );
  AOI22_X1 U20528 ( .A1(n17248), .A2(n19464), .B1(n20434), .B2(n17249), .ZN(
        U361) );
  INV_X1 U20529 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19462) );
  INV_X1 U20530 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20433) );
  AOI22_X1 U20531 ( .A1(n17248), .A2(n19462), .B1(n20433), .B2(n17249), .ZN(
        U362) );
  INV_X1 U20532 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19460) );
  INV_X1 U20533 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20431) );
  AOI22_X1 U20534 ( .A1(n17248), .A2(n19460), .B1(n20431), .B2(n17249), .ZN(
        U363) );
  INV_X1 U20535 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19458) );
  INV_X1 U20536 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20430) );
  AOI22_X1 U20537 ( .A1(n17248), .A2(n19458), .B1(n20430), .B2(n17249), .ZN(
        U364) );
  INV_X1 U20538 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19425) );
  INV_X1 U20539 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20398) );
  AOI22_X1 U20540 ( .A1(n17248), .A2(n19425), .B1(n20398), .B2(n17249), .ZN(
        U365) );
  INV_X1 U20541 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19456) );
  INV_X1 U20542 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20428) );
  AOI22_X1 U20543 ( .A1(n17248), .A2(n19456), .B1(n20428), .B2(n17249), .ZN(
        U366) );
  INV_X1 U20544 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19454) );
  INV_X1 U20545 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20426) );
  AOI22_X1 U20546 ( .A1(n17248), .A2(n19454), .B1(n20426), .B2(n17249), .ZN(
        U367) );
  INV_X1 U20547 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19452) );
  INV_X1 U20548 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20424) );
  AOI22_X1 U20549 ( .A1(n17248), .A2(n19452), .B1(n20424), .B2(n17249), .ZN(
        U368) );
  INV_X1 U20550 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19449) );
  INV_X1 U20551 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20421) );
  AOI22_X1 U20552 ( .A1(n17248), .A2(n19449), .B1(n20421), .B2(n17249), .ZN(
        U369) );
  INV_X1 U20553 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19448) );
  INV_X1 U20554 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20419) );
  AOI22_X1 U20555 ( .A1(n17248), .A2(n19448), .B1(n20419), .B2(n17249), .ZN(
        U370) );
  INV_X1 U20556 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19446) );
  INV_X1 U20557 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n21122) );
  AOI22_X1 U20558 ( .A1(n17250), .A2(n19446), .B1(n21122), .B2(n17249), .ZN(
        U371) );
  INV_X1 U20559 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19444) );
  INV_X1 U20560 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20418) );
  AOI22_X1 U20561 ( .A1(n17250), .A2(n19444), .B1(n20418), .B2(n17249), .ZN(
        U372) );
  INV_X1 U20562 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19443) );
  INV_X1 U20563 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20416) );
  AOI22_X1 U20564 ( .A1(n17250), .A2(n19443), .B1(n20416), .B2(n17249), .ZN(
        U373) );
  INV_X1 U20565 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n21149) );
  INV_X1 U20566 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20415) );
  AOI22_X1 U20567 ( .A1(n17250), .A2(n21149), .B1(n20415), .B2(n17249), .ZN(
        U374) );
  INV_X1 U20568 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19441) );
  INV_X1 U20569 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20413) );
  AOI22_X1 U20570 ( .A1(n17250), .A2(n19441), .B1(n20413), .B2(n17249), .ZN(
        U375) );
  INV_X1 U20571 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19422) );
  INV_X1 U20572 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20397) );
  AOI22_X1 U20573 ( .A1(n17250), .A2(n19422), .B1(n20397), .B2(n17249), .ZN(
        U376) );
  INV_X1 U20574 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19421) );
  NAND2_X1 U20575 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19421), .ZN(n19407) );
  AOI21_X1 U20576 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19489), .ZN(n17251) );
  INV_X1 U20577 ( .A(n17251), .ZN(P3_U2633) );
  OAI21_X1 U20578 ( .B1(n17259), .B2(n18123), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17252) );
  OAI21_X1 U20579 ( .B1(n17253), .B2(n19396), .A(n17252), .ZN(P3_U2634) );
  AOI21_X1 U20580 ( .B1(n19419), .B2(n19421), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17254) );
  AOI22_X1 U20581 ( .A1(n19484), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17254), 
        .B2(n19548), .ZN(P3_U2635) );
  NOR2_X1 U20582 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n17255) );
  OAI21_X1 U20583 ( .B1(n17255), .B2(BS16), .A(n19489), .ZN(n19487) );
  OAI21_X1 U20584 ( .B1(n19489), .B2(n19538), .A(n19487), .ZN(P3_U2636) );
  INV_X1 U20585 ( .A(n17256), .ZN(n17258) );
  NOR3_X1 U20586 ( .A1(n17259), .A2(n17258), .A3(n17257), .ZN(n19327) );
  NOR2_X1 U20587 ( .A1(n19327), .A2(n19391), .ZN(n19532) );
  OAI21_X1 U20588 ( .B1(n19532), .B2(n18881), .A(n17260), .ZN(P3_U2637) );
  NOR2_X1 U20589 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21288) );
  AOI211_X1 U20590 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_16__SCAN_IN), .B(
        P3_DATAWIDTH_REG_20__SCAN_IN), .ZN(n17261) );
  INV_X1 U20591 ( .A(P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n21145) );
  INV_X1 U20592 ( .A(P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n21166) );
  NAND4_X1 U20593 ( .A1(n21288), .A2(n17261), .A3(n21145), .A4(n21166), .ZN(
        n17269) );
  OR4_X1 U20594 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n17268) );
  OR4_X1 U20595 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n17267) );
  NOR4_X1 U20596 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n17265) );
  NOR4_X1 U20597 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n17264) );
  NOR4_X1 U20598 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_26__SCAN_IN), .A3(P3_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(n17263) );
  NOR4_X1 U20599 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_23__SCAN_IN), .A3(P3_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17262) );
  NAND4_X1 U20600 ( .A1(n17265), .A2(n17264), .A3(n17263), .A4(n17262), .ZN(
        n17266) );
  INV_X1 U20601 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19483) );
  NOR3_X1 U20602 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17271) );
  OAI21_X1 U20603 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17271), .A(n19530), .ZN(
        n17270) );
  OAI21_X1 U20604 ( .B1(n19530), .B2(n19483), .A(n17270), .ZN(P3_U2638) );
  INV_X1 U20605 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19488) );
  AOI21_X1 U20606 ( .B1(n19423), .B2(n19488), .A(n17271), .ZN(n17273) );
  INV_X1 U20607 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17272) );
  INV_X1 U20608 ( .A(n19530), .ZN(n19527) );
  AOI22_X1 U20609 ( .A1(n19530), .A2(n17273), .B1(n17272), .B2(n19527), .ZN(
        P3_U2639) );
  NOR2_X1 U20610 ( .A1(n17615), .A2(n17274), .ZN(n17293) );
  INV_X1 U20611 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17633) );
  INV_X1 U20612 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19479) );
  NAND4_X1 U20613 ( .A1(n17298), .A2(P3_REIP_REG_29__SCAN_IN), .A3(
        P3_REIP_REG_28__SCAN_IN), .A4(P3_REIP_REG_27__SCAN_IN), .ZN(n17279) );
  NOR3_X1 U20614 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19479), .A3(n17279), 
        .ZN(n17278) );
  INV_X1 U20615 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n17275) );
  OAI22_X1 U20616 ( .A1(n17276), .A2(n17605), .B1(n17275), .B2(n17608), .ZN(
        n17277) );
  AOI211_X1 U20617 ( .C1(n17293), .C2(n17633), .A(n17278), .B(n17277), .ZN(
        n17283) );
  NOR2_X1 U20618 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17279), .ZN(n17289) );
  INV_X1 U20619 ( .A(n17287), .ZN(n17280) );
  OAI21_X1 U20620 ( .B1(n17289), .B2(n17280), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n17282) );
  NAND4_X1 U20621 ( .A1(n17547), .A2(n17591), .A3(n17284), .A4(n17285), .ZN(
        n17281) );
  NAND3_X1 U20622 ( .A1(n17283), .A2(n17282), .A3(n17281), .ZN(P3_U2640) );
  XNOR2_X1 U20623 ( .A(n17286), .B(n17285), .ZN(n17292) );
  OAI22_X1 U20624 ( .A1(n17288), .A2(n17605), .B1(n19479), .B2(n17287), .ZN(
        n17290) );
  AOI21_X1 U20625 ( .B1(n17292), .B2(n17591), .A(n17291), .ZN(n17295) );
  OAI21_X1 U20626 ( .B1(n17617), .B2(n17293), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17294) );
  OAI211_X1 U20627 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17296), .A(n17295), .B(
        n17294), .ZN(P3_U2641) );
  NAND2_X1 U20628 ( .A1(n17298), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17307) );
  AOI22_X1 U20629 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17598), .B1(
        n17617), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17306) );
  NAND2_X1 U20630 ( .A1(n17619), .A2(n17297), .ZN(n17324) );
  INV_X1 U20631 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19469) );
  NAND2_X1 U20632 ( .A1(n17298), .A2(n19469), .ZN(n17310) );
  NAND2_X1 U20633 ( .A1(n17324), .A2(n17310), .ZN(n17304) );
  AOI211_X1 U20634 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17313), .A(n17299), .B(
        n17615), .ZN(n17303) );
  AOI211_X1 U20635 ( .C1(n18194), .C2(n17301), .A(n17300), .B(n19399), .ZN(
        n17302) );
  AOI211_X1 U20636 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17304), .A(n17303), 
        .B(n17302), .ZN(n17305) );
  OAI211_X1 U20637 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17307), .A(n17306), 
        .B(n17305), .ZN(P3_U2643) );
  AOI211_X1 U20638 ( .C1(n18203), .C2(n17309), .A(n17308), .B(n19399), .ZN(
        n17312) );
  OAI21_X1 U20639 ( .B1(n17671), .B2(n17608), .A(n17310), .ZN(n17311) );
  AOI211_X1 U20640 ( .C1(n17598), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17312), .B(n17311), .ZN(n17315) );
  OAI211_X1 U20641 ( .C1(n17317), .C2(n17671), .A(n17616), .B(n17313), .ZN(
        n17314) );
  OAI211_X1 U20642 ( .C1(n17324), .C2(n19469), .A(n17315), .B(n17314), .ZN(
        P3_U2644) );
  NOR2_X1 U20643 ( .A1(n17609), .A2(n17316), .ZN(n17331) );
  AOI21_X1 U20644 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n17331), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20645 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17598), .B1(
        n17617), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17323) );
  AOI211_X1 U20646 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17332), .A(n17317), .B(
        n17615), .ZN(n17321) );
  AOI211_X1 U20647 ( .C1(n18217), .C2(n17319), .A(n17318), .B(n19399), .ZN(
        n17320) );
  NOR2_X1 U20648 ( .A1(n17321), .A2(n17320), .ZN(n17322) );
  OAI211_X1 U20649 ( .C1(n17325), .C2(n17324), .A(n17323), .B(n17322), .ZN(
        P3_U2645) );
  INV_X1 U20650 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19463) );
  OAI21_X1 U20651 ( .B1(n17337), .B2(n17609), .A(n17620), .ZN(n17346) );
  AOI21_X1 U20652 ( .B1(n17600), .B2(n19463), .A(n17346), .ZN(n17335) );
  AOI211_X1 U20653 ( .C1(n18227), .C2(n17327), .A(n17326), .B(n19399), .ZN(
        n17330) );
  OAI22_X1 U20654 ( .A1(n17328), .A2(n17605), .B1(n17608), .B2(n17624), .ZN(
        n17329) );
  AOI211_X1 U20655 ( .C1(n17331), .C2(n19465), .A(n17330), .B(n17329), .ZN(
        n17334) );
  OAI211_X1 U20656 ( .C1(n17338), .C2(n17624), .A(n17616), .B(n17332), .ZN(
        n17333) );
  OAI211_X1 U20657 ( .C1(n17335), .C2(n19465), .A(n17334), .B(n17333), .ZN(
        P3_U2646) );
  NOR2_X1 U20658 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17609), .ZN(n17336) );
  AOI22_X1 U20659 ( .A1(n17617), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17337), 
        .B2(n17336), .ZN(n17344) );
  AOI211_X1 U20660 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17351), .A(n17338), .B(
        n17615), .ZN(n17342) );
  AOI211_X1 U20661 ( .C1(n18240), .C2(n17340), .A(n17339), .B(n19399), .ZN(
        n17341) );
  AOI211_X1 U20662 ( .C1(n17346), .C2(P3_REIP_REG_24__SCAN_IN), .A(n17342), 
        .B(n17341), .ZN(n17343) );
  OAI211_X1 U20663 ( .C1(n18244), .C2(n17605), .A(n17344), .B(n17343), .ZN(
        P3_U2647) );
  AOI21_X1 U20664 ( .B1(n17600), .B2(n17345), .A(P3_REIP_REG_23__SCAN_IN), 
        .ZN(n17355) );
  INV_X1 U20665 ( .A(n17346), .ZN(n17354) );
  AOI211_X1 U20666 ( .C1(n18257), .C2(n17347), .A(n9808), .B(n19399), .ZN(
        n17350) );
  OAI22_X1 U20667 ( .A1(n17348), .A2(n17605), .B1(n17608), .B2(n17626), .ZN(
        n17349) );
  NOR2_X1 U20668 ( .A1(n17350), .A2(n17349), .ZN(n17353) );
  OAI211_X1 U20669 ( .C1(n17356), .C2(n17626), .A(n17616), .B(n17351), .ZN(
        n17352) );
  OAI211_X1 U20670 ( .C1(n17355), .C2(n17354), .A(n17353), .B(n17352), .ZN(
        P3_U2648) );
  AOI21_X1 U20671 ( .B1(n17600), .B2(n17359), .A(n17604), .ZN(n17372) );
  AOI211_X1 U20672 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17369), .A(n17356), .B(
        n17615), .ZN(n17363) );
  AOI211_X1 U20673 ( .C1(n18273), .C2(n17358), .A(n17357), .B(n19399), .ZN(
        n17362) );
  NOR3_X1 U20674 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17609), .A3(n17359), 
        .ZN(n17361) );
  OAI22_X1 U20675 ( .A1(n18270), .A2(n17605), .B1(n17608), .B2(n17625), .ZN(
        n17360) );
  NOR4_X1 U20676 ( .A1(n17363), .A2(n17362), .A3(n17361), .A4(n17360), .ZN(
        n17364) );
  OAI21_X1 U20677 ( .B1(n19459), .B2(n17372), .A(n17364), .ZN(P3_U2649) );
  NAND2_X1 U20678 ( .A1(n17600), .A2(n17376), .ZN(n17436) );
  NOR2_X1 U20679 ( .A1(n17377), .A2(n17436), .ZN(n17405) );
  AOI21_X1 U20680 ( .B1(n17378), .B2(n17405), .A(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n17373) );
  AOI211_X1 U20681 ( .C1(n18289), .C2(n17366), .A(n17365), .B(n19399), .ZN(
        n17368) );
  OAI22_X1 U20682 ( .A1(n18286), .A2(n17605), .B1(n17608), .B2(n17703), .ZN(
        n17367) );
  NOR2_X1 U20683 ( .A1(n17368), .A2(n17367), .ZN(n17371) );
  OAI211_X1 U20684 ( .C1(n17374), .C2(n17703), .A(n17616), .B(n17369), .ZN(
        n17370) );
  OAI211_X1 U20685 ( .C1(n17373), .C2(n17372), .A(n17371), .B(n17370), .ZN(
        P3_U2650) );
  AOI211_X1 U20686 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17391), .A(n17374), .B(
        n17615), .ZN(n17375) );
  AOI21_X1 U20687 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17617), .A(n17375), .ZN(
        n17386) );
  NAND2_X1 U20688 ( .A1(n17376), .A2(n17620), .ZN(n17439) );
  NOR2_X1 U20689 ( .A1(n17377), .A2(n17439), .ZN(n17387) );
  AOI21_X1 U20690 ( .B1(n17378), .B2(n17387), .A(n19455), .ZN(n17384) );
  AOI211_X1 U20691 ( .C1(n17381), .C2(n17380), .A(n17379), .B(n19399), .ZN(
        n17383) );
  NAND2_X1 U20692 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n17405), .ZN(n17398) );
  NOR3_X1 U20693 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n19453), .A3(n17398), 
        .ZN(n17382) );
  AOI211_X1 U20694 ( .C1(n17384), .C2(n17619), .A(n17383), .B(n17382), .ZN(
        n17385) );
  OAI211_X1 U20695 ( .C1(n21230), .C2(n17605), .A(n17386), .B(n17385), .ZN(
        P3_U2651) );
  NOR2_X1 U20696 ( .A1(n17388), .A2(n17387), .ZN(n17416) );
  AOI21_X1 U20697 ( .B1(n17405), .B2(n19451), .A(n17416), .ZN(n17397) );
  AOI211_X1 U20698 ( .C1(n18308), .C2(n17390), .A(n17389), .B(n19399), .ZN(
        n17395) );
  OAI211_X1 U20699 ( .C1(n17399), .C2(n17393), .A(n17616), .B(n17391), .ZN(
        n17392) );
  OAI211_X1 U20700 ( .C1(n17608), .C2(n17393), .A(n18833), .B(n17392), .ZN(
        n17394) );
  AOI211_X1 U20701 ( .C1(n17598), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n17395), .B(n17394), .ZN(n17396) );
  OAI221_X1 U20702 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(n17398), .C1(n19453), 
        .C2(n17397), .A(n17396), .ZN(P3_U2652) );
  AOI211_X1 U20703 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17410), .A(n17399), .B(
        n17615), .ZN(n17400) );
  AOI211_X1 U20704 ( .C1(n17617), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18828), .B(
        n17400), .ZN(n17407) );
  AOI211_X1 U20705 ( .C1(n17403), .C2(n17402), .A(n17401), .B(n19399), .ZN(
        n17404) );
  AOI221_X1 U20706 ( .B1(n17416), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n17405), 
        .C2(n19451), .A(n17404), .ZN(n17406) );
  OAI211_X1 U20707 ( .C1(n18327), .C2(n17605), .A(n17407), .B(n17406), .ZN(
        P3_U2653) );
  INV_X1 U20708 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19447) );
  INV_X1 U20709 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n21323) );
  OR2_X1 U20710 ( .A1(n21323), .A2(n17436), .ZN(n17425) );
  INV_X1 U20711 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19450) );
  OAI21_X1 U20712 ( .B1(n19447), .B2(n17425), .A(n19450), .ZN(n17415) );
  AOI211_X1 U20713 ( .C1(n18339), .C2(n17409), .A(n17408), .B(n19399), .ZN(
        n17414) );
  OAI211_X1 U20714 ( .C1(n17419), .C2(n17412), .A(n17616), .B(n17410), .ZN(
        n17411) );
  OAI21_X1 U20715 ( .B1(n17412), .B2(n17608), .A(n17411), .ZN(n17413) );
  AOI211_X1 U20716 ( .C1(n17416), .C2(n17415), .A(n17414), .B(n17413), .ZN(
        n17417) );
  OAI211_X1 U20717 ( .C1(n18337), .C2(n17605), .A(n17417), .B(n18833), .ZN(
        P3_U2654) );
  OAI21_X1 U20718 ( .B1(n21323), .B2(n17439), .A(n17619), .ZN(n17437) );
  AOI211_X1 U20719 ( .C1(n18348), .C2(n10325), .A(n17418), .B(n19399), .ZN(
        n17423) );
  AOI211_X1 U20720 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17430), .A(n17419), .B(
        n17615), .ZN(n17422) );
  AOI22_X1 U20721 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17598), .B1(
        n17617), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n17420) );
  INV_X1 U20722 ( .A(n17420), .ZN(n17421) );
  NOR4_X1 U20723 ( .A1(n18828), .A2(n17423), .A3(n17422), .A4(n17421), .ZN(
        n17424) );
  OAI221_X1 U20724 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n17425), .C1(n19447), 
        .C2(n17437), .A(n17424), .ZN(P3_U2655) );
  OAI21_X1 U20725 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18347), .A(
        n17426), .ZN(n18357) );
  INV_X1 U20726 ( .A(n18357), .ZN(n17429) );
  NOR2_X1 U20727 ( .A1(n19399), .A2(n17547), .ZN(n17560) );
  INV_X1 U20728 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17607) );
  AOI21_X1 U20729 ( .B1(n18347), .B2(n17607), .A(n18357), .ZN(n17427) );
  NOR2_X1 U20730 ( .A1(n17427), .A2(n19399), .ZN(n17428) );
  OAI22_X1 U20731 ( .A1(n10325), .A2(n17429), .B1(n17560), .B2(n17428), .ZN(
        n17433) );
  OAI211_X1 U20732 ( .C1(n17438), .C2(n17431), .A(n17616), .B(n17430), .ZN(
        n17432) );
  OAI211_X1 U20733 ( .C1(n17605), .C2(n18360), .A(n17433), .B(n17432), .ZN(
        n17434) );
  AOI211_X1 U20734 ( .C1(n17617), .C2(P3_EBX_REG_15__SCAN_IN), .A(n18828), .B(
        n17434), .ZN(n17435) );
  OAI221_X1 U20735 ( .B1(n17437), .B2(n21323), .C1(n17437), .C2(n17436), .A(
        n17435), .ZN(P3_U2656) );
  AOI211_X1 U20736 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17452), .A(n17438), .B(
        n17615), .ZN(n17445) );
  INV_X1 U20737 ( .A(n17439), .ZN(n17443) );
  NOR2_X1 U20738 ( .A1(n17609), .A2(n17440), .ZN(n17447) );
  AOI22_X1 U20739 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17447), .B1(
        P3_REIP_REG_14__SCAN_IN), .B2(n17619), .ZN(n17442) );
  NOR2_X1 U20740 ( .A1(n18387), .A2(n18548), .ZN(n18386) );
  INV_X1 U20741 ( .A(n18386), .ZN(n17463) );
  AOI221_X1 U20742 ( .B1(n18389), .B2(n21325), .C1(n17463), .C2(n21325), .A(
        n18347), .ZN(n18373) );
  NOR2_X1 U20743 ( .A1(n18548), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17592) );
  INV_X1 U20744 ( .A(n17592), .ZN(n17567) );
  OAI21_X1 U20745 ( .B1(n18387), .B2(n17567), .A(n17547), .ZN(n17464) );
  INV_X1 U20746 ( .A(n17464), .ZN(n17466) );
  AOI21_X1 U20747 ( .B1(n18389), .B2(n17547), .A(n17466), .ZN(n17451) );
  XOR2_X1 U20748 ( .A(n18373), .B(n17451), .Z(n17441) );
  OAI22_X1 U20749 ( .A1(n17443), .A2(n17442), .B1(n19399), .B2(n17441), .ZN(
        n17444) );
  AOI211_X1 U20750 ( .C1(n17598), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17445), .B(n17444), .ZN(n17446) );
  OAI211_X1 U20751 ( .C1(n17608), .C2(n17812), .A(n17446), .B(n18833), .ZN(
        P3_U2657) );
  AOI22_X1 U20752 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17598), .B1(
        n17447), .B2(n21324), .ZN(n17459) );
  INV_X1 U20753 ( .A(n17448), .ZN(n17460) );
  AOI21_X1 U20754 ( .B1(n17600), .B2(n17460), .A(n17604), .ZN(n17477) );
  OAI21_X1 U20755 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17609), .A(n17477), 
        .ZN(n17457) );
  INV_X1 U20756 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18405) );
  NOR2_X1 U20757 ( .A1(n18405), .A2(n17463), .ZN(n17462) );
  OAI22_X1 U20758 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17462), .B1(
        n17463), .B2(n18389), .ZN(n18392) );
  INV_X1 U20759 ( .A(n17560), .ZN(n17595) );
  NOR2_X1 U20760 ( .A1(n18387), .A2(n17567), .ZN(n17449) );
  OAI221_X1 U20761 ( .B1(n18392), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C1(
        n18392), .C2(n17449), .A(n17591), .ZN(n17450) );
  AOI22_X1 U20762 ( .A1(n17451), .A2(n18392), .B1(n17595), .B2(n17450), .ZN(
        n17456) );
  OAI211_X1 U20763 ( .C1(n17467), .C2(n17454), .A(n17616), .B(n17452), .ZN(
        n17453) );
  OAI21_X1 U20764 ( .B1(n17454), .B2(n17608), .A(n17453), .ZN(n17455) );
  AOI211_X1 U20765 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17457), .A(n17456), 
        .B(n17455), .ZN(n17458) );
  NAND3_X1 U20766 ( .A1(n17459), .A2(n17458), .A3(n18833), .ZN(P3_U2658) );
  INV_X1 U20767 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19442) );
  NOR3_X1 U20768 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17609), .A3(n17460), 
        .ZN(n17461) );
  AOI211_X1 U20769 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17598), .A(
        n18828), .B(n17461), .ZN(n17471) );
  AOI21_X1 U20770 ( .B1(n18405), .B2(n17463), .A(n17462), .ZN(n18400) );
  INV_X1 U20771 ( .A(n18400), .ZN(n17465) );
  AOI221_X1 U20772 ( .B1(n18400), .B2(n17466), .C1(n17465), .C2(n17464), .A(
        n19399), .ZN(n17469) );
  AOI211_X1 U20773 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17480), .A(n17467), .B(
        n17615), .ZN(n17468) );
  AOI211_X1 U20774 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17617), .A(n17469), .B(
        n17468), .ZN(n17470) );
  OAI211_X1 U20775 ( .C1(n19442), .C2(n17477), .A(n17471), .B(n17470), .ZN(
        P3_U2659) );
  INV_X1 U20776 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17484) );
  NOR2_X1 U20777 ( .A1(n17609), .A2(n17485), .ZN(n17541) );
  INV_X1 U20778 ( .A(n17541), .ZN(n17521) );
  NOR2_X1 U20779 ( .A1(n17486), .A2(n17521), .ZN(n17500) );
  AOI21_X1 U20780 ( .B1(n17472), .B2(n17500), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17478) );
  NOR2_X1 U20781 ( .A1(n18481), .A2(n18548), .ZN(n17546) );
  INV_X1 U20782 ( .A(n17546), .ZN(n17537) );
  NOR2_X1 U20783 ( .A1(n18492), .A2(n17537), .ZN(n17536) );
  AND2_X1 U20784 ( .A1(n17504), .A2(n17536), .ZN(n17512) );
  NAND2_X1 U20785 ( .A1(n17473), .A2(n17512), .ZN(n17487) );
  OAI21_X1 U20786 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17487), .A(
        n17547), .ZN(n17475) );
  AOI21_X1 U20787 ( .B1(n17484), .B2(n17487), .A(n18386), .ZN(n17474) );
  INV_X1 U20788 ( .A(n17474), .ZN(n18416) );
  XNOR2_X1 U20789 ( .A(n17475), .B(n18416), .ZN(n17476) );
  OAI22_X1 U20790 ( .A1(n17478), .A2(n17477), .B1(n19399), .B2(n17476), .ZN(
        n17479) );
  AOI211_X1 U20791 ( .C1(n17617), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18828), .B(
        n17479), .ZN(n17483) );
  OAI211_X1 U20792 ( .C1(n17490), .C2(n17481), .A(n17616), .B(n17480), .ZN(
        n17482) );
  OAI211_X1 U20793 ( .C1(n17605), .C2(n17484), .A(n17483), .B(n17482), .ZN(
        P3_U2660) );
  AOI21_X1 U20794 ( .B1(n17485), .B2(n17600), .A(n17604), .ZN(n17550) );
  INV_X1 U20795 ( .A(n17550), .ZN(n17540) );
  AOI21_X1 U20796 ( .B1(n17600), .B2(n17486), .A(n17540), .ZN(n17516) );
  NAND2_X1 U20797 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17512), .ZN(
        n17503) );
  OAI21_X1 U20798 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17503), .A(
        n17547), .ZN(n17506) );
  INV_X1 U20799 ( .A(n17503), .ZN(n17488) );
  OAI21_X1 U20800 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17488), .A(
        n17487), .ZN(n18439) );
  OAI21_X1 U20801 ( .B1(n17506), .B2(n18439), .A(n17591), .ZN(n17489) );
  AOI21_X1 U20802 ( .B1(n17506), .B2(n18439), .A(n17489), .ZN(n17495) );
  AOI211_X1 U20803 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17491), .A(n17490), .B(
        n17615), .ZN(n17494) );
  AOI22_X1 U20804 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17598), .B1(
        n17617), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n17492) );
  INV_X1 U20805 ( .A(n17492), .ZN(n17493) );
  NOR4_X1 U20806 ( .A1(n18828), .A2(n17495), .A3(n17494), .A4(n17493), .ZN(
        n17498) );
  OAI211_X1 U20807 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n17500), .B(n17496), .ZN(n17497) );
  OAI211_X1 U20808 ( .C1(n17516), .C2(n19439), .A(n17498), .B(n17497), .ZN(
        P3_U2661) );
  AOI21_X1 U20809 ( .B1(n17616), .B2(n17502), .A(n17617), .ZN(n17499) );
  INV_X1 U20810 ( .A(n17499), .ZN(n17501) );
  AOI22_X1 U20811 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17501), .B1(n17500), .B2(
        n19437), .ZN(n17510) );
  NOR2_X1 U20812 ( .A1(n17502), .A2(n17615), .ZN(n17514) );
  OAI21_X1 U20813 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17512), .A(
        n17503), .ZN(n18444) );
  INV_X1 U20814 ( .A(n17511), .ZN(n18471) );
  NOR2_X1 U20815 ( .A1(n18471), .A2(n17567), .ZN(n17538) );
  OAI221_X1 U20816 ( .B1(n18444), .B2(n17504), .C1(n18444), .C2(n17538), .A(
        n17591), .ZN(n17505) );
  AOI22_X1 U20817 ( .A1(n17506), .A2(n18444), .B1(n17595), .B2(n17505), .ZN(
        n17508) );
  INV_X1 U20818 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18431) );
  OAI21_X1 U20819 ( .B1(n18431), .B2(n17605), .A(n18833), .ZN(n17507) );
  AOI211_X1 U20820 ( .C1(n17514), .C2(n17854), .A(n17508), .B(n17507), .ZN(
        n17509) );
  OAI211_X1 U20821 ( .C1(n17516), .C2(n19437), .A(n17510), .B(n17509), .ZN(
        P3_U2662) );
  NAND3_X1 U20822 ( .A1(n17511), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17522) );
  AOI21_X1 U20823 ( .B1(n18457), .B2(n17522), .A(n17512), .ZN(n18453) );
  OAI21_X1 U20824 ( .B1(n17522), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n17547), .ZN(n17524) );
  XOR2_X1 U20825 ( .A(n18453), .B(n17524), .Z(n17520) );
  INV_X1 U20826 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19434) );
  INV_X1 U20827 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19432) );
  NOR4_X1 U20828 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n19434), .A3(n19432), .A4(
        n17521), .ZN(n17518) );
  INV_X1 U20829 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n21222) );
  NAND2_X1 U20830 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17529), .ZN(n17513) );
  AOI22_X1 U20831 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17598), .B1(
        n17514), .B2(n17513), .ZN(n17515) );
  OAI211_X1 U20832 ( .C1(n17516), .C2(n21222), .A(n17515), .B(n18833), .ZN(
        n17517) );
  AOI211_X1 U20833 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17617), .A(n17518), .B(
        n17517), .ZN(n17519) );
  OAI21_X1 U20834 ( .B1(n19399), .B2(n17520), .A(n17519), .ZN(P3_U2663) );
  OAI21_X1 U20835 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n17521), .A(n17550), .ZN(
        n17528) );
  OAI21_X1 U20836 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17536), .A(
        n17522), .ZN(n18480) );
  OAI21_X1 U20837 ( .B1(n17538), .B2(n18480), .A(n17591), .ZN(n17523) );
  AOI22_X1 U20838 ( .A1(n18480), .A2(n17524), .B1(n17595), .B2(n17523), .ZN(
        n17527) );
  NAND3_X1 U20839 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17541), .A3(n19434), 
        .ZN(n17525) );
  OAI211_X1 U20840 ( .C1(n17608), .C2(n17530), .A(n18833), .B(n17525), .ZN(
        n17526) );
  AOI211_X1 U20841 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n17528), .A(n17527), .B(
        n17526), .ZN(n17532) );
  OAI211_X1 U20842 ( .C1(n17533), .C2(n17530), .A(n17616), .B(n17529), .ZN(
        n17531) );
  OAI211_X1 U20843 ( .C1(n17605), .C2(n18469), .A(n17532), .B(n17531), .ZN(
        P3_U2664) );
  AOI211_X1 U20844 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17552), .A(n17533), .B(
        n17615), .ZN(n17535) );
  OAI22_X1 U20845 ( .A1(n18492), .A2(n17605), .B1(n17608), .B2(n17890), .ZN(
        n17534) );
  NOR3_X1 U20846 ( .A1(n18828), .A2(n17535), .A3(n17534), .ZN(n17545) );
  AOI21_X1 U20847 ( .B1(n18492), .B2(n17537), .A(n17536), .ZN(n18489) );
  NAND2_X1 U20848 ( .A1(n17547), .A2(n17591), .ZN(n17606) );
  NOR3_X1 U20849 ( .A1(n18489), .A2(n17538), .A3(n17606), .ZN(n17539) );
  AOI221_X1 U20850 ( .B1(n17541), .B2(n19432), .C1(n17540), .C2(
        P3_REIP_REG_6__SCAN_IN), .A(n17539), .ZN(n17544) );
  NOR2_X1 U20851 ( .A1(n10186), .A2(n17607), .ZN(n17542) );
  NOR2_X1 U20852 ( .A1(n17542), .A2(n19399), .ZN(n17612) );
  OAI211_X1 U20853 ( .C1(n17546), .C2(n10186), .A(n18489), .B(n17612), .ZN(
        n17543) );
  NAND3_X1 U20854 ( .A1(n17545), .A2(n17544), .A3(n17543), .ZN(P3_U2665) );
  INV_X1 U20855 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17556) );
  AND2_X1 U20856 ( .A1(n17600), .A2(n17573), .ZN(n17559) );
  AOI21_X1 U20857 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17559), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17549) );
  NAND2_X1 U20858 ( .A1(n18493), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17557) );
  AOI21_X1 U20859 ( .B1(n17556), .B2(n17557), .A(n17546), .ZN(n18501) );
  OAI21_X1 U20860 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17557), .A(
        n17547), .ZN(n17568) );
  XOR2_X1 U20861 ( .A(n18501), .B(n17568), .Z(n17548) );
  OAI22_X1 U20862 ( .A1(n17550), .A2(n17549), .B1(n19399), .B2(n17548), .ZN(
        n17551) );
  AOI211_X1 U20863 ( .C1(n17617), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18828), .B(
        n17551), .ZN(n17555) );
  OAI211_X1 U20864 ( .C1(n17561), .C2(n17553), .A(n17616), .B(n17552), .ZN(
        n17554) );
  OAI211_X1 U20865 ( .C1(n17605), .C2(n17556), .A(n17555), .B(n17554), .ZN(
        P3_U2666) );
  NAND2_X1 U20866 ( .A1(n9836), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17578) );
  INV_X1 U20867 ( .A(n17557), .ZN(n17558) );
  AOI21_X1 U20868 ( .B1(n17566), .B2(n17578), .A(n17558), .ZN(n18510) );
  INV_X1 U20869 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19428) );
  AOI22_X1 U20870 ( .A1(n17560), .A2(n18510), .B1(n17559), .B2(n19428), .ZN(
        n17572) );
  AOI211_X1 U20871 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17582), .A(n17561), .B(
        n17615), .ZN(n17565) );
  NOR2_X1 U20872 ( .A1(n17562), .A2(n19551), .ZN(n17618) );
  OAI21_X1 U20873 ( .B1(n17763), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n17618), .ZN(n17563) );
  OAI211_X1 U20874 ( .C1(n17566), .C2(n17605), .A(n18833), .B(n17563), .ZN(
        n17564) );
  AOI211_X1 U20875 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17617), .A(n17565), .B(
        n17564), .ZN(n17571) );
  NAND2_X1 U20876 ( .A1(n9836), .A2(n17566), .ZN(n18518) );
  OAI22_X1 U20877 ( .A1(n18510), .A2(n17568), .B1(n17567), .B2(n18518), .ZN(
        n17569) );
  OAI21_X1 U20878 ( .B1(n17573), .B2(n17609), .A(n17620), .ZN(n17580) );
  AOI22_X1 U20879 ( .A1(n17591), .A2(n17569), .B1(P3_REIP_REG_4__SCAN_IN), 
        .B2(n17580), .ZN(n17570) );
  NAND3_X1 U20880 ( .A1(n17572), .A2(n17571), .A3(n17570), .ZN(P3_U2667) );
  AOI22_X1 U20881 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17598), .B1(
        n17617), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n17586) );
  NOR2_X1 U20882 ( .A1(n17573), .A2(n17609), .ZN(n17575) );
  NOR2_X1 U20883 ( .A1(n19515), .A2(n12306), .ZN(n19339) );
  INV_X1 U20884 ( .A(n19339), .ZN(n19348) );
  NOR2_X1 U20885 ( .A1(n19522), .A2(n19348), .ZN(n19338) );
  INV_X1 U20886 ( .A(n19338), .ZN(n17574) );
  AOI21_X1 U20887 ( .B1(n19499), .B2(n17574), .A(n17763), .ZN(n19495) );
  AOI22_X1 U20888 ( .A1(n17576), .A2(n17575), .B1(n17618), .B2(n19495), .ZN(
        n17585) );
  NAND2_X1 U20889 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17589) );
  INV_X1 U20890 ( .A(n17589), .ZN(n17579) );
  AOI21_X1 U20891 ( .B1(n17579), .B2(n17607), .A(n10186), .ZN(n17590) );
  OAI21_X1 U20892 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17579), .A(
        n17578), .ZN(n18530) );
  XNOR2_X1 U20893 ( .A(n17590), .B(n18530), .ZN(n17581) );
  AOI22_X1 U20894 ( .A1(n17591), .A2(n17581), .B1(P3_REIP_REG_3__SCAN_IN), 
        .B2(n17580), .ZN(n17584) );
  OAI211_X1 U20895 ( .C1(n17587), .C2(n17906), .A(n17616), .B(n17582), .ZN(
        n17583) );
  NAND4_X1 U20896 ( .A1(n17586), .A2(n17585), .A3(n17584), .A4(n17583), .ZN(
        P3_U2668) );
  INV_X1 U20897 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17923) );
  INV_X1 U20898 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17917) );
  NAND2_X1 U20899 ( .A1(n17923), .A2(n17917), .ZN(n17588) );
  AOI211_X1 U20900 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17588), .A(n17587), .B(
        n17615), .ZN(n17597) );
  OAI21_X1 U20901 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17589), .ZN(n18537) );
  AOI21_X1 U20902 ( .B1(n12306), .B2(n19355), .A(n19338), .ZN(n19506) );
  AOI22_X1 U20903 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n17604), .B1(n19506), 
        .B2(n17618), .ZN(n17594) );
  OAI211_X1 U20904 ( .C1(n17592), .C2(n18537), .A(n17591), .B(n17590), .ZN(
        n17593) );
  OAI211_X1 U20905 ( .C1(n17595), .C2(n18537), .A(n17594), .B(n17593), .ZN(
        n17596) );
  AOI211_X1 U20906 ( .C1(n17598), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17597), .B(n17596), .ZN(n17602) );
  OAI211_X1 U20907 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17600), .B(n17599), .ZN(n17601) );
  OAI211_X1 U20908 ( .C1(n17910), .C2(n17608), .A(n17602), .B(n17601), .ZN(
        P3_U2669) );
  OAI21_X1 U20909 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17912), .ZN(n17919) );
  NAND2_X1 U20910 ( .A1(n19355), .A2(n17603), .ZN(n19362) );
  INV_X1 U20911 ( .A(n19362), .ZN(n19512) );
  AOI22_X1 U20912 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17604), .B1(n19512), 
        .B2(n17618), .ZN(n17614) );
  OAI21_X1 U20913 ( .B1(n17607), .B2(n17606), .A(n17605), .ZN(n17611) );
  OAI22_X1 U20914 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17609), .B1(n17608), 
        .B2(n17917), .ZN(n17610) );
  AOI221_X1 U20915 ( .B1(n17612), .B2(n18548), .C1(n17611), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17610), .ZN(n17613) );
  OAI211_X1 U20916 ( .C1(n17615), .C2(n17919), .A(n17614), .B(n17613), .ZN(
        P3_U2670) );
  NOR2_X1 U20917 ( .A1(n17617), .A2(n17616), .ZN(n17623) );
  AOI22_X1 U20918 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17619), .B1(n17618), 
        .B2(n19522), .ZN(n17622) );
  NAND3_X1 U20919 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19497), .A3(
        n17620), .ZN(n17621) );
  OAI211_X1 U20920 ( .C1(n17623), .C2(n17923), .A(n17622), .B(n17621), .ZN(
        P3_U2671) );
  INV_X1 U20921 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17675) );
  NOR2_X1 U20922 ( .A1(n17675), .A2(n17624), .ZN(n17629) );
  NOR4_X1 U20923 ( .A1(n17659), .A2(n17627), .A3(n17626), .A4(n17625), .ZN(
        n17628) );
  NAND4_X1 U20924 ( .A1(n9786), .A2(n17629), .A3(n17660), .A4(n17628), .ZN(
        n17632) );
  NAND2_X1 U20925 ( .A1(n17916), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17631) );
  NAND2_X1 U20926 ( .A1(n17658), .A2(n18929), .ZN(n17630) );
  OAI22_X1 U20927 ( .A1(n17658), .A2(n17631), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17630), .ZN(P3_U2672) );
  NAND2_X1 U20928 ( .A1(n17633), .A2(n17632), .ZN(n17634) );
  NAND2_X1 U20929 ( .A1(n17634), .A2(n17916), .ZN(n17657) );
  AOI22_X1 U20930 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17644) );
  AOI22_X1 U20931 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17643) );
  AOI22_X1 U20932 ( .A1(n16556), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17635) );
  OAI21_X1 U20933 ( .B1(n17877), .B2(n21187), .A(n17635), .ZN(n17641) );
  AOI22_X1 U20934 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17639) );
  AOI22_X1 U20935 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17763), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17638) );
  AOI22_X1 U20936 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17637) );
  AOI22_X1 U20937 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17636) );
  NAND4_X1 U20938 ( .A1(n17639), .A2(n17638), .A3(n17637), .A4(n17636), .ZN(
        n17640) );
  AOI211_X1 U20939 ( .C1(n17879), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17641), .B(n17640), .ZN(n17642) );
  NAND3_X1 U20940 ( .A1(n17644), .A2(n17643), .A3(n17642), .ZN(n17656) );
  AOI22_X1 U20941 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17648) );
  AOI22_X1 U20942 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17647) );
  AOI22_X1 U20943 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17646) );
  AOI22_X1 U20944 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12130), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17645) );
  NAND4_X1 U20945 ( .A1(n17648), .A2(n17647), .A3(n17646), .A4(n17645), .ZN(
        n17654) );
  AOI22_X1 U20946 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17652) );
  AOI22_X1 U20947 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17651) );
  AOI22_X1 U20948 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U20949 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17649) );
  NAND4_X1 U20950 ( .A1(n17652), .A2(n17651), .A3(n17650), .A4(n17649), .ZN(
        n17653) );
  NOR2_X1 U20951 ( .A1(n17654), .A2(n17653), .ZN(n17663) );
  NOR3_X1 U20952 ( .A1(n17663), .A2(n17661), .A3(n17662), .ZN(n17655) );
  XNOR2_X1 U20953 ( .A(n17656), .B(n17655), .ZN(n17930) );
  OAI22_X1 U20954 ( .A1(n17658), .A2(n17657), .B1(n17930), .B2(n17916), .ZN(
        P3_U2673) );
  NAND2_X1 U20955 ( .A1(n17660), .A2(n17659), .ZN(n17667) );
  NOR2_X1 U20956 ( .A1(n17662), .A2(n17661), .ZN(n17664) );
  XNOR2_X1 U20957 ( .A(n17664), .B(n17663), .ZN(n17934) );
  OAI21_X1 U20958 ( .B1(n17672), .B2(n17667), .A(n17666), .ZN(P3_U2674) );
  AOI21_X1 U20959 ( .B1(n17669), .B2(n17947), .A(n17668), .ZN(n17943) );
  NAND2_X1 U20960 ( .A1(n17921), .A2(n17943), .ZN(n17670) );
  OAI221_X1 U20961 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17672), .C1(n17671), 
        .C2(n17674), .A(n17670), .ZN(P3_U2676) );
  NAND2_X1 U20962 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17684), .ZN(n17677) );
  OAI211_X1 U20963 ( .C1(n17949), .C2(n17948), .A(n17921), .B(n17947), .ZN(
        n17673) );
  OAI221_X1 U20964 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17677), .C1(n17675), 
        .C2(n17674), .A(n17673), .ZN(P3_U2677) );
  XNOR2_X1 U20965 ( .A(n17676), .B(n17680), .ZN(n17958) );
  OAI211_X1 U20966 ( .C1(n17684), .C2(P3_EBX_REG_25__SCAN_IN), .A(n17916), .B(
        n17677), .ZN(n17678) );
  OAI21_X1 U20967 ( .B1(n17958), .B2(n17916), .A(n17678), .ZN(P3_U2678) );
  INV_X1 U20968 ( .A(n17679), .ZN(n17689) );
  AOI21_X1 U20969 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17916), .A(n17689), .ZN(
        n17683) );
  OAI21_X1 U20970 ( .B1(n17682), .B2(n17681), .A(n17680), .ZN(n17963) );
  OAI22_X1 U20971 ( .A1(n17684), .A2(n17683), .B1(n17916), .B2(n17963), .ZN(
        P3_U2679) );
  AOI21_X1 U20972 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17916), .A(n17685), .ZN(
        n17688) );
  XNOR2_X1 U20973 ( .A(n17687), .B(n17686), .ZN(n17968) );
  OAI22_X1 U20974 ( .A1(n17689), .A2(n17688), .B1(n17916), .B2(n17968), .ZN(
        P3_U2680) );
  AOI22_X1 U20975 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17693) );
  AOI22_X1 U20976 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17692) );
  AOI22_X1 U20977 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17691) );
  AOI22_X1 U20978 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17690) );
  NAND4_X1 U20979 ( .A1(n17693), .A2(n17692), .A3(n17691), .A4(n17690), .ZN(
        n17699) );
  AOI22_X1 U20980 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17697) );
  AOI22_X1 U20981 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17696) );
  AOI22_X1 U20982 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17695) );
  AOI22_X1 U20983 ( .A1(n12105), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17694) );
  NAND4_X1 U20984 ( .A1(n17697), .A2(n17696), .A3(n17695), .A4(n17694), .ZN(
        n17698) );
  NOR2_X1 U20985 ( .A1(n17699), .A2(n17698), .ZN(n17970) );
  NAND3_X1 U20986 ( .A1(n17701), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17916), 
        .ZN(n17700) );
  OAI221_X1 U20987 ( .B1(n17701), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17916), 
        .C2(n17970), .A(n17700), .ZN(P3_U2681) );
  AOI21_X1 U20988 ( .B1(n17703), .B2(n17702), .A(n17921), .ZN(n17704) );
  INV_X1 U20989 ( .A(n17704), .ZN(n17715) );
  AOI22_X1 U20990 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17708) );
  AOI22_X1 U20991 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17763), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17707) );
  AOI22_X1 U20992 ( .A1(n9698), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17706) );
  AOI22_X1 U20993 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17705) );
  NAND4_X1 U20994 ( .A1(n17708), .A2(n17707), .A3(n17706), .A4(n17705), .ZN(
        n17714) );
  AOI22_X1 U20995 ( .A1(n17857), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17712) );
  AOI22_X1 U20996 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17711) );
  AOI22_X1 U20997 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17710) );
  AOI22_X1 U20998 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17709) );
  NAND4_X1 U20999 ( .A1(n17712), .A2(n17711), .A3(n17710), .A4(n17709), .ZN(
        n17713) );
  NOR2_X1 U21000 ( .A1(n17714), .A2(n17713), .ZN(n17976) );
  OAI22_X1 U21001 ( .A1(n9786), .A2(n17715), .B1(n17976), .B2(n17916), .ZN(
        P3_U2682) );
  NAND2_X1 U21002 ( .A1(n18929), .A2(n17716), .ZN(n17728) );
  NOR2_X1 U21003 ( .A1(n17921), .A2(n17716), .ZN(n17740) );
  AOI22_X1 U21004 ( .A1(n12105), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17726) );
  AOI22_X1 U21005 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17725) );
  INV_X1 U21006 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n21152) );
  AOI22_X1 U21007 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17717) );
  OAI21_X1 U21008 ( .B1(n9754), .B2(n21152), .A(n17717), .ZN(n17723) );
  AOI22_X1 U21009 ( .A1(n17820), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17721) );
  AOI22_X1 U21010 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17720) );
  AOI22_X1 U21011 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9698), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17719) );
  AOI22_X1 U21012 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12130), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17718) );
  NAND4_X1 U21013 ( .A1(n17721), .A2(n17720), .A3(n17719), .A4(n17718), .ZN(
        n17722) );
  AOI211_X1 U21014 ( .C1(n17859), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n17723), .B(n17722), .ZN(n17724) );
  NAND3_X1 U21015 ( .A1(n17726), .A2(n17725), .A3(n17724), .ZN(n17980) );
  AOI22_X1 U21016 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17740), .B1(n17921), 
        .B2(n17980), .ZN(n17727) );
  OAI21_X1 U21017 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17728), .A(n17727), .ZN(
        P3_U2683) );
  AOI22_X1 U21018 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17820), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17732) );
  AOI22_X1 U21019 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17731) );
  AOI22_X1 U21020 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17730) );
  AOI22_X1 U21021 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9695), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17729) );
  NAND4_X1 U21022 ( .A1(n17732), .A2(n17731), .A3(n17730), .A4(n17729), .ZN(
        n17738) );
  AOI22_X1 U21023 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17736) );
  AOI22_X1 U21024 ( .A1(n12105), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17735) );
  AOI22_X1 U21025 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17734) );
  AOI22_X1 U21026 ( .A1(n17879), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17733) );
  NAND4_X1 U21027 ( .A1(n17736), .A2(n17735), .A3(n17734), .A4(n17733), .ZN(
        n17737) );
  NOR2_X1 U21028 ( .A1(n17738), .A2(n17737), .ZN(n17988) );
  INV_X1 U21029 ( .A(n17739), .ZN(n17741) );
  OAI21_X1 U21030 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17741), .A(n17740), .ZN(
        n17742) );
  OAI21_X1 U21031 ( .B1(n17988), .B2(n17916), .A(n17742), .ZN(P3_U2684) );
  NAND2_X1 U21032 ( .A1(n18929), .A2(n17743), .ZN(n17757) );
  NOR2_X1 U21033 ( .A1(n17921), .A2(n17743), .ZN(n17770) );
  AOI22_X1 U21034 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17755) );
  AOI22_X1 U21035 ( .A1(n12105), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17826), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17754) );
  AOI22_X1 U21036 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17744) );
  OAI21_X1 U21037 ( .B1(n17745), .B2(n21247), .A(n17744), .ZN(n17751) );
  AOI22_X1 U21038 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U21039 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17857), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17748) );
  AOI22_X1 U21040 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17747) );
  AOI22_X1 U21041 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17746) );
  NAND4_X1 U21042 ( .A1(n17749), .A2(n17748), .A3(n17747), .A4(n17746), .ZN(
        n17750) );
  AOI211_X1 U21043 ( .C1(n17752), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n17751), .B(n17750), .ZN(n17753) );
  NAND3_X1 U21044 ( .A1(n17755), .A2(n17754), .A3(n17753), .ZN(n17989) );
  AOI22_X1 U21045 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17770), .B1(n17921), 
        .B2(n17989), .ZN(n17756) );
  OAI21_X1 U21046 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17757), .A(n17756), .ZN(
        P3_U2685) );
  AOI22_X1 U21047 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n16556), .ZN(n17762) );
  AOI22_X1 U21048 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12128), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17761) );
  AOI22_X1 U21049 ( .A1(n9698), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17857), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17760) );
  AOI22_X1 U21050 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12130), .B1(
        n17758), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17759) );
  NAND4_X1 U21051 ( .A1(n17762), .A2(n17761), .A3(n17760), .A4(n17759), .ZN(
        n17769) );
  AOI22_X1 U21052 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12175), .B1(
        n17875), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17767) );
  AOI22_X1 U21053 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n9696), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17766) );
  AOI22_X1 U21054 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12093), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17765) );
  AOI22_X1 U21055 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17763), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17860), .ZN(n17764) );
  NAND4_X1 U21056 ( .A1(n17767), .A2(n17766), .A3(n17765), .A4(n17764), .ZN(
        n17768) );
  NOR2_X1 U21057 ( .A1(n17769), .A2(n17768), .ZN(n17999) );
  OAI21_X1 U21058 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n10032), .A(n17770), .ZN(
        n17771) );
  OAI21_X1 U21059 ( .B1(n17999), .B2(n17916), .A(n17771), .ZN(P3_U2686) );
  AOI22_X1 U21060 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9698), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17775) );
  AOI22_X1 U21061 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17857), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17774) );
  AOI22_X1 U21062 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17773) );
  AOI22_X1 U21063 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17772) );
  NAND4_X1 U21064 ( .A1(n17775), .A2(n17774), .A3(n17773), .A4(n17772), .ZN(
        n17781) );
  AOI22_X1 U21065 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17779) );
  AOI22_X1 U21066 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17778) );
  AOI22_X1 U21067 ( .A1(n17820), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17777) );
  AOI22_X1 U21068 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17826), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17776) );
  NAND4_X1 U21069 ( .A1(n17779), .A2(n17778), .A3(n17777), .A4(n17776), .ZN(
        n17780) );
  NOR2_X1 U21070 ( .A1(n17781), .A2(n17780), .ZN(n18005) );
  OAI21_X1 U21071 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17796), .A(n17782), .ZN(
        n17783) );
  AOI22_X1 U21072 ( .A1(n17921), .A2(n18005), .B1(n17783), .B2(n17916), .ZN(
        P3_U2687) );
  OAI21_X1 U21073 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17784), .A(n17916), .ZN(
        n17795) );
  AOI22_X1 U21074 ( .A1(n17752), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17788) );
  AOI22_X1 U21075 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17826), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17787) );
  AOI22_X1 U21076 ( .A1(n17844), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17786) );
  AOI22_X1 U21077 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17785) );
  NAND4_X1 U21078 ( .A1(n17788), .A2(n17787), .A3(n17786), .A4(n17785), .ZN(
        n17794) );
  AOI22_X1 U21079 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17857), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17792) );
  AOI22_X1 U21080 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17797), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17791) );
  AOI22_X1 U21081 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17820), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17790) );
  AOI22_X1 U21082 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17789) );
  NAND4_X1 U21083 ( .A1(n17792), .A2(n17791), .A3(n17790), .A4(n17789), .ZN(
        n17793) );
  NOR2_X1 U21084 ( .A1(n17794), .A2(n17793), .ZN(n18009) );
  OAI22_X1 U21085 ( .A1(n17796), .A2(n17795), .B1(n18009), .B2(n17916), .ZN(
        P3_U2688) );
  AOI22_X1 U21086 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17820), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17807) );
  AOI22_X1 U21087 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17806) );
  AOI22_X1 U21088 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17857), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17798) );
  OAI21_X1 U21089 ( .B1(n17877), .B2(n18925), .A(n17798), .ZN(n17804) );
  AOI22_X1 U21090 ( .A1(n16555), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17802) );
  AOI22_X1 U21091 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17801) );
  AOI22_X1 U21092 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17800) );
  AOI22_X1 U21093 ( .A1(n12175), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17826), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17799) );
  NAND4_X1 U21094 ( .A1(n17802), .A2(n17801), .A3(n17800), .A4(n17799), .ZN(
        n17803) );
  AOI211_X1 U21095 ( .C1(n17859), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n17804), .B(n17803), .ZN(n17805) );
  NAND3_X1 U21096 ( .A1(n17807), .A2(n17806), .A3(n17805), .ZN(n18010) );
  NOR3_X1 U21097 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17969), .A3(n17808), .ZN(
        n17809) );
  AOI21_X1 U21098 ( .B1(n17921), .B2(n18010), .A(n17809), .ZN(n17810) );
  OAI21_X1 U21099 ( .B1(n17812), .B2(n17811), .A(n17810), .ZN(P3_U2689) );
  AOI22_X1 U21100 ( .A1(n12105), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17855), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17823) );
  AOI22_X1 U21101 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16556), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17822) );
  INV_X1 U21102 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n21173) );
  AOI22_X1 U21103 ( .A1(n17826), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17813) );
  OAI21_X1 U21104 ( .B1(n17877), .B2(n21173), .A(n17813), .ZN(n17819) );
  AOI22_X1 U21105 ( .A1(n9698), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17817) );
  AOI22_X1 U21106 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17816) );
  AOI22_X1 U21107 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17857), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17815) );
  AOI22_X1 U21108 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17814) );
  NAND4_X1 U21109 ( .A1(n17817), .A2(n17816), .A3(n17815), .A4(n17814), .ZN(
        n17818) );
  AOI211_X1 U21110 ( .C1(n17820), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n17819), .B(n17818), .ZN(n17821) );
  NAND3_X1 U21111 ( .A1(n17823), .A2(n17822), .A3(n17821), .ZN(n18018) );
  INV_X1 U21112 ( .A(n18018), .ZN(n17825) );
  OAI21_X1 U21113 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17838), .A(n9784), .ZN(
        n17824) );
  AOI22_X1 U21114 ( .A1(n17921), .A2(n17825), .B1(n17824), .B2(n17916), .ZN(
        P3_U2691) );
  OAI21_X1 U21115 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17852), .A(n17916), .ZN(
        n17837) );
  AOI22_X1 U21116 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17857), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17830) );
  AOI22_X1 U21117 ( .A1(n17758), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17829) );
  AOI22_X1 U21118 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12130), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17828) );
  AOI22_X1 U21119 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17826), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17827) );
  NAND4_X1 U21120 ( .A1(n17830), .A2(n17829), .A3(n17828), .A4(n17827), .ZN(
        n17836) );
  AOI22_X1 U21121 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17834) );
  AOI22_X1 U21122 ( .A1(n17820), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17833) );
  AOI22_X1 U21123 ( .A1(n12105), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17832) );
  AOI22_X1 U21124 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17831) );
  NAND4_X1 U21125 ( .A1(n17834), .A2(n17833), .A3(n17832), .A4(n17831), .ZN(
        n17835) );
  NOR2_X1 U21126 ( .A1(n17836), .A2(n17835), .ZN(n18022) );
  OAI22_X1 U21127 ( .A1(n17838), .A2(n17837), .B1(n18022), .B2(n17916), .ZN(
        P3_U2692) );
  AOI22_X1 U21128 ( .A1(n18929), .A2(n17853), .B1(P3_EBX_REG_10__SCAN_IN), 
        .B2(n17916), .ZN(n17851) );
  AOI22_X1 U21129 ( .A1(n17879), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17843) );
  AOI22_X1 U21130 ( .A1(n17856), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17842) );
  AOI22_X1 U21131 ( .A1(n12128), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17841) );
  AOI22_X1 U21132 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17839), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17840) );
  NAND4_X1 U21133 ( .A1(n17843), .A2(n17842), .A3(n17841), .A4(n17840), .ZN(
        n17850) );
  AOI22_X1 U21134 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17844), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17848) );
  AOI22_X1 U21135 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17847) );
  AOI22_X1 U21136 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17846) );
  AOI22_X1 U21137 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17845) );
  NAND4_X1 U21138 ( .A1(n17848), .A2(n17847), .A3(n17846), .A4(n17845), .ZN(
        n17849) );
  NOR2_X1 U21139 ( .A1(n17850), .A2(n17849), .ZN(n18029) );
  OAI22_X1 U21140 ( .A1(n17852), .A2(n17851), .B1(n18029), .B2(n17916), .ZN(
        P3_U2693) );
  INV_X1 U21141 ( .A(n17853), .ZN(n17871) );
  AOI21_X1 U21142 ( .B1(n17854), .B2(n17891), .A(n17921), .ZN(n17870) );
  AOI22_X1 U21143 ( .A1(n17855), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n9696), .ZN(n17869) );
  AOI22_X1 U21144 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17873), .B1(
        n17856), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17868) );
  AOI22_X1 U21145 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17857), .B1(
        n17752), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17858) );
  OAI21_X1 U21146 ( .B1(n21120), .B2(n12221), .A(n17858), .ZN(n17866) );
  AOI22_X1 U21147 ( .A1(n17839), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n9697), .ZN(n17864) );
  AOI22_X1 U21148 ( .A1(n17859), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n16555), .ZN(n17863) );
  AOI22_X1 U21149 ( .A1(n17820), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17862) );
  AOI22_X1 U21150 ( .A1(n17797), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17860), .ZN(n17861) );
  NAND4_X1 U21151 ( .A1(n17864), .A2(n17863), .A3(n17862), .A4(n17861), .ZN(
        n17865) );
  AOI211_X1 U21152 ( .C1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .C2(n17826), .A(
        n17866), .B(n17865), .ZN(n17867) );
  NAND3_X1 U21153 ( .A1(n17869), .A2(n17868), .A3(n17867), .ZN(n18030) );
  AOI22_X1 U21154 ( .A1(n17871), .A2(n17870), .B1(n18030), .B2(n17921), .ZN(
        n17872) );
  INV_X1 U21155 ( .A(n17872), .ZN(P3_U2694) );
  AOI22_X1 U21156 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17873), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17889) );
  AOI22_X1 U21157 ( .A1(n17875), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17874), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17888) );
  AOI22_X1 U21158 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16555), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17876) );
  OAI21_X1 U21159 ( .B1(n17877), .B2(n18897), .A(n17876), .ZN(n17886) );
  AOI22_X1 U21160 ( .A1(n17758), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12216), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17884) );
  AOI22_X1 U21161 ( .A1(n17878), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12175), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17883) );
  AOI22_X1 U21162 ( .A1(n17763), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17879), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17882) );
  AOI22_X1 U21163 ( .A1(n17880), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12093), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17881) );
  NAND4_X1 U21164 ( .A1(n17884), .A2(n17883), .A3(n17882), .A4(n17881), .ZN(
        n17885) );
  AOI211_X1 U21165 ( .C1(n17826), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n17886), .B(n17885), .ZN(n17887) );
  NAND3_X1 U21166 ( .A1(n17889), .A2(n17888), .A3(n17887), .ZN(n18033) );
  INV_X1 U21167 ( .A(n18033), .ZN(n17893) );
  NOR3_X1 U21168 ( .A1(n17969), .A2(n17890), .A3(n17896), .ZN(n17898) );
  OAI221_X1 U21169 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(P3_EBX_REG_7__SCAN_IN), 
        .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17898), .A(n17891), .ZN(n17892) );
  AOI22_X1 U21170 ( .A1(n17921), .A2(n17893), .B1(n17892), .B2(n17916), .ZN(
        P3_U2695) );
  AOI21_X1 U21171 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17916), .A(n17898), .ZN(
        n17894) );
  INV_X1 U21172 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18932) );
  OAI22_X1 U21173 ( .A1(n17895), .A2(n17894), .B1(n18932), .B2(n17916), .ZN(
        P3_U2696) );
  NOR2_X1 U21174 ( .A1(n17969), .A2(n17896), .ZN(n17901) );
  AOI21_X1 U21175 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17916), .A(n17901), .ZN(
        n17897) );
  OAI22_X1 U21176 ( .A1(n17898), .A2(n17897), .B1(n18925), .B2(n17916), .ZN(
        P3_U2697) );
  OAI21_X1 U21177 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17899), .A(n17916), .ZN(
        n17900) );
  INV_X1 U21178 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18920) );
  OAI22_X1 U21179 ( .A1(n17901), .A2(n17900), .B1(n18920), .B2(n17916), .ZN(
        P3_U2698) );
  NAND2_X1 U21180 ( .A1(n17902), .A2(n17920), .ZN(n17913) );
  NOR2_X1 U21181 ( .A1(n17906), .A2(n17913), .ZN(n17909) );
  AOI21_X1 U21182 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17916), .A(n17909), .ZN(
        n17905) );
  NOR2_X1 U21183 ( .A1(n17903), .A2(n17918), .ZN(n17904) );
  OAI22_X1 U21184 ( .A1(n17905), .A2(n17904), .B1(n21173), .B2(n17916), .ZN(
        P3_U2699) );
  OAI21_X1 U21185 ( .B1(n17906), .B2(n17921), .A(n17913), .ZN(n17907) );
  INV_X1 U21186 ( .A(n17907), .ZN(n17908) );
  INV_X1 U21187 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18912) );
  OAI22_X1 U21188 ( .A1(n17909), .A2(n17908), .B1(n18912), .B2(n17916), .ZN(
        P3_U2700) );
  OAI221_X1 U21189 ( .B1(n17912), .B2(n17911), .C1(n18929), .C2(n17911), .A(
        n17910), .ZN(n17914) );
  OAI211_X1 U21190 ( .C1(n17916), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17914), .B(n17913), .ZN(n17915) );
  INV_X1 U21191 ( .A(n17915), .ZN(P3_U2701) );
  INV_X1 U21192 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18902) );
  OAI222_X1 U21193 ( .A1(n17919), .A2(n17918), .B1(n17917), .B2(n17924), .C1(
        n18902), .C2(n17916), .ZN(P3_U2702) );
  AOI22_X1 U21194 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17921), .B1(
        n17920), .B2(n17923), .ZN(n17922) );
  OAI21_X1 U21195 ( .B1(n17924), .B2(n17923), .A(n17922), .ZN(P3_U2703) );
  INV_X1 U21196 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18080) );
  INV_X1 U21197 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n21123) );
  INV_X1 U21198 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n21203) );
  INV_X1 U21199 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18177) );
  INV_X1 U21200 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n21139) );
  NAND3_X1 U21201 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n18040) );
  NAND4_X1 U21202 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_5__SCAN_IN), .ZN(n17925) );
  INV_X1 U21203 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18098) );
  INV_X1 U21204 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18138) );
  INV_X1 U21205 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18148) );
  OR2_X1 U21206 ( .A1(n17935), .A2(n18148), .ZN(n17929) );
  NAND2_X1 U21207 ( .A1(n17926), .A2(n18063), .ZN(n17994) );
  NAND2_X1 U21208 ( .A1(n18060), .A2(n17935), .ZN(n17933) );
  OAI21_X1 U21209 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18064), .A(n17933), .ZN(
        n17927) );
  AOI22_X1 U21210 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18000), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17927), .ZN(n17928) );
  OAI21_X1 U21211 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17929), .A(n17928), .ZN(
        P3_U2704) );
  NAND2_X1 U21212 ( .A1(n18917), .A2(n18063), .ZN(n17975) );
  OAI22_X1 U21213 ( .A1(n17930), .A2(n18052), .B1(n19894), .B2(n17994), .ZN(
        n17931) );
  AOI21_X1 U21214 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18001), .A(n17931), .ZN(
        n17932) );
  OAI221_X1 U21215 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17935), .C1(n18148), 
        .C2(n17933), .A(n17932), .ZN(P3_U2705) );
  AOI22_X1 U21216 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18000), .B1(n17934), .B2(
        n18067), .ZN(n17938) );
  OAI211_X1 U21217 ( .C1(n17936), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18060), .B(
        n17935), .ZN(n17937) );
  OAI211_X1 U21218 ( .C1(n17975), .C2(n21221), .A(n17938), .B(n17937), .ZN(
        P3_U2706) );
  INV_X1 U21219 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18170) );
  AOI22_X1 U21220 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18000), .B1(n17939), .B2(
        n18067), .ZN(n17942) );
  OAI211_X1 U21221 ( .C1(n9787), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18060), .B(
        n17940), .ZN(n17941) );
  OAI211_X1 U21222 ( .C1(n17975), .C2(n18170), .A(n17942), .B(n17941), .ZN(
        P3_U2707) );
  INV_X1 U21223 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n21078) );
  AOI22_X1 U21224 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18001), .B1(n17943), .B2(
        n18067), .ZN(n17946) );
  AOI211_X1 U21225 ( .C1(n18080), .C2(n17950), .A(n9787), .B(n18063), .ZN(
        n17944) );
  INV_X1 U21226 ( .A(n17944), .ZN(n17945) );
  OAI211_X1 U21227 ( .C1(n17994), .C2(n21078), .A(n17946), .B(n17945), .ZN(
        P3_U2708) );
  OAI21_X1 U21228 ( .B1(n17949), .B2(n17948), .A(n17947), .ZN(n17953) );
  AOI22_X1 U21229 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18001), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18000), .ZN(n17952) );
  OAI211_X1 U21230 ( .C1(n17954), .C2(P3_EAX_REG_26__SCAN_IN), .A(n18060), .B(
        n17950), .ZN(n17951) );
  OAI211_X1 U21231 ( .C1(n18052), .C2(n17953), .A(n17952), .B(n17951), .ZN(
        P3_U2709) );
  AOI22_X1 U21232 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18001), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18000), .ZN(n17957) );
  AOI211_X1 U21233 ( .C1(n21123), .C2(n17959), .A(n17954), .B(n18063), .ZN(
        n17955) );
  INV_X1 U21234 ( .A(n17955), .ZN(n17956) );
  OAI211_X1 U21235 ( .C1(n18052), .C2(n17958), .A(n17957), .B(n17956), .ZN(
        P3_U2710) );
  AOI22_X1 U21236 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18001), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18000), .ZN(n17962) );
  OAI211_X1 U21237 ( .C1(n17960), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18060), .B(
        n17959), .ZN(n17961) );
  OAI211_X1 U21238 ( .C1(n18052), .C2(n17963), .A(n17962), .B(n17961), .ZN(
        P3_U2711) );
  AOI22_X1 U21239 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18001), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18000), .ZN(n17967) );
  OAI211_X1 U21240 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17965), .A(n18060), .B(
        n17964), .ZN(n17966) );
  OAI211_X1 U21241 ( .C1(n18052), .C2(n17968), .A(n17967), .B(n17966), .ZN(
        P3_U2712) );
  INV_X1 U21242 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18131) );
  INV_X1 U21243 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18129) );
  NAND2_X1 U21244 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17990), .ZN(n17985) );
  NAND2_X1 U21245 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17981), .ZN(n17979) );
  NAND2_X1 U21246 ( .A1(n18060), .A2(n17979), .ZN(n17984) );
  OAI21_X1 U21247 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18064), .A(n17984), .ZN(
        n17972) );
  OAI22_X1 U21248 ( .A1(n17970), .A2(n18052), .B1(n16122), .B2(n17994), .ZN(
        n17971) );
  AOI21_X1 U21249 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n17972), .A(n17971), .ZN(
        n17974) );
  INV_X1 U21250 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18136) );
  OR3_X1 U21251 ( .A1(n18136), .A2(n17979), .A3(P3_EAX_REG_22__SCAN_IN), .ZN(
        n17973) );
  OAI211_X1 U21252 ( .C1(n17975), .C2(n18921), .A(n17974), .B(n17973), .ZN(
        P3_U2713) );
  OAI22_X1 U21253 ( .A1(n17976), .A2(n18052), .B1(n16133), .B2(n17994), .ZN(
        n17977) );
  AOI21_X1 U21254 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n18001), .A(n17977), .ZN(
        n17978) );
  OAI221_X1 U21255 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17979), .C1(n18136), 
        .C2(n17984), .A(n17978), .ZN(P3_U2714) );
  INV_X1 U21256 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18134) );
  AOI22_X1 U21257 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18000), .B1(n18067), .B2(
        n17980), .ZN(n17983) );
  AOI22_X1 U21258 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18001), .B1(n17981), .B2(
        n18134), .ZN(n17982) );
  OAI211_X1 U21259 ( .C1(n18134), .C2(n17984), .A(n17983), .B(n17982), .ZN(
        P3_U2715) );
  AOI22_X1 U21260 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18001), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18000), .ZN(n17987) );
  OAI211_X1 U21261 ( .C1(n17990), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18060), .B(
        n17985), .ZN(n17986) );
  OAI211_X1 U21262 ( .C1(n17988), .C2(n18052), .A(n17987), .B(n17986), .ZN(
        P3_U2716) );
  AOI22_X1 U21263 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18001), .B1(n18067), .B2(
        n17989), .ZN(n17993) );
  AOI211_X1 U21264 ( .C1(n18131), .C2(n17995), .A(n17990), .B(n18063), .ZN(
        n17991) );
  INV_X1 U21265 ( .A(n17991), .ZN(n17992) );
  OAI211_X1 U21266 ( .C1(n17994), .C2(n16157), .A(n17993), .B(n17992), .ZN(
        P3_U2717) );
  AOI22_X1 U21267 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18001), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18000), .ZN(n17998) );
  INV_X1 U21268 ( .A(n18002), .ZN(n17996) );
  OAI211_X1 U21269 ( .C1(n17996), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18060), .B(
        n17995), .ZN(n17997) );
  OAI211_X1 U21270 ( .C1(n17999), .C2(n18052), .A(n17998), .B(n17997), .ZN(
        P3_U2718) );
  AOI22_X1 U21271 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18001), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18000), .ZN(n18004) );
  OAI211_X1 U21272 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18006), .A(n18060), .B(
        n18002), .ZN(n18003) );
  OAI211_X1 U21273 ( .C1(n18005), .C2(n18052), .A(n18004), .B(n18003), .ZN(
        P3_U2719) );
  AOI21_X1 U21274 ( .B1(n18177), .B2(n18011), .A(n18006), .ZN(n18007) );
  AOI22_X1 U21275 ( .A1(n18068), .A2(BUF2_REG_15__SCAN_IN), .B1(n18007), .B2(
        n18060), .ZN(n18008) );
  OAI21_X1 U21276 ( .B1(n18009), .B2(n18052), .A(n18008), .ZN(P3_U2720) );
  AOI22_X1 U21277 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18068), .B1(n18067), .B2(
        n18010), .ZN(n18014) );
  OAI211_X1 U21278 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n18012), .A(n18060), .B(
        n18011), .ZN(n18013) );
  NAND2_X1 U21279 ( .A1(n18014), .A2(n18013), .ZN(P3_U2721) );
  INV_X1 U21280 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18164) );
  NAND4_X1 U21281 ( .A1(n18929), .A2(P3_EAX_REG_7__SCAN_IN), .A3(n18043), .A4(
        P3_EAX_REG_8__SCAN_IN), .ZN(n18032) );
  OR2_X1 U21282 ( .A1(n18164), .A2(n18032), .ZN(n18026) );
  NOR2_X1 U21283 ( .A1(n21139), .A2(n18026), .ZN(n18025) );
  NAND3_X1 U21284 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(n18025), .ZN(n18017) );
  NAND2_X1 U21285 ( .A1(n18060), .A2(n18017), .ZN(n18020) );
  AOI22_X1 U21286 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18068), .B1(n18067), .B2(
        n18015), .ZN(n18016) );
  OAI221_X1 U21287 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18017), .C1(n18098), 
        .C2(n18020), .A(n18016), .ZN(P3_U2722) );
  NAND2_X1 U21288 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18025), .ZN(n18021) );
  INV_X1 U21289 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18100) );
  AOI22_X1 U21290 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18068), .B1(n18067), .B2(
        n18018), .ZN(n18019) );
  OAI221_X1 U21291 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18021), .C1(n18100), 
        .C2(n18020), .A(n18019), .ZN(P3_U2723) );
  INV_X1 U21292 ( .A(n18068), .ZN(n18055) );
  INV_X1 U21293 ( .A(n18021), .ZN(n18024) );
  AOI21_X1 U21294 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18060), .A(n18025), .ZN(
        n18023) );
  OAI222_X1 U21295 ( .A1(n18055), .A2(n18168), .B1(n18024), .B2(n18023), .C1(
        n18052), .C2(n18022), .ZN(P3_U2724) );
  AOI21_X1 U21296 ( .B1(n21139), .B2(n18026), .A(n18025), .ZN(n18027) );
  AOI22_X1 U21297 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18068), .B1(n18027), .B2(
        n18060), .ZN(n18028) );
  OAI21_X1 U21298 ( .B1(n18029), .B2(n18052), .A(n18028), .ZN(P3_U2725) );
  NAND2_X1 U21299 ( .A1(n18060), .A2(n18032), .ZN(n18035) );
  AOI22_X1 U21300 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18068), .B1(n18067), .B2(
        n18030), .ZN(n18031) );
  OAI221_X1 U21301 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18032), .C1(n18164), 
        .C2(n18035), .A(n18031), .ZN(P3_U2726) );
  INV_X1 U21302 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18107) );
  AOI22_X1 U21303 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18068), .B1(n18067), .B2(
        n18033), .ZN(n18034) );
  OAI221_X1 U21304 ( .B1(n18035), .B2(n18037), .C1(n18035), .C2(n18107), .A(
        n18034), .ZN(P3_U2727) );
  AOI22_X1 U21305 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18068), .B1(n18067), .B2(
        n18036), .ZN(n18039) );
  OAI211_X1 U21306 ( .C1(P3_EAX_REG_7__SCAN_IN), .C2(n18043), .A(n18060), .B(
        n18037), .ZN(n18038) );
  NAND2_X1 U21307 ( .A1(n18039), .A2(n18038), .ZN(P3_U2728) );
  INV_X1 U21308 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21047) );
  INV_X1 U21309 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18115) );
  NOR2_X1 U21310 ( .A1(n18040), .A2(n18064), .ZN(n18050) );
  INV_X1 U21311 ( .A(n18050), .ZN(n18059) );
  NOR3_X1 U21312 ( .A1(n21047), .A2(n18115), .A3(n18059), .ZN(n18049) );
  AND2_X1 U21313 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18049), .ZN(n18046) );
  AOI21_X1 U21314 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18060), .A(n18046), .ZN(
        n18042) );
  OAI222_X1 U21315 ( .A1(n18055), .A2(n18921), .B1(n18043), .B2(n18042), .C1(
        n18052), .C2(n18041), .ZN(P3_U2729) );
  AOI21_X1 U21316 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18060), .A(n18049), .ZN(
        n18045) );
  OAI222_X1 U21317 ( .A1(n21293), .A2(n18055), .B1(n18046), .B2(n18045), .C1(
        n18052), .C2(n18044), .ZN(P3_U2730) );
  INV_X1 U21318 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18913) );
  AOI22_X1 U21319 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18060), .B1(
        P3_EAX_REG_3__SCAN_IN), .B2(n18050), .ZN(n18048) );
  OAI222_X1 U21320 ( .A1(n18913), .A2(n18055), .B1(n18049), .B2(n18048), .C1(
        n18052), .C2(n18047), .ZN(P3_U2731) );
  NOR2_X1 U21321 ( .A1(n18115), .A2(n18059), .ZN(n18054) );
  AOI21_X1 U21322 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18060), .A(n18050), .ZN(
        n18053) );
  OAI222_X1 U21323 ( .A1(n18908), .A2(n18055), .B1(n18054), .B2(n18053), .C1(
        n18052), .C2(n18051), .ZN(P3_U2732) );
  AOI22_X1 U21324 ( .A1(n18068), .A2(BUF2_REG_2__SCAN_IN), .B1(n18067), .B2(
        n18056), .ZN(n18062) );
  NAND2_X1 U21325 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n18057) );
  NOR2_X1 U21326 ( .A1(n18058), .A2(n18057), .ZN(n18071) );
  OAI211_X1 U21327 ( .C1(P3_EAX_REG_2__SCAN_IN), .C2(n18071), .A(n18060), .B(
        n18059), .ZN(n18061) );
  NAND2_X1 U21328 ( .A1(n18062), .A2(n18061), .ZN(P3_U2733) );
  INV_X1 U21329 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18152) );
  AOI221_X1 U21330 ( .B1(n18152), .B2(n18150), .C1(n18152), .C2(n18064), .A(
        n18063), .ZN(n18065) );
  INV_X1 U21331 ( .A(n18065), .ZN(n18070) );
  AOI22_X1 U21332 ( .A1(n18068), .A2(BUF2_REG_1__SCAN_IN), .B1(n18067), .B2(
        n18066), .ZN(n18069) );
  OAI21_X1 U21333 ( .B1(n18071), .B2(n18070), .A(n18069), .ZN(P3_U2734) );
  NAND2_X1 U21334 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18384), .ZN(n18102) );
  NOR2_X1 U21335 ( .A1(n18085), .A2(n18073), .ZN(P3_U2736) );
  NOR2_X1 U21336 ( .A1(n18121), .A2(n18893), .ZN(n18083) );
  INV_X1 U21337 ( .A(n18083), .ZN(n18094) );
  AOI22_X1 U21338 ( .A1(n18119), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18074) );
  OAI21_X1 U21339 ( .B1(n18148), .B2(n18094), .A(n18074), .ZN(P3_U2737) );
  INV_X1 U21340 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18076) );
  AOI22_X1 U21341 ( .A1(n18119), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18075) );
  OAI21_X1 U21342 ( .B1(n18076), .B2(n18094), .A(n18075), .ZN(P3_U2738) );
  INV_X1 U21343 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18078) );
  AOI22_X1 U21344 ( .A1(n18119), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18077) );
  OAI21_X1 U21345 ( .B1(n18078), .B2(n18094), .A(n18077), .ZN(P3_U2739) );
  AOI22_X1 U21346 ( .A1(n18119), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18079) );
  OAI21_X1 U21347 ( .B1(n18080), .B2(n18094), .A(n18079), .ZN(P3_U2740) );
  INV_X1 U21348 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n21237) );
  AOI22_X1 U21349 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18083), .B1(n18119), 
        .B2(P3_UWORD_REG_10__SCAN_IN), .ZN(n18081) );
  OAI21_X1 U21350 ( .B1(n21237), .B2(n18085), .A(n18081), .ZN(P3_U2741) );
  AOI22_X1 U21351 ( .A1(n18119), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18082) );
  OAI21_X1 U21352 ( .B1(n21123), .B2(n18094), .A(n18082), .ZN(P3_U2742) );
  INV_X1 U21353 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n21106) );
  AOI22_X1 U21354 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18083), .B1(n18119), 
        .B2(P3_UWORD_REG_8__SCAN_IN), .ZN(n18084) );
  OAI21_X1 U21355 ( .B1(n21106), .B2(n18085), .A(n18084), .ZN(P3_U2743) );
  INV_X1 U21356 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18140) );
  AOI22_X1 U21357 ( .A1(n18119), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18086) );
  OAI21_X1 U21358 ( .B1(n18140), .B2(n18094), .A(n18086), .ZN(P3_U2744) );
  AOI22_X1 U21359 ( .A1(n18119), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18087) );
  OAI21_X1 U21360 ( .B1(n18138), .B2(n18094), .A(n18087), .ZN(P3_U2745) );
  AOI22_X1 U21361 ( .A1(n18119), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18088) );
  OAI21_X1 U21362 ( .B1(n18136), .B2(n18094), .A(n18088), .ZN(P3_U2746) );
  AOI22_X1 U21363 ( .A1(n18119), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18089) );
  OAI21_X1 U21364 ( .B1(n18134), .B2(n18094), .A(n18089), .ZN(P3_U2747) );
  AOI22_X1 U21365 ( .A1(n18119), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18090) );
  OAI21_X1 U21366 ( .B1(n21203), .B2(n18094), .A(n18090), .ZN(P3_U2748) );
  AOI22_X1 U21367 ( .A1(n18119), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18091) );
  OAI21_X1 U21368 ( .B1(n18131), .B2(n18094), .A(n18091), .ZN(P3_U2749) );
  AOI22_X1 U21369 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(n18118), .B1(n18119), 
        .B2(P3_UWORD_REG_1__SCAN_IN), .ZN(n18092) );
  OAI21_X1 U21370 ( .B1(n18129), .B2(n18094), .A(n18092), .ZN(P3_U2750) );
  INV_X1 U21371 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18127) );
  AOI22_X1 U21372 ( .A1(n18119), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18093) );
  OAI21_X1 U21373 ( .B1(n18127), .B2(n18094), .A(n18093), .ZN(P3_U2751) );
  INV_X1 U21374 ( .A(P3_LWORD_REG_15__SCAN_IN), .ZN(n21067) );
  AOI22_X1 U21375 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n18104), .B1(n18118), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18095) );
  OAI21_X1 U21376 ( .B1(n21067), .B2(n18102), .A(n18095), .ZN(P3_U2752) );
  INV_X1 U21377 ( .A(P3_LWORD_REG_14__SCAN_IN), .ZN(n21054) );
  AOI22_X1 U21378 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18104), .B1(n18118), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18096) );
  OAI21_X1 U21379 ( .B1(n21054), .B2(n18102), .A(n18096), .ZN(P3_U2753) );
  AOI22_X1 U21380 ( .A1(n18119), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18097) );
  OAI21_X1 U21381 ( .B1(n18098), .B2(n18121), .A(n18097), .ZN(P3_U2754) );
  AOI22_X1 U21382 ( .A1(n18119), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18099) );
  OAI21_X1 U21383 ( .B1(n18100), .B2(n18121), .A(n18099), .ZN(P3_U2755) );
  INV_X1 U21384 ( .A(P3_LWORD_REG_11__SCAN_IN), .ZN(n21097) );
  AOI22_X1 U21385 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18104), .B1(n18118), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18101) );
  OAI21_X1 U21386 ( .B1(n21097), .B2(n18102), .A(n18101), .ZN(P3_U2756) );
  AOI22_X1 U21387 ( .A1(n18119), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18103) );
  OAI21_X1 U21388 ( .B1(n21139), .B2(n18121), .A(n18103), .ZN(P3_U2757) );
  AOI222_X1 U21389 ( .A1(P3_LWORD_REG_9__SCAN_IN), .A2(n18119), .B1(n18118), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .C1(P3_EAX_REG_9__SCAN_IN), .C2(n18104), 
        .ZN(n18105) );
  INV_X1 U21390 ( .A(n18105), .ZN(P3_U2758) );
  AOI22_X1 U21391 ( .A1(n18119), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18106) );
  OAI21_X1 U21392 ( .B1(n18107), .B2(n18121), .A(n18106), .ZN(P3_U2759) );
  INV_X1 U21393 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18160) );
  AOI22_X1 U21394 ( .A1(n18119), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18108) );
  OAI21_X1 U21395 ( .B1(n18160), .B2(n18121), .A(n18108), .ZN(P3_U2760) );
  INV_X1 U21396 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18110) );
  AOI22_X1 U21397 ( .A1(n18119), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18109) );
  OAI21_X1 U21398 ( .B1(n18110), .B2(n18121), .A(n18109), .ZN(P3_U2761) );
  INV_X1 U21399 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18112) );
  AOI22_X1 U21400 ( .A1(n18119), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18111) );
  OAI21_X1 U21401 ( .B1(n18112), .B2(n18121), .A(n18111), .ZN(P3_U2762) );
  AOI22_X1 U21402 ( .A1(n18119), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18113) );
  OAI21_X1 U21403 ( .B1(n21047), .B2(n18121), .A(n18113), .ZN(P3_U2763) );
  AOI22_X1 U21404 ( .A1(n18119), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18114) );
  OAI21_X1 U21405 ( .B1(n18115), .B2(n18121), .A(n18114), .ZN(P3_U2764) );
  INV_X1 U21406 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18154) );
  AOI22_X1 U21407 ( .A1(n18119), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18116) );
  OAI21_X1 U21408 ( .B1(n18154), .B2(n18121), .A(n18116), .ZN(P3_U2765) );
  AOI22_X1 U21409 ( .A1(n18119), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18117) );
  OAI21_X1 U21410 ( .B1(n18152), .B2(n18121), .A(n18117), .ZN(P3_U2766) );
  AOI22_X1 U21411 ( .A1(n18119), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18118), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18120) );
  OAI21_X1 U21412 ( .B1(n18150), .B2(n18121), .A(n18120), .ZN(P3_U2767) );
  NAND2_X1 U21413 ( .A1(n19539), .A2(n18122), .ZN(n19384) );
  NOR2_X2 U21414 ( .A1(n18123), .A2(n19384), .ZN(n18173) );
  AOI211_X1 U21415 ( .C1(n18125), .C2(n19411), .A(n18124), .B(n18123), .ZN(
        n18178) );
  NAND2_X1 U21416 ( .A1(n18125), .A2(n18178), .ZN(n18180) );
  AOI22_X1 U21417 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18174), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18171), .ZN(n18126) );
  OAI21_X1 U21418 ( .B1(n18127), .B2(n18176), .A(n18126), .ZN(P3_U2768) );
  AOI22_X1 U21419 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18174), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18171), .ZN(n18128) );
  OAI21_X1 U21420 ( .B1(n18129), .B2(n18176), .A(n18128), .ZN(P3_U2769) );
  AOI22_X1 U21421 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18174), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18171), .ZN(n18130) );
  OAI21_X1 U21422 ( .B1(n18131), .B2(n18176), .A(n18130), .ZN(P3_U2770) );
  AOI22_X1 U21423 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18174), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18171), .ZN(n18132) );
  OAI21_X1 U21424 ( .B1(n21203), .B2(n18176), .A(n18132), .ZN(P3_U2771) );
  AOI22_X1 U21425 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18174), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18171), .ZN(n18133) );
  OAI21_X1 U21426 ( .B1(n18134), .B2(n18176), .A(n18133), .ZN(P3_U2772) );
  AOI22_X1 U21427 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18174), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18171), .ZN(n18135) );
  OAI21_X1 U21428 ( .B1(n18136), .B2(n18176), .A(n18135), .ZN(P3_U2773) );
  AOI22_X1 U21429 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18174), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18171), .ZN(n18137) );
  OAI21_X1 U21430 ( .B1(n18138), .B2(n18176), .A(n18137), .ZN(P3_U2774) );
  AOI22_X1 U21431 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18174), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18171), .ZN(n18139) );
  OAI21_X1 U21432 ( .B1(n18140), .B2(n18176), .A(n18139), .ZN(P3_U2775) );
  AOI22_X1 U21433 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18173), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18171), .ZN(n18141) );
  OAI21_X1 U21434 ( .B1(n18162), .B2(n18180), .A(n18141), .ZN(P3_U2776) );
  AOI22_X1 U21435 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18174), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18171), .ZN(n18142) );
  OAI21_X1 U21436 ( .B1(n21123), .B2(n18176), .A(n18142), .ZN(P3_U2777) );
  INV_X1 U21437 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18166) );
  AOI22_X1 U21438 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18173), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18171), .ZN(n18143) );
  OAI21_X1 U21439 ( .B1(n18166), .B2(n18180), .A(n18143), .ZN(P3_U2778) );
  AOI22_X1 U21440 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n18173), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18171), .ZN(n18144) );
  OAI21_X1 U21441 ( .B1(n18168), .B2(n18180), .A(n18144), .ZN(P3_U2779) );
  AOI22_X1 U21442 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18173), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18171), .ZN(n18145) );
  OAI21_X1 U21443 ( .B1(n18170), .B2(n18180), .A(n18145), .ZN(P3_U2780) );
  AOI22_X1 U21444 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18173), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18171), .ZN(n18146) );
  OAI21_X1 U21445 ( .B1(n21221), .B2(n18180), .A(n18146), .ZN(P3_U2781) );
  AOI22_X1 U21446 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18174), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18171), .ZN(n18147) );
  OAI21_X1 U21447 ( .B1(n18148), .B2(n18176), .A(n18147), .ZN(P3_U2782) );
  AOI22_X1 U21448 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18174), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18171), .ZN(n18149) );
  OAI21_X1 U21449 ( .B1(n18150), .B2(n18176), .A(n18149), .ZN(P3_U2783) );
  AOI22_X1 U21450 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18174), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18171), .ZN(n18151) );
  OAI21_X1 U21451 ( .B1(n18152), .B2(n18176), .A(n18151), .ZN(P3_U2784) );
  AOI22_X1 U21452 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18174), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18171), .ZN(n18153) );
  OAI21_X1 U21453 ( .B1(n18154), .B2(n18176), .A(n18153), .ZN(P3_U2785) );
  AOI22_X1 U21454 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18173), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18171), .ZN(n18155) );
  OAI21_X1 U21455 ( .B1(n18908), .B2(n18180), .A(n18155), .ZN(P3_U2786) );
  AOI22_X1 U21456 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18173), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18171), .ZN(n18156) );
  OAI21_X1 U21457 ( .B1(n18913), .B2(n18180), .A(n18156), .ZN(P3_U2787) );
  AOI22_X1 U21458 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18173), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18171), .ZN(n18157) );
  OAI21_X1 U21459 ( .B1(n21293), .B2(n18180), .A(n18157), .ZN(P3_U2788) );
  AOI22_X1 U21460 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18173), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18171), .ZN(n18158) );
  OAI21_X1 U21461 ( .B1(n18921), .B2(n18180), .A(n18158), .ZN(P3_U2789) );
  AOI22_X1 U21462 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18174), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18171), .ZN(n18159) );
  OAI21_X1 U21463 ( .B1(n18160), .B2(n18176), .A(n18159), .ZN(P3_U2790) );
  AOI22_X1 U21464 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18173), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18171), .ZN(n18161) );
  OAI21_X1 U21465 ( .B1(n18162), .B2(n18180), .A(n18161), .ZN(P3_U2791) );
  AOI22_X1 U21466 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18174), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18171), .ZN(n18163) );
  OAI21_X1 U21467 ( .B1(n18164), .B2(n18176), .A(n18163), .ZN(P3_U2792) );
  AOI22_X1 U21468 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18173), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18171), .ZN(n18165) );
  OAI21_X1 U21469 ( .B1(n18166), .B2(n18180), .A(n18165), .ZN(P3_U2793) );
  AOI22_X1 U21470 ( .A1(P3_LWORD_REG_11__SCAN_IN), .A2(n18171), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n18173), .ZN(n18167) );
  OAI21_X1 U21471 ( .B1(n18168), .B2(n18180), .A(n18167), .ZN(P3_U2794) );
  AOI22_X1 U21472 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18173), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18171), .ZN(n18169) );
  OAI21_X1 U21473 ( .B1(n18170), .B2(n18180), .A(n18169), .ZN(P3_U2795) );
  AOI22_X1 U21474 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18173), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18171), .ZN(n18172) );
  OAI21_X1 U21475 ( .B1(n21221), .B2(n18180), .A(n18172), .ZN(P3_U2796) );
  AOI22_X1 U21476 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18174), .B1(
        P3_EAX_REG_14__SCAN_IN), .B2(n18173), .ZN(n18175) );
  OAI21_X1 U21477 ( .B1(n18178), .B2(n21054), .A(n18175), .ZN(P3_U2797) );
  OAI222_X1 U21478 ( .A1(n18180), .A2(n18179), .B1(n21067), .B2(n18178), .C1(
        n18177), .C2(n18176), .ZN(P3_U2798) );
  NOR2_X1 U21479 ( .A1(n18309), .A2(n18629), .ZN(n18628) );
  INV_X1 U21480 ( .A(n18628), .ZN(n18564) );
  NOR3_X1 U21481 ( .A1(n18636), .A2(n18356), .A3(n18564), .ZN(n18264) );
  INV_X1 U21482 ( .A(n18264), .ZN(n18251) );
  AOI211_X1 U21483 ( .C1(n18183), .C2(n18182), .A(n18181), .B(n18399), .ZN(
        n18193) );
  INV_X1 U21484 ( .A(n18388), .ZN(n18266) );
  NAND2_X1 U21485 ( .A1(n18184), .A2(n18266), .ZN(n18190) );
  NOR3_X1 U21486 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18388), .A3(
        n10179), .ZN(n18208) );
  OAI21_X1 U21487 ( .B1(n18185), .B2(n18509), .A(n18554), .ZN(n18186) );
  AOI21_X1 U21488 ( .B1(n18384), .B2(n18187), .A(n18186), .ZN(n18211) );
  OAI21_X1 U21489 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18256), .A(
        n18211), .ZN(n18209) );
  OAI21_X1 U21490 ( .B1(n18208), .B2(n18209), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18189) );
  OAI211_X1 U21491 ( .C1(n18191), .C2(n18190), .A(n18189), .B(n18188), .ZN(
        n18192) );
  AOI211_X1 U21492 ( .C1(n18194), .C2(n18401), .A(n18193), .B(n18192), .ZN(
        n18198) );
  NAND2_X1 U21493 ( .A1(n18560), .A2(n18467), .ZN(n18294) );
  AOI22_X1 U21494 ( .A1(n18547), .A2(n18195), .B1(n18396), .B2(n18572), .ZN(
        n18224) );
  NAND2_X1 U21495 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18224), .ZN(
        n18196) );
  NAND3_X1 U21496 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18294), .A3(
        n18196), .ZN(n18197) );
  OAI211_X1 U21497 ( .C1(n18199), .C2(n18251), .A(n18198), .B(n18197), .ZN(
        P3_U2802) );
  NAND2_X1 U21498 ( .A1(n18201), .A2(n18200), .ZN(n18202) );
  XOR2_X1 U21499 ( .A(n18202), .B(n18382), .Z(n18578) );
  AOI22_X1 U21500 ( .A1(n18869), .A2(P3_REIP_REG_27__SCAN_IN), .B1(n18401), 
        .B2(n18203), .ZN(n18204) );
  OAI221_X1 U21501 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18206), 
        .C1(n18205), .C2(n18224), .A(n18204), .ZN(n18207) );
  AOI211_X1 U21502 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n18209), .A(
        n18208), .B(n18207), .ZN(n18210) );
  OAI21_X1 U21503 ( .B1(n18578), .B2(n18399), .A(n18210), .ZN(P3_U2803) );
  NAND2_X1 U21504 ( .A1(n18869), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18583) );
  INV_X1 U21505 ( .A(n18583), .ZN(n18215) );
  INV_X2 U21506 ( .A(n19265), .ZN(n18999) );
  AOI221_X1 U21507 ( .B1(n18999), .B2(n18213), .C1(n18212), .C2(n18213), .A(
        n18211), .ZN(n18214) );
  AOI211_X1 U21508 ( .C1(n18217), .C2(n18216), .A(n18215), .B(n18214), .ZN(
        n18223) );
  OAI21_X1 U21509 ( .B1(n18219), .B2(n18585), .A(n18218), .ZN(n18581) );
  NOR2_X1 U21510 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18251), .ZN(
        n18220) );
  AOI22_X1 U21511 ( .A1(n18464), .A2(n18581), .B1(n18221), .B2(n18220), .ZN(
        n18222) );
  OAI211_X1 U21512 ( .C1(n18224), .C2(n18585), .A(n18223), .B(n18222), .ZN(
        P3_U2804) );
  OAI21_X1 U21513 ( .B1(n18234), .B2(n18999), .A(n18554), .ZN(n18225) );
  AOI21_X1 U21514 ( .B1(n18384), .B2(n18226), .A(n18225), .ZN(n18261) );
  OAI21_X1 U21515 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18256), .A(
        n18261), .ZN(n18243) );
  AOI22_X1 U21516 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18243), .B1(
        n18401), .B2(n18227), .ZN(n18239) );
  XOR2_X1 U21517 ( .A(n18228), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18598) );
  XOR2_X1 U21518 ( .A(n18229), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18600) );
  OAI21_X1 U21519 ( .B1(n18463), .B2(n18231), .A(n18230), .ZN(n18232) );
  XOR2_X1 U21520 ( .A(n18232), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18596) );
  OAI22_X1 U21521 ( .A1(n18560), .A2(n18600), .B1(n18399), .B2(n18596), .ZN(
        n18233) );
  AOI21_X1 U21522 ( .B1(n18396), .B2(n18598), .A(n18233), .ZN(n18238) );
  NAND2_X1 U21523 ( .A1(n18828), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18594) );
  NOR2_X1 U21524 ( .A1(n18388), .A2(n18235), .ZN(n18245) );
  OAI211_X1 U21525 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18245), .B(n18236), .ZN(n18237) );
  NAND4_X1 U21526 ( .A1(n18239), .A2(n18238), .A3(n18594), .A4(n18237), .ZN(
        P3_U2805) );
  NAND2_X1 U21527 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18609), .ZN(
        n18616) );
  INV_X1 U21528 ( .A(n18240), .ZN(n18241) );
  NAND2_X1 U21529 ( .A1(n18869), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18613) );
  OAI21_X1 U21530 ( .B1(n18241), .B2(n18393), .A(n18613), .ZN(n18242) );
  AOI221_X1 U21531 ( .B1(n18245), .B2(n18244), .C1(n18243), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18242), .ZN(n18250) );
  NOR2_X1 U21532 ( .A1(n18697), .A2(n18246), .ZN(n18604) );
  NOR2_X1 U21533 ( .A1(n18623), .A2(n18246), .ZN(n18602) );
  OAI22_X1 U21534 ( .A1(n18604), .A2(n18467), .B1(n18602), .B2(n18560), .ZN(
        n18263) );
  OAI21_X1 U21535 ( .B1(n18248), .B2(n18609), .A(n18247), .ZN(n18612) );
  AOI22_X1 U21536 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18263), .B1(
        n18464), .B2(n18612), .ZN(n18249) );
  OAI211_X1 U21537 ( .C1(n18251), .C2(n18616), .A(n18250), .B(n18249), .ZN(
        P3_U2806) );
  OAI22_X1 U21538 ( .A1(n18463), .A2(n18636), .B1(n18252), .B2(n18275), .ZN(
        n18253) );
  NOR2_X1 U21539 ( .A1(n18253), .A2(n18302), .ZN(n18254) );
  XOR2_X1 U21540 ( .A(n18254), .B(n21089), .Z(n18621) );
  AOI21_X1 U21541 ( .B1(n18255), .B2(n19265), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18260) );
  OAI21_X1 U21542 ( .B1(n18401), .B2(n18296), .A(n18257), .ZN(n18259) );
  NAND2_X1 U21543 ( .A1(n18869), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18258) );
  OAI211_X1 U21544 ( .C1(n18261), .C2(n18260), .A(n18259), .B(n18258), .ZN(
        n18262) );
  AOI221_X1 U21545 ( .B1(n18264), .B2(n21089), .C1(n18263), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n18262), .ZN(n18265) );
  OAI21_X1 U21546 ( .B1(n18399), .B2(n18621), .A(n18265), .ZN(P3_U2807) );
  NAND2_X1 U21547 ( .A1(n18340), .A2(n18628), .ZN(n18280) );
  NAND2_X1 U21548 ( .A1(n18269), .A2(n18266), .ZN(n18287) );
  AOI221_X1 U21549 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n18286), .C2(n18270), .A(
        n18287), .ZN(n18272) );
  OR2_X1 U21550 ( .A1(n18555), .A2(n18267), .ZN(n18268) );
  OAI211_X1 U21551 ( .C1(n18269), .C2(n18509), .A(n18554), .B(n18268), .ZN(
        n18301) );
  AOI21_X1 U21552 ( .B1(n18296), .B2(n21230), .A(n18301), .ZN(n18285) );
  OAI22_X1 U21553 ( .A1(n18285), .A2(n18270), .B1(n18833), .B2(n19459), .ZN(
        n18271) );
  AOI211_X1 U21554 ( .C1(n18273), .C2(n18401), .A(n18272), .B(n18271), .ZN(
        n18279) );
  AOI22_X1 U21555 ( .A1(n18547), .A2(n18623), .B1(n18396), .B2(n18697), .ZN(
        n18355) );
  INV_X1 U21556 ( .A(n18355), .ZN(n18329) );
  AOI21_X1 U21557 ( .B1(n18294), .B2(n18564), .A(n18329), .ZN(n18274) );
  INV_X1 U21558 ( .A(n18274), .ZN(n18291) );
  INV_X1 U21559 ( .A(n18275), .ZN(n18276) );
  AOI221_X1 U21560 ( .B1(n18344), .B2(n18276), .C1(n18564), .C2(n18276), .A(
        n18302), .ZN(n18277) );
  XOR2_X1 U21561 ( .A(n18277), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n18622) );
  AOI22_X1 U21562 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18291), .B1(
        n18464), .B2(n18622), .ZN(n18278) );
  OAI211_X1 U21563 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18280), .A(
        n18279), .B(n18278), .ZN(P3_U2808) );
  NAND3_X1 U21564 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18463), .A3(
        n18281), .ZN(n18310) );
  INV_X1 U21565 ( .A(n18322), .ZN(n18311) );
  OAI22_X1 U21566 ( .A1(n18290), .A2(n18310), .B1(n18311), .B2(n18282), .ZN(
        n18283) );
  XNOR2_X1 U21567 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18283), .ZN(
        n18647) );
  NAND2_X1 U21568 ( .A1(n18828), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18284) );
  OAI221_X1 U21569 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18287), .C1(
        n18286), .C2(n18285), .A(n18284), .ZN(n18288) );
  AOI21_X1 U21570 ( .B1(n18401), .B2(n18289), .A(n18288), .ZN(n18293) );
  NOR3_X1 U21571 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18309), .A3(
        n18290), .ZN(n18637) );
  AOI22_X1 U21572 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18291), .B1(
        n18340), .B2(n18637), .ZN(n18292) );
  OAI211_X1 U21573 ( .C1(n18647), .C2(n18399), .A(n18293), .B(n18292), .ZN(
        P3_U2809) );
  INV_X1 U21574 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18313) );
  NOR2_X1 U21575 ( .A1(n18309), .A2(n18313), .ZN(n18651) );
  INV_X1 U21576 ( .A(n18651), .ZN(n18624) );
  AOI21_X1 U21577 ( .B1(n18294), .B2(n18624), .A(n18329), .ZN(n18314) );
  OAI21_X1 U21578 ( .B1(n18999), .B2(n18295), .A(n21230), .ZN(n18300) );
  NOR2_X1 U21579 ( .A1(n18833), .A2(n19455), .ZN(n18299) );
  AOI21_X1 U21580 ( .B1(n18393), .B2(n18256), .A(n18297), .ZN(n18298) );
  AOI211_X1 U21581 ( .C1(n18301), .C2(n18300), .A(n18299), .B(n18298), .ZN(
        n18305) );
  AOI221_X1 U21582 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18310), 
        .C1(n18313), .C2(n18320), .A(n18302), .ZN(n18303) );
  XOR2_X1 U21583 ( .A(n18303), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n18649) );
  NOR2_X1 U21584 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18624), .ZN(
        n18648) );
  AOI22_X1 U21585 ( .A1(n18464), .A2(n18649), .B1(n18340), .B2(n18648), .ZN(
        n18304) );
  OAI211_X1 U21586 ( .C1(n18314), .C2(n18306), .A(n18305), .B(n18304), .ZN(
        P3_U2810) );
  OAI21_X1 U21587 ( .B1(n18526), .B2(n18316), .A(n18549), .ZN(n18335) );
  OAI21_X1 U21588 ( .B1(n18307), .B2(n18555), .A(n18335), .ZN(n18326) );
  AOI22_X1 U21589 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18326), .B1(
        n18401), .B2(n18308), .ZN(n18319) );
  NOR2_X1 U21590 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18309), .ZN(
        n18655) );
  OAI21_X1 U21591 ( .B1(n18320), .B2(n18311), .A(n18310), .ZN(n18312) );
  XOR2_X1 U21592 ( .A(n18312), .B(n18313), .Z(n18660) );
  OAI22_X1 U21593 ( .A1(n18660), .A2(n18399), .B1(n18314), .B2(n18313), .ZN(
        n18315) );
  AOI21_X1 U21594 ( .B1(n18340), .B2(n18655), .A(n18315), .ZN(n18318) );
  NAND2_X1 U21595 ( .A1(n18828), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18658) );
  NOR2_X1 U21596 ( .A1(n18388), .A2(n18316), .ZN(n18328) );
  OAI221_X1 U21597 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C1(n21075), .C2(n18327), .A(
        n18328), .ZN(n18317) );
  NAND4_X1 U21598 ( .A1(n18319), .A2(n18318), .A3(n18658), .A4(n18317), .ZN(
        P3_U2811) );
  OAI21_X1 U21599 ( .B1(n18382), .B2(n18321), .A(n18320), .ZN(n18323) );
  XOR2_X1 U21600 ( .A(n18323), .B(n18322), .Z(n18676) );
  NAND2_X1 U21601 ( .A1(n18869), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18674) );
  OAI21_X1 U21602 ( .B1(n18324), .B2(n18393), .A(n18674), .ZN(n18325) );
  AOI221_X1 U21603 ( .B1(n18328), .B2(n18327), .C1(n18326), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18325), .ZN(n18332) );
  AOI21_X1 U21604 ( .B1(n18662), .B2(n18340), .A(n18329), .ZN(n18330) );
  INV_X1 U21605 ( .A(n18330), .ZN(n18341) );
  NOR2_X1 U21606 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18662), .ZN(
        n18672) );
  AOI22_X1 U21607 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18341), .B1(
        n18340), .B2(n18672), .ZN(n18331) );
  OAI211_X1 U21608 ( .C1(n18399), .C2(n18676), .A(n18332), .B(n18331), .ZN(
        P3_U2812) );
  AOI21_X1 U21609 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18334), .A(
        n18333), .ZN(n18683) );
  AOI221_X1 U21610 ( .B1(n18999), .B2(n18337), .C1(n18336), .C2(n18337), .A(
        n18335), .ZN(n18338) );
  NOR2_X1 U21611 ( .A1(n18833), .A2(n19450), .ZN(n18680) );
  AOI211_X1 U21612 ( .C1(n18339), .C2(n18216), .A(n18338), .B(n18680), .ZN(
        n18343) );
  NOR2_X1 U21613 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18692), .ZN(
        n18678) );
  AOI22_X1 U21614 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18341), .B1(
        n18340), .B2(n18678), .ZN(n18342) );
  OAI211_X1 U21615 ( .C1(n18683), .C2(n18399), .A(n18343), .B(n18342), .ZN(
        P3_U2813) );
  NOR2_X1 U21616 ( .A1(n18382), .A2(n18729), .ZN(n18441) );
  AOI22_X1 U21617 ( .A1(n18441), .A2(n18345), .B1(n18344), .B2(n18382), .ZN(
        n18346) );
  XOR2_X1 U21618 ( .A(n18692), .B(n18346), .Z(n18694) );
  OAI21_X1 U21619 ( .B1(n18526), .B2(n18349), .A(n18549), .ZN(n18370) );
  OAI21_X1 U21620 ( .B1(n18347), .B2(n18555), .A(n18370), .ZN(n18359) );
  AOI22_X1 U21621 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18359), .B1(
        n18401), .B2(n18348), .ZN(n18352) );
  NOR2_X1 U21622 ( .A1(n18388), .A2(n18349), .ZN(n18361) );
  OAI221_X1 U21623 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n18360), .C2(n18350), .A(
        n18361), .ZN(n18351) );
  OAI211_X1 U21624 ( .C1(n19447), .C2(n18833), .A(n18352), .B(n18351), .ZN(
        n18353) );
  AOI21_X1 U21625 ( .B1(n18464), .B2(n18694), .A(n18353), .ZN(n18354) );
  OAI221_X1 U21626 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18356), 
        .C1(n18692), .C2(n18355), .A(n18354), .ZN(P3_U2814) );
  NOR2_X1 U21627 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18374), .ZN(
        n18698) );
  NAND2_X1 U21628 ( .A1(n18396), .A2(n18697), .ZN(n18366) );
  OAI22_X1 U21629 ( .A1(n18833), .A2(n21323), .B1(n18393), .B2(n18357), .ZN(
        n18358) );
  AOI221_X1 U21630 ( .B1(n18361), .B2(n18360), .C1(n18359), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18358), .ZN(n18365) );
  NAND2_X1 U21631 ( .A1(n18732), .A2(n18441), .ZN(n18375) );
  NOR2_X1 U21632 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18749), .ZN(
        n18737) );
  AOI221_X1 U21633 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18375), 
        .C1(n18721), .C2(n9785), .A(n18737), .ZN(n18362) );
  XOR2_X1 U21634 ( .A(n18362), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n18708) );
  NOR2_X1 U21635 ( .A1(n18705), .A2(n18560), .ZN(n18363) );
  NAND2_X1 U21636 ( .A1(n18367), .A2(n18699), .ZN(n18706) );
  AOI22_X1 U21637 ( .A1(n18464), .A2(n18708), .B1(n18363), .B2(n18706), .ZN(
        n18364) );
  OAI211_X1 U21638 ( .C1(n18698), .C2(n18366), .A(n18365), .B(n18364), .ZN(
        P3_U2815) );
  OAI21_X1 U21639 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18368), .A(
        n18367), .ZN(n18728) );
  INV_X1 U21640 ( .A(n18389), .ZN(n18369) );
  NOR2_X1 U21641 ( .A1(n18999), .A2(n18387), .ZN(n18418) );
  AOI21_X1 U21642 ( .B1(n18369), .B2(n18418), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18371) );
  OAI22_X1 U21643 ( .A1(n18371), .A2(n18370), .B1(n18833), .B2(n19445), .ZN(
        n18372) );
  AOI21_X1 U21644 ( .B1(n18373), .B2(n18216), .A(n18372), .ZN(n18378) );
  AOI221_X1 U21645 ( .B1(n18718), .B2(n18721), .C1(n18729), .C2(n18721), .A(
        n18374), .ZN(n18724) );
  AOI21_X1 U21646 ( .B1(n18375), .B2(n9785), .A(n18737), .ZN(n18376) );
  XOR2_X1 U21647 ( .A(n18376), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18723) );
  AOI22_X1 U21648 ( .A1(n18396), .A2(n18724), .B1(n18464), .B2(n18723), .ZN(
        n18377) );
  OAI211_X1 U21649 ( .C1(n18560), .C2(n18728), .A(n18378), .B(n18377), .ZN(
        P3_U2816) );
  INV_X1 U21650 ( .A(n18379), .ZN(n18380) );
  AOI22_X1 U21651 ( .A1(n18380), .A2(n18732), .B1(n18749), .B2(n18382), .ZN(
        n18381) );
  AOI21_X1 U21652 ( .B1(n18382), .B2(n18403), .A(n18381), .ZN(n18383) );
  XNOR2_X1 U21653 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18383), .ZN(
        n18741) );
  AOI21_X1 U21654 ( .B1(n18452), .B2(n18387), .A(n18384), .ZN(n18385) );
  OAI21_X1 U21655 ( .B1(n18386), .B2(n18385), .A(n18554), .ZN(n18402) );
  NOR2_X1 U21656 ( .A1(n18388), .A2(n18387), .ZN(n18406) );
  OAI211_X1 U21657 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18406), .B(n18389), .ZN(n18391) );
  NAND2_X1 U21658 ( .A1(n18828), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18390) );
  OAI211_X1 U21659 ( .C1(n18393), .C2(n18392), .A(n18391), .B(n18390), .ZN(
        n18394) );
  AOI21_X1 U21660 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18402), .A(
        n18394), .ZN(n18398) );
  INV_X1 U21661 ( .A(n18395), .ZN(n18451) );
  AOI22_X1 U21662 ( .A1(n18547), .A2(n18731), .B1(n18396), .B2(n18729), .ZN(
        n18450) );
  OAI21_X1 U21663 ( .B1(n18732), .B2(n18451), .A(n18450), .ZN(n18407) );
  NOR2_X1 U21664 ( .A1(n18451), .A2(n18736), .ZN(n18408) );
  AOI22_X1 U21665 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18407), .B1(
        n18737), .B2(n18408), .ZN(n18397) );
  OAI211_X1 U21666 ( .C1(n18399), .C2(n18741), .A(n18398), .B(n18397), .ZN(
        P3_U2817) );
  AOI22_X1 U21667 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18402), .B1(
        n18401), .B2(n18400), .ZN(n18411) );
  NAND2_X1 U21668 ( .A1(n18756), .A2(n18441), .ZN(n18412) );
  OAI21_X1 U21669 ( .B1(n18413), .B2(n18412), .A(n18403), .ZN(n18404) );
  XOR2_X1 U21670 ( .A(n18404), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18746) );
  AOI22_X1 U21671 ( .A1(n18464), .A2(n18746), .B1(n18406), .B2(n18405), .ZN(
        n18410) );
  NAND2_X1 U21672 ( .A1(n18828), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18747) );
  OAI21_X1 U21673 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18408), .A(
        n18407), .ZN(n18409) );
  NAND4_X1 U21674 ( .A1(n18411), .A2(n18410), .A3(n18747), .A4(n18409), .ZN(
        P3_U2818) );
  NAND2_X1 U21675 ( .A1(n18756), .A2(n18413), .ZN(n18762) );
  INV_X1 U21676 ( .A(n18412), .ZN(n18427) );
  NOR2_X1 U21677 ( .A1(n18427), .A2(n9805), .ZN(n18414) );
  XOR2_X1 U21678 ( .A(n18414), .B(n18413), .Z(n18750) );
  NOR2_X1 U21679 ( .A1(n18833), .A2(n21135), .ZN(n18420) );
  NOR4_X1 U21680 ( .A1(n18999), .A2(n18471), .A3(n18469), .A4(n18457), .ZN(
        n18443) );
  INV_X1 U21681 ( .A(n18443), .ZN(n18430) );
  NOR2_X1 U21682 ( .A1(n18415), .A2(n18430), .ZN(n18433) );
  AOI21_X1 U21683 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18549), .A(
        n18433), .ZN(n18417) );
  OAI22_X1 U21684 ( .A1(n18418), .A2(n18417), .B1(n18538), .B2(n18416), .ZN(
        n18419) );
  AOI211_X1 U21685 ( .C1(n18464), .C2(n18750), .A(n18420), .B(n18419), .ZN(
        n18422) );
  NOR2_X1 U21686 ( .A1(n18756), .A2(n18451), .ZN(n18428) );
  INV_X1 U21687 ( .A(n18450), .ZN(n18429) );
  OAI21_X1 U21688 ( .B1(n18428), .B2(n18429), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18421) );
  OAI211_X1 U21689 ( .C1(n18451), .C2(n18762), .A(n18422), .B(n18421), .ZN(
        P3_U2819) );
  NOR4_X1 U21690 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18463), .A3(
        n18424), .A4(n18423), .ZN(n18426) );
  AOI221_X1 U21691 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18441), .C1(
        n18776), .C2(n18440), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18425) );
  NOR3_X1 U21692 ( .A1(n18427), .A2(n18426), .A3(n18425), .ZN(n18767) );
  AOI21_X1 U21693 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18429), .A(
        n18428), .ZN(n18434) );
  NOR2_X1 U21694 ( .A1(n18431), .A2(n18430), .ZN(n18446) );
  AOI21_X1 U21695 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18549), .A(
        n18446), .ZN(n18432) );
  OAI22_X1 U21696 ( .A1(n18435), .A2(n18434), .B1(n18433), .B2(n18432), .ZN(
        n18436) );
  AOI21_X1 U21697 ( .B1(n18464), .B2(n18767), .A(n18436), .ZN(n18438) );
  NAND2_X1 U21698 ( .A1(n18828), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18437) );
  OAI211_X1 U21699 ( .C1(n18538), .C2(n18439), .A(n18438), .B(n18437), .ZN(
        P3_U2820) );
  NOR2_X1 U21700 ( .A1(n18441), .A2(n18440), .ZN(n18442) );
  XOR2_X1 U21701 ( .A(n18442), .B(n18776), .Z(n18773) );
  NOR2_X1 U21702 ( .A1(n18833), .A2(n19437), .ZN(n18448) );
  AOI21_X1 U21703 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18549), .A(
        n18443), .ZN(n18445) );
  OAI22_X1 U21704 ( .A1(n18446), .A2(n18445), .B1(n18538), .B2(n18444), .ZN(
        n18447) );
  AOI211_X1 U21705 ( .C1(n18464), .C2(n18773), .A(n18448), .B(n18447), .ZN(
        n18449) );
  OAI221_X1 U21706 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18451), .C1(
        n18776), .C2(n18450), .A(n18449), .ZN(P3_U2821) );
  NOR3_X1 U21707 ( .A1(n18999), .A2(n18471), .A3(n18469), .ZN(n18458) );
  AOI21_X1 U21708 ( .B1(n18452), .B2(n18471), .A(n18526), .ZN(n18468) );
  OAI21_X1 U21709 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18999), .A(
        n18468), .ZN(n18456) );
  AOI22_X1 U21710 ( .A1(n18216), .A2(n18453), .B1(n18869), .B2(
        P3_REIP_REG_8__SCAN_IN), .ZN(n18454) );
  INV_X1 U21711 ( .A(n18454), .ZN(n18455) );
  AOI221_X1 U21712 ( .B1(n18458), .B2(n18457), .C1(n18456), .C2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(n18455), .ZN(n18466) );
  AOI21_X1 U21713 ( .B1(n18460), .B2(n21202), .A(n18459), .ZN(n18789) );
  OAI21_X1 U21714 ( .B1(n18463), .B2(n18462), .A(n18461), .ZN(n18787) );
  AOI22_X1 U21715 ( .A1(n18547), .A2(n18789), .B1(n18464), .B2(n18787), .ZN(
        n18465) );
  OAI211_X1 U21716 ( .C1(n18467), .C2(n18793), .A(n18466), .B(n18465), .ZN(
        P3_U2822) );
  NAND2_X1 U21717 ( .A1(n19265), .A2(n18469), .ZN(n18470) );
  OAI22_X1 U21718 ( .A1(n18471), .A2(n18470), .B1(n18469), .B2(n18468), .ZN(
        n18478) );
  NAND2_X1 U21719 ( .A1(n18473), .A2(n18472), .ZN(n18474) );
  XOR2_X1 U21720 ( .A(n18474), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18796) );
  INV_X1 U21721 ( .A(n18502), .ZN(n18558) );
  OAI21_X1 U21722 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18476), .A(
        n18475), .ZN(n18795) );
  OAI22_X1 U21723 ( .A1(n18560), .A2(n18796), .B1(n18558), .B2(n18795), .ZN(
        n18477) );
  AOI211_X1 U21724 ( .C1(n18828), .C2(P3_REIP_REG_7__SCAN_IN), .A(n18478), .B(
        n18477), .ZN(n18479) );
  OAI21_X1 U21725 ( .B1(n18538), .B2(n18480), .A(n18479), .ZN(P3_U2823) );
  OAI21_X1 U21726 ( .B1(n18481), .B2(n18999), .A(n18549), .ZN(n18505) );
  OR2_X1 U21727 ( .A1(n18999), .A2(n18481), .ZN(n18485) );
  OAI21_X1 U21728 ( .B1(n18484), .B2(n18483), .A(n18482), .ZN(n18804) );
  OAI22_X1 U21729 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18485), .B1(
        n18558), .B2(n18804), .ZN(n18486) );
  AOI21_X1 U21730 ( .B1(n18828), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18486), .ZN(
        n18491) );
  AOI21_X1 U21731 ( .B1(n18488), .B2(n18808), .A(n18487), .ZN(n18806) );
  AOI22_X1 U21732 ( .A1(n18547), .A2(n18806), .B1(n18489), .B2(n18216), .ZN(
        n18490) );
  OAI211_X1 U21733 ( .C1(n18492), .C2(n18505), .A(n18491), .B(n18490), .ZN(
        P3_U2824) );
  AOI21_X1 U21734 ( .B1(n18493), .B2(n18554), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18506) );
  AOI21_X1 U21735 ( .B1(n18496), .B2(n18495), .A(n18494), .ZN(n18813) );
  AOI22_X1 U21736 ( .A1(n18547), .A2(n18813), .B1(n18828), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18504) );
  AOI21_X1 U21737 ( .B1(n18499), .B2(n18498), .A(n18497), .ZN(n18500) );
  XOR2_X1 U21738 ( .A(n18500), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18810) );
  AOI22_X1 U21739 ( .A1(n18502), .A2(n18810), .B1(n18501), .B2(n18216), .ZN(
        n18503) );
  OAI211_X1 U21740 ( .C1(n18506), .C2(n18505), .A(n18504), .B(n18503), .ZN(
        P3_U2825) );
  AOI21_X1 U21741 ( .B1(n18811), .B2(n18508), .A(n18507), .ZN(n18827) );
  AOI22_X1 U21742 ( .A1(n18547), .A2(n18827), .B1(n18869), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n18517) );
  OAI21_X1 U21743 ( .B1(n9836), .B2(n18509), .A(n18554), .ZN(n18527) );
  INV_X1 U21744 ( .A(n18510), .ZN(n18514) );
  OAI21_X1 U21745 ( .B1(n18513), .B2(n18512), .A(n18511), .ZN(n18831) );
  OAI22_X1 U21746 ( .A1(n18538), .A2(n18514), .B1(n18558), .B2(n18831), .ZN(
        n18515) );
  AOI21_X1 U21747 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18527), .A(
        n18515), .ZN(n18516) );
  OAI211_X1 U21748 ( .C1(n18999), .C2(n18518), .A(n18517), .B(n18516), .ZN(
        P3_U2826) );
  AOI21_X1 U21749 ( .B1(n18521), .B2(n18520), .A(n18519), .ZN(n18835) );
  OAI21_X1 U21750 ( .B1(n18524), .B2(n18523), .A(n18522), .ZN(n18832) );
  OAI22_X1 U21751 ( .A1(n18558), .A2(n18832), .B1(n18833), .B2(n19426), .ZN(
        n18525) );
  AOI21_X1 U21752 ( .B1(n18547), .B2(n18835), .A(n18525), .ZN(n18529) );
  INV_X1 U21753 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18542) );
  NOR2_X1 U21754 ( .A1(n18526), .A2(n18542), .ZN(n18543) );
  OAI21_X1 U21755 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18543), .A(
        n18527), .ZN(n18528) );
  OAI211_X1 U21756 ( .C1(n18538), .C2(n18530), .A(n18529), .B(n18528), .ZN(
        P3_U2827) );
  AOI21_X1 U21757 ( .B1(n18533), .B2(n18532), .A(n18531), .ZN(n18848) );
  NAND2_X1 U21758 ( .A1(n18869), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18855) );
  INV_X1 U21759 ( .A(n18855), .ZN(n18540) );
  OAI21_X1 U21760 ( .B1(n18536), .B2(n18535), .A(n18534), .ZN(n18857) );
  OAI22_X1 U21761 ( .A1(n18538), .A2(n18537), .B1(n18558), .B2(n18857), .ZN(
        n18539) );
  AOI211_X1 U21762 ( .C1(n18547), .C2(n18848), .A(n18540), .B(n18539), .ZN(
        n18541) );
  OAI221_X1 U21763 ( .B1(n18543), .B2(n18999), .C1(n18543), .C2(n18542), .A(
        n18541), .ZN(P3_U2828) );
  OAI21_X1 U21764 ( .B1(n18545), .B2(n18552), .A(n18544), .ZN(n18860) );
  NAND2_X1 U21765 ( .A1(n19519), .A2(n18553), .ZN(n18546) );
  XNOR2_X1 U21766 ( .A(n18546), .B(n18545), .ZN(n18863) );
  AOI22_X1 U21767 ( .A1(n18547), .A2(n18863), .B1(n18828), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18551) );
  AOI22_X1 U21768 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18549), .B1(
        n18216), .B2(n18548), .ZN(n18550) );
  OAI211_X1 U21769 ( .C1(n18558), .C2(n18860), .A(n18551), .B(n18550), .ZN(
        P3_U2829) );
  AOI21_X1 U21770 ( .B1(n18553), .B2(n19519), .A(n18552), .ZN(n18879) );
  INV_X1 U21771 ( .A(n18879), .ZN(n18559) );
  NAND3_X1 U21772 ( .A1(n19503), .A2(n18555), .A3(n18554), .ZN(n18556) );
  AOI22_X1 U21773 ( .A1(n18869), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18556), .ZN(n18557) );
  OAI221_X1 U21774 ( .B1(n18879), .B2(n18560), .C1(n18559), .C2(n18558), .A(
        n18557), .ZN(P3_U2830) );
  NOR2_X1 U21775 ( .A1(n18561), .A2(n18564), .ZN(n18633) );
  NAND2_X1 U21776 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18633), .ZN(
        n18617) );
  NOR2_X1 U21777 ( .A1(n18562), .A2(n18617), .ZN(n18574) );
  NOR2_X1 U21778 ( .A1(n19331), .A2(n19358), .ZN(n18846) );
  INV_X1 U21779 ( .A(n18846), .ZN(n18821) );
  OAI21_X1 U21780 ( .B1(n18636), .B2(n19358), .A(n18563), .ZN(n18630) );
  OAI21_X1 U21781 ( .B1(n18625), .B2(n18564), .A(n19331), .ZN(n18565) );
  OAI21_X1 U21782 ( .B1(n18846), .B2(n18630), .A(n18565), .ZN(n18606) );
  AOI21_X1 U21783 ( .B1(n18566), .B2(n18821), .A(n18606), .ZN(n18591) );
  AOI21_X1 U21784 ( .B1(n18568), .B2(n18821), .A(n18567), .ZN(n18569) );
  OAI211_X1 U21785 ( .C1(n18570), .C2(n18601), .A(n18591), .B(n18569), .ZN(
        n18571) );
  AOI21_X1 U21786 ( .B1(n18730), .B2(n18572), .A(n18571), .ZN(n18579) );
  INV_X1 U21787 ( .A(n18579), .ZN(n18573) );
  MUX2_X1 U21788 ( .A(n18574), .B(n18573), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n18575) );
  AOI22_X1 U21789 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18873), .B1(
        n18854), .B2(n18575), .ZN(n18577) );
  NAND2_X1 U21790 ( .A1(n18869), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18576) );
  OAI211_X1 U21791 ( .C1(n18578), .C2(n18740), .A(n18577), .B(n18576), .ZN(
        P3_U2835) );
  AOI221_X1 U21792 ( .B1(n18580), .B2(n18585), .C1(n18617), .C2(n18585), .A(
        n18579), .ZN(n18582) );
  AOI22_X1 U21793 ( .A1(n18854), .A2(n18582), .B1(n18788), .B2(n18581), .ZN(
        n18584) );
  OAI211_X1 U21794 ( .C1(n18841), .C2(n18585), .A(n18584), .B(n18583), .ZN(
        P3_U2836) );
  INV_X1 U21795 ( .A(n18586), .ZN(n18589) );
  AOI221_X1 U21796 ( .B1(n18589), .B2(n18588), .C1(n18587), .C2(n18588), .A(
        n18871), .ZN(n18593) );
  NAND3_X1 U21797 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18591), .A3(
        n18590), .ZN(n18592) );
  AOI22_X1 U21798 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18873), .B1(
        n18593), .B2(n18592), .ZN(n18595) );
  OAI211_X1 U21799 ( .C1(n18596), .C2(n18740), .A(n18595), .B(n18594), .ZN(
        n18597) );
  AOI21_X1 U21800 ( .B1(n18725), .B2(n18598), .A(n18597), .ZN(n18599) );
  OAI21_X1 U21801 ( .B1(n18878), .B2(n18600), .A(n18599), .ZN(P3_U2837) );
  OAI22_X1 U21802 ( .A1(n18604), .A2(n18603), .B1(n18602), .B2(n18601), .ZN(
        n18605) );
  NOR3_X1 U21803 ( .A1(n18873), .A2(n18606), .A3(n18605), .ZN(n18610) );
  AOI21_X1 U21804 ( .B1(n19334), .B2(n18607), .A(n21089), .ZN(n18608) );
  AOI21_X1 U21805 ( .B1(n18610), .B2(n18608), .A(n18828), .ZN(n18619) );
  AOI21_X1 U21806 ( .B1(n18783), .B2(n18610), .A(n18609), .ZN(n18611) );
  AOI22_X1 U21807 ( .A1(n18788), .A2(n18612), .B1(n18619), .B2(n18611), .ZN(
        n18614) );
  OAI211_X1 U21808 ( .C1(n18616), .C2(n18615), .A(n18614), .B(n18613), .ZN(
        P3_U2838) );
  OAI21_X1 U21809 ( .B1(n18873), .B2(n18617), .A(n21089), .ZN(n18618) );
  AOI22_X1 U21810 ( .A1(n18869), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18619), 
        .B2(n18618), .ZN(n18620) );
  OAI21_X1 U21811 ( .B1(n18740), .B2(n18621), .A(n18620), .ZN(P3_U2839) );
  AOI22_X1 U21812 ( .A1(n18869), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n18788), 
        .B2(n18622), .ZN(n18635) );
  AOI22_X1 U21813 ( .A1(n19320), .A2(n18623), .B1(n18730), .B2(n18697), .ZN(
        n18639) );
  OAI21_X1 U21814 ( .B1(n18625), .B2(n18624), .A(n19331), .ZN(n18626) );
  OAI221_X1 U21815 ( .B1(n19353), .B2(n18638), .C1(n19353), .C2(n18627), .A(
        n18626), .ZN(n18640) );
  NOR2_X1 U21816 ( .A1(n19320), .A2(n18730), .ZN(n18755) );
  OAI22_X1 U21817 ( .A1(n19360), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18628), .B2(n18755), .ZN(n18644) );
  AOI211_X1 U21818 ( .C1(n18763), .C2(n18629), .A(n18640), .B(n18644), .ZN(
        n18631) );
  NAND3_X1 U21819 ( .A1(n18639), .A2(n18631), .A3(n18630), .ZN(n18632) );
  OAI211_X1 U21820 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18633), .A(
        n18854), .B(n18632), .ZN(n18634) );
  OAI211_X1 U21821 ( .C1(n18841), .C2(n18636), .A(n18635), .B(n18634), .ZN(
        P3_U2840) );
  AOI22_X1 U21822 ( .A1(n18869), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18656), 
        .B2(n18637), .ZN(n18646) );
  NOR2_X1 U21823 ( .A1(n19334), .A2(n19358), .ZN(n18859) );
  AOI21_X1 U21824 ( .B1(n18638), .B2(n18686), .A(n19345), .ZN(n18641) );
  NAND2_X1 U21825 ( .A1(n18854), .A2(n18639), .ZN(n18691) );
  NOR3_X1 U21826 ( .A1(n18641), .A2(n18691), .A3(n18640), .ZN(n18650) );
  OAI21_X1 U21827 ( .B1(n18642), .B2(n18859), .A(n18650), .ZN(n18643) );
  OAI211_X1 U21828 ( .C1(n18644), .C2(n18643), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18833), .ZN(n18645) );
  OAI211_X1 U21829 ( .C1(n18647), .C2(n18740), .A(n18646), .B(n18645), .ZN(
        P3_U2841) );
  AOI22_X1 U21830 ( .A1(n18788), .A2(n18649), .B1(n18656), .B2(n18648), .ZN(
        n18654) );
  AOI221_X1 U21831 ( .B1(n18651), .B2(n18650), .C1(n18755), .C2(n18650), .A(
        n18869), .ZN(n18657) );
  NOR3_X1 U21832 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18859), .A3(
        n19393), .ZN(n18652) );
  OAI21_X1 U21833 ( .B1(n18657), .B2(n18652), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18653) );
  OAI211_X1 U21834 ( .C1(n19455), .C2(n18833), .A(n18654), .B(n18653), .ZN(
        P3_U2842) );
  AOI22_X1 U21835 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18657), .B1(
        n18656), .B2(n18655), .ZN(n18659) );
  OAI211_X1 U21836 ( .C1(n18660), .C2(n18740), .A(n18659), .B(n18658), .ZN(
        P3_U2843) );
  NOR2_X1 U21837 ( .A1(n19345), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18781) );
  INV_X1 U21838 ( .A(n18781), .ZN(n18845) );
  NAND3_X1 U21839 ( .A1(n18661), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18845), .ZN(n18666) );
  AOI21_X1 U21840 ( .B1(n19334), .B2(n18663), .A(n18662), .ZN(n18664) );
  AOI21_X1 U21841 ( .B1(n18755), .B2(n19353), .A(n18664), .ZN(n18665) );
  AOI211_X1 U21842 ( .C1(n18821), .C2(n18666), .A(n18665), .B(n18691), .ZN(
        n18677) );
  AOI221_X1 U21843 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18677), 
        .C1(n18846), .C2(n18677), .A(n18869), .ZN(n18673) );
  INV_X1 U21844 ( .A(n18667), .ZN(n18670) );
  OAI22_X1 U21845 ( .A1(n18844), .A2(n19353), .B1(n18852), .B2(n18820), .ZN(
        n18837) );
  INV_X1 U21846 ( .A(n18837), .ZN(n18819) );
  NOR2_X1 U21847 ( .A1(n18819), .A2(n18668), .ZN(n18794) );
  NAND2_X1 U21848 ( .A1(n18669), .A2(n18794), .ZN(n18717) );
  NAND2_X1 U21849 ( .A1(n18670), .A2(n18717), .ZN(n18742) );
  NAND2_X1 U21850 ( .A1(n18854), .A2(n18742), .ZN(n18777) );
  NOR2_X1 U21851 ( .A1(n18671), .A2(n18777), .ZN(n18693) );
  AOI22_X1 U21852 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18673), .B1(
        n18693), .B2(n18672), .ZN(n18675) );
  OAI211_X1 U21853 ( .C1(n18740), .C2(n18676), .A(n18675), .B(n18674), .ZN(
        P3_U2844) );
  NOR2_X1 U21854 ( .A1(n18828), .A2(n18677), .ZN(n18679) );
  AOI22_X1 U21855 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18679), .B1(
        n18693), .B2(n18678), .ZN(n18682) );
  INV_X1 U21856 ( .A(n18680), .ZN(n18681) );
  OAI211_X1 U21857 ( .C1(n18683), .C2(n18740), .A(n18682), .B(n18681), .ZN(
        P3_U2845) );
  AOI22_X1 U21858 ( .A1(n19334), .A2(n18685), .B1(n19331), .B2(n18684), .ZN(
        n18752) );
  INV_X1 U21859 ( .A(n18686), .ZN(n18687) );
  OAI21_X1 U21860 ( .B1(n18699), .B2(n19358), .A(n18687), .ZN(n18688) );
  OAI211_X1 U21861 ( .C1(n18758), .C2(n18689), .A(n18752), .B(n18688), .ZN(
        n18702) );
  OAI221_X1 U21862 ( .B1(n18691), .B2(n18690), .C1(n18691), .C2(n18702), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18696) );
  AOI22_X1 U21863 ( .A1(n18788), .A2(n18694), .B1(n18693), .B2(n18692), .ZN(
        n18695) );
  OAI221_X1 U21864 ( .B1(n18828), .B2(n18696), .C1(n18833), .C2(n19447), .A(
        n18695), .ZN(P3_U2846) );
  AND2_X1 U21865 ( .A1(n18697), .A2(n18730), .ZN(n18704) );
  INV_X1 U21866 ( .A(n18698), .ZN(n18703) );
  OAI21_X1 U21867 ( .B1(n18700), .B2(n18717), .A(n18699), .ZN(n18701) );
  AOI22_X1 U21868 ( .A1(n18704), .A2(n18703), .B1(n18702), .B2(n18701), .ZN(
        n18711) );
  AOI22_X1 U21869 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18873), .B1(
        n18869), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18710) );
  NOR2_X1 U21870 ( .A1(n18705), .A2(n18878), .ZN(n18707) );
  AOI22_X1 U21871 ( .A1(n18788), .A2(n18708), .B1(n18707), .B2(n18706), .ZN(
        n18709) );
  OAI211_X1 U21872 ( .C1(n18711), .C2(n18871), .A(n18710), .B(n18709), .ZN(
        P3_U2847) );
  AOI22_X1 U21873 ( .A1(n19345), .A2(n18752), .B1(n18732), .B2(n18712), .ZN(
        n18734) );
  INV_X1 U21874 ( .A(n18718), .ZN(n18713) );
  OAI22_X1 U21875 ( .A1(n19360), .A2(n18713), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18859), .ZN(n18714) );
  INV_X1 U21876 ( .A(n18714), .ZN(n18715) );
  OAI211_X1 U21877 ( .C1(n18732), .C2(n19353), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18715), .ZN(n18716) );
  OAI21_X1 U21878 ( .B1(n18734), .B2(n18716), .A(n18854), .ZN(n18720) );
  OR2_X1 U21879 ( .A1(n18718), .A2(n18717), .ZN(n18719) );
  AOI222_X1 U21880 ( .A1(n18721), .A2(n18720), .B1(n18721), .B2(n18719), .C1(
        n18720), .C2(n18841), .ZN(n18722) );
  AOI21_X1 U21881 ( .B1(n18828), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18722), 
        .ZN(n18727) );
  AOI22_X1 U21882 ( .A1(n18725), .A2(n18724), .B1(n18788), .B2(n18723), .ZN(
        n18726) );
  OAI211_X1 U21883 ( .C1(n18878), .C2(n18728), .A(n18727), .B(n18726), .ZN(
        P3_U2848) );
  AOI22_X1 U21884 ( .A1(n19320), .A2(n18731), .B1(n18730), .B2(n18729), .ZN(
        n18751) );
  OAI21_X1 U21885 ( .B1(n18732), .B2(n18755), .A(n18751), .ZN(n18733) );
  AOI211_X1 U21886 ( .C1(n18763), .C2(n18736), .A(n18734), .B(n18733), .ZN(
        n18744) );
  OAI211_X1 U21887 ( .C1(n18758), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18854), .B(n18744), .ZN(n18735) );
  OAI221_X1 U21888 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n18833), .C1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18828), .A(n18735), .ZN(
        n18739) );
  INV_X1 U21889 ( .A(n18736), .ZN(n18757) );
  NAND4_X1 U21890 ( .A1(n18854), .A2(n18757), .A3(n18737), .A4(n18742), .ZN(
        n18738) );
  OAI211_X1 U21891 ( .C1(n18741), .C2(n18740), .A(n18739), .B(n18738), .ZN(
        P3_U2849) );
  NAND2_X1 U21892 ( .A1(n18757), .A2(n18742), .ZN(n18743) );
  AOI221_X1 U21893 ( .B1(n18744), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), 
        .C1(n18743), .C2(n18749), .A(n18871), .ZN(n18745) );
  AOI21_X1 U21894 ( .B1(n18788), .B2(n18746), .A(n18745), .ZN(n18748) );
  OAI211_X1 U21895 ( .C1(n18841), .C2(n18749), .A(n18748), .B(n18747), .ZN(
        P3_U2850) );
  AOI22_X1 U21896 ( .A1(n18869), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18788), 
        .B2(n18750), .ZN(n18761) );
  NAND2_X1 U21897 ( .A1(n18854), .A2(n18751), .ZN(n18772) );
  INV_X1 U21898 ( .A(n18772), .ZN(n18754) );
  NAND2_X1 U21899 ( .A1(n19345), .A2(n18752), .ZN(n18770) );
  OAI21_X1 U21900 ( .B1(n18771), .B2(n18776), .A(n18770), .ZN(n18753) );
  OAI211_X1 U21901 ( .C1(n18756), .C2(n18755), .A(n18754), .B(n18753), .ZN(
        n18764) );
  OAI22_X1 U21902 ( .A1(n18758), .A2(n18757), .B1(n19345), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18759) );
  OAI211_X1 U21903 ( .C1(n18764), .C2(n18759), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18833), .ZN(n18760) );
  OAI211_X1 U21904 ( .C1(n18762), .C2(n18777), .A(n18761), .B(n18760), .ZN(
        P3_U2851) );
  OAI221_X1 U21905 ( .B1(n18764), .B2(n18763), .C1(n18764), .C2(n18776), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18769) );
  INV_X1 U21906 ( .A(n18777), .ZN(n18766) );
  NOR2_X1 U21907 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18776), .ZN(
        n18765) );
  AOI22_X1 U21908 ( .A1(n18788), .A2(n18767), .B1(n18766), .B2(n18765), .ZN(
        n18768) );
  OAI221_X1 U21909 ( .B1(n18828), .B2(n18769), .C1(n18833), .C2(n19439), .A(
        n18768), .ZN(P3_U2852) );
  OAI221_X1 U21910 ( .B1(n18772), .B2(n18771), .C1(n18772), .C2(n18770), .A(
        n18833), .ZN(n18775) );
  AOI22_X1 U21911 ( .A1(n18869), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18788), 
        .B2(n18773), .ZN(n18774) );
  OAI221_X1 U21912 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18777), .C1(
        n18776), .C2(n18775), .A(n18774), .ZN(P3_U2853) );
  NAND2_X1 U21913 ( .A1(n18854), .A2(n18794), .ZN(n18809) );
  NOR3_X1 U21914 ( .A1(n21225), .A2(n18808), .A3(n18809), .ZN(n18786) );
  OAI22_X1 U21915 ( .A1(n18779), .A2(n19353), .B1(n18846), .B2(n18778), .ZN(
        n18780) );
  NOR2_X1 U21916 ( .A1(n18781), .A2(n18780), .ZN(n18802) );
  OAI211_X1 U21917 ( .C1(n18783), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18802), .ZN(n18782) );
  NAND2_X1 U21918 ( .A1(n18854), .A2(n18782), .ZN(n18800) );
  OAI21_X1 U21919 ( .B1(n18783), .B2(n18800), .A(n18841), .ZN(n18785) );
  NOR2_X1 U21920 ( .A1(n18833), .A2(n21222), .ZN(n18784) );
  AOI221_X1 U21921 ( .B1(n18786), .B2(n21202), .C1(n18785), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18784), .ZN(n18791) );
  AOI22_X1 U21922 ( .A1(n18864), .A2(n18789), .B1(n18788), .B2(n18787), .ZN(
        n18790) );
  OAI211_X1 U21923 ( .C1(n18793), .C2(n18792), .A(n18791), .B(n18790), .ZN(
        P3_U2854) );
  AOI21_X1 U21924 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18794), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18801) );
  NOR2_X1 U21925 ( .A1(n18833), .A2(n19434), .ZN(n18798) );
  INV_X1 U21926 ( .A(n18868), .ZN(n18861) );
  OAI22_X1 U21927 ( .A1(n18878), .A2(n18796), .B1(n18861), .B2(n18795), .ZN(
        n18797) );
  AOI211_X1 U21928 ( .C1(n18873), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18798), .B(n18797), .ZN(n18799) );
  OAI21_X1 U21929 ( .B1(n18801), .B2(n18800), .A(n18799), .ZN(P3_U2855) );
  AOI21_X1 U21930 ( .B1(n18854), .B2(n18802), .A(n18828), .ZN(n18803) );
  INV_X1 U21931 ( .A(n18803), .ZN(n18816) );
  OAI22_X1 U21932 ( .A1(n18833), .A2(n19432), .B1(n18861), .B2(n18804), .ZN(
        n18805) );
  AOI21_X1 U21933 ( .B1(n18864), .B2(n18806), .A(n18805), .ZN(n18807) );
  OAI221_X1 U21934 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18809), .C1(
        n18808), .C2(n18816), .A(n18807), .ZN(P3_U2856) );
  AOI22_X1 U21935 ( .A1(n18869), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18868), 
        .B2(n18810), .ZN(n18815) );
  NOR4_X1 U21936 ( .A1(n18819), .A2(n18811), .A3(n18840), .A4(n18871), .ZN(
        n18812) );
  AOI22_X1 U21937 ( .A1(n18813), .A2(n18864), .B1(n18812), .B2(n18817), .ZN(
        n18814) );
  OAI211_X1 U21938 ( .C1(n18817), .C2(n18816), .A(n18815), .B(n18814), .ZN(
        P3_U2857) );
  NAND2_X1 U21939 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18854), .ZN(
        n18818) );
  NOR2_X1 U21940 ( .A1(n18819), .A2(n18818), .ZN(n18825) );
  AOI22_X1 U21941 ( .A1(n19334), .A2(n18844), .B1(n18821), .B2(n18820), .ZN(
        n18822) );
  NAND3_X1 U21942 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18822), .A3(
        n18845), .ZN(n18836) );
  AOI21_X1 U21943 ( .B1(n18858), .B2(n18836), .A(n18873), .ZN(n18823) );
  INV_X1 U21944 ( .A(n18823), .ZN(n18824) );
  MUX2_X1 U21945 ( .A(n18825), .B(n18824), .S(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n18826) );
  AOI21_X1 U21946 ( .B1(n18864), .B2(n18827), .A(n18826), .ZN(n18830) );
  NAND2_X1 U21947 ( .A1(n18828), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18829) );
  OAI211_X1 U21948 ( .C1(n18831), .C2(n18861), .A(n18830), .B(n18829), .ZN(
        P3_U2858) );
  OAI22_X1 U21949 ( .A1(n18833), .A2(n19426), .B1(n18861), .B2(n18832), .ZN(
        n18834) );
  AOI21_X1 U21950 ( .B1(n18864), .B2(n18835), .A(n18834), .ZN(n18839) );
  OAI211_X1 U21951 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18837), .A(
        n18854), .B(n18836), .ZN(n18838) );
  OAI211_X1 U21952 ( .C1(n18841), .C2(n18840), .A(n18839), .B(n18838), .ZN(
        P3_U2859) );
  NAND2_X1 U21953 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18842), .ZN(
        n18851) );
  INV_X1 U21954 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19504) );
  NOR2_X1 U21955 ( .A1(n19519), .A2(n19504), .ZN(n18843) );
  OAI221_X1 U21956 ( .B1(n18844), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18844), .C2(n18843), .A(n19334), .ZN(n18850) );
  OAI21_X1 U21957 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18846), .A(
        n18845), .ZN(n18847) );
  AOI22_X1 U21958 ( .A1(n19320), .A2(n18848), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18847), .ZN(n18849) );
  OAI211_X1 U21959 ( .C1(n18852), .C2(n18851), .A(n18850), .B(n18849), .ZN(
        n18853) );
  AOI22_X1 U21960 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18873), .B1(
        n18854), .B2(n18853), .ZN(n18856) );
  OAI211_X1 U21961 ( .C1(n18857), .C2(n18861), .A(n18856), .B(n18855), .ZN(
        P3_U2860) );
  OAI21_X1 U21962 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19331), .A(
        n18858), .ZN(n18867) );
  NOR2_X1 U21963 ( .A1(n18859), .A2(n18871), .ZN(n18870) );
  AOI21_X1 U21964 ( .B1(n18870), .B2(n19519), .A(n18873), .ZN(n18866) );
  OAI22_X1 U21965 ( .A1(n18833), .A2(n19423), .B1(n18861), .B2(n18860), .ZN(
        n18862) );
  AOI21_X1 U21966 ( .B1(n18864), .B2(n18863), .A(n18862), .ZN(n18865) );
  OAI221_X1 U21967 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18867), .C1(
        n19504), .C2(n18866), .A(n18865), .ZN(P3_U2861) );
  AOI22_X1 U21968 ( .A1(n18869), .A2(P3_REIP_REG_0__SCAN_IN), .B1(n18868), 
        .B2(n18879), .ZN(n18877) );
  INV_X1 U21969 ( .A(n18870), .ZN(n18875) );
  NOR2_X1 U21970 ( .A1(n19360), .A2(n18871), .ZN(n18872) );
  NOR2_X1 U21971 ( .A1(n18873), .A2(n18872), .ZN(n18874) );
  MUX2_X1 U21972 ( .A(n18875), .B(n18874), .S(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n18876) );
  OAI211_X1 U21973 ( .C1(n18879), .C2(n18878), .A(n18877), .B(n18876), .ZN(
        P3_U2862) );
  AOI211_X1 U21974 ( .C1(n18881), .C2(n18880), .A(n19393), .B(n19503), .ZN(
        n19386) );
  OAI21_X1 U21975 ( .B1(n19386), .B2(n18934), .A(n18886), .ZN(n18882) );
  OAI221_X1 U21976 ( .B1(n19364), .B2(n19534), .C1(n19364), .C2(n18886), .A(
        n18882), .ZN(P3_U2863) );
  INV_X1 U21977 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19374) );
  NOR2_X1 U21978 ( .A1(n19371), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19071) );
  NOR2_X1 U21979 ( .A1(n19374), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19160) );
  NOR2_X1 U21980 ( .A1(n19071), .A2(n19160), .ZN(n18884) );
  OAI22_X1 U21981 ( .A1(n18885), .A2(n19374), .B1(n18884), .B2(n18883), .ZN(
        P3_U2866) );
  NOR2_X1 U21982 ( .A1(n19375), .A2(n18886), .ZN(P3_U2867) );
  NOR2_X1 U21983 ( .A1(n19374), .A2(n19047), .ZN(n19263) );
  NAND2_X1 U21984 ( .A1(n19263), .A2(n19364), .ZN(n19252) );
  INV_X1 U21985 ( .A(n19252), .ZN(n19254) );
  NOR3_X1 U21986 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19371), .A3(
        n19374), .ZN(n19264) );
  NAND2_X1 U21987 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19264), .ZN(
        n19299) );
  INV_X1 U21988 ( .A(n19299), .ZN(n19309) );
  NOR2_X1 U21989 ( .A1(n19254), .A2(n19309), .ZN(n19226) );
  NAND2_X1 U21990 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19263), .ZN(
        n19307) );
  INV_X1 U21991 ( .A(n19307), .ZN(n19313) );
  NAND2_X1 U21992 ( .A1(n19366), .A2(n19364), .ZN(n19367) );
  NOR2_X1 U21993 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18978) );
  INV_X1 U21994 ( .A(n18978), .ZN(n18957) );
  NOR2_X2 U21995 ( .A1(n19367), .A2(n18957), .ZN(n18991) );
  NOR2_X1 U21996 ( .A1(n19313), .A2(n18991), .ZN(n18958) );
  INV_X1 U21997 ( .A(n18887), .ZN(n18888) );
  OAI22_X1 U21998 ( .A1(n19227), .A2(n19226), .B1(n18958), .B2(n18888), .ZN(
        n18889) );
  AND2_X1 U21999 ( .A1(n18889), .A2(n19230), .ZN(n18933) );
  NAND2_X1 U22000 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19265), .ZN(n19234) );
  INV_X1 U22001 ( .A(n19234), .ZN(n19261) );
  NOR2_X2 U22002 ( .A1(n19001), .A2(n18890), .ZN(n19260) );
  INV_X1 U22003 ( .A(n19259), .ZN(n19394) );
  NOR2_X1 U22004 ( .A1(n19394), .A2(n18958), .ZN(n18927) );
  AOI22_X1 U22005 ( .A1(n19261), .A2(n19309), .B1(n19260), .B2(n18927), .ZN(
        n18896) );
  NAND2_X1 U22006 ( .A1(n18892), .A2(n18891), .ZN(n18928) );
  NOR2_X1 U22007 ( .A1(n18893), .A2(n18928), .ZN(n19231) );
  INV_X1 U22008 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18894) );
  NOR2_X2 U22009 ( .A1(n18999), .A2(n18894), .ZN(n19266) );
  AOI22_X1 U22010 ( .A1(n19231), .A2(n18991), .B1(n19266), .B2(n19254), .ZN(
        n18895) );
  OAI211_X1 U22011 ( .C1(n18933), .C2(n18897), .A(n18896), .B(n18895), .ZN(
        P3_U2868) );
  INV_X1 U22012 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18898) );
  NOR2_X2 U22013 ( .A1(n18999), .A2(n18898), .ZN(n19271) );
  NOR2_X2 U22014 ( .A1(n19001), .A2(n18899), .ZN(n19270) );
  AOI22_X1 U22015 ( .A1(n19271), .A2(n19254), .B1(n19270), .B2(n18927), .ZN(
        n18901) );
  NOR2_X1 U22016 ( .A1(n18928), .A2(n19539), .ZN(n18937) );
  AND2_X1 U22017 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19265), .ZN(n19272) );
  AOI22_X1 U22018 ( .A1(n18937), .A2(n18991), .B1(n19272), .B2(n19309), .ZN(
        n18900) );
  OAI211_X1 U22019 ( .C1(n18933), .C2(n18902), .A(n18901), .B(n18900), .ZN(
        P3_U2869) );
  INV_X1 U22020 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18907) );
  NOR2_X2 U22021 ( .A1(n18999), .A2(n16157), .ZN(n19277) );
  NOR2_X2 U22022 ( .A1(n19001), .A2(n18903), .ZN(n19276) );
  AOI22_X1 U22023 ( .A1(n19277), .A2(n19254), .B1(n19276), .B2(n18927), .ZN(
        n18906) );
  NOR2_X1 U22024 ( .A1(n18928), .A2(n18904), .ZN(n18940) );
  AND2_X1 U22025 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19265), .ZN(n19278) );
  AOI22_X1 U22026 ( .A1(n18940), .A2(n18991), .B1(n19278), .B2(n19309), .ZN(
        n18905) );
  OAI211_X1 U22027 ( .C1(n18933), .C2(n18907), .A(n18906), .B(n18905), .ZN(
        P3_U2870) );
  NOR2_X1 U22028 ( .A1(n21078), .A2(n18999), .ZN(n19239) );
  NOR2_X2 U22029 ( .A1(n19001), .A2(n18908), .ZN(n19283) );
  AOI22_X1 U22030 ( .A1(n19239), .A2(n19309), .B1(n19283), .B2(n18927), .ZN(
        n18911) );
  NOR2_X2 U22031 ( .A1(n18909), .A2(n18928), .ZN(n19284) );
  NAND2_X1 U22032 ( .A1(n19265), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19242) );
  INV_X1 U22033 ( .A(n19242), .ZN(n19282) );
  AOI22_X1 U22034 ( .A1(n19284), .A2(n18991), .B1(n19282), .B2(n19254), .ZN(
        n18910) );
  OAI211_X1 U22035 ( .C1(n18933), .C2(n18912), .A(n18911), .B(n18910), .ZN(
        P3_U2871) );
  NOR2_X2 U22036 ( .A1(n18999), .A2(n16139), .ZN(n19289) );
  NOR2_X2 U22037 ( .A1(n19001), .A2(n18913), .ZN(n19288) );
  AOI22_X1 U22038 ( .A1(n19289), .A2(n19254), .B1(n19288), .B2(n18927), .ZN(
        n18916) );
  NOR2_X1 U22039 ( .A1(n18928), .A2(n18914), .ZN(n18945) );
  INV_X1 U22040 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21208) );
  NOR2_X2 U22041 ( .A1(n21208), .A2(n18999), .ZN(n19290) );
  AOI22_X1 U22042 ( .A1(n18945), .A2(n18991), .B1(n19290), .B2(n19309), .ZN(
        n18915) );
  OAI211_X1 U22043 ( .C1(n18933), .C2(n21173), .A(n18916), .B(n18915), .ZN(
        P3_U2872) );
  NOR2_X2 U22044 ( .A1(n19001), .A2(n21293), .ZN(n19294) );
  NAND2_X1 U22045 ( .A1(n19265), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19300) );
  INV_X1 U22046 ( .A(n19300), .ZN(n19245) );
  AOI22_X1 U22047 ( .A1(n19294), .A2(n18927), .B1(n19245), .B2(n19254), .ZN(
        n18919) );
  NAND2_X1 U22048 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19265), .ZN(n19248) );
  INV_X1 U22049 ( .A(n19248), .ZN(n19295) );
  NOR2_X2 U22050 ( .A1(n18917), .A2(n18928), .ZN(n19296) );
  AOI22_X1 U22051 ( .A1(n19295), .A2(n19309), .B1(n19296), .B2(n18991), .ZN(
        n18918) );
  OAI211_X1 U22052 ( .C1(n18933), .C2(n18920), .A(n18919), .B(n18918), .ZN(
        P3_U2873) );
  NOR2_X2 U22053 ( .A1(n16122), .A2(n18999), .ZN(n19302) );
  NOR2_X2 U22054 ( .A1(n18921), .A2(n19001), .ZN(n19301) );
  AOI22_X1 U22055 ( .A1(n19302), .A2(n19254), .B1(n19301), .B2(n18927), .ZN(
        n18924) );
  NOR2_X1 U22056 ( .A1(n18928), .A2(n18922), .ZN(n18950) );
  NOR2_X2 U22057 ( .A1(n19894), .A2(n18999), .ZN(n19304) );
  AOI22_X1 U22058 ( .A1(n18950), .A2(n18991), .B1(n19304), .B2(n19309), .ZN(
        n18923) );
  OAI211_X1 U22059 ( .C1(n18933), .C2(n18925), .A(n18924), .B(n18923), .ZN(
        P3_U2874) );
  NOR2_X2 U22060 ( .A1(n18926), .A2(n19001), .ZN(n19312) );
  NAND2_X1 U22061 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19265), .ZN(n19225) );
  INV_X1 U22062 ( .A(n19225), .ZN(n19310) );
  AOI22_X1 U22063 ( .A1(n19312), .A2(n18927), .B1(n19310), .B2(n19254), .ZN(
        n18931) );
  NOR2_X1 U22064 ( .A1(n18999), .A2(n19901), .ZN(n19221) );
  NOR2_X2 U22065 ( .A1(n18929), .A2(n18928), .ZN(n19314) );
  AOI22_X1 U22066 ( .A1(n19221), .A2(n19309), .B1(n19314), .B2(n18991), .ZN(
        n18930) );
  OAI211_X1 U22067 ( .C1(n18933), .C2(n18932), .A(n18931), .B(n18930), .ZN(
        P3_U2875) );
  NAND2_X1 U22068 ( .A1(n19366), .A2(n19259), .ZN(n19113) );
  NOR2_X1 U22069 ( .A1(n18957), .A2(n19113), .ZN(n18953) );
  AOI22_X1 U22070 ( .A1(n19260), .A2(n18953), .B1(n19266), .B2(n19313), .ZN(
        n18936) );
  NOR2_X1 U22071 ( .A1(n19001), .A2(n18934), .ZN(n19262) );
  AND2_X1 U22072 ( .A1(n19366), .A2(n19262), .ZN(n19114) );
  AOI22_X1 U22073 ( .A1(n19265), .A2(n19263), .B1(n18978), .B2(n19114), .ZN(
        n18954) );
  NAND2_X1 U22074 ( .A1(n19366), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19024) );
  INV_X1 U22075 ( .A(n19024), .ZN(n19116) );
  NAND2_X1 U22076 ( .A1(n19116), .A2(n18978), .ZN(n19023) );
  INV_X1 U22077 ( .A(n19023), .ZN(n19015) );
  AOI22_X1 U22078 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18954), .B1(
        n19231), .B2(n19015), .ZN(n18935) );
  OAI211_X1 U22079 ( .C1(n19234), .C2(n19252), .A(n18936), .B(n18935), .ZN(
        P3_U2876) );
  INV_X1 U22080 ( .A(n18937), .ZN(n19275) );
  AOI22_X1 U22081 ( .A1(n19270), .A2(n18953), .B1(n19272), .B2(n19254), .ZN(
        n18939) );
  AOI22_X1 U22082 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18954), .B1(
        n19271), .B2(n19313), .ZN(n18938) );
  OAI211_X1 U22083 ( .C1(n19275), .C2(n19023), .A(n18939), .B(n18938), .ZN(
        P3_U2877) );
  AOI22_X1 U22084 ( .A1(n19277), .A2(n19313), .B1(n19276), .B2(n18953), .ZN(
        n18942) );
  AOI22_X1 U22085 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18954), .B1(
        n19278), .B2(n19254), .ZN(n18941) );
  OAI211_X1 U22086 ( .C1(n19281), .C2(n19023), .A(n18942), .B(n18941), .ZN(
        P3_U2878) );
  INV_X1 U22087 ( .A(n19239), .ZN(n19287) );
  AOI22_X1 U22088 ( .A1(n19283), .A2(n18953), .B1(n19282), .B2(n19313), .ZN(
        n18944) );
  AOI22_X1 U22089 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18954), .B1(
        n19284), .B2(n19015), .ZN(n18943) );
  OAI211_X1 U22090 ( .C1(n19287), .C2(n19252), .A(n18944), .B(n18943), .ZN(
        P3_U2879) );
  INV_X1 U22091 ( .A(n18945), .ZN(n19293) );
  AOI22_X1 U22092 ( .A1(n19290), .A2(n19254), .B1(n19288), .B2(n18953), .ZN(
        n18947) );
  AOI22_X1 U22093 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18954), .B1(
        n19289), .B2(n19313), .ZN(n18946) );
  OAI211_X1 U22094 ( .C1(n19293), .C2(n19023), .A(n18947), .B(n18946), .ZN(
        P3_U2880) );
  AOI22_X1 U22095 ( .A1(n19295), .A2(n19254), .B1(n19294), .B2(n18953), .ZN(
        n18949) );
  AOI22_X1 U22096 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18954), .B1(
        n19296), .B2(n19015), .ZN(n18948) );
  OAI211_X1 U22097 ( .C1(n19300), .C2(n19307), .A(n18949), .B(n18948), .ZN(
        P3_U2881) );
  INV_X1 U22098 ( .A(n18950), .ZN(n19308) );
  AOI22_X1 U22099 ( .A1(n19304), .A2(n19254), .B1(n19301), .B2(n18953), .ZN(
        n18952) );
  AOI22_X1 U22100 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18954), .B1(
        n19302), .B2(n19313), .ZN(n18951) );
  OAI211_X1 U22101 ( .C1(n19308), .C2(n19023), .A(n18952), .B(n18951), .ZN(
        P3_U2882) );
  INV_X1 U22102 ( .A(n19221), .ZN(n19319) );
  AOI22_X1 U22103 ( .A1(n19312), .A2(n18953), .B1(n19310), .B2(n19313), .ZN(
        n18956) );
  AOI22_X1 U22104 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18954), .B1(
        n19314), .B2(n19015), .ZN(n18955) );
  OAI211_X1 U22105 ( .C1(n19319), .C2(n19252), .A(n18956), .B(n18955), .ZN(
        P3_U2883) );
  INV_X1 U22106 ( .A(n19231), .ZN(n19269) );
  NOR2_X1 U22107 ( .A1(n19366), .A2(n18957), .ZN(n19026) );
  NAND2_X1 U22108 ( .A1(n19026), .A2(n19364), .ZN(n19046) );
  INV_X1 U22109 ( .A(n19046), .ZN(n19039) );
  NOR2_X1 U22110 ( .A1(n19015), .A2(n19039), .ZN(n19000) );
  NOR2_X1 U22111 ( .A1(n19394), .A2(n19000), .ZN(n18974) );
  AOI22_X1 U22112 ( .A1(n19261), .A2(n19313), .B1(n19260), .B2(n18974), .ZN(
        n18961) );
  OAI21_X1 U22113 ( .B1(n18958), .B2(n19227), .A(n19000), .ZN(n18959) );
  OAI211_X1 U22114 ( .C1(n19039), .C2(n19492), .A(n19230), .B(n18959), .ZN(
        n18975) );
  AOI22_X1 U22115 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18975), .B1(
        n19266), .B2(n18991), .ZN(n18960) );
  OAI211_X1 U22116 ( .C1(n19269), .C2(n19046), .A(n18961), .B(n18960), .ZN(
        P3_U2884) );
  AOI22_X1 U22117 ( .A1(n19271), .A2(n18991), .B1(n19270), .B2(n18974), .ZN(
        n18963) );
  AOI22_X1 U22118 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18975), .B1(
        n19272), .B2(n19313), .ZN(n18962) );
  OAI211_X1 U22119 ( .C1(n19275), .C2(n19046), .A(n18963), .B(n18962), .ZN(
        P3_U2885) );
  AOI22_X1 U22120 ( .A1(n19277), .A2(n18991), .B1(n19276), .B2(n18974), .ZN(
        n18965) );
  AOI22_X1 U22121 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18975), .B1(
        n19278), .B2(n19313), .ZN(n18964) );
  OAI211_X1 U22122 ( .C1(n19281), .C2(n19046), .A(n18965), .B(n18964), .ZN(
        P3_U2886) );
  INV_X1 U22123 ( .A(n18991), .ZN(n18998) );
  AOI22_X1 U22124 ( .A1(n19239), .A2(n19313), .B1(n19283), .B2(n18974), .ZN(
        n18967) );
  AOI22_X1 U22125 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18975), .B1(
        n19284), .B2(n19039), .ZN(n18966) );
  OAI211_X1 U22126 ( .C1(n19242), .C2(n18998), .A(n18967), .B(n18966), .ZN(
        P3_U2887) );
  AOI22_X1 U22127 ( .A1(n19289), .A2(n18991), .B1(n19288), .B2(n18974), .ZN(
        n18969) );
  AOI22_X1 U22128 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18975), .B1(
        n19290), .B2(n19313), .ZN(n18968) );
  OAI211_X1 U22129 ( .C1(n19293), .C2(n19046), .A(n18969), .B(n18968), .ZN(
        P3_U2888) );
  AOI22_X1 U22130 ( .A1(n19295), .A2(n19313), .B1(n19294), .B2(n18974), .ZN(
        n18971) );
  AOI22_X1 U22131 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18975), .B1(
        n19296), .B2(n19039), .ZN(n18970) );
  OAI211_X1 U22132 ( .C1(n19300), .C2(n18998), .A(n18971), .B(n18970), .ZN(
        P3_U2889) );
  AOI22_X1 U22133 ( .A1(n19304), .A2(n19313), .B1(n19301), .B2(n18974), .ZN(
        n18973) );
  AOI22_X1 U22134 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18975), .B1(
        n19302), .B2(n18991), .ZN(n18972) );
  OAI211_X1 U22135 ( .C1(n19308), .C2(n19046), .A(n18973), .B(n18972), .ZN(
        P3_U2890) );
  AOI22_X1 U22136 ( .A1(n19221), .A2(n19313), .B1(n19312), .B2(n18974), .ZN(
        n18977) );
  AOI22_X1 U22137 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18975), .B1(
        n19314), .B2(n19039), .ZN(n18976) );
  OAI211_X1 U22138 ( .C1(n19225), .C2(n18998), .A(n18977), .B(n18976), .ZN(
        P3_U2891) );
  NAND2_X1 U22139 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19026), .ZN(
        n19069) );
  INV_X1 U22140 ( .A(n19069), .ZN(n19062) );
  AOI21_X1 U22141 ( .B1(n19366), .B2(n19227), .A(n19001), .ZN(n19070) );
  OAI211_X1 U22142 ( .C1(n19062), .C2(n19492), .A(n18978), .B(n19070), .ZN(
        n18995) );
  AND2_X1 U22143 ( .A1(n19259), .A2(n19026), .ZN(n18994) );
  AOI22_X1 U22144 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18995), .B1(
        n19260), .B2(n18994), .ZN(n18980) );
  AOI22_X1 U22145 ( .A1(n19062), .A2(n19231), .B1(n19266), .B2(n19015), .ZN(
        n18979) );
  OAI211_X1 U22146 ( .C1(n19234), .C2(n18998), .A(n18980), .B(n18979), .ZN(
        P3_U2892) );
  AOI22_X1 U22147 ( .A1(n19270), .A2(n18994), .B1(n19272), .B2(n18991), .ZN(
        n18982) );
  AOI22_X1 U22148 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18995), .B1(
        n19271), .B2(n19015), .ZN(n18981) );
  OAI211_X1 U22149 ( .C1(n19069), .C2(n19275), .A(n18982), .B(n18981), .ZN(
        P3_U2893) );
  AOI22_X1 U22150 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18995), .B1(
        n19276), .B2(n18994), .ZN(n18984) );
  AOI22_X1 U22151 ( .A1(n19277), .A2(n19015), .B1(n19278), .B2(n18991), .ZN(
        n18983) );
  OAI211_X1 U22152 ( .C1(n19069), .C2(n19281), .A(n18984), .B(n18983), .ZN(
        P3_U2894) );
  AOI22_X1 U22153 ( .A1(n19239), .A2(n18991), .B1(n19283), .B2(n18994), .ZN(
        n18986) );
  AOI22_X1 U22154 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18995), .B1(
        n19062), .B2(n19284), .ZN(n18985) );
  OAI211_X1 U22155 ( .C1(n19242), .C2(n19023), .A(n18986), .B(n18985), .ZN(
        P3_U2895) );
  AOI22_X1 U22156 ( .A1(n19289), .A2(n19015), .B1(n19288), .B2(n18994), .ZN(
        n18988) );
  AOI22_X1 U22157 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18995), .B1(
        n19290), .B2(n18991), .ZN(n18987) );
  OAI211_X1 U22158 ( .C1(n19069), .C2(n19293), .A(n18988), .B(n18987), .ZN(
        P3_U2896) );
  AOI22_X1 U22159 ( .A1(n19295), .A2(n18991), .B1(n19294), .B2(n18994), .ZN(
        n18990) );
  AOI22_X1 U22160 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18995), .B1(
        n19062), .B2(n19296), .ZN(n18989) );
  OAI211_X1 U22161 ( .C1(n19300), .C2(n19023), .A(n18990), .B(n18989), .ZN(
        P3_U2897) );
  AOI22_X1 U22162 ( .A1(n19302), .A2(n19015), .B1(n19301), .B2(n18994), .ZN(
        n18993) );
  AOI22_X1 U22163 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18995), .B1(
        n19304), .B2(n18991), .ZN(n18992) );
  OAI211_X1 U22164 ( .C1(n19069), .C2(n19308), .A(n18993), .B(n18992), .ZN(
        P3_U2898) );
  AOI22_X1 U22165 ( .A1(n19312), .A2(n18994), .B1(n19310), .B2(n19015), .ZN(
        n18997) );
  AOI22_X1 U22166 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18995), .B1(
        n19062), .B2(n19314), .ZN(n18996) );
  OAI211_X1 U22167 ( .C1(n19319), .C2(n18998), .A(n18997), .B(n18996), .ZN(
        P3_U2899) );
  INV_X1 U22168 ( .A(n19071), .ZN(n19025) );
  INV_X1 U22169 ( .A(n9689), .ZN(n19018) );
  NOR2_X1 U22170 ( .A1(n9689), .A2(n19062), .ZN(n19048) );
  NOR2_X1 U22171 ( .A1(n19394), .A2(n19048), .ZN(n19019) );
  AOI22_X1 U22172 ( .A1(n19261), .A2(n19015), .B1(n19260), .B2(n19019), .ZN(
        n19004) );
  OAI22_X1 U22173 ( .A1(n19048), .A2(n19001), .B1(n19000), .B2(n18999), .ZN(
        n19002) );
  OAI21_X1 U22174 ( .B1(n9689), .B2(n19492), .A(n19002), .ZN(n19020) );
  AOI22_X1 U22175 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19020), .B1(
        n19266), .B2(n19039), .ZN(n19003) );
  OAI211_X1 U22176 ( .C1(n19018), .C2(n19269), .A(n19004), .B(n19003), .ZN(
        P3_U2900) );
  AOI22_X1 U22177 ( .A1(n19271), .A2(n19039), .B1(n19270), .B2(n19019), .ZN(
        n19006) );
  AOI22_X1 U22178 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19020), .B1(
        n19272), .B2(n19015), .ZN(n19005) );
  OAI211_X1 U22179 ( .C1(n19018), .C2(n19275), .A(n19006), .B(n19005), .ZN(
        P3_U2901) );
  AOI22_X1 U22180 ( .A1(n19278), .A2(n19015), .B1(n19276), .B2(n19019), .ZN(
        n19008) );
  AOI22_X1 U22181 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19020), .B1(
        n19277), .B2(n19039), .ZN(n19007) );
  OAI211_X1 U22182 ( .C1(n19018), .C2(n19281), .A(n19008), .B(n19007), .ZN(
        P3_U2902) );
  AOI22_X1 U22183 ( .A1(n19239), .A2(n19015), .B1(n19283), .B2(n19019), .ZN(
        n19010) );
  AOI22_X1 U22184 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19020), .B1(
        n9689), .B2(n19284), .ZN(n19009) );
  OAI211_X1 U22185 ( .C1(n19242), .C2(n19046), .A(n19010), .B(n19009), .ZN(
        P3_U2903) );
  AOI22_X1 U22186 ( .A1(n19289), .A2(n19039), .B1(n19288), .B2(n19019), .ZN(
        n19012) );
  AOI22_X1 U22187 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19020), .B1(
        n19290), .B2(n19015), .ZN(n19011) );
  OAI211_X1 U22188 ( .C1(n19018), .C2(n19293), .A(n19012), .B(n19011), .ZN(
        P3_U2904) );
  AOI22_X1 U22189 ( .A1(n19294), .A2(n19019), .B1(n19245), .B2(n19039), .ZN(
        n19014) );
  AOI22_X1 U22190 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19020), .B1(
        n9689), .B2(n19296), .ZN(n19013) );
  OAI211_X1 U22191 ( .C1(n19248), .C2(n19023), .A(n19014), .B(n19013), .ZN(
        P3_U2905) );
  AOI22_X1 U22192 ( .A1(n19302), .A2(n19039), .B1(n19301), .B2(n19019), .ZN(
        n19017) );
  AOI22_X1 U22193 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19020), .B1(
        n19304), .B2(n19015), .ZN(n19016) );
  OAI211_X1 U22194 ( .C1(n19018), .C2(n19308), .A(n19017), .B(n19016), .ZN(
        P3_U2906) );
  AOI22_X1 U22195 ( .A1(n19312), .A2(n19019), .B1(n19310), .B2(n19039), .ZN(
        n19022) );
  AOI22_X1 U22196 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19020), .B1(
        n9689), .B2(n19314), .ZN(n19021) );
  OAI211_X1 U22197 ( .C1(n19319), .C2(n19023), .A(n19022), .B(n19021), .ZN(
        P3_U2907) );
  NOR2_X2 U22198 ( .A1(n19024), .A2(n19025), .ZN(n19105) );
  INV_X1 U22199 ( .A(n19105), .ZN(n19112) );
  NOR2_X1 U22200 ( .A1(n19025), .A2(n19113), .ZN(n19042) );
  AOI22_X1 U22201 ( .A1(n19062), .A2(n19266), .B1(n19260), .B2(n19042), .ZN(
        n19028) );
  AOI22_X1 U22202 ( .A1(n19265), .A2(n19026), .B1(n19071), .B2(n19114), .ZN(
        n19043) );
  AOI22_X1 U22203 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19043), .B1(
        n19261), .B2(n19039), .ZN(n19027) );
  OAI211_X1 U22204 ( .C1(n19112), .C2(n19269), .A(n19028), .B(n19027), .ZN(
        P3_U2908) );
  AOI22_X1 U22205 ( .A1(n19062), .A2(n19271), .B1(n19270), .B2(n19042), .ZN(
        n19030) );
  AOI22_X1 U22206 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19043), .B1(
        n19272), .B2(n19039), .ZN(n19029) );
  OAI211_X1 U22207 ( .C1(n19112), .C2(n19275), .A(n19030), .B(n19029), .ZN(
        P3_U2909) );
  AOI22_X1 U22208 ( .A1(n19062), .A2(n19277), .B1(n19276), .B2(n19042), .ZN(
        n19032) );
  AOI22_X1 U22209 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19043), .B1(
        n19278), .B2(n19039), .ZN(n19031) );
  OAI211_X1 U22210 ( .C1(n19112), .C2(n19281), .A(n19032), .B(n19031), .ZN(
        P3_U2910) );
  AOI22_X1 U22211 ( .A1(n19239), .A2(n19039), .B1(n19283), .B2(n19042), .ZN(
        n19034) );
  AOI22_X1 U22212 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19043), .B1(
        n19105), .B2(n19284), .ZN(n19033) );
  OAI211_X1 U22213 ( .C1(n19069), .C2(n19242), .A(n19034), .B(n19033), .ZN(
        P3_U2911) );
  AOI22_X1 U22214 ( .A1(n19290), .A2(n19039), .B1(n19288), .B2(n19042), .ZN(
        n19036) );
  AOI22_X1 U22215 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19043), .B1(
        n19062), .B2(n19289), .ZN(n19035) );
  OAI211_X1 U22216 ( .C1(n19112), .C2(n19293), .A(n19036), .B(n19035), .ZN(
        P3_U2912) );
  AOI22_X1 U22217 ( .A1(n19062), .A2(n19245), .B1(n19294), .B2(n19042), .ZN(
        n19038) );
  AOI22_X1 U22218 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19043), .B1(
        n19105), .B2(n19296), .ZN(n19037) );
  OAI211_X1 U22219 ( .C1(n19248), .C2(n19046), .A(n19038), .B(n19037), .ZN(
        P3_U2913) );
  AOI22_X1 U22220 ( .A1(n19062), .A2(n19302), .B1(n19301), .B2(n19042), .ZN(
        n19041) );
  AOI22_X1 U22221 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19043), .B1(
        n19304), .B2(n19039), .ZN(n19040) );
  OAI211_X1 U22222 ( .C1(n19112), .C2(n19308), .A(n19041), .B(n19040), .ZN(
        P3_U2914) );
  AOI22_X1 U22223 ( .A1(n19062), .A2(n19310), .B1(n19312), .B2(n19042), .ZN(
        n19045) );
  AOI22_X1 U22224 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19043), .B1(
        n19105), .B2(n19314), .ZN(n19044) );
  OAI211_X1 U22225 ( .C1(n19319), .C2(n19046), .A(n19045), .B(n19044), .ZN(
        P3_U2915) );
  NOR2_X1 U22226 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19047), .ZN(
        n19115) );
  NAND2_X1 U22227 ( .A1(n19115), .A2(n19364), .ZN(n19136) );
  AOI21_X1 U22228 ( .B1(n19136), .B2(n19112), .A(n19394), .ZN(n19065) );
  AOI22_X1 U22229 ( .A1(n9689), .A2(n19266), .B1(n19260), .B2(n19065), .ZN(
        n19051) );
  INV_X1 U22230 ( .A(n19136), .ZN(n19129) );
  AOI221_X1 U22231 ( .B1(n19048), .B2(n19112), .C1(n19227), .C2(n19112), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19049) );
  OAI21_X1 U22232 ( .B1(n19129), .B2(n19049), .A(n19230), .ZN(n19066) );
  AOI22_X1 U22233 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19066), .B1(
        n19129), .B2(n19231), .ZN(n19050) );
  OAI211_X1 U22234 ( .C1(n19069), .C2(n19234), .A(n19051), .B(n19050), .ZN(
        P3_U2916) );
  AOI22_X1 U22235 ( .A1(n19062), .A2(n19272), .B1(n19065), .B2(n19270), .ZN(
        n19053) );
  AOI22_X1 U22236 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19066), .B1(
        n9689), .B2(n19271), .ZN(n19052) );
  OAI211_X1 U22237 ( .C1(n19136), .C2(n19275), .A(n19053), .B(n19052), .ZN(
        P3_U2917) );
  AOI22_X1 U22238 ( .A1(n19062), .A2(n19278), .B1(n19065), .B2(n19276), .ZN(
        n19055) );
  AOI22_X1 U22239 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19066), .B1(
        n9689), .B2(n19277), .ZN(n19054) );
  OAI211_X1 U22240 ( .C1(n19136), .C2(n19281), .A(n19055), .B(n19054), .ZN(
        P3_U2918) );
  AOI22_X1 U22241 ( .A1(n9689), .A2(n19282), .B1(n19065), .B2(n19283), .ZN(
        n19057) );
  AOI22_X1 U22242 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19066), .B1(
        n19129), .B2(n19284), .ZN(n19056) );
  OAI211_X1 U22243 ( .C1(n19069), .C2(n19287), .A(n19057), .B(n19056), .ZN(
        P3_U2919) );
  AOI22_X1 U22244 ( .A1(n19062), .A2(n19290), .B1(n19065), .B2(n19288), .ZN(
        n19059) );
  AOI22_X1 U22245 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19066), .B1(
        n9689), .B2(n19289), .ZN(n19058) );
  OAI211_X1 U22246 ( .C1(n19136), .C2(n19293), .A(n19059), .B(n19058), .ZN(
        P3_U2920) );
  AOI22_X1 U22247 ( .A1(n9689), .A2(n19245), .B1(n19065), .B2(n19294), .ZN(
        n19061) );
  AOI22_X1 U22248 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19066), .B1(
        n19129), .B2(n19296), .ZN(n19060) );
  OAI211_X1 U22249 ( .C1(n19069), .C2(n19248), .A(n19061), .B(n19060), .ZN(
        P3_U2921) );
  AOI22_X1 U22250 ( .A1(n19062), .A2(n19304), .B1(n19065), .B2(n19301), .ZN(
        n19064) );
  AOI22_X1 U22251 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19066), .B1(
        n9689), .B2(n19302), .ZN(n19063) );
  OAI211_X1 U22252 ( .C1(n19136), .C2(n19308), .A(n19064), .B(n19063), .ZN(
        P3_U2922) );
  AOI22_X1 U22253 ( .A1(n9689), .A2(n19310), .B1(n19065), .B2(n19312), .ZN(
        n19068) );
  AOI22_X1 U22254 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19066), .B1(
        n19129), .B2(n19314), .ZN(n19067) );
  OAI211_X1 U22255 ( .C1(n19069), .C2(n19319), .A(n19068), .B(n19067), .ZN(
        P3_U2923) );
  NAND2_X1 U22256 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19115), .ZN(
        n19152) );
  AND2_X1 U22257 ( .A1(n19259), .A2(n19115), .ZN(n19087) );
  AOI22_X1 U22258 ( .A1(n19105), .A2(n19266), .B1(n19260), .B2(n19087), .ZN(
        n19073) );
  INV_X1 U22259 ( .A(n19152), .ZN(n19156) );
  OAI211_X1 U22260 ( .C1(n19156), .C2(n19492), .A(n19071), .B(n19070), .ZN(
        n19088) );
  AOI22_X1 U22261 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19088), .B1(
        n9689), .B2(n19261), .ZN(n19072) );
  OAI211_X1 U22262 ( .C1(n19269), .C2(n19152), .A(n19073), .B(n19072), .ZN(
        P3_U2924) );
  AOI22_X1 U22263 ( .A1(n9689), .A2(n19272), .B1(n19270), .B2(n19087), .ZN(
        n19075) );
  AOI22_X1 U22264 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19088), .B1(
        n19105), .B2(n19271), .ZN(n19074) );
  OAI211_X1 U22265 ( .C1(n19275), .C2(n19152), .A(n19075), .B(n19074), .ZN(
        P3_U2925) );
  AOI22_X1 U22266 ( .A1(n9689), .A2(n19278), .B1(n19276), .B2(n19087), .ZN(
        n19077) );
  AOI22_X1 U22267 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19088), .B1(
        n19105), .B2(n19277), .ZN(n19076) );
  OAI211_X1 U22268 ( .C1(n19281), .C2(n19152), .A(n19077), .B(n19076), .ZN(
        P3_U2926) );
  AOI22_X1 U22269 ( .A1(n9689), .A2(n19239), .B1(n19283), .B2(n19087), .ZN(
        n19079) );
  AOI22_X1 U22270 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19088), .B1(
        n19284), .B2(n19156), .ZN(n19078) );
  OAI211_X1 U22271 ( .C1(n19112), .C2(n19242), .A(n19079), .B(n19078), .ZN(
        P3_U2927) );
  AOI22_X1 U22272 ( .A1(n19105), .A2(n19289), .B1(n19288), .B2(n19087), .ZN(
        n19081) );
  AOI22_X1 U22273 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19088), .B1(
        n9689), .B2(n19290), .ZN(n19080) );
  OAI211_X1 U22274 ( .C1(n19293), .C2(n19152), .A(n19081), .B(n19080), .ZN(
        P3_U2928) );
  AOI22_X1 U22275 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19088), .B1(
        n19294), .B2(n19087), .ZN(n19083) );
  AOI22_X1 U22276 ( .A1(n9689), .A2(n19295), .B1(n19296), .B2(n19156), .ZN(
        n19082) );
  OAI211_X1 U22277 ( .C1(n19112), .C2(n19300), .A(n19083), .B(n19082), .ZN(
        P3_U2929) );
  AOI22_X1 U22278 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19088), .B1(
        n19301), .B2(n19087), .ZN(n19086) );
  AOI22_X1 U22279 ( .A1(n19105), .A2(n19302), .B1(n9689), .B2(n19304), .ZN(
        n19085) );
  OAI211_X1 U22280 ( .C1(n19308), .C2(n19152), .A(n19086), .B(n19085), .ZN(
        P3_U2930) );
  AOI22_X1 U22281 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19088), .B1(
        n19312), .B2(n19087), .ZN(n19090) );
  AOI22_X1 U22282 ( .A1(n9689), .A2(n19221), .B1(n19314), .B2(n19156), .ZN(
        n19089) );
  OAI211_X1 U22283 ( .C1(n19112), .C2(n19225), .A(n19090), .B(n19089), .ZN(
        P3_U2931) );
  INV_X1 U22284 ( .A(n19160), .ZN(n19137) );
  NOR2_X2 U22285 ( .A1(n19367), .A2(n19137), .ZN(n19177) );
  NOR2_X1 U22286 ( .A1(n19156), .A2(n19177), .ZN(n19138) );
  NOR2_X1 U22287 ( .A1(n19394), .A2(n19138), .ZN(n19108) );
  AOI22_X1 U22288 ( .A1(n19129), .A2(n19266), .B1(n19260), .B2(n19108), .ZN(
        n19094) );
  NOR2_X1 U22289 ( .A1(n19129), .A2(n19105), .ZN(n19091) );
  OAI21_X1 U22290 ( .B1(n19091), .B2(n19227), .A(n19138), .ZN(n19092) );
  OAI211_X1 U22291 ( .C1(n19177), .C2(n19492), .A(n19230), .B(n19092), .ZN(
        n19109) );
  AOI22_X1 U22292 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19109), .B1(
        n19231), .B2(n19177), .ZN(n19093) );
  OAI211_X1 U22293 ( .C1(n19112), .C2(n19234), .A(n19094), .B(n19093), .ZN(
        P3_U2932) );
  INV_X1 U22294 ( .A(n19177), .ZN(n19173) );
  AOI22_X1 U22295 ( .A1(n19105), .A2(n19272), .B1(n19270), .B2(n19108), .ZN(
        n19096) );
  AOI22_X1 U22296 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19109), .B1(
        n19129), .B2(n19271), .ZN(n19095) );
  OAI211_X1 U22297 ( .C1(n19275), .C2(n19173), .A(n19096), .B(n19095), .ZN(
        P3_U2933) );
  AOI22_X1 U22298 ( .A1(n19129), .A2(n19277), .B1(n19276), .B2(n19108), .ZN(
        n19098) );
  AOI22_X1 U22299 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19109), .B1(
        n19105), .B2(n19278), .ZN(n19097) );
  OAI211_X1 U22300 ( .C1(n19281), .C2(n19173), .A(n19098), .B(n19097), .ZN(
        P3_U2934) );
  AOI22_X1 U22301 ( .A1(n19129), .A2(n19282), .B1(n19283), .B2(n19108), .ZN(
        n19100) );
  AOI22_X1 U22302 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19109), .B1(
        n19284), .B2(n19177), .ZN(n19099) );
  OAI211_X1 U22303 ( .C1(n19112), .C2(n19287), .A(n19100), .B(n19099), .ZN(
        P3_U2935) );
  AOI22_X1 U22304 ( .A1(n19129), .A2(n19289), .B1(n19288), .B2(n19108), .ZN(
        n19102) );
  AOI22_X1 U22305 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19109), .B1(
        n19105), .B2(n19290), .ZN(n19101) );
  OAI211_X1 U22306 ( .C1(n19293), .C2(n19173), .A(n19102), .B(n19101), .ZN(
        P3_U2936) );
  AOI22_X1 U22307 ( .A1(n19129), .A2(n19245), .B1(n19294), .B2(n19108), .ZN(
        n19104) );
  AOI22_X1 U22308 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19109), .B1(
        n19296), .B2(n19177), .ZN(n19103) );
  OAI211_X1 U22309 ( .C1(n19112), .C2(n19248), .A(n19104), .B(n19103), .ZN(
        P3_U2937) );
  AOI22_X1 U22310 ( .A1(n19105), .A2(n19304), .B1(n19301), .B2(n19108), .ZN(
        n19107) );
  AOI22_X1 U22311 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19109), .B1(
        n19129), .B2(n19302), .ZN(n19106) );
  OAI211_X1 U22312 ( .C1(n19308), .C2(n19173), .A(n19107), .B(n19106), .ZN(
        P3_U2938) );
  AOI22_X1 U22313 ( .A1(n19129), .A2(n19310), .B1(n19312), .B2(n19108), .ZN(
        n19111) );
  AOI22_X1 U22314 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19109), .B1(
        n19314), .B2(n19177), .ZN(n19110) );
  OAI211_X1 U22315 ( .C1(n19112), .C2(n19319), .A(n19111), .B(n19110), .ZN(
        P3_U2939) );
  NOR2_X1 U22316 ( .A1(n19113), .A2(n19137), .ZN(n19132) );
  AOI22_X1 U22317 ( .A1(n19260), .A2(n19132), .B1(n19266), .B2(n19156), .ZN(
        n19118) );
  AOI22_X1 U22318 ( .A1(n19265), .A2(n19115), .B1(n19114), .B2(n19160), .ZN(
        n19133) );
  NAND2_X1 U22319 ( .A1(n19116), .A2(n19160), .ZN(n19202) );
  INV_X1 U22320 ( .A(n19202), .ZN(n19195) );
  AOI22_X1 U22321 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19133), .B1(
        n19231), .B2(n19195), .ZN(n19117) );
  OAI211_X1 U22322 ( .C1(n19136), .C2(n19234), .A(n19118), .B(n19117), .ZN(
        P3_U2940) );
  AOI22_X1 U22323 ( .A1(n19129), .A2(n19272), .B1(n19270), .B2(n19132), .ZN(
        n19120) );
  AOI22_X1 U22324 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19133), .B1(
        n19271), .B2(n19156), .ZN(n19119) );
  OAI211_X1 U22325 ( .C1(n19275), .C2(n19202), .A(n19120), .B(n19119), .ZN(
        P3_U2941) );
  AOI22_X1 U22326 ( .A1(n19129), .A2(n19278), .B1(n19276), .B2(n19132), .ZN(
        n19122) );
  AOI22_X1 U22327 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19133), .B1(
        n19277), .B2(n19156), .ZN(n19121) );
  OAI211_X1 U22328 ( .C1(n19281), .C2(n19202), .A(n19122), .B(n19121), .ZN(
        P3_U2942) );
  AOI22_X1 U22329 ( .A1(n19129), .A2(n19239), .B1(n19283), .B2(n19132), .ZN(
        n19124) );
  AOI22_X1 U22330 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19133), .B1(
        n19284), .B2(n19195), .ZN(n19123) );
  OAI211_X1 U22331 ( .C1(n19242), .C2(n19152), .A(n19124), .B(n19123), .ZN(
        P3_U2943) );
  AOI22_X1 U22332 ( .A1(n19289), .A2(n19156), .B1(n19288), .B2(n19132), .ZN(
        n19126) );
  AOI22_X1 U22333 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19133), .B1(
        n19129), .B2(n19290), .ZN(n19125) );
  OAI211_X1 U22334 ( .C1(n19293), .C2(n19202), .A(n19126), .B(n19125), .ZN(
        P3_U2944) );
  AOI22_X1 U22335 ( .A1(n19294), .A2(n19132), .B1(n19245), .B2(n19156), .ZN(
        n19128) );
  AOI22_X1 U22336 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19133), .B1(
        n19296), .B2(n19195), .ZN(n19127) );
  OAI211_X1 U22337 ( .C1(n19136), .C2(n19248), .A(n19128), .B(n19127), .ZN(
        P3_U2945) );
  AOI22_X1 U22338 ( .A1(n19129), .A2(n19304), .B1(n19301), .B2(n19132), .ZN(
        n19131) );
  AOI22_X1 U22339 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19133), .B1(
        n19302), .B2(n19156), .ZN(n19130) );
  OAI211_X1 U22340 ( .C1(n19308), .C2(n19202), .A(n19131), .B(n19130), .ZN(
        P3_U2946) );
  AOI22_X1 U22341 ( .A1(n19312), .A2(n19132), .B1(n19310), .B2(n19156), .ZN(
        n19135) );
  AOI22_X1 U22342 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19133), .B1(
        n19314), .B2(n19195), .ZN(n19134) );
  OAI211_X1 U22343 ( .C1(n19136), .C2(n19319), .A(n19135), .B(n19134), .ZN(
        P3_U2947) );
  NOR2_X1 U22344 ( .A1(n19366), .A2(n19137), .ZN(n19203) );
  NAND2_X1 U22345 ( .A1(n19364), .A2(n19203), .ZN(n19216) );
  INV_X1 U22346 ( .A(n19216), .ZN(n19220) );
  NOR2_X1 U22347 ( .A1(n19195), .A2(n19220), .ZN(n19181) );
  NOR2_X1 U22348 ( .A1(n19394), .A2(n19181), .ZN(n19155) );
  AOI22_X1 U22349 ( .A1(n19260), .A2(n19155), .B1(n19266), .B2(n19177), .ZN(
        n19141) );
  OAI21_X1 U22350 ( .B1(n19138), .B2(n19227), .A(n19181), .ZN(n19139) );
  OAI211_X1 U22351 ( .C1(n19220), .C2(n19492), .A(n19230), .B(n19139), .ZN(
        n19157) );
  AOI22_X1 U22352 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19157), .B1(
        n19231), .B2(n19220), .ZN(n19140) );
  OAI211_X1 U22353 ( .C1(n19234), .C2(n19152), .A(n19141), .B(n19140), .ZN(
        P3_U2948) );
  AOI22_X1 U22354 ( .A1(n19271), .A2(n19177), .B1(n19270), .B2(n19155), .ZN(
        n19143) );
  AOI22_X1 U22355 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19157), .B1(
        n19272), .B2(n19156), .ZN(n19142) );
  OAI211_X1 U22356 ( .C1(n19275), .C2(n19216), .A(n19143), .B(n19142), .ZN(
        P3_U2949) );
  AOI22_X1 U22357 ( .A1(n19277), .A2(n19177), .B1(n19276), .B2(n19155), .ZN(
        n19145) );
  AOI22_X1 U22358 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19157), .B1(
        n19278), .B2(n19156), .ZN(n19144) );
  OAI211_X1 U22359 ( .C1(n19281), .C2(n19216), .A(n19145), .B(n19144), .ZN(
        P3_U2950) );
  AOI22_X1 U22360 ( .A1(n19239), .A2(n19156), .B1(n19283), .B2(n19155), .ZN(
        n19147) );
  AOI22_X1 U22361 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19157), .B1(
        n19284), .B2(n19220), .ZN(n19146) );
  OAI211_X1 U22362 ( .C1(n19242), .C2(n19173), .A(n19147), .B(n19146), .ZN(
        P3_U2951) );
  AOI22_X1 U22363 ( .A1(n19290), .A2(n19156), .B1(n19288), .B2(n19155), .ZN(
        n19149) );
  AOI22_X1 U22364 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19157), .B1(
        n19289), .B2(n19177), .ZN(n19148) );
  OAI211_X1 U22365 ( .C1(n19293), .C2(n19216), .A(n19149), .B(n19148), .ZN(
        P3_U2952) );
  AOI22_X1 U22366 ( .A1(n19294), .A2(n19155), .B1(n19245), .B2(n19177), .ZN(
        n19151) );
  AOI22_X1 U22367 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19157), .B1(
        n19296), .B2(n19220), .ZN(n19150) );
  OAI211_X1 U22368 ( .C1(n19248), .C2(n19152), .A(n19151), .B(n19150), .ZN(
        P3_U2953) );
  AOI22_X1 U22369 ( .A1(n19302), .A2(n19177), .B1(n19301), .B2(n19155), .ZN(
        n19154) );
  AOI22_X1 U22370 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19157), .B1(
        n19304), .B2(n19156), .ZN(n19153) );
  OAI211_X1 U22371 ( .C1(n19308), .C2(n19216), .A(n19154), .B(n19153), .ZN(
        P3_U2954) );
  AOI22_X1 U22372 ( .A1(n19221), .A2(n19156), .B1(n19312), .B2(n19155), .ZN(
        n19159) );
  AOI22_X1 U22373 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19157), .B1(
        n19314), .B2(n19220), .ZN(n19158) );
  OAI211_X1 U22374 ( .C1(n19225), .C2(n19173), .A(n19159), .B(n19158), .ZN(
        P3_U2955) );
  AND2_X1 U22375 ( .A1(n19259), .A2(n19203), .ZN(n19176) );
  AOI22_X1 U22376 ( .A1(n19260), .A2(n19176), .B1(n19266), .B2(n19195), .ZN(
        n19162) );
  AOI22_X1 U22377 ( .A1(n19265), .A2(n19160), .B1(n19262), .B2(n19203), .ZN(
        n19178) );
  NAND2_X1 U22378 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19203), .ZN(
        n19258) );
  INV_X1 U22379 ( .A(n19258), .ZN(n19249) );
  AOI22_X1 U22380 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19178), .B1(
        n19231), .B2(n19249), .ZN(n19161) );
  OAI211_X1 U22381 ( .C1(n19234), .C2(n19173), .A(n19162), .B(n19161), .ZN(
        P3_U2956) );
  AOI22_X1 U22382 ( .A1(n19270), .A2(n19176), .B1(n19272), .B2(n19177), .ZN(
        n19164) );
  AOI22_X1 U22383 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19178), .B1(
        n19271), .B2(n19195), .ZN(n19163) );
  OAI211_X1 U22384 ( .C1(n19275), .C2(n19258), .A(n19164), .B(n19163), .ZN(
        P3_U2957) );
  AOI22_X1 U22385 ( .A1(n19278), .A2(n19177), .B1(n19276), .B2(n19176), .ZN(
        n19166) );
  AOI22_X1 U22386 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19178), .B1(
        n19277), .B2(n19195), .ZN(n19165) );
  OAI211_X1 U22387 ( .C1(n19281), .C2(n19258), .A(n19166), .B(n19165), .ZN(
        P3_U2958) );
  AOI22_X1 U22388 ( .A1(n19283), .A2(n19176), .B1(n19282), .B2(n19195), .ZN(
        n19168) );
  AOI22_X1 U22389 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19178), .B1(
        n19284), .B2(n19249), .ZN(n19167) );
  OAI211_X1 U22390 ( .C1(n19287), .C2(n19173), .A(n19168), .B(n19167), .ZN(
        P3_U2959) );
  AOI22_X1 U22391 ( .A1(n19290), .A2(n19177), .B1(n19288), .B2(n19176), .ZN(
        n19170) );
  AOI22_X1 U22392 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19178), .B1(
        n19289), .B2(n19195), .ZN(n19169) );
  OAI211_X1 U22393 ( .C1(n19293), .C2(n19258), .A(n19170), .B(n19169), .ZN(
        P3_U2960) );
  AOI22_X1 U22394 ( .A1(n19294), .A2(n19176), .B1(n19245), .B2(n19195), .ZN(
        n19172) );
  AOI22_X1 U22395 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19178), .B1(
        n19296), .B2(n19249), .ZN(n19171) );
  OAI211_X1 U22396 ( .C1(n19248), .C2(n19173), .A(n19172), .B(n19171), .ZN(
        P3_U2961) );
  AOI22_X1 U22397 ( .A1(n19304), .A2(n19177), .B1(n19301), .B2(n19176), .ZN(
        n19175) );
  AOI22_X1 U22398 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19178), .B1(
        n19302), .B2(n19195), .ZN(n19174) );
  OAI211_X1 U22399 ( .C1(n19308), .C2(n19258), .A(n19175), .B(n19174), .ZN(
        P3_U2962) );
  AOI22_X1 U22400 ( .A1(n19221), .A2(n19177), .B1(n19312), .B2(n19176), .ZN(
        n19180) );
  AOI22_X1 U22401 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19178), .B1(
        n19314), .B2(n19249), .ZN(n19179) );
  OAI211_X1 U22402 ( .C1(n19225), .C2(n19202), .A(n19180), .B(n19179), .ZN(
        P3_U2963) );
  NAND2_X1 U22403 ( .A1(n19264), .A2(n19364), .ZN(n19318) );
  INV_X1 U22404 ( .A(n19318), .ZN(n19303) );
  NOR2_X1 U22405 ( .A1(n19249), .A2(n19303), .ZN(n19228) );
  NOR2_X1 U22406 ( .A1(n19394), .A2(n19228), .ZN(n19198) );
  AOI22_X1 U22407 ( .A1(n19260), .A2(n19198), .B1(n19266), .B2(n19220), .ZN(
        n19184) );
  OAI21_X1 U22408 ( .B1(n19181), .B2(n19227), .A(n19228), .ZN(n19182) );
  OAI211_X1 U22409 ( .C1(n19303), .C2(n19492), .A(n19230), .B(n19182), .ZN(
        n19199) );
  AOI22_X1 U22410 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19199), .B1(
        n19261), .B2(n19195), .ZN(n19183) );
  OAI211_X1 U22411 ( .C1(n19269), .C2(n19318), .A(n19184), .B(n19183), .ZN(
        P3_U2964) );
  AOI22_X1 U22412 ( .A1(n19270), .A2(n19198), .B1(n19272), .B2(n19195), .ZN(
        n19186) );
  AOI22_X1 U22413 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19199), .B1(
        n19271), .B2(n19220), .ZN(n19185) );
  OAI211_X1 U22414 ( .C1(n19275), .C2(n19318), .A(n19186), .B(n19185), .ZN(
        P3_U2965) );
  AOI22_X1 U22415 ( .A1(n19278), .A2(n19195), .B1(n19276), .B2(n19198), .ZN(
        n19188) );
  AOI22_X1 U22416 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19199), .B1(
        n19277), .B2(n19220), .ZN(n19187) );
  OAI211_X1 U22417 ( .C1(n19281), .C2(n19318), .A(n19188), .B(n19187), .ZN(
        P3_U2966) );
  AOI22_X1 U22418 ( .A1(n19283), .A2(n19198), .B1(n19282), .B2(n19220), .ZN(
        n19190) );
  AOI22_X1 U22419 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19199), .B1(
        n19284), .B2(n19303), .ZN(n19189) );
  OAI211_X1 U22420 ( .C1(n19287), .C2(n19202), .A(n19190), .B(n19189), .ZN(
        P3_U2967) );
  AOI22_X1 U22421 ( .A1(n19290), .A2(n19195), .B1(n19288), .B2(n19198), .ZN(
        n19192) );
  AOI22_X1 U22422 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19199), .B1(
        n19289), .B2(n19220), .ZN(n19191) );
  OAI211_X1 U22423 ( .C1(n19293), .C2(n19318), .A(n19192), .B(n19191), .ZN(
        P3_U2968) );
  AOI22_X1 U22424 ( .A1(n19295), .A2(n19195), .B1(n19294), .B2(n19198), .ZN(
        n19194) );
  AOI22_X1 U22425 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19199), .B1(
        n19296), .B2(n19303), .ZN(n19193) );
  OAI211_X1 U22426 ( .C1(n19300), .C2(n19216), .A(n19194), .B(n19193), .ZN(
        P3_U2969) );
  AOI22_X1 U22427 ( .A1(n19302), .A2(n19220), .B1(n19301), .B2(n19198), .ZN(
        n19197) );
  AOI22_X1 U22428 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19199), .B1(
        n19304), .B2(n19195), .ZN(n19196) );
  OAI211_X1 U22429 ( .C1(n19308), .C2(n19318), .A(n19197), .B(n19196), .ZN(
        P3_U2970) );
  AOI22_X1 U22430 ( .A1(n19312), .A2(n19198), .B1(n19310), .B2(n19220), .ZN(
        n19201) );
  AOI22_X1 U22431 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19199), .B1(
        n19314), .B2(n19303), .ZN(n19200) );
  OAI211_X1 U22432 ( .C1(n19319), .C2(n19202), .A(n19201), .B(n19200), .ZN(
        P3_U2971) );
  AND2_X1 U22433 ( .A1(n19259), .A2(n19264), .ZN(n19219) );
  AOI22_X1 U22434 ( .A1(n19261), .A2(n19220), .B1(n19260), .B2(n19219), .ZN(
        n19205) );
  AOI22_X1 U22435 ( .A1(n19265), .A2(n19203), .B1(n19264), .B2(n19262), .ZN(
        n19222) );
  AOI22_X1 U22436 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19222), .B1(
        n19266), .B2(n19249), .ZN(n19204) );
  OAI211_X1 U22437 ( .C1(n19269), .C2(n19299), .A(n19205), .B(n19204), .ZN(
        P3_U2972) );
  AOI22_X1 U22438 ( .A1(n19271), .A2(n19249), .B1(n19270), .B2(n19219), .ZN(
        n19207) );
  AOI22_X1 U22439 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19222), .B1(
        n19272), .B2(n19220), .ZN(n19206) );
  OAI211_X1 U22440 ( .C1(n19275), .C2(n19299), .A(n19207), .B(n19206), .ZN(
        P3_U2973) );
  AOI22_X1 U22441 ( .A1(n19278), .A2(n19220), .B1(n19276), .B2(n19219), .ZN(
        n19209) );
  AOI22_X1 U22442 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19222), .B1(
        n19277), .B2(n19249), .ZN(n19208) );
  OAI211_X1 U22443 ( .C1(n19281), .C2(n19299), .A(n19209), .B(n19208), .ZN(
        P3_U2974) );
  AOI22_X1 U22444 ( .A1(n19239), .A2(n19220), .B1(n19283), .B2(n19219), .ZN(
        n19211) );
  AOI22_X1 U22445 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19222), .B1(
        n19284), .B2(n19309), .ZN(n19210) );
  OAI211_X1 U22446 ( .C1(n19242), .C2(n19258), .A(n19211), .B(n19210), .ZN(
        P3_U2975) );
  AOI22_X1 U22447 ( .A1(n19290), .A2(n19220), .B1(n19288), .B2(n19219), .ZN(
        n19213) );
  AOI22_X1 U22448 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19222), .B1(
        n19289), .B2(n19249), .ZN(n19212) );
  OAI211_X1 U22449 ( .C1(n19293), .C2(n19299), .A(n19213), .B(n19212), .ZN(
        P3_U2976) );
  AOI22_X1 U22450 ( .A1(n19294), .A2(n19219), .B1(n19245), .B2(n19249), .ZN(
        n19215) );
  AOI22_X1 U22451 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19222), .B1(
        n19296), .B2(n19309), .ZN(n19214) );
  OAI211_X1 U22452 ( .C1(n19248), .C2(n19216), .A(n19215), .B(n19214), .ZN(
        P3_U2977) );
  AOI22_X1 U22453 ( .A1(n19302), .A2(n19249), .B1(n19301), .B2(n19219), .ZN(
        n19218) );
  AOI22_X1 U22454 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19222), .B1(
        n19304), .B2(n19220), .ZN(n19217) );
  OAI211_X1 U22455 ( .C1(n19308), .C2(n19299), .A(n19218), .B(n19217), .ZN(
        P3_U2978) );
  AOI22_X1 U22456 ( .A1(n19221), .A2(n19220), .B1(n19312), .B2(n19219), .ZN(
        n19224) );
  AOI22_X1 U22457 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19222), .B1(
        n19314), .B2(n19309), .ZN(n19223) );
  OAI211_X1 U22458 ( .C1(n19225), .C2(n19258), .A(n19224), .B(n19223), .ZN(
        P3_U2979) );
  NOR2_X1 U22459 ( .A1(n19394), .A2(n19226), .ZN(n19253) );
  AOI22_X1 U22460 ( .A1(n19260), .A2(n19253), .B1(n19266), .B2(n19303), .ZN(
        n19233) );
  OAI21_X1 U22461 ( .B1(n19228), .B2(n19227), .A(n19226), .ZN(n19229) );
  OAI211_X1 U22462 ( .C1(n19254), .C2(n19492), .A(n19230), .B(n19229), .ZN(
        n19255) );
  AOI22_X1 U22463 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19255), .B1(
        n19231), .B2(n19254), .ZN(n19232) );
  OAI211_X1 U22464 ( .C1(n19234), .C2(n19258), .A(n19233), .B(n19232), .ZN(
        P3_U2980) );
  AOI22_X1 U22465 ( .A1(n19271), .A2(n19303), .B1(n19270), .B2(n19253), .ZN(
        n19236) );
  AOI22_X1 U22466 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19255), .B1(
        n19272), .B2(n19249), .ZN(n19235) );
  OAI211_X1 U22467 ( .C1(n19275), .C2(n19252), .A(n19236), .B(n19235), .ZN(
        P3_U2981) );
  AOI22_X1 U22468 ( .A1(n19278), .A2(n19249), .B1(n19276), .B2(n19253), .ZN(
        n19238) );
  AOI22_X1 U22469 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19255), .B1(
        n19277), .B2(n19303), .ZN(n19237) );
  OAI211_X1 U22470 ( .C1(n19281), .C2(n19252), .A(n19238), .B(n19237), .ZN(
        P3_U2982) );
  AOI22_X1 U22471 ( .A1(n19239), .A2(n19249), .B1(n19283), .B2(n19253), .ZN(
        n19241) );
  AOI22_X1 U22472 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19255), .B1(
        n19284), .B2(n19254), .ZN(n19240) );
  OAI211_X1 U22473 ( .C1(n19242), .C2(n19318), .A(n19241), .B(n19240), .ZN(
        P3_U2983) );
  AOI22_X1 U22474 ( .A1(n19290), .A2(n19249), .B1(n19288), .B2(n19253), .ZN(
        n19244) );
  AOI22_X1 U22475 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19255), .B1(
        n19289), .B2(n19303), .ZN(n19243) );
  OAI211_X1 U22476 ( .C1(n19293), .C2(n19252), .A(n19244), .B(n19243), .ZN(
        P3_U2984) );
  AOI22_X1 U22477 ( .A1(n19294), .A2(n19253), .B1(n19245), .B2(n19303), .ZN(
        n19247) );
  AOI22_X1 U22478 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19255), .B1(
        n19296), .B2(n19254), .ZN(n19246) );
  OAI211_X1 U22479 ( .C1(n19248), .C2(n19258), .A(n19247), .B(n19246), .ZN(
        P3_U2985) );
  AOI22_X1 U22480 ( .A1(n19304), .A2(n19249), .B1(n19301), .B2(n19253), .ZN(
        n19251) );
  AOI22_X1 U22481 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19255), .B1(
        n19302), .B2(n19303), .ZN(n19250) );
  OAI211_X1 U22482 ( .C1(n19308), .C2(n19252), .A(n19251), .B(n19250), .ZN(
        P3_U2986) );
  AOI22_X1 U22483 ( .A1(n19312), .A2(n19253), .B1(n19310), .B2(n19303), .ZN(
        n19257) );
  AOI22_X1 U22484 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19255), .B1(
        n19314), .B2(n19254), .ZN(n19256) );
  OAI211_X1 U22485 ( .C1(n19319), .C2(n19258), .A(n19257), .B(n19256), .ZN(
        P3_U2987) );
  AND2_X1 U22486 ( .A1(n19259), .A2(n19263), .ZN(n19311) );
  AOI22_X1 U22487 ( .A1(n19261), .A2(n19303), .B1(n19260), .B2(n19311), .ZN(
        n19268) );
  AOI22_X1 U22488 ( .A1(n19265), .A2(n19264), .B1(n19263), .B2(n19262), .ZN(
        n19315) );
  AOI22_X1 U22489 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19315), .B1(
        n19266), .B2(n19309), .ZN(n19267) );
  OAI211_X1 U22490 ( .C1(n19269), .C2(n19307), .A(n19268), .B(n19267), .ZN(
        P3_U2988) );
  AOI22_X1 U22491 ( .A1(n19271), .A2(n19309), .B1(n19270), .B2(n19311), .ZN(
        n19274) );
  AOI22_X1 U22492 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19315), .B1(
        n19272), .B2(n19303), .ZN(n19273) );
  OAI211_X1 U22493 ( .C1(n19275), .C2(n19307), .A(n19274), .B(n19273), .ZN(
        P3_U2989) );
  AOI22_X1 U22494 ( .A1(n19277), .A2(n19309), .B1(n19276), .B2(n19311), .ZN(
        n19280) );
  AOI22_X1 U22495 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19315), .B1(
        n19278), .B2(n19303), .ZN(n19279) );
  OAI211_X1 U22496 ( .C1(n19281), .C2(n19307), .A(n19280), .B(n19279), .ZN(
        P3_U2990) );
  AOI22_X1 U22497 ( .A1(n19283), .A2(n19311), .B1(n19282), .B2(n19309), .ZN(
        n19286) );
  AOI22_X1 U22498 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19315), .B1(
        n19284), .B2(n19313), .ZN(n19285) );
  OAI211_X1 U22499 ( .C1(n19287), .C2(n19318), .A(n19286), .B(n19285), .ZN(
        P3_U2991) );
  AOI22_X1 U22500 ( .A1(n19289), .A2(n19309), .B1(n19288), .B2(n19311), .ZN(
        n19292) );
  AOI22_X1 U22501 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19315), .B1(
        n19290), .B2(n19303), .ZN(n19291) );
  OAI211_X1 U22502 ( .C1(n19293), .C2(n19307), .A(n19292), .B(n19291), .ZN(
        P3_U2992) );
  AOI22_X1 U22503 ( .A1(n19295), .A2(n19303), .B1(n19294), .B2(n19311), .ZN(
        n19298) );
  AOI22_X1 U22504 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19315), .B1(
        n19296), .B2(n19313), .ZN(n19297) );
  OAI211_X1 U22505 ( .C1(n19300), .C2(n19299), .A(n19298), .B(n19297), .ZN(
        P3_U2993) );
  AOI22_X1 U22506 ( .A1(n19302), .A2(n19309), .B1(n19301), .B2(n19311), .ZN(
        n19306) );
  AOI22_X1 U22507 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19315), .B1(
        n19304), .B2(n19303), .ZN(n19305) );
  OAI211_X1 U22508 ( .C1(n19308), .C2(n19307), .A(n19306), .B(n19305), .ZN(
        P3_U2994) );
  AOI22_X1 U22509 ( .A1(n19312), .A2(n19311), .B1(n19310), .B2(n19309), .ZN(
        n19317) );
  AOI22_X1 U22510 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19315), .B1(
        n19314), .B2(n19313), .ZN(n19316) );
  OAI211_X1 U22511 ( .C1(n19319), .C2(n19318), .A(n19317), .B(n19316), .ZN(
        P3_U2995) );
  NOR2_X1 U22512 ( .A1(n19334), .A2(n19320), .ZN(n19322) );
  OAI222_X1 U22513 ( .A1(n19326), .A2(n19325), .B1(n19324), .B2(n19323), .C1(
        n19322), .C2(n19321), .ZN(n19533) );
  OAI21_X1 U22514 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19327), .ZN(n19328) );
  OAI211_X1 U22515 ( .C1(n19330), .C2(n19357), .A(n19329), .B(n19328), .ZN(
        n19380) );
  NAND2_X1 U22516 ( .A1(n12306), .A2(n19355), .ZN(n19333) );
  NOR2_X1 U22517 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19331), .ZN(
        n19361) );
  INV_X1 U22518 ( .A(n19361), .ZN(n19332) );
  AOI22_X1 U22519 ( .A1(n19334), .A2(n19333), .B1(n19339), .B2(n19332), .ZN(
        n19493) );
  NOR2_X1 U22520 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19493), .ZN(
        n19342) );
  AOI21_X1 U22521 ( .B1(n19337), .B2(n19336), .A(n19335), .ZN(n19344) );
  OAI22_X1 U22522 ( .A1(n19360), .A2(n19339), .B1(n19344), .B2(n19338), .ZN(
        n19340) );
  AOI21_X1 U22523 ( .B1(n12306), .B2(n19355), .A(n19340), .ZN(n19496) );
  NAND2_X1 U22524 ( .A1(n19357), .A2(n19496), .ZN(n19341) );
  AOI22_X1 U22525 ( .A1(n19357), .A2(n19342), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19341), .ZN(n19378) );
  INV_X1 U22526 ( .A(n19357), .ZN(n19369) );
  AOI221_X1 U22527 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19344), 
        .C1(n19343), .C2(n19344), .A(n12306), .ZN(n19356) );
  NOR2_X1 U22528 ( .A1(n19345), .A2(n19522), .ZN(n19347) );
  OAI211_X1 U22529 ( .C1(n19347), .C2(n19346), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n12306), .ZN(n19352) );
  OAI211_X1 U22530 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n19350), .A(
        n19349), .B(n19348), .ZN(n19351) );
  OAI211_X1 U22531 ( .C1(n19506), .C2(n19353), .A(n19352), .B(n19351), .ZN(
        n19354) );
  AOI21_X1 U22532 ( .B1(n19356), .B2(n19355), .A(n19354), .ZN(n19502) );
  AOI22_X1 U22533 ( .A1(n19369), .A2(n12306), .B1(n19502), .B2(n19357), .ZN(
        n19373) );
  NOR2_X1 U22534 ( .A1(n19359), .A2(n19358), .ZN(n19363) );
  AOI22_X1 U22535 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19360), .B1(
        n19363), .B2(n19522), .ZN(n19517) );
  OAI22_X1 U22536 ( .A1(n19363), .A2(n19362), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19361), .ZN(n19513) );
  OR3_X1 U22537 ( .A1(n19517), .A2(n19366), .A3(n19364), .ZN(n19365) );
  AOI22_X1 U22538 ( .A1(n19517), .A2(n19366), .B1(n19513), .B2(n19365), .ZN(
        n19368) );
  OAI21_X1 U22539 ( .B1(n19369), .B2(n19368), .A(n19367), .ZN(n19372) );
  AND2_X1 U22540 ( .A1(n19373), .A2(n19372), .ZN(n19370) );
  OAI221_X1 U22541 ( .B1(n19373), .B2(n19372), .C1(n19371), .C2(n19370), .A(
        n19375), .ZN(n19377) );
  AOI21_X1 U22542 ( .B1(n19375), .B2(n19374), .A(n19373), .ZN(n19376) );
  AOI222_X1 U22543 ( .A1(n19378), .A2(n19377), .B1(n19378), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n19377), .C2(n19376), .ZN(
        n19379) );
  NOR4_X1 U22544 ( .A1(n19381), .A2(n19533), .A3(n19380), .A4(n19379), .ZN(
        n19392) );
  INV_X1 U22545 ( .A(n19382), .ZN(n19516) );
  NAND2_X1 U22546 ( .A1(n19503), .A2(n19393), .ZN(n19402) );
  INV_X1 U22547 ( .A(n19402), .ZN(n19543) );
  AOI22_X1 U22548 ( .A1(n19516), .A2(n19543), .B1(n19411), .B2(n18119), .ZN(
        n19383) );
  INV_X1 U22549 ( .A(n19383), .ZN(n19388) );
  OAI211_X1 U22550 ( .C1(n19385), .C2(n19384), .A(n19535), .B(n19392), .ZN(
        n19491) );
  OAI21_X1 U22551 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19540), .A(n19491), 
        .ZN(n19395) );
  NOR2_X1 U22552 ( .A1(n19386), .A2(n19395), .ZN(n19387) );
  MUX2_X1 U22553 ( .A(n19388), .B(n19387), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19390) );
  OAI211_X1 U22554 ( .C1(n19392), .C2(n19391), .A(n19390), .B(n19389), .ZN(
        P3_U2996) );
  NAND2_X1 U22555 ( .A1(n19411), .A2(n18119), .ZN(n19398) );
  NAND4_X1 U22556 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n19411), .A4(n19393), .ZN(n19400) );
  OR3_X1 U22557 ( .A1(n19396), .A2(n19395), .A3(n19394), .ZN(n19397) );
  NAND4_X1 U22558 ( .A1(n19399), .A2(n19398), .A3(n19400), .A4(n19397), .ZN(
        P3_U2997) );
  AND4_X1 U22559 ( .A1(n19402), .A2(n19401), .A3(n19400), .A4(n19490), .ZN(
        P3_U2998) );
  INV_X1 U22560 ( .A(n19489), .ZN(n19403) );
  AND2_X1 U22561 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19403), .ZN(
        P3_U2999) );
  INV_X1 U22562 ( .A(P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n21066) );
  NOR2_X1 U22563 ( .A1(n21066), .A2(n19489), .ZN(P3_U3000) );
  AND2_X1 U22564 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19403), .ZN(
        P3_U3001) );
  AND2_X1 U22565 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19403), .ZN(
        P3_U3002) );
  NOR2_X1 U22566 ( .A1(n21145), .A2(n19489), .ZN(P3_U3003) );
  AND2_X1 U22567 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19403), .ZN(
        P3_U3004) );
  AND2_X1 U22568 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19403), .ZN(
        P3_U3005) );
  AND2_X1 U22569 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19403), .ZN(
        P3_U3006) );
  AND2_X1 U22570 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19403), .ZN(
        P3_U3007) );
  AND2_X1 U22571 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19403), .ZN(
        P3_U3008) );
  AND2_X1 U22572 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19403), .ZN(
        P3_U3009) );
  INV_X1 U22573 ( .A(P3_DATAWIDTH_REG_20__SCAN_IN), .ZN(n21243) );
  NOR2_X1 U22574 ( .A1(n21243), .A2(n19489), .ZN(P3_U3010) );
  INV_X1 U22575 ( .A(P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21210) );
  NOR2_X1 U22576 ( .A1(n21210), .A2(n19489), .ZN(P3_U3011) );
  AND2_X1 U22577 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19403), .ZN(
        P3_U3012) );
  AND2_X1 U22578 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19403), .ZN(
        P3_U3013) );
  INV_X1 U22579 ( .A(P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(n21211) );
  NOR2_X1 U22580 ( .A1(n21211), .A2(n19489), .ZN(P3_U3014) );
  AND2_X1 U22581 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19403), .ZN(
        P3_U3015) );
  NOR2_X1 U22582 ( .A1(n21166), .A2(n19489), .ZN(P3_U3016) );
  AND2_X1 U22583 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19403), .ZN(
        P3_U3017) );
  AND2_X1 U22584 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19403), .ZN(
        P3_U3018) );
  AND2_X1 U22585 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19403), .ZN(
        P3_U3019) );
  AND2_X1 U22586 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19403), .ZN(
        P3_U3020) );
  AND2_X1 U22587 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19403), .ZN(P3_U3021) );
  AND2_X1 U22588 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19403), .ZN(P3_U3022) );
  AND2_X1 U22589 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19403), .ZN(P3_U3023) );
  AND2_X1 U22590 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19403), .ZN(P3_U3024) );
  AND2_X1 U22591 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19403), .ZN(P3_U3025) );
  AND2_X1 U22592 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19403), .ZN(P3_U3026) );
  AND2_X1 U22593 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19403), .ZN(P3_U3027) );
  AND2_X1 U22594 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19403), .ZN(P3_U3028) );
  INV_X1 U22595 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19408) );
  NOR2_X1 U22596 ( .A1(n19421), .A2(n20938), .ZN(n19417) );
  INV_X1 U22597 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19404) );
  NOR2_X1 U22598 ( .A1(n19417), .A2(n19404), .ZN(n19410) );
  OAI21_X1 U22599 ( .B1(n19408), .B2(n20938), .A(n19410), .ZN(n19405) );
  AOI22_X1 U22600 ( .A1(n19419), .A2(n19421), .B1(n19548), .B2(n19405), .ZN(
        n19406) );
  NAND3_X1 U22601 ( .A1(NA), .A2(n19419), .A3(n19408), .ZN(n19414) );
  OAI211_X1 U22602 ( .C1(n19540), .C2(n19407), .A(n19406), .B(n19414), .ZN(
        P3_U3029) );
  NOR2_X1 U22603 ( .A1(n19408), .A2(n20938), .ZN(n19409) );
  AOI22_X1 U22604 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19410), .B1(n19409), 
        .B2(n19421), .ZN(n19412) );
  NAND2_X1 U22605 ( .A1(n19411), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19415) );
  NAND3_X1 U22606 ( .A1(n19412), .A2(n19537), .A3(n19415), .ZN(P3_U3030) );
  INV_X1 U22607 ( .A(n19415), .ZN(n19413) );
  AOI21_X1 U22608 ( .B1(n19419), .B2(n19414), .A(n19413), .ZN(n19420) );
  OAI22_X1 U22609 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19415), .ZN(n19416) );
  OAI22_X1 U22610 ( .A1(n19417), .A2(n19416), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19418) );
  OAI22_X1 U22611 ( .A1(n19420), .A2(n19421), .B1(n19419), .B2(n19418), .ZN(
        P3_U3031) );
  OAI222_X1 U22612 ( .A1(n19423), .A2(n19474), .B1(n19422), .B2(n19484), .C1(
        n19424), .C2(n19471), .ZN(P3_U3032) );
  OAI222_X1 U22613 ( .A1(n19471), .A2(n19426), .B1(n19425), .B2(n19484), .C1(
        n19424), .C2(n19474), .ZN(P3_U3033) );
  OAI222_X1 U22614 ( .A1(n19471), .A2(n19428), .B1(n19427), .B2(n19484), .C1(
        n19426), .C2(n19474), .ZN(P3_U3034) );
  INV_X1 U22615 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19431) );
  OAI222_X1 U22616 ( .A1(n19471), .A2(n19431), .B1(n19429), .B2(n19484), .C1(
        n19428), .C2(n19474), .ZN(P3_U3035) );
  OAI222_X1 U22617 ( .A1(n19431), .A2(n19474), .B1(n19430), .B2(n19484), .C1(
        n19432), .C2(n19471), .ZN(P3_U3036) );
  OAI222_X1 U22618 ( .A1(n19471), .A2(n19434), .B1(n19433), .B2(n19484), .C1(
        n19432), .C2(n19474), .ZN(P3_U3037) );
  OAI222_X1 U22619 ( .A1(n19471), .A2(n21222), .B1(n19435), .B2(n19484), .C1(
        n19434), .C2(n19474), .ZN(P3_U3038) );
  OAI222_X1 U22620 ( .A1(n21222), .A2(n19474), .B1(n19436), .B2(n19484), .C1(
        n19437), .C2(n19471), .ZN(P3_U3039) );
  OAI222_X1 U22621 ( .A1(n19471), .A2(n19439), .B1(n19438), .B2(n19484), .C1(
        n19437), .C2(n19474), .ZN(P3_U3040) );
  OAI222_X1 U22622 ( .A1(n19471), .A2(n21135), .B1(n19440), .B2(n19484), .C1(
        n19439), .C2(n19474), .ZN(P3_U3041) );
  OAI222_X1 U22623 ( .A1(n19471), .A2(n19442), .B1(n19441), .B2(n19484), .C1(
        n21135), .C2(n19474), .ZN(P3_U3042) );
  OAI222_X1 U22624 ( .A1(n19471), .A2(n21324), .B1(n21149), .B2(n19484), .C1(
        n19442), .C2(n19474), .ZN(P3_U3043) );
  OAI222_X1 U22625 ( .A1(n21324), .A2(n19474), .B1(n19443), .B2(n19484), .C1(
        n19445), .C2(n19471), .ZN(P3_U3044) );
  OAI222_X1 U22626 ( .A1(n19445), .A2(n19474), .B1(n19444), .B2(n19484), .C1(
        n21323), .C2(n19471), .ZN(P3_U3045) );
  OAI222_X1 U22627 ( .A1(n21323), .A2(n19474), .B1(n19446), .B2(n19484), .C1(
        n19447), .C2(n19471), .ZN(P3_U3046) );
  OAI222_X1 U22628 ( .A1(n19471), .A2(n19450), .B1(n19448), .B2(n19484), .C1(
        n19447), .C2(n19474), .ZN(P3_U3047) );
  OAI222_X1 U22629 ( .A1(n19450), .A2(n19474), .B1(n19449), .B2(n19484), .C1(
        n19451), .C2(n19471), .ZN(P3_U3048) );
  OAI222_X1 U22630 ( .A1(n19471), .A2(n19453), .B1(n19452), .B2(n19484), .C1(
        n19451), .C2(n19480), .ZN(P3_U3049) );
  OAI222_X1 U22631 ( .A1(n19471), .A2(n19455), .B1(n19454), .B2(n19484), .C1(
        n19453), .C2(n19480), .ZN(P3_U3050) );
  INV_X1 U22632 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19457) );
  OAI222_X1 U22633 ( .A1(n19471), .A2(n19457), .B1(n19456), .B2(n19484), .C1(
        n19455), .C2(n19480), .ZN(P3_U3051) );
  OAI222_X1 U22634 ( .A1(n19471), .A2(n19459), .B1(n19458), .B2(n19484), .C1(
        n19457), .C2(n19480), .ZN(P3_U3052) );
  INV_X1 U22635 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19461) );
  OAI222_X1 U22636 ( .A1(n19471), .A2(n19461), .B1(n19460), .B2(n19484), .C1(
        n19459), .C2(n19480), .ZN(P3_U3053) );
  OAI222_X1 U22637 ( .A1(n19471), .A2(n19463), .B1(n19462), .B2(n19484), .C1(
        n19461), .C2(n19480), .ZN(P3_U3054) );
  OAI222_X1 U22638 ( .A1(n19471), .A2(n19465), .B1(n19464), .B2(n19484), .C1(
        n19463), .C2(n19480), .ZN(P3_U3055) );
  OAI222_X1 U22639 ( .A1(n19471), .A2(n19468), .B1(n19466), .B2(n19484), .C1(
        n19465), .C2(n19480), .ZN(P3_U3056) );
  OAI222_X1 U22640 ( .A1(n19468), .A2(n19474), .B1(n19467), .B2(n19484), .C1(
        n19469), .C2(n19471), .ZN(P3_U3057) );
  INV_X1 U22641 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19472) );
  OAI222_X1 U22642 ( .A1(n19471), .A2(n19472), .B1(n19470), .B2(n19484), .C1(
        n19469), .C2(n19480), .ZN(P3_U3058) );
  OAI222_X1 U22643 ( .A1(n19471), .A2(n19475), .B1(n19473), .B2(n19484), .C1(
        n19472), .C2(n19474), .ZN(P3_U3059) );
  OAI222_X1 U22644 ( .A1(n19471), .A2(n19479), .B1(n19476), .B2(n19484), .C1(
        n19475), .C2(n19474), .ZN(P3_U3060) );
  OAI222_X1 U22645 ( .A1(n19480), .A2(n19479), .B1(n19478), .B2(n19484), .C1(
        n19477), .C2(n19471), .ZN(P3_U3061) );
  OAI22_X1 U22646 ( .A1(n19548), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19484), .ZN(n19481) );
  INV_X1 U22647 ( .A(n19481), .ZN(P3_U3274) );
  OAI22_X1 U22648 ( .A1(n19548), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19484), .ZN(n19482) );
  INV_X1 U22649 ( .A(n19482), .ZN(P3_U3275) );
  INV_X1 U22650 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n21228) );
  AOI22_X1 U22651 ( .A1(n19484), .A2(n19483), .B1(n21228), .B2(n19548), .ZN(
        P3_U3276) );
  OAI22_X1 U22652 ( .A1(n19548), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19484), .ZN(n19485) );
  INV_X1 U22653 ( .A(n19485), .ZN(P3_U3277) );
  OAI21_X1 U22654 ( .B1(n19489), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19487), 
        .ZN(n19486) );
  INV_X1 U22655 ( .A(n19486), .ZN(P3_U3280) );
  OAI21_X1 U22656 ( .B1(n19489), .B2(n19488), .A(n19487), .ZN(P3_U3281) );
  OAI221_X1 U22657 ( .B1(n19492), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19492), 
        .C2(n19491), .A(n19490), .ZN(P3_U3282) );
  NOR3_X1 U22658 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19493), .A3(
        n19497), .ZN(n19494) );
  AOI21_X1 U22659 ( .B1(n19495), .B2(n19516), .A(n19494), .ZN(n19501) );
  OAI21_X1 U22660 ( .B1(n19497), .B2(n19496), .A(n19520), .ZN(n19498) );
  INV_X1 U22661 ( .A(n19498), .ZN(n19500) );
  OAI22_X1 U22662 ( .A1(n19523), .A2(n19501), .B1(n19500), .B2(n19499), .ZN(
        P3_U3285) );
  INV_X1 U22663 ( .A(n19502), .ZN(n19508) );
  NOR2_X1 U22664 ( .A1(n19503), .A2(n19519), .ZN(n19510) );
  OAI22_X1 U22665 ( .A1(n19505), .A2(n19504), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19511) );
  INV_X1 U22666 ( .A(n19511), .ZN(n19507) );
  AOI222_X1 U22667 ( .A1(n19508), .A2(n19518), .B1(n19510), .B2(n19507), .C1(
        n19516), .C2(n19506), .ZN(n19509) );
  AOI22_X1 U22668 ( .A1(n19523), .A2(n12306), .B1(n19509), .B2(n19520), .ZN(
        P3_U3288) );
  AOI222_X1 U22669 ( .A1(n19513), .A2(n19518), .B1(n19516), .B2(n19512), .C1(
        n19511), .C2(n19510), .ZN(n19514) );
  AOI22_X1 U22670 ( .A1(n19523), .A2(n19515), .B1(n19514), .B2(n19520), .ZN(
        P3_U3289) );
  AOI222_X1 U22671 ( .A1(n19519), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19518), 
        .B2(n19517), .C1(n19522), .C2(n19516), .ZN(n19521) );
  AOI22_X1 U22672 ( .A1(n19523), .A2(n19522), .B1(n19521), .B2(n19520), .ZN(
        P3_U3290) );
  AOI211_X1 U22673 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19524) );
  AOI21_X1 U22674 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19524), .ZN(n19526) );
  INV_X1 U22675 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19525) );
  AOI22_X1 U22676 ( .A1(n19530), .A2(n19526), .B1(n19525), .B2(n19527), .ZN(
        P3_U3292) );
  NOR2_X1 U22677 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n19529) );
  INV_X1 U22678 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19528) );
  AOI22_X1 U22679 ( .A1(n19530), .A2(n19529), .B1(n19528), .B2(n19527), .ZN(
        P3_U3293) );
  INV_X1 U22680 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19531) );
  AOI22_X1 U22681 ( .A1(n19484), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19531), 
        .B2(n19548), .ZN(P3_U3294) );
  MUX2_X1 U22682 ( .A(P3_MORE_REG_SCAN_IN), .B(n19533), .S(n19532), .Z(
        P3_U3295) );
  OAI21_X1 U22683 ( .B1(n19535), .B2(n19534), .A(n19551), .ZN(n19536) );
  AOI21_X1 U22684 ( .B1(n18119), .B2(n19540), .A(n19536), .ZN(n19547) );
  AOI21_X1 U22685 ( .B1(n19539), .B2(n19538), .A(n19537), .ZN(n19541) );
  OAI211_X1 U22686 ( .C1(n19542), .C2(n19541), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19540), .ZN(n19544) );
  AOI21_X1 U22687 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19544), .A(n19543), 
        .ZN(n19546) );
  NAND2_X1 U22688 ( .A1(n19547), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19545) );
  OAI21_X1 U22689 ( .B1(n19547), .B2(n19546), .A(n19545), .ZN(P3_U3296) );
  MUX2_X1 U22690 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .B(P3_M_IO_N_REG_SCAN_IN), 
        .S(n19548), .Z(P3_U3297) );
  OAI21_X1 U22691 ( .B1(n19552), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19551), 
        .ZN(n19549) );
  OAI21_X1 U22692 ( .B1(n19551), .B2(n19550), .A(n19549), .ZN(P3_U3298) );
  NOR2_X1 U22693 ( .A1(n19552), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19554)
         );
  OAI21_X1 U22694 ( .B1(n19555), .B2(n19554), .A(n19553), .ZN(P3_U3299) );
  INV_X1 U22695 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20389) );
  NAND2_X1 U22696 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20395), .ZN(n20382) );
  NAND2_X1 U22697 ( .A1(n20389), .A2(n20374), .ZN(n20378) );
  OAI21_X1 U22698 ( .B1(n20389), .B2(n20382), .A(n20378), .ZN(n20453) );
  AOI21_X1 U22699 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20453), .ZN(n19556) );
  INV_X1 U22700 ( .A(n19556), .ZN(P2_U2815) );
  INV_X1 U22701 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19559) );
  OAI22_X1 U22702 ( .A1(n19558), .A2(n20133), .B1(n19557), .B2(n19559), .ZN(
        P2_U2816) );
  OR2_X1 U22703 ( .A1(n20374), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n20505) );
  INV_X1 U22704 ( .A(n20505), .ZN(n20494) );
  AOI22_X1 U22705 ( .A1(n20494), .A2(n19559), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n20505), .ZN(n19560) );
  OAI21_X1 U22706 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n20378), .A(n19560), 
        .ZN(P2_U2817) );
  OAI21_X1 U22707 ( .B1(n20387), .B2(BS16), .A(n20453), .ZN(n20452) );
  OAI21_X1 U22708 ( .B1(n20453), .B2(n21150), .A(n20452), .ZN(P2_U2818) );
  NOR2_X1 U22709 ( .A1(n19562), .A2(n19561), .ZN(n20503) );
  OAI21_X1 U22710 ( .B1(n20503), .B2(n19564), .A(n19563), .ZN(P2_U2819) );
  NOR4_X1 U22711 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19568) );
  NOR4_X1 U22712 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19567) );
  NOR4_X1 U22713 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19566) );
  NOR4_X1 U22714 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19565) );
  NAND4_X1 U22715 ( .A1(n19568), .A2(n19567), .A3(n19566), .A4(n19565), .ZN(
        n19574) );
  NOR4_X1 U22716 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19572) );
  AOI211_X1 U22717 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19571) );
  NOR4_X1 U22718 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19570) );
  NOR4_X1 U22719 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19569) );
  NAND4_X1 U22720 ( .A1(n19572), .A2(n19571), .A3(n19570), .A4(n19569), .ZN(
        n19573) );
  NOR2_X1 U22721 ( .A1(n19574), .A2(n19573), .ZN(n19585) );
  INV_X1 U22722 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19576) );
  OAI21_X1 U22723 ( .B1(P2_REIP_REG_0__SCAN_IN), .B2(P2_REIP_REG_1__SCAN_IN), 
        .A(n19585), .ZN(n19575) );
  OAI21_X1 U22724 ( .B1(n19585), .B2(n19576), .A(n19575), .ZN(P2_U2820) );
  INV_X1 U22725 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19578) );
  NOR3_X1 U22726 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19581) );
  OAI21_X1 U22727 ( .B1(P2_REIP_REG_1__SCAN_IN), .B2(n19581), .A(n19585), .ZN(
        n19577) );
  OAI21_X1 U22728 ( .B1(n19585), .B2(n19578), .A(n19577), .ZN(P2_U2821) );
  AOI21_X1 U22729 ( .B1(P2_REIP_REG_0__SCAN_IN), .B2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19579) );
  OAI22_X1 U22730 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(n20396), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19579), .ZN(n19580) );
  INV_X1 U22731 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20448) );
  INV_X1 U22732 ( .A(n19585), .ZN(n19582) );
  AOI22_X1 U22733 ( .A1(n19585), .A2(n19580), .B1(n20448), .B2(n19582), .ZN(
        P2_U2822) );
  INV_X1 U22734 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21188) );
  AOI21_X1 U22735 ( .B1(n20396), .B2(n21188), .A(n19581), .ZN(n19584) );
  INV_X1 U22736 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19583) );
  AOI22_X1 U22737 ( .A1(n19585), .A2(n19584), .B1(n19583), .B2(n19582), .ZN(
        P2_U2823) );
  NOR2_X1 U22738 ( .A1(n19656), .A2(n19586), .ZN(n19588) );
  XOR2_X1 U22739 ( .A(n19588), .B(n19587), .Z(n19597) );
  AOI22_X1 U22740 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n19678), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19672), .ZN(n19589) );
  OAI21_X1 U22741 ( .B1(n19590), .B2(n19692), .A(n19589), .ZN(n19591) );
  AOI211_X1 U22742 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19697), .A(n19825), 
        .B(n19591), .ZN(n19596) );
  INV_X1 U22743 ( .A(n19592), .ZN(n19594) );
  AOI22_X1 U22744 ( .A1(n19594), .A2(n19698), .B1(n19593), .B2(n19671), .ZN(
        n19595) );
  OAI211_X1 U22745 ( .C1(n19704), .C2(n19597), .A(n19596), .B(n19595), .ZN(
        P2_U2837) );
  NOR2_X1 U22746 ( .A1(n19656), .A2(n19598), .ZN(n19600) );
  XOR2_X1 U22747 ( .A(n19600), .B(n19599), .Z(n19608) );
  AOI22_X1 U22748 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(n19678), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19672), .ZN(n19601) );
  OAI21_X1 U22749 ( .B1(n19602), .B2(n19692), .A(n19601), .ZN(n19603) );
  AOI211_X1 U22750 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19697), .A(n19825), 
        .B(n19603), .ZN(n19607) );
  AOI22_X1 U22751 ( .A1(n19605), .A2(n19698), .B1(n19604), .B2(n19671), .ZN(
        n19606) );
  OAI211_X1 U22752 ( .C1(n19704), .C2(n19608), .A(n19607), .B(n19606), .ZN(
        P2_U2839) );
  AOI22_X1 U22753 ( .A1(n19609), .A2(n19679), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19672), .ZN(n19610) );
  OAI211_X1 U22754 ( .C1(n20417), .C2(n19676), .A(n19610), .B(n19856), .ZN(
        n19611) );
  AOI21_X1 U22755 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n19678), .A(n19611), .ZN(
        n19617) );
  NOR2_X1 U22756 ( .A1(n19656), .A2(n19612), .ZN(n19614) );
  XNOR2_X1 U22757 ( .A(n19614), .B(n19613), .ZN(n19615) );
  AOI22_X1 U22758 ( .A1(n19724), .A2(n19671), .B1(n19684), .B2(n19615), .ZN(
        n19616) );
  OAI211_X1 U22759 ( .C1(n19618), .C2(n19687), .A(n19617), .B(n19616), .ZN(
        P2_U2841) );
  OAI21_X1 U22760 ( .B1(n20414), .B2(n19676), .A(n19838), .ZN(n19621) );
  OAI22_X1 U22761 ( .A1(n19619), .A2(n19692), .B1(n11077), .B2(n19694), .ZN(
        n19620) );
  AOI211_X1 U22762 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n19672), .A(
        n19621), .B(n19620), .ZN(n19626) );
  NOR2_X1 U22763 ( .A1(n19656), .A2(n19632), .ZN(n19623) );
  XNOR2_X1 U22764 ( .A(n19623), .B(n19622), .ZN(n19624) );
  AOI22_X1 U22765 ( .A1(n19624), .A2(n19684), .B1(n19671), .B2(n19729), .ZN(
        n19625) );
  OAI211_X1 U22766 ( .C1(n19627), .C2(n19687), .A(n19626), .B(n19625), .ZN(
        P2_U2843) );
  INV_X1 U22767 ( .A(n19634), .ZN(n19640) );
  AOI22_X1 U22768 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n19678), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19672), .ZN(n19628) );
  OAI211_X1 U22769 ( .C1(n19703), .C2(n19734), .A(n19628), .B(n19838), .ZN(
        n19631) );
  NOR2_X1 U22770 ( .A1(n19629), .A2(n19692), .ZN(n19630) );
  AOI211_X1 U22771 ( .C1(n19697), .C2(P2_REIP_REG_11__SCAN_IN), .A(n19631), 
        .B(n19630), .ZN(n19639) );
  AOI21_X1 U22772 ( .B1(n19634), .B2(n19633), .A(n19632), .ZN(n19635) );
  AOI22_X1 U22773 ( .A1(n19637), .A2(n19698), .B1(n19636), .B2(n19635), .ZN(
        n19638) );
  OAI211_X1 U22774 ( .C1(n19640), .C2(n19710), .A(n19639), .B(n19638), .ZN(
        P2_U2844) );
  INV_X1 U22775 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21194) );
  OAI22_X1 U22776 ( .A1(n19641), .A2(n19692), .B1(n19690), .B2(n21194), .ZN(
        n19642) );
  AOI211_X1 U22777 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19697), .A(n19825), 
        .B(n19642), .ZN(n19651) );
  NOR2_X1 U22778 ( .A1(n19656), .A2(n19643), .ZN(n19644) );
  XNOR2_X1 U22779 ( .A(n19645), .B(n19644), .ZN(n19649) );
  INV_X1 U22780 ( .A(n19646), .ZN(n19647) );
  OAI22_X1 U22781 ( .A1(n19736), .A2(n19703), .B1(n19647), .B2(n19687), .ZN(
        n19648) );
  AOI21_X1 U22782 ( .B1(n19649), .B2(n19684), .A(n19648), .ZN(n19650) );
  OAI211_X1 U22783 ( .C1(n19694), .C2(n10104), .A(n19651), .B(n19650), .ZN(
        P2_U2845) );
  AOI22_X1 U22784 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n19678), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19672), .ZN(n19652) );
  OAI21_X1 U22785 ( .B1(n19653), .B2(n19692), .A(n19652), .ZN(n19654) );
  AOI211_X1 U22786 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19697), .A(n19825), .B(
        n19654), .ZN(n19661) );
  NOR2_X1 U22787 ( .A1(n19656), .A2(n19655), .ZN(n19658) );
  XNOR2_X1 U22788 ( .A(n19658), .B(n19657), .ZN(n19659) );
  AOI22_X1 U22789 ( .A1(n19659), .A2(n19684), .B1(n19671), .B2(n19739), .ZN(
        n19660) );
  OAI211_X1 U22790 ( .C1(n19662), .C2(n19687), .A(n19661), .B(n19660), .ZN(
        P2_U2847) );
  NOR2_X1 U22791 ( .A1(n19656), .A2(n19663), .ZN(n19664) );
  XNOR2_X1 U22792 ( .A(n19833), .B(n19664), .ZN(n19685) );
  INV_X1 U22793 ( .A(n19665), .ZN(n19670) );
  INV_X1 U22794 ( .A(n19666), .ZN(n19667) );
  OAI21_X1 U22795 ( .B1(n11865), .B2(n19668), .A(n19667), .ZN(n19669) );
  NAND2_X1 U22796 ( .A1(n19670), .A2(n19669), .ZN(n19761) );
  NAND2_X1 U22797 ( .A1(n19671), .A2(n19759), .ZN(n19675) );
  AND2_X1 U22798 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19672), .ZN(
        n19673) );
  NOR2_X1 U22799 ( .A1(n19825), .A2(n19673), .ZN(n19674) );
  OAI211_X1 U22800 ( .C1(n19676), .C2(n20400), .A(n19675), .B(n19674), .ZN(
        n19677) );
  AOI21_X1 U22801 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n19678), .A(n19677), .ZN(
        n19682) );
  NAND2_X1 U22802 ( .A1(n19680), .A2(n19679), .ZN(n19681) );
  OAI211_X1 U22803 ( .C1(n19761), .C2(n19688), .A(n19682), .B(n19681), .ZN(
        n19683) );
  AOI21_X1 U22804 ( .B1(n19685), .B2(n19684), .A(n19683), .ZN(n19686) );
  OAI21_X1 U22805 ( .B1(n19687), .B2(n19826), .A(n19686), .ZN(P2_U2851) );
  INV_X1 U22806 ( .A(n19688), .ZN(n19708) );
  OAI22_X1 U22807 ( .A1(n19692), .A2(n19691), .B1(n19690), .B2(n19689), .ZN(
        n19696) );
  NOR2_X1 U22808 ( .A1(n19694), .A2(n19693), .ZN(n19695) );
  AOI211_X1 U22809 ( .C1(n19697), .C2(P2_REIP_REG_1__SCAN_IN), .A(n19696), .B(
        n19695), .ZN(n19701) );
  NAND2_X1 U22810 ( .A1(n9706), .A2(n19698), .ZN(n19700) );
  OAI211_X1 U22811 ( .C1(n19703), .C2(n19702), .A(n19701), .B(n19700), .ZN(
        n19707) );
  NOR2_X1 U22812 ( .A1(n19705), .A2(n19704), .ZN(n19706) );
  AOI211_X1 U22813 ( .C1(n19708), .C2(n20478), .A(n19707), .B(n19706), .ZN(
        n19709) );
  OAI21_X1 U22814 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19710), .A(
        n19709), .ZN(P2_U2854) );
  INV_X1 U22815 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19711) );
  OAI22_X1 U22816 ( .A1(n19761), .A2(n19713), .B1(n19712), .B2(n19711), .ZN(
        n19714) );
  INV_X1 U22817 ( .A(n19714), .ZN(n19715) );
  OAI21_X1 U22818 ( .B1(n19716), .B2(n19826), .A(n19715), .ZN(P2_U2883) );
  AOI22_X1 U22819 ( .A1(n19718), .A2(n19772), .B1(n19717), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19721) );
  AOI22_X1 U22820 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19771), .B1(n19719), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19720) );
  NAND2_X1 U22821 ( .A1(n19721), .A2(n19720), .ZN(P2_U2888) );
  OAI222_X1 U22822 ( .A1(n19723), .A2(n19758), .B1(n19787), .B2(n19744), .C1(
        n19722), .C2(n19779), .ZN(P2_U2904) );
  INV_X1 U22823 ( .A(n19724), .ZN(n19726) );
  AOI22_X1 U22824 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19771), .B1(n19818), 
        .B2(n19746), .ZN(n19725) );
  OAI21_X1 U22825 ( .B1(n19758), .B2(n19726), .A(n19725), .ZN(P2_U2905) );
  INV_X1 U22826 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19792) );
  OAI222_X1 U22827 ( .A1(n19728), .A2(n19758), .B1(n19792), .B2(n19744), .C1(
        n19779), .C2(n19727), .ZN(P2_U2906) );
  INV_X1 U22828 ( .A(n19729), .ZN(n19732) );
  AOI22_X1 U22829 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19771), .B1(n19730), 
        .B2(n19746), .ZN(n19731) );
  OAI21_X1 U22830 ( .B1(n19758), .B2(n19732), .A(n19731), .ZN(P2_U2907) );
  OAI222_X1 U22831 ( .A1(n19734), .A2(n19758), .B1(n12657), .B2(n19744), .C1(
        n19779), .C2(n19733), .ZN(P2_U2908) );
  OAI222_X1 U22832 ( .A1(n19736), .A2(n19758), .B1(n12633), .B2(n19744), .C1(
        n19779), .C2(n19735), .ZN(P2_U2909) );
  INV_X1 U22833 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19799) );
  OAI222_X1 U22834 ( .A1(n19738), .A2(n19758), .B1(n19799), .B2(n19744), .C1(
        n19779), .C2(n19737), .ZN(P2_U2910) );
  INV_X1 U22835 ( .A(n19739), .ZN(n19742) );
  AOI22_X1 U22836 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19771), .B1(n19740), .B2(
        n19746), .ZN(n19741) );
  OAI21_X1 U22837 ( .B1(n19758), .B2(n19742), .A(n19741), .ZN(P2_U2911) );
  OAI222_X1 U22838 ( .A1(n19743), .A2(n19758), .B1(n12665), .B2(n19744), .C1(
        n19779), .C2(n19908), .ZN(P2_U2912) );
  INV_X1 U22839 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19804) );
  OAI222_X1 U22840 ( .A1(n19745), .A2(n19758), .B1(n19804), .B2(n19744), .C1(
        n19779), .C2(n19897), .ZN(P2_U2913) );
  AOI22_X1 U22841 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19771), .B1(n19747), .B2(
        n19746), .ZN(n19756) );
  NAND2_X1 U22842 ( .A1(n19749), .A2(n19748), .ZN(n19753) );
  XNOR2_X1 U22843 ( .A(n19749), .B(n20459), .ZN(n19767) );
  NAND2_X1 U22844 ( .A1(n19750), .A2(n20466), .ZN(n19752) );
  NAND2_X1 U22845 ( .A1(n19752), .A2(n19751), .ZN(n19766) );
  NAND2_X1 U22846 ( .A1(n19767), .A2(n19766), .ZN(n19765) );
  AOI21_X1 U22847 ( .B1(n19753), .B2(n19765), .A(n19759), .ZN(n19760) );
  OR3_X1 U22848 ( .A1(n19760), .A2(n19761), .A3(n19754), .ZN(n19755) );
  OAI211_X1 U22849 ( .C1(n19758), .C2(n19757), .A(n19756), .B(n19755), .ZN(
        P2_U2914) );
  AOI22_X1 U22850 ( .A1(n19772), .A2(n19759), .B1(n19771), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19764) );
  XOR2_X1 U22851 ( .A(n19761), .B(n19760), .Z(n19762) );
  NAND2_X1 U22852 ( .A1(n19762), .A2(n19773), .ZN(n19763) );
  OAI211_X1 U22853 ( .C1(n19891), .C2(n19779), .A(n19764), .B(n19763), .ZN(
        P2_U2915) );
  OAI21_X1 U22854 ( .B1(n19767), .B2(n19766), .A(n19765), .ZN(n19768) );
  NAND2_X1 U22855 ( .A1(n19768), .A2(n19773), .ZN(n19770) );
  AOI22_X1 U22856 ( .A1(n20459), .A2(n19772), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19771), .ZN(n19769) );
  OAI211_X1 U22857 ( .C1(n19886), .C2(n19779), .A(n19770), .B(n19769), .ZN(
        P2_U2916) );
  AOI22_X1 U22858 ( .A1(n19772), .A2(n19775), .B1(n19771), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19778) );
  OAI211_X1 U22859 ( .C1(n19776), .C2(n19775), .A(n19774), .B(n19773), .ZN(
        n19777) );
  OAI211_X1 U22860 ( .C1(n19780), .C2(n19779), .A(n19778), .B(n19777), .ZN(
        P2_U2919) );
  NOR2_X1 U22861 ( .A1(n19791), .A2(n19781), .ZN(P2_U2920) );
  INV_X1 U22862 ( .A(n19782), .ZN(n19783) );
  AOI22_X1 U22863 ( .A1(n19783), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n19814), .ZN(n19784) );
  OAI21_X1 U22864 ( .B1(n19791), .B2(n19785), .A(n19784), .ZN(P2_U2921) );
  OAI222_X1 U22865 ( .A1(n19791), .A2(n21246), .B1(n19816), .B2(n19787), .C1(
        n19793), .C2(n19786), .ZN(P2_U2936) );
  INV_X1 U22866 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19789) );
  AOI22_X1 U22867 ( .A1(n19814), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19788) );
  OAI21_X1 U22868 ( .B1(n19789), .B2(n19816), .A(n19788), .ZN(P2_U2937) );
  OAI222_X1 U22869 ( .A1(n19793), .A2(n12705), .B1(n19816), .B2(n19792), .C1(
        n19791), .C2(n19790), .ZN(P2_U2938) );
  AOI22_X1 U22870 ( .A1(n19814), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19794) );
  OAI21_X1 U22871 ( .B1(n19795), .B2(n19816), .A(n19794), .ZN(P2_U2939) );
  AOI22_X1 U22872 ( .A1(n19814), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19796) );
  OAI21_X1 U22873 ( .B1(n12657), .B2(n19816), .A(n19796), .ZN(P2_U2940) );
  AOI22_X1 U22874 ( .A1(n19814), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19797) );
  OAI21_X1 U22875 ( .B1(n12633), .B2(n19816), .A(n19797), .ZN(P2_U2941) );
  AOI22_X1 U22876 ( .A1(n19814), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19798) );
  OAI21_X1 U22877 ( .B1(n19799), .B2(n19816), .A(n19798), .ZN(P2_U2942) );
  AOI22_X1 U22878 ( .A1(n19814), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19800) );
  OAI21_X1 U22879 ( .B1(n19801), .B2(n19816), .A(n19800), .ZN(P2_U2943) );
  AOI22_X1 U22880 ( .A1(n19814), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19802) );
  OAI21_X1 U22881 ( .B1(n12665), .B2(n19816), .A(n19802), .ZN(P2_U2944) );
  AOI22_X1 U22882 ( .A1(n19814), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19803) );
  OAI21_X1 U22883 ( .B1(n19804), .B2(n19816), .A(n19803), .ZN(P2_U2945) );
  INV_X1 U22884 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19806) );
  AOI22_X1 U22885 ( .A1(n19814), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19805) );
  OAI21_X1 U22886 ( .B1(n19806), .B2(n19816), .A(n19805), .ZN(P2_U2946) );
  AOI22_X1 U22887 ( .A1(n19814), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19807) );
  OAI21_X1 U22888 ( .B1(n12649), .B2(n19816), .A(n19807), .ZN(P2_U2947) );
  AOI22_X1 U22889 ( .A1(n19814), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19808) );
  OAI21_X1 U22890 ( .B1(n12636), .B2(n19816), .A(n19808), .ZN(P2_U2948) );
  INV_X1 U22891 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19810) );
  AOI22_X1 U22892 ( .A1(n19814), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19809) );
  OAI21_X1 U22893 ( .B1(n19810), .B2(n19816), .A(n19809), .ZN(P2_U2949) );
  INV_X1 U22894 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19812) );
  AOI22_X1 U22895 ( .A1(n19814), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19811) );
  OAI21_X1 U22896 ( .B1(n19812), .B2(n19816), .A(n19811), .ZN(P2_U2950) );
  AOI22_X1 U22897 ( .A1(n19814), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19813), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19815) );
  OAI21_X1 U22898 ( .B1(n19817), .B2(n19816), .A(n19815), .ZN(P2_U2951) );
  AOI22_X1 U22899 ( .A1(n19822), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19821), .ZN(n19820) );
  NAND2_X1 U22900 ( .A1(n19819), .A2(n19818), .ZN(n19823) );
  NAND2_X1 U22901 ( .A1(n19820), .A2(n19823), .ZN(P2_U2966) );
  AOI22_X1 U22902 ( .A1(n19822), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19821), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n19824) );
  NAND2_X1 U22903 ( .A1(n19824), .A2(n19823), .ZN(P2_U2981) );
  AOI22_X1 U22904 ( .A1(n19837), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19825), .ZN(n19832) );
  INV_X1 U22905 ( .A(n19826), .ZN(n19829) );
  AOI222_X1 U22906 ( .A1(n19830), .A2(n11531), .B1(n19848), .B2(n19829), .C1(
        n19828), .C2(n19827), .ZN(n19831) );
  OAI211_X1 U22907 ( .C1(n19840), .C2(n19833), .A(n19832), .B(n19831), .ZN(
        P2_U3010) );
  AOI21_X1 U22908 ( .B1(n19836), .B2(n19835), .A(n19834), .ZN(n19855) );
  AOI22_X1 U22909 ( .A1(n19855), .A2(n11531), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19837), .ZN(n19850) );
  OAI22_X1 U22910 ( .A1(n19840), .A2(n19839), .B1(n19857), .B2(n19838), .ZN(
        n19847) );
  NAND2_X1 U22911 ( .A1(n19842), .A2(n19841), .ZN(n19843) );
  NAND2_X1 U22912 ( .A1(n19844), .A2(n19843), .ZN(n19864) );
  NOR2_X1 U22913 ( .A1(n19864), .A2(n19845), .ZN(n19846) );
  AOI211_X1 U22914 ( .C1(n19848), .C2(n10541), .A(n19847), .B(n19846), .ZN(
        n19849) );
  NAND2_X1 U22915 ( .A1(n19850), .A2(n19849), .ZN(P2_U3012) );
  AOI221_X1 U22916 ( .B1(n19853), .B2(n19862), .C1(n19863), .C2(n19852), .A(
        n19851), .ZN(n19877) );
  NAND2_X1 U22917 ( .A1(n20468), .A2(n19854), .ZN(n19874) );
  INV_X1 U22918 ( .A(n19855), .ZN(n19858) );
  OAI22_X1 U22919 ( .A1(n19859), .A2(n19858), .B1(n19857), .B2(n19856), .ZN(
        n19860) );
  NOR2_X1 U22920 ( .A1(n19861), .A2(n19860), .ZN(n19873) );
  NAND3_X1 U22921 ( .A1(n19863), .A2(n19862), .A3(n19876), .ZN(n19868) );
  INV_X1 U22922 ( .A(n19864), .ZN(n19865) );
  NAND2_X1 U22923 ( .A1(n19866), .A2(n19865), .ZN(n19867) );
  AND2_X1 U22924 ( .A1(n19868), .A2(n19867), .ZN(n19872) );
  OR2_X1 U22925 ( .A1(n19870), .A2(n19869), .ZN(n19871) );
  AND4_X1 U22926 ( .A1(n19874), .A2(n19873), .A3(n19872), .A4(n19871), .ZN(
        n19875) );
  OAI21_X1 U22927 ( .B1(n19877), .B2(n19876), .A(n19875), .ZN(P2_U3044) );
  AOI22_X1 U22928 ( .A1(n19907), .A2(n20322), .B1(n20314), .B2(n19906), .ZN(
        n19879) );
  AOI22_X1 U22929 ( .A1(n13231), .A2(n19911), .B1(n19937), .B2(n20173), .ZN(
        n19878) );
  OAI211_X1 U22930 ( .C1(n19914), .C2(n11767), .A(n19879), .B(n19878), .ZN(
        P2_U3048) );
  AOI22_X1 U22931 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19909), .ZN(n20182) );
  AND2_X1 U22932 ( .A1(n19880), .A2(n19904), .ZN(n20331) );
  AOI22_X1 U22933 ( .A1(n19907), .A2(n20333), .B1(n19906), .B2(n20331), .ZN(
        n19883) );
  NOR2_X2 U22934 ( .A1(n19881), .A2(n20074), .ZN(n20332) );
  AOI22_X1 U22935 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19909), .ZN(n20336) );
  AOI22_X1 U22936 ( .A1(n20332), .A2(n19911), .B1(n19937), .B2(n20288), .ZN(
        n19882) );
  OAI211_X1 U22937 ( .C1(n19914), .C2(n19884), .A(n19883), .B(n19882), .ZN(
        P2_U3050) );
  NOR2_X2 U22938 ( .A1(n10470), .A2(n19890), .ZN(n20337) );
  AOI22_X1 U22939 ( .A1(n20339), .A2(n19907), .B1(n19906), .B2(n20337), .ZN(
        n19888) );
  NOR2_X2 U22940 ( .A1(n19886), .A2(n20074), .ZN(n20338) );
  AOI22_X1 U22941 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19909), .ZN(n20342) );
  AOI22_X1 U22942 ( .A1(n20338), .A2(n19911), .B1(n19937), .B2(n20291), .ZN(
        n19887) );
  OAI211_X1 U22943 ( .C1(n19914), .C2(n11842), .A(n19888), .B(n19887), .ZN(
        P2_U3051) );
  OAI22_X1 U22944 ( .A1(n19889), .A2(n19902), .B1(n21208), .B2(n19900), .ZN(
        n20345) );
  AOI22_X1 U22945 ( .A1(n20345), .A2(n19907), .B1(n19906), .B2(n20343), .ZN(
        n19893) );
  NOR2_X2 U22946 ( .A1(n19891), .A2(n20074), .ZN(n20344) );
  AOI22_X1 U22947 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19909), .ZN(n20348) );
  AOI22_X1 U22948 ( .A1(n20344), .A2(n19911), .B1(n19937), .B2(n20294), .ZN(
        n19892) );
  OAI211_X1 U22949 ( .C1(n19914), .C2(n11865), .A(n19893), .B(n19892), .ZN(
        P2_U3052) );
  OAI22_X2 U22950 ( .A1(n19895), .A2(n19902), .B1(n19894), .B2(n19900), .ZN(
        n20357) );
  AND2_X1 U22951 ( .A1(n19896), .A2(n19904), .ZN(n20355) );
  AOI22_X1 U22952 ( .A1(n20357), .A2(n19907), .B1(n19906), .B2(n20355), .ZN(
        n19899) );
  NOR2_X2 U22953 ( .A1(n19897), .A2(n20074), .ZN(n20356) );
  AOI22_X1 U22954 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19909), .ZN(n20360) );
  INV_X1 U22955 ( .A(n20360), .ZN(n20300) );
  AOI22_X1 U22956 ( .A1(n20356), .A2(n19911), .B1(n19937), .B2(n20300), .ZN(
        n19898) );
  OAI211_X1 U22957 ( .C1(n19914), .C2(n13317), .A(n19899), .B(n19898), .ZN(
        P2_U3054) );
  OAI22_X1 U22958 ( .A1(n19903), .A2(n19902), .B1(n19901), .B2(n19900), .ZN(
        n20365) );
  AND2_X1 U22959 ( .A1(n19905), .A2(n19904), .ZN(n20362) );
  AOI22_X1 U22960 ( .A1(n20365), .A2(n19907), .B1(n19906), .B2(n20362), .ZN(
        n19913) );
  NOR2_X2 U22961 ( .A1(n19908), .A2(n20074), .ZN(n20363) );
  AOI22_X1 U22962 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19910), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19909), .ZN(n20371) );
  AOI22_X1 U22963 ( .A1(n20363), .A2(n19911), .B1(n19937), .B2(n20304), .ZN(
        n19912) );
  OAI211_X1 U22964 ( .C1(n19914), .C2(n21174), .A(n19913), .B(n19912), .ZN(
        P2_U3055) );
  INV_X1 U22965 ( .A(n10778), .ZN(n19915) );
  NOR2_X1 U22966 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20492), .ZN(
        n20131) );
  AND2_X1 U22967 ( .A1(n20131), .A2(n19941), .ZN(n19935) );
  OAI21_X1 U22968 ( .B1(n19915), .B2(n19935), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19916) );
  OAI21_X1 U22969 ( .B1(n19917), .B2(n20133), .A(n19916), .ZN(n19936) );
  AOI22_X1 U22970 ( .A1(n19936), .A2(n13231), .B1(n20314), .B2(n19935), .ZN(
        n19922) );
  OAI21_X1 U22971 ( .B1(n20072), .B2(n20132), .A(n19917), .ZN(n19920) );
  INV_X1 U22972 ( .A(n19935), .ZN(n19918) );
  OAI211_X1 U22973 ( .C1(n10778), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19918), 
        .B(n20133), .ZN(n19919) );
  NAND3_X1 U22974 ( .A1(n19920), .A2(n20320), .A3(n19919), .ZN(n19938) );
  AOI22_X1 U22975 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19938), .B1(
        n19937), .B2(n20322), .ZN(n19921) );
  OAI211_X1 U22976 ( .C1(n20325), .C2(n19968), .A(n19922), .B(n19921), .ZN(
        P2_U3056) );
  AOI22_X1 U22977 ( .A1(n19936), .A2(n14253), .B1(n20326), .B2(n19935), .ZN(
        n19924) );
  AOI22_X1 U22978 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19938), .B1(
        n19937), .B2(n20327), .ZN(n19923) );
  OAI211_X1 U22979 ( .C1(n20330), .C2(n19968), .A(n19924), .B(n19923), .ZN(
        P2_U3057) );
  AOI22_X1 U22980 ( .A1(n19936), .A2(n20332), .B1(n20331), .B2(n19935), .ZN(
        n19926) );
  AOI22_X1 U22981 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19938), .B1(
        n19937), .B2(n20333), .ZN(n19925) );
  OAI211_X1 U22982 ( .C1(n20336), .C2(n19968), .A(n19926), .B(n19925), .ZN(
        P2_U3058) );
  AOI22_X1 U22983 ( .A1(n19936), .A2(n20338), .B1(n20337), .B2(n19935), .ZN(
        n19928) );
  AOI22_X1 U22984 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19938), .B1(
        n19937), .B2(n20339), .ZN(n19927) );
  OAI211_X1 U22985 ( .C1(n20342), .C2(n19968), .A(n19928), .B(n19927), .ZN(
        P2_U3059) );
  AOI22_X1 U22986 ( .A1(n19936), .A2(n20344), .B1(n20343), .B2(n19935), .ZN(
        n19930) );
  AOI22_X1 U22987 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19938), .B1(
        n19937), .B2(n20345), .ZN(n19929) );
  OAI211_X1 U22988 ( .C1(n20348), .C2(n19968), .A(n19930), .B(n19929), .ZN(
        P2_U3060) );
  AOI22_X1 U22989 ( .A1(n19936), .A2(n20350), .B1(n20349), .B2(n19935), .ZN(
        n19932) );
  AOI22_X1 U22990 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19938), .B1(
        n19937), .B2(n20351), .ZN(n19931) );
  OAI211_X1 U22991 ( .C1(n20354), .C2(n19968), .A(n19932), .B(n19931), .ZN(
        P2_U3061) );
  AOI22_X1 U22992 ( .A1(n19936), .A2(n20356), .B1(n20355), .B2(n19935), .ZN(
        n19934) );
  AOI22_X1 U22993 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19938), .B1(
        n19937), .B2(n20357), .ZN(n19933) );
  OAI211_X1 U22994 ( .C1(n20360), .C2(n19968), .A(n19934), .B(n19933), .ZN(
        P2_U3062) );
  AOI22_X1 U22995 ( .A1(n19936), .A2(n20363), .B1(n20362), .B2(n19935), .ZN(
        n19940) );
  AOI22_X1 U22996 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19938), .B1(
        n19937), .B2(n20365), .ZN(n19939) );
  OAI211_X1 U22997 ( .C1(n20371), .C2(n19968), .A(n19940), .B(n19939), .ZN(
        P2_U3063) );
  NOR2_X1 U22998 ( .A1(n20481), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20163) );
  NAND2_X1 U22999 ( .A1(n20163), .A2(n19941), .ZN(n19945) );
  AND2_X1 U23000 ( .A1(n10760), .A2(n19945), .ZN(n19943) );
  NAND3_X1 U23001 ( .A1(n20458), .A2(n19942), .A3(n19941), .ZN(n19944) );
  OAI21_X1 U23002 ( .B1(n19943), .B2(n20312), .A(n19944), .ZN(n19964) );
  INV_X1 U23003 ( .A(n19945), .ZN(n19963) );
  AOI22_X1 U23004 ( .A1(n19964), .A2(n13231), .B1(n20314), .B2(n19963), .ZN(
        n19950) );
  OAI221_X1 U23005 ( .B1(n21150), .B2(n19989), .C1(n21150), .C2(n19968), .A(
        n19944), .ZN(n19947) );
  OAI21_X1 U23006 ( .B1(n10760), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19945), 
        .ZN(n19946) );
  MUX2_X1 U23007 ( .A(n19947), .B(n19946), .S(n20133), .Z(n19948) );
  NAND2_X1 U23008 ( .A1(n19948), .A2(n20320), .ZN(n19965) );
  AOI22_X1 U23009 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19965), .B1(
        n19981), .B2(n20173), .ZN(n19949) );
  OAI211_X1 U23010 ( .C1(n20176), .C2(n19968), .A(n19950), .B(n19949), .ZN(
        P2_U3064) );
  AOI22_X1 U23011 ( .A1(n19964), .A2(n14253), .B1(n20326), .B2(n19963), .ZN(
        n19952) );
  AOI22_X1 U23012 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19965), .B1(
        n19981), .B2(n20285), .ZN(n19951) );
  OAI211_X1 U23013 ( .C1(n20179), .C2(n19968), .A(n19952), .B(n19951), .ZN(
        P2_U3065) );
  AOI22_X1 U23014 ( .A1(n19964), .A2(n20332), .B1(n20331), .B2(n19963), .ZN(
        n19954) );
  AOI22_X1 U23015 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19965), .B1(
        n19981), .B2(n20288), .ZN(n19953) );
  OAI211_X1 U23016 ( .C1(n20182), .C2(n19968), .A(n19954), .B(n19953), .ZN(
        P2_U3066) );
  AOI22_X1 U23017 ( .A1(n19964), .A2(n20338), .B1(n20337), .B2(n19963), .ZN(
        n19956) );
  AOI22_X1 U23018 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19965), .B1(
        n19981), .B2(n20291), .ZN(n19955) );
  OAI211_X1 U23019 ( .C1(n20185), .C2(n19968), .A(n19956), .B(n19955), .ZN(
        P2_U3067) );
  INV_X1 U23020 ( .A(n20345), .ZN(n20188) );
  AOI22_X1 U23021 ( .A1(n19964), .A2(n20344), .B1(n20343), .B2(n19963), .ZN(
        n19958) );
  AOI22_X1 U23022 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19965), .B1(
        n19981), .B2(n20294), .ZN(n19957) );
  OAI211_X1 U23023 ( .C1(n20188), .C2(n19968), .A(n19958), .B(n19957), .ZN(
        P2_U3068) );
  AOI22_X1 U23024 ( .A1(n19964), .A2(n20350), .B1(n20349), .B2(n19963), .ZN(
        n19960) );
  AOI22_X1 U23025 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19965), .B1(
        n19981), .B2(n20297), .ZN(n19959) );
  OAI211_X1 U23026 ( .C1(n20191), .C2(n19968), .A(n19960), .B(n19959), .ZN(
        P2_U3069) );
  INV_X1 U23027 ( .A(n20357), .ZN(n20194) );
  AOI22_X1 U23028 ( .A1(n19964), .A2(n20356), .B1(n20355), .B2(n19963), .ZN(
        n19962) );
  AOI22_X1 U23029 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19965), .B1(
        n19981), .B2(n20300), .ZN(n19961) );
  OAI211_X1 U23030 ( .C1(n20194), .C2(n19968), .A(n19962), .B(n19961), .ZN(
        P2_U3070) );
  INV_X1 U23031 ( .A(n20365), .ZN(n20201) );
  AOI22_X1 U23032 ( .A1(n19964), .A2(n20363), .B1(n20362), .B2(n19963), .ZN(
        n19967) );
  AOI22_X1 U23033 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19965), .B1(
        n19981), .B2(n20304), .ZN(n19966) );
  OAI211_X1 U23034 ( .C1(n20201), .C2(n19968), .A(n19967), .B(n19966), .ZN(
        P2_U3071) );
  AOI22_X1 U23035 ( .A1(n20327), .A2(n19981), .B1(n20326), .B2(n19984), .ZN(
        n19970) );
  AOI22_X1 U23036 ( .A1(n14253), .A2(n19985), .B1(n20011), .B2(n20285), .ZN(
        n19969) );
  OAI211_X1 U23037 ( .C1(n19974), .C2(n10608), .A(n19970), .B(n19969), .ZN(
        P2_U3073) );
  INV_X1 U23038 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n19973) );
  AOI22_X1 U23039 ( .A1(n19981), .A2(n20333), .B1(n19984), .B2(n20331), .ZN(
        n19972) );
  AOI22_X1 U23040 ( .A1(n20332), .A2(n19985), .B1(n20011), .B2(n20288), .ZN(
        n19971) );
  OAI211_X1 U23041 ( .C1(n19974), .C2(n19973), .A(n19972), .B(n19971), .ZN(
        P2_U3074) );
  AOI22_X1 U23042 ( .A1(n20291), .A2(n20011), .B1(n19984), .B2(n20337), .ZN(
        n19976) );
  AOI22_X1 U23043 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19986), .B1(
        n20338), .B2(n19985), .ZN(n19975) );
  OAI211_X1 U23044 ( .C1(n20185), .C2(n19989), .A(n19976), .B(n19975), .ZN(
        P2_U3075) );
  AOI22_X1 U23045 ( .A1(n20294), .A2(n20011), .B1(n19984), .B2(n20343), .ZN(
        n19978) );
  AOI22_X1 U23046 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19986), .B1(
        n20344), .B2(n19985), .ZN(n19977) );
  OAI211_X1 U23047 ( .C1(n20188), .C2(n19989), .A(n19978), .B(n19977), .ZN(
        P2_U3076) );
  AOI22_X1 U23048 ( .A1(n19981), .A2(n20351), .B1(n20349), .B2(n19984), .ZN(
        n19980) );
  AOI22_X1 U23049 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19986), .B1(
        n20350), .B2(n19985), .ZN(n19979) );
  OAI211_X1 U23050 ( .C1(n20354), .C2(n20019), .A(n19980), .B(n19979), .ZN(
        P2_U3077) );
  AOI22_X1 U23051 ( .A1(n20357), .A2(n19981), .B1(n19984), .B2(n20355), .ZN(
        n19983) );
  AOI22_X1 U23052 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19986), .B1(
        n20356), .B2(n19985), .ZN(n19982) );
  OAI211_X1 U23053 ( .C1(n20360), .C2(n20019), .A(n19983), .B(n19982), .ZN(
        P2_U3078) );
  AOI22_X1 U23054 ( .A1(n20304), .A2(n20011), .B1(n19984), .B2(n20362), .ZN(
        n19988) );
  AOI22_X1 U23055 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19986), .B1(
        n20363), .B2(n19985), .ZN(n19987) );
  OAI211_X1 U23056 ( .C1(n20201), .C2(n19989), .A(n19988), .B(n19987), .ZN(
        P2_U3079) );
  NAND2_X1 U23057 ( .A1(n19990), .A2(n20463), .ZN(n19997) );
  INV_X1 U23058 ( .A(n19991), .ZN(n19994) );
  NOR2_X1 U23059 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19992), .ZN(
        n20014) );
  OAI21_X1 U23060 ( .B1(n19994), .B2(n20014), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19993) );
  OAI21_X1 U23061 ( .B1(n19997), .B2(n20133), .A(n19993), .ZN(n20015) );
  AOI22_X1 U23062 ( .A1(n20015), .A2(n13231), .B1(n20314), .B2(n20014), .ZN(
        n20000) );
  OAI21_X1 U23063 ( .B1(n20011), .B2(n20022), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19996) );
  AOI211_X1 U23064 ( .C1(n19994), .C2(n20101), .A(n20014), .B(n20458), .ZN(
        n19995) );
  AOI211_X1 U23065 ( .C1(n19997), .C2(n19996), .A(n20074), .B(n19995), .ZN(
        n19998) );
  AOI22_X1 U23066 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20016), .B1(
        n20022), .B2(n20173), .ZN(n19999) );
  OAI211_X1 U23067 ( .C1(n20176), .C2(n20019), .A(n20000), .B(n19999), .ZN(
        P2_U3080) );
  AOI22_X1 U23068 ( .A1(n20015), .A2(n14253), .B1(n20326), .B2(n20014), .ZN(
        n20002) );
  AOI22_X1 U23069 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20016), .B1(
        n20022), .B2(n20285), .ZN(n20001) );
  OAI211_X1 U23070 ( .C1(n20179), .C2(n20019), .A(n20002), .B(n20001), .ZN(
        P2_U3081) );
  AOI22_X1 U23071 ( .A1(n20015), .A2(n20332), .B1(n20331), .B2(n20014), .ZN(
        n20004) );
  AOI22_X1 U23072 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20016), .B1(
        n20022), .B2(n20288), .ZN(n20003) );
  OAI211_X1 U23073 ( .C1(n20182), .C2(n20019), .A(n20004), .B(n20003), .ZN(
        P2_U3082) );
  AOI22_X1 U23074 ( .A1(n20015), .A2(n20338), .B1(n20337), .B2(n20014), .ZN(
        n20006) );
  AOI22_X1 U23075 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20016), .B1(
        n20022), .B2(n20291), .ZN(n20005) );
  OAI211_X1 U23076 ( .C1(n20185), .C2(n20019), .A(n20006), .B(n20005), .ZN(
        P2_U3083) );
  AOI22_X1 U23077 ( .A1(n20015), .A2(n20344), .B1(n20343), .B2(n20014), .ZN(
        n20008) );
  AOI22_X1 U23078 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20016), .B1(
        n20022), .B2(n20294), .ZN(n20007) );
  OAI211_X1 U23079 ( .C1(n20188), .C2(n20019), .A(n20008), .B(n20007), .ZN(
        P2_U3084) );
  AOI22_X1 U23080 ( .A1(n20015), .A2(n20350), .B1(n20349), .B2(n20014), .ZN(
        n20010) );
  AOI22_X1 U23081 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20016), .B1(
        n20011), .B2(n20351), .ZN(n20009) );
  OAI211_X1 U23082 ( .C1(n20354), .C2(n20038), .A(n20010), .B(n20009), .ZN(
        P2_U3085) );
  AOI22_X1 U23083 ( .A1(n20015), .A2(n20356), .B1(n20355), .B2(n20014), .ZN(
        n20013) );
  AOI22_X1 U23084 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20016), .B1(
        n20011), .B2(n20357), .ZN(n20012) );
  OAI211_X1 U23085 ( .C1(n20360), .C2(n20038), .A(n20013), .B(n20012), .ZN(
        P2_U3086) );
  AOI22_X1 U23086 ( .A1(n20015), .A2(n20363), .B1(n20362), .B2(n20014), .ZN(
        n20018) );
  AOI22_X1 U23087 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20016), .B1(
        n20022), .B2(n20304), .ZN(n20017) );
  OAI211_X1 U23088 ( .C1(n20201), .C2(n20019), .A(n20018), .B(n20017), .ZN(
        P2_U3087) );
  INV_X1 U23089 ( .A(n20066), .ZN(n20033) );
  AOI22_X1 U23090 ( .A1(n20033), .A2(n20285), .B1(n20326), .B2(n20044), .ZN(
        n20021) );
  AOI22_X1 U23091 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20035), .B1(
        n14253), .B2(n20034), .ZN(n20020) );
  OAI211_X1 U23092 ( .C1(n20179), .C2(n20038), .A(n20021), .B(n20020), .ZN(
        P2_U3089) );
  AOI22_X1 U23093 ( .A1(n20022), .A2(n20333), .B1(n20044), .B2(n20331), .ZN(
        n20024) );
  AOI22_X1 U23094 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20035), .B1(
        n20332), .B2(n20034), .ZN(n20023) );
  OAI211_X1 U23095 ( .C1(n20336), .C2(n20066), .A(n20024), .B(n20023), .ZN(
        P2_U3090) );
  AOI22_X1 U23096 ( .A1(n20033), .A2(n20291), .B1(n20044), .B2(n20337), .ZN(
        n20026) );
  AOI22_X1 U23097 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20035), .B1(
        n20338), .B2(n20034), .ZN(n20025) );
  OAI211_X1 U23098 ( .C1(n20185), .C2(n20038), .A(n20026), .B(n20025), .ZN(
        P2_U3091) );
  AOI22_X1 U23099 ( .A1(n20033), .A2(n20294), .B1(n20044), .B2(n20343), .ZN(
        n20028) );
  AOI22_X1 U23100 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20035), .B1(
        n20344), .B2(n20034), .ZN(n20027) );
  OAI211_X1 U23101 ( .C1(n20188), .C2(n20038), .A(n20028), .B(n20027), .ZN(
        P2_U3092) );
  AOI22_X1 U23102 ( .A1(n20297), .A2(n20033), .B1(n20349), .B2(n20044), .ZN(
        n20030) );
  AOI22_X1 U23103 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20035), .B1(
        n20350), .B2(n20034), .ZN(n20029) );
  OAI211_X1 U23104 ( .C1(n20191), .C2(n20038), .A(n20030), .B(n20029), .ZN(
        P2_U3093) );
  AOI22_X1 U23105 ( .A1(n20300), .A2(n20033), .B1(n20044), .B2(n20355), .ZN(
        n20032) );
  AOI22_X1 U23106 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20035), .B1(
        n20356), .B2(n20034), .ZN(n20031) );
  OAI211_X1 U23107 ( .C1(n20194), .C2(n20038), .A(n20032), .B(n20031), .ZN(
        P2_U3094) );
  AOI22_X1 U23108 ( .A1(n20033), .A2(n20304), .B1(n20044), .B2(n20362), .ZN(
        n20037) );
  AOI22_X1 U23109 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20035), .B1(
        n20363), .B2(n20034), .ZN(n20036) );
  OAI211_X1 U23110 ( .C1(n20201), .C2(n20038), .A(n20037), .B(n20036), .ZN(
        P2_U3095) );
  NOR2_X1 U23111 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20071), .ZN(
        n20061) );
  NOR2_X1 U23112 ( .A1(n20044), .A2(n20061), .ZN(n20040) );
  INV_X1 U23113 ( .A(n10773), .ZN(n20039) );
  NOR3_X1 U23114 ( .A1(n20039), .A2(n20061), .A3(n20312), .ZN(n20045) );
  AOI211_X2 U23115 ( .C1(n20040), .C2(n20312), .A(n20070), .B(n20045), .ZN(
        n20062) );
  AOI22_X1 U23116 ( .A1(n20062), .A2(n13231), .B1(n20314), .B2(n20061), .ZN(
        n20048) );
  INV_X1 U23117 ( .A(n20093), .ZN(n20042) );
  AOI21_X1 U23118 ( .B1(n20066), .B2(n20042), .A(n21150), .ZN(n20043) );
  AOI221_X1 U23119 ( .B1(n20101), .B2(n20044), .C1(n20101), .C2(n20043), .A(
        n20061), .ZN(n20046) );
  AOI22_X1 U23120 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20063), .B1(
        n20093), .B2(n20173), .ZN(n20047) );
  OAI211_X1 U23121 ( .C1(n20176), .C2(n20066), .A(n20048), .B(n20047), .ZN(
        P2_U3096) );
  AOI22_X1 U23122 ( .A1(n20062), .A2(n14253), .B1(n20326), .B2(n20061), .ZN(
        n20050) );
  AOI22_X1 U23123 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20063), .B1(
        n20093), .B2(n20285), .ZN(n20049) );
  OAI211_X1 U23124 ( .C1(n20179), .C2(n20066), .A(n20050), .B(n20049), .ZN(
        P2_U3097) );
  AOI22_X1 U23125 ( .A1(n20062), .A2(n20332), .B1(n20331), .B2(n20061), .ZN(
        n20052) );
  AOI22_X1 U23126 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20063), .B1(
        n20093), .B2(n20288), .ZN(n20051) );
  OAI211_X1 U23127 ( .C1(n20182), .C2(n20066), .A(n20052), .B(n20051), .ZN(
        P2_U3098) );
  AOI22_X1 U23128 ( .A1(n20062), .A2(n20338), .B1(n20337), .B2(n20061), .ZN(
        n20054) );
  AOI22_X1 U23129 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20063), .B1(
        n20093), .B2(n20291), .ZN(n20053) );
  OAI211_X1 U23130 ( .C1(n20185), .C2(n20066), .A(n20054), .B(n20053), .ZN(
        P2_U3099) );
  AOI22_X1 U23131 ( .A1(n20062), .A2(n20344), .B1(n20343), .B2(n20061), .ZN(
        n20056) );
  AOI22_X1 U23132 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20063), .B1(
        n20093), .B2(n20294), .ZN(n20055) );
  OAI211_X1 U23133 ( .C1(n20188), .C2(n20066), .A(n20056), .B(n20055), .ZN(
        P2_U3100) );
  AOI22_X1 U23134 ( .A1(n20062), .A2(n20350), .B1(n20349), .B2(n20061), .ZN(
        n20058) );
  AOI22_X1 U23135 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20063), .B1(
        n20093), .B2(n20297), .ZN(n20057) );
  OAI211_X1 U23136 ( .C1(n20191), .C2(n20066), .A(n20058), .B(n20057), .ZN(
        P2_U3101) );
  AOI22_X1 U23137 ( .A1(n20062), .A2(n20356), .B1(n20355), .B2(n20061), .ZN(
        n20060) );
  AOI22_X1 U23138 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20063), .B1(
        n20093), .B2(n20300), .ZN(n20059) );
  OAI211_X1 U23139 ( .C1(n20194), .C2(n20066), .A(n20060), .B(n20059), .ZN(
        P2_U3102) );
  AOI22_X1 U23140 ( .A1(n20062), .A2(n20363), .B1(n20362), .B2(n20061), .ZN(
        n20065) );
  AOI22_X1 U23141 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20063), .B1(
        n20093), .B2(n20304), .ZN(n20064) );
  OAI211_X1 U23142 ( .C1(n20201), .C2(n20066), .A(n20065), .B(n20064), .ZN(
        P2_U3103) );
  INV_X1 U23143 ( .A(n10759), .ZN(n20069) );
  NOR3_X1 U23144 ( .A1(n20069), .A2(n20091), .A3(n20312), .ZN(n20073) );
  AOI211_X2 U23145 ( .C1(n20071), .C2(n20312), .A(n20070), .B(n20073), .ZN(
        n20092) );
  AOI22_X1 U23146 ( .A1(n20092), .A2(n13231), .B1(n20314), .B2(n20091), .ZN(
        n20078) );
  INV_X1 U23147 ( .A(n20071), .ZN(n20076) );
  NOR2_X1 U23148 ( .A1(n20072), .A2(n20316), .ZN(n20457) );
  INV_X1 U23149 ( .A(n20091), .ZN(n20104) );
  AOI211_X1 U23150 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20104), .A(n20074), 
        .B(n20073), .ZN(n20075) );
  OAI21_X1 U23151 ( .B1(n20076), .B2(n20457), .A(n20075), .ZN(n20094) );
  AOI22_X1 U23152 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20094), .B1(
        n20093), .B2(n20322), .ZN(n20077) );
  OAI211_X1 U23153 ( .C1(n20325), .C2(n20129), .A(n20078), .B(n20077), .ZN(
        P2_U3104) );
  AOI22_X1 U23154 ( .A1(n20092), .A2(n14253), .B1(n20326), .B2(n20091), .ZN(
        n20080) );
  AOI22_X1 U23155 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20094), .B1(
        n20093), .B2(n20327), .ZN(n20079) );
  OAI211_X1 U23156 ( .C1(n20330), .C2(n20129), .A(n20080), .B(n20079), .ZN(
        P2_U3105) );
  AOI22_X1 U23157 ( .A1(n20092), .A2(n20332), .B1(n20331), .B2(n20091), .ZN(
        n20082) );
  AOI22_X1 U23158 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20094), .B1(
        n20093), .B2(n20333), .ZN(n20081) );
  OAI211_X1 U23159 ( .C1(n20336), .C2(n20129), .A(n20082), .B(n20081), .ZN(
        P2_U3106) );
  AOI22_X1 U23160 ( .A1(n20092), .A2(n20338), .B1(n20337), .B2(n20091), .ZN(
        n20084) );
  AOI22_X1 U23161 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20094), .B1(
        n20093), .B2(n20339), .ZN(n20083) );
  OAI211_X1 U23162 ( .C1(n20342), .C2(n20129), .A(n20084), .B(n20083), .ZN(
        P2_U3107) );
  AOI22_X1 U23163 ( .A1(n20092), .A2(n20344), .B1(n20343), .B2(n20091), .ZN(
        n20086) );
  AOI22_X1 U23164 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20094), .B1(
        n20093), .B2(n20345), .ZN(n20085) );
  OAI211_X1 U23165 ( .C1(n20348), .C2(n20129), .A(n20086), .B(n20085), .ZN(
        P2_U3108) );
  AOI22_X1 U23166 ( .A1(n20092), .A2(n20350), .B1(n20349), .B2(n20091), .ZN(
        n20088) );
  AOI22_X1 U23167 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20094), .B1(
        n20093), .B2(n20351), .ZN(n20087) );
  OAI211_X1 U23168 ( .C1(n20354), .C2(n20129), .A(n20088), .B(n20087), .ZN(
        P2_U3109) );
  AOI22_X1 U23169 ( .A1(n20092), .A2(n20356), .B1(n20355), .B2(n20091), .ZN(
        n20090) );
  AOI22_X1 U23170 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20094), .B1(
        n20093), .B2(n20357), .ZN(n20089) );
  OAI211_X1 U23171 ( .C1(n20360), .C2(n20129), .A(n20090), .B(n20089), .ZN(
        P2_U3110) );
  AOI22_X1 U23172 ( .A1(n20092), .A2(n20363), .B1(n20362), .B2(n20091), .ZN(
        n20096) );
  AOI22_X1 U23173 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20094), .B1(
        n20093), .B2(n20365), .ZN(n20095) );
  OAI211_X1 U23174 ( .C1(n20371), .C2(n20129), .A(n20096), .B(n20095), .ZN(
        P2_U3111) );
  INV_X1 U23175 ( .A(n20166), .ZN(n20098) );
  NAND2_X1 U23176 ( .A1(n20470), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20202) );
  NOR2_X1 U23177 ( .A1(n20202), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20135) );
  INV_X1 U23178 ( .A(n20135), .ZN(n20139) );
  NOR2_X1 U23179 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20139), .ZN(
        n20124) );
  AOI22_X1 U23180 ( .A1(n20153), .A2(n20173), .B1(n20314), .B2(n20124), .ZN(
        n20111) );
  AOI21_X1 U23181 ( .B1(n20161), .B2(n20129), .A(n21150), .ZN(n20099) );
  NOR2_X1 U23182 ( .A1(n20099), .A2(n20133), .ZN(n20105) );
  INV_X1 U23183 ( .A(n20100), .ZN(n20107) );
  OAI21_X1 U23184 ( .B1(n20107), .B2(n20312), .A(n20101), .ZN(n20102) );
  AOI21_X1 U23185 ( .B1(n20105), .B2(n20104), .A(n20102), .ZN(n20103) );
  INV_X1 U23186 ( .A(n20104), .ZN(n20106) );
  OAI21_X1 U23187 ( .B1(n20124), .B2(n20106), .A(n20105), .ZN(n20109) );
  OAI21_X1 U23188 ( .B1(n20107), .B2(n20124), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20108) );
  NAND2_X1 U23189 ( .A1(n20109), .A2(n20108), .ZN(n20125) );
  AOI22_X1 U23190 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20126), .B1(
        n13231), .B2(n20125), .ZN(n20110) );
  OAI211_X1 U23191 ( .C1(n20176), .C2(n20129), .A(n20111), .B(n20110), .ZN(
        P2_U3112) );
  AOI22_X1 U23192 ( .A1(n20153), .A2(n20285), .B1(n20326), .B2(n20124), .ZN(
        n20113) );
  AOI22_X1 U23193 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20126), .B1(
        n20125), .B2(n14253), .ZN(n20112) );
  OAI211_X1 U23194 ( .C1(n20179), .C2(n20129), .A(n20113), .B(n20112), .ZN(
        P2_U3113) );
  AOI22_X1 U23195 ( .A1(n20153), .A2(n20288), .B1(n20331), .B2(n20124), .ZN(
        n20115) );
  AOI22_X1 U23196 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20126), .B1(
        n20125), .B2(n20332), .ZN(n20114) );
  OAI211_X1 U23197 ( .C1(n20182), .C2(n20129), .A(n20115), .B(n20114), .ZN(
        P2_U3114) );
  AOI22_X1 U23198 ( .A1(n20153), .A2(n20291), .B1(n20337), .B2(n20124), .ZN(
        n20117) );
  AOI22_X1 U23199 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20126), .B1(
        n20125), .B2(n20338), .ZN(n20116) );
  OAI211_X1 U23200 ( .C1(n20185), .C2(n20129), .A(n20117), .B(n20116), .ZN(
        P2_U3115) );
  AOI22_X1 U23201 ( .A1(n20153), .A2(n20294), .B1(n20343), .B2(n20124), .ZN(
        n20119) );
  AOI22_X1 U23202 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20126), .B1(
        n20125), .B2(n20344), .ZN(n20118) );
  OAI211_X1 U23203 ( .C1(n20188), .C2(n20129), .A(n20119), .B(n20118), .ZN(
        P2_U3116) );
  AOI22_X1 U23204 ( .A1(n20153), .A2(n20297), .B1(n20349), .B2(n20124), .ZN(
        n20121) );
  AOI22_X1 U23205 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20126), .B1(
        n20125), .B2(n20350), .ZN(n20120) );
  OAI211_X1 U23206 ( .C1(n20191), .C2(n20129), .A(n20121), .B(n20120), .ZN(
        P2_U3117) );
  AOI22_X1 U23207 ( .A1(n20153), .A2(n20300), .B1(n20355), .B2(n20124), .ZN(
        n20123) );
  AOI22_X1 U23208 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20126), .B1(
        n20125), .B2(n20356), .ZN(n20122) );
  OAI211_X1 U23209 ( .C1(n20194), .C2(n20129), .A(n20123), .B(n20122), .ZN(
        P2_U3118) );
  AOI22_X1 U23210 ( .A1(n20153), .A2(n20304), .B1(n20362), .B2(n20124), .ZN(
        n20128) );
  AOI22_X1 U23211 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20126), .B1(
        n20125), .B2(n20363), .ZN(n20127) );
  OAI211_X1 U23212 ( .C1(n20201), .C2(n20129), .A(n20128), .B(n20127), .ZN(
        P2_U3119) );
  INV_X1 U23213 ( .A(n20202), .ZN(n20206) );
  NAND2_X1 U23214 ( .A1(n20131), .A2(n20206), .ZN(n20170) );
  INV_X1 U23215 ( .A(n20170), .ZN(n20156) );
  AOI22_X1 U23216 ( .A1(n20167), .A2(n20173), .B1(n20314), .B2(n20156), .ZN(
        n20142) );
  NAND2_X1 U23217 ( .A1(n20460), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20317) );
  OAI21_X1 U23218 ( .B1(n20317), .B2(n20132), .A(n20458), .ZN(n20140) );
  OAI211_X1 U23219 ( .C1(n20136), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20170), 
        .B(n20133), .ZN(n20134) );
  OAI211_X1 U23220 ( .C1(n20140), .C2(n20135), .A(n20320), .B(n20134), .ZN(
        n20158) );
  INV_X1 U23221 ( .A(n20136), .ZN(n20137) );
  OAI21_X1 U23222 ( .B1(n20137), .B2(n20156), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20138) );
  OAI21_X1 U23223 ( .B1(n20140), .B2(n20139), .A(n20138), .ZN(n20157) );
  AOI22_X1 U23224 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20158), .B1(
        n13231), .B2(n20157), .ZN(n20141) );
  OAI211_X1 U23225 ( .C1(n20176), .C2(n20161), .A(n20142), .B(n20141), .ZN(
        P2_U3120) );
  AOI22_X1 U23226 ( .A1(n20153), .A2(n20327), .B1(n20326), .B2(n20156), .ZN(
        n20144) );
  AOI22_X1 U23227 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20158), .B1(
        n14253), .B2(n20157), .ZN(n20143) );
  OAI211_X1 U23228 ( .C1(n20330), .C2(n20200), .A(n20144), .B(n20143), .ZN(
        P2_U3121) );
  AOI22_X1 U23229 ( .A1(n20153), .A2(n20333), .B1(n20331), .B2(n20156), .ZN(
        n20146) );
  AOI22_X1 U23230 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20158), .B1(
        n20332), .B2(n20157), .ZN(n20145) );
  OAI211_X1 U23231 ( .C1(n20336), .C2(n20200), .A(n20146), .B(n20145), .ZN(
        P2_U3122) );
  AOI22_X1 U23232 ( .A1(n20339), .A2(n20153), .B1(n20337), .B2(n20156), .ZN(
        n20148) );
  AOI22_X1 U23233 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20158), .B1(
        n20338), .B2(n20157), .ZN(n20147) );
  OAI211_X1 U23234 ( .C1(n20342), .C2(n20200), .A(n20148), .B(n20147), .ZN(
        P2_U3123) );
  AOI22_X1 U23235 ( .A1(n20167), .A2(n20294), .B1(n20343), .B2(n20156), .ZN(
        n20150) );
  AOI22_X1 U23236 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20158), .B1(
        n20344), .B2(n20157), .ZN(n20149) );
  OAI211_X1 U23237 ( .C1(n20188), .C2(n20161), .A(n20150), .B(n20149), .ZN(
        P2_U3124) );
  AOI22_X1 U23238 ( .A1(n20153), .A2(n20351), .B1(n20349), .B2(n20156), .ZN(
        n20152) );
  AOI22_X1 U23239 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20158), .B1(
        n20350), .B2(n20157), .ZN(n20151) );
  OAI211_X1 U23240 ( .C1(n20354), .C2(n20200), .A(n20152), .B(n20151), .ZN(
        P2_U3125) );
  AOI22_X1 U23241 ( .A1(n20357), .A2(n20153), .B1(n20355), .B2(n20156), .ZN(
        n20155) );
  AOI22_X1 U23242 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20158), .B1(
        n20356), .B2(n20157), .ZN(n20154) );
  OAI211_X1 U23243 ( .C1(n20360), .C2(n20200), .A(n20155), .B(n20154), .ZN(
        P2_U3126) );
  AOI22_X1 U23244 ( .A1(n20167), .A2(n20304), .B1(n20362), .B2(n20156), .ZN(
        n20160) );
  AOI22_X1 U23245 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20158), .B1(
        n20363), .B2(n20157), .ZN(n20159) );
  OAI211_X1 U23246 ( .C1(n20201), .C2(n20161), .A(n20160), .B(n20159), .ZN(
        P2_U3127) );
  INV_X1 U23247 ( .A(n20162), .ZN(n20168) );
  AND2_X1 U23248 ( .A1(n20163), .A2(n20206), .ZN(n20195) );
  OAI21_X1 U23249 ( .B1(n20168), .B2(n20195), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20164) );
  OAI21_X1 U23250 ( .B1(n20202), .B2(n20165), .A(n20164), .ZN(n20196) );
  AOI22_X1 U23251 ( .A1(n20196), .A2(n13231), .B1(n20314), .B2(n20195), .ZN(
        n20175) );
  OAI21_X1 U23252 ( .B1(n20167), .B2(n20229), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20171) );
  OAI21_X1 U23253 ( .B1(n20168), .B2(n20312), .A(n20101), .ZN(n20169) );
  AOI21_X1 U23254 ( .B1(n20171), .B2(n20170), .A(n20169), .ZN(n20172) );
  AOI22_X1 U23255 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20197), .B1(
        n20229), .B2(n20173), .ZN(n20174) );
  OAI211_X1 U23256 ( .C1(n20176), .C2(n20200), .A(n20175), .B(n20174), .ZN(
        P2_U3128) );
  AOI22_X1 U23257 ( .A1(n20196), .A2(n14253), .B1(n20326), .B2(n20195), .ZN(
        n20178) );
  AOI22_X1 U23258 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20197), .B1(
        n20229), .B2(n20285), .ZN(n20177) );
  OAI211_X1 U23259 ( .C1(n20179), .C2(n20200), .A(n20178), .B(n20177), .ZN(
        P2_U3129) );
  AOI22_X1 U23260 ( .A1(n20196), .A2(n20332), .B1(n20331), .B2(n20195), .ZN(
        n20181) );
  AOI22_X1 U23261 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20197), .B1(
        n20229), .B2(n20288), .ZN(n20180) );
  OAI211_X1 U23262 ( .C1(n20182), .C2(n20200), .A(n20181), .B(n20180), .ZN(
        P2_U3130) );
  AOI22_X1 U23263 ( .A1(n20196), .A2(n20338), .B1(n20337), .B2(n20195), .ZN(
        n20184) );
  AOI22_X1 U23264 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20197), .B1(
        n20229), .B2(n20291), .ZN(n20183) );
  OAI211_X1 U23265 ( .C1(n20185), .C2(n20200), .A(n20184), .B(n20183), .ZN(
        P2_U3131) );
  AOI22_X1 U23266 ( .A1(n20196), .A2(n20344), .B1(n20343), .B2(n20195), .ZN(
        n20187) );
  AOI22_X1 U23267 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20197), .B1(
        n20229), .B2(n20294), .ZN(n20186) );
  OAI211_X1 U23268 ( .C1(n20188), .C2(n20200), .A(n20187), .B(n20186), .ZN(
        P2_U3132) );
  AOI22_X1 U23269 ( .A1(n20196), .A2(n20350), .B1(n20349), .B2(n20195), .ZN(
        n20190) );
  AOI22_X1 U23270 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20197), .B1(
        n20229), .B2(n20297), .ZN(n20189) );
  OAI211_X1 U23271 ( .C1(n20191), .C2(n20200), .A(n20190), .B(n20189), .ZN(
        P2_U3133) );
  AOI22_X1 U23272 ( .A1(n20196), .A2(n20356), .B1(n20355), .B2(n20195), .ZN(
        n20193) );
  AOI22_X1 U23273 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20197), .B1(
        n20229), .B2(n20300), .ZN(n20192) );
  OAI211_X1 U23274 ( .C1(n20194), .C2(n20200), .A(n20193), .B(n20192), .ZN(
        P2_U3134) );
  AOI22_X1 U23275 ( .A1(n20196), .A2(n20363), .B1(n20362), .B2(n20195), .ZN(
        n20199) );
  AOI22_X1 U23276 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20197), .B1(
        n20229), .B2(n20304), .ZN(n20198) );
  OAI211_X1 U23277 ( .C1(n20201), .C2(n20200), .A(n20199), .B(n20198), .ZN(
        P2_U3135) );
  NOR2_X1 U23278 ( .A1(n20203), .A2(n20202), .ZN(n20227) );
  NOR2_X1 U23279 ( .A1(n20227), .A2(n20312), .ZN(n20204) );
  NAND2_X1 U23280 ( .A1(n20205), .A2(n20204), .ZN(n20210) );
  NAND2_X1 U23281 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20206), .ZN(
        n20208) );
  OAI21_X1 U23282 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20208), .A(n20312), 
        .ZN(n20207) );
  AND2_X1 U23283 ( .A1(n20210), .A2(n20207), .ZN(n20228) );
  AOI22_X1 U23284 ( .A1(n20228), .A2(n13231), .B1(n20314), .B2(n20227), .ZN(
        n20214) );
  OAI21_X1 U23285 ( .B1(n20317), .B2(n20209), .A(n20208), .ZN(n20211) );
  AND2_X1 U23286 ( .A1(n20211), .A2(n20210), .ZN(n20212) );
  OAI211_X1 U23287 ( .C1(n20227), .C2(n20101), .A(n20212), .B(n20320), .ZN(
        n20230) );
  AOI22_X1 U23288 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20230), .B1(
        n20229), .B2(n20322), .ZN(n20213) );
  OAI211_X1 U23289 ( .C1(n20325), .C2(n20233), .A(n20214), .B(n20213), .ZN(
        P2_U3136) );
  AOI22_X1 U23290 ( .A1(n20228), .A2(n14253), .B1(n20326), .B2(n20227), .ZN(
        n20216) );
  AOI22_X1 U23291 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20230), .B1(
        n20229), .B2(n20327), .ZN(n20215) );
  OAI211_X1 U23292 ( .C1(n20330), .C2(n20233), .A(n20216), .B(n20215), .ZN(
        P2_U3137) );
  AOI22_X1 U23293 ( .A1(n20228), .A2(n20332), .B1(n20331), .B2(n20227), .ZN(
        n20218) );
  AOI22_X1 U23294 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20230), .B1(
        n20229), .B2(n20333), .ZN(n20217) );
  OAI211_X1 U23295 ( .C1(n20336), .C2(n20233), .A(n20218), .B(n20217), .ZN(
        P2_U3138) );
  AOI22_X1 U23296 ( .A1(n20228), .A2(n20338), .B1(n20337), .B2(n20227), .ZN(
        n20220) );
  AOI22_X1 U23297 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20230), .B1(
        n20229), .B2(n20339), .ZN(n20219) );
  OAI211_X1 U23298 ( .C1(n20342), .C2(n20233), .A(n20220), .B(n20219), .ZN(
        P2_U3139) );
  AOI22_X1 U23299 ( .A1(n20228), .A2(n20344), .B1(n20343), .B2(n20227), .ZN(
        n20222) );
  AOI22_X1 U23300 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20230), .B1(
        n20229), .B2(n20345), .ZN(n20221) );
  OAI211_X1 U23301 ( .C1(n20348), .C2(n20233), .A(n20222), .B(n20221), .ZN(
        P2_U3140) );
  AOI22_X1 U23302 ( .A1(n20228), .A2(n20350), .B1(n20349), .B2(n20227), .ZN(
        n20224) );
  AOI22_X1 U23303 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20230), .B1(
        n20229), .B2(n20351), .ZN(n20223) );
  OAI211_X1 U23304 ( .C1(n20354), .C2(n20233), .A(n20224), .B(n20223), .ZN(
        P2_U3141) );
  AOI22_X1 U23305 ( .A1(n20228), .A2(n20356), .B1(n20355), .B2(n20227), .ZN(
        n20226) );
  AOI22_X1 U23306 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20230), .B1(
        n20229), .B2(n20357), .ZN(n20225) );
  OAI211_X1 U23307 ( .C1(n20360), .C2(n20233), .A(n20226), .B(n20225), .ZN(
        P2_U3142) );
  AOI22_X1 U23308 ( .A1(n20228), .A2(n20363), .B1(n20362), .B2(n20227), .ZN(
        n20232) );
  AOI22_X1 U23309 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20230), .B1(
        n20229), .B2(n20365), .ZN(n20231) );
  OAI211_X1 U23310 ( .C1(n20371), .C2(n20233), .A(n20232), .B(n20231), .ZN(
        P2_U3143) );
  INV_X1 U23311 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n20236) );
  AOI22_X1 U23312 ( .A1(n20249), .A2(n14253), .B1(n20326), .B2(n20248), .ZN(
        n20235) );
  AOI22_X1 U23313 ( .A1(n20280), .A2(n20285), .B1(n20250), .B2(n20327), .ZN(
        n20234) );
  OAI211_X1 U23314 ( .C1(n20254), .C2(n20236), .A(n20235), .B(n20234), .ZN(
        P2_U3145) );
  INV_X1 U23315 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20239) );
  AOI22_X1 U23316 ( .A1(n20249), .A2(n20332), .B1(n20248), .B2(n20331), .ZN(
        n20238) );
  AOI22_X1 U23317 ( .A1(n20280), .A2(n20288), .B1(n20250), .B2(n20333), .ZN(
        n20237) );
  OAI211_X1 U23318 ( .C1(n20254), .C2(n20239), .A(n20238), .B(n20237), .ZN(
        P2_U3146) );
  AOI22_X1 U23319 ( .A1(n20249), .A2(n20338), .B1(n20248), .B2(n20337), .ZN(
        n20241) );
  AOI22_X1 U23320 ( .A1(n20280), .A2(n20291), .B1(n20250), .B2(n20339), .ZN(
        n20240) );
  OAI211_X1 U23321 ( .C1(n20254), .C2(n21045), .A(n20241), .B(n20240), .ZN(
        P2_U3147) );
  AOI22_X1 U23322 ( .A1(n20249), .A2(n20344), .B1(n20248), .B2(n20343), .ZN(
        n20243) );
  AOI22_X1 U23323 ( .A1(n20280), .A2(n20294), .B1(n20250), .B2(n20345), .ZN(
        n20242) );
  OAI211_X1 U23324 ( .C1(n20254), .C2(n10724), .A(n20243), .B(n20242), .ZN(
        P2_U3148) );
  AOI22_X1 U23325 ( .A1(n20249), .A2(n20350), .B1(n20349), .B2(n20248), .ZN(
        n20245) );
  AOI22_X1 U23326 ( .A1(n20280), .A2(n20297), .B1(n20250), .B2(n20351), .ZN(
        n20244) );
  OAI211_X1 U23327 ( .C1(n20254), .C2(n10775), .A(n20245), .B(n20244), .ZN(
        P2_U3149) );
  AOI22_X1 U23328 ( .A1(n20249), .A2(n20356), .B1(n20248), .B2(n20355), .ZN(
        n20247) );
  AOI22_X1 U23329 ( .A1(n20280), .A2(n20300), .B1(n20250), .B2(n20357), .ZN(
        n20246) );
  OAI211_X1 U23330 ( .C1(n20254), .C2(n11733), .A(n20247), .B(n20246), .ZN(
        P2_U3150) );
  INV_X1 U23331 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n20253) );
  AOI22_X1 U23332 ( .A1(n20249), .A2(n20363), .B1(n20248), .B2(n20362), .ZN(
        n20252) );
  AOI22_X1 U23333 ( .A1(n20280), .A2(n20304), .B1(n20250), .B2(n20365), .ZN(
        n20251) );
  OAI211_X1 U23334 ( .C1(n20254), .C2(n20253), .A(n20252), .B(n20251), .ZN(
        P2_U3151) );
  INV_X1 U23335 ( .A(n20278), .ZN(n20255) );
  AND2_X1 U23336 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20255), .ZN(n20256) );
  NAND2_X1 U23337 ( .A1(n20257), .A2(n20256), .ZN(n20261) );
  OAI21_X1 U23338 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20259), .A(n20312), 
        .ZN(n20258) );
  AOI22_X1 U23339 ( .A1(n20279), .A2(n13231), .B1(n20314), .B2(n20278), .ZN(
        n20265) );
  OAI21_X1 U23340 ( .B1(n20317), .B2(n20260), .A(n20259), .ZN(n20262) );
  AND2_X1 U23341 ( .A1(n20262), .A2(n20261), .ZN(n20263) );
  OAI211_X1 U23342 ( .C1(n20278), .C2(n20101), .A(n20263), .B(n20320), .ZN(
        n20281) );
  AOI22_X1 U23343 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20322), .ZN(n20264) );
  OAI211_X1 U23344 ( .C1(n20325), .C2(n20284), .A(n20265), .B(n20264), .ZN(
        P2_U3152) );
  AOI22_X1 U23345 ( .A1(n20279), .A2(n14253), .B1(n20326), .B2(n20278), .ZN(
        n20267) );
  AOI22_X1 U23346 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20327), .ZN(n20266) );
  OAI211_X1 U23347 ( .C1(n20330), .C2(n20284), .A(n20267), .B(n20266), .ZN(
        P2_U3153) );
  AOI22_X1 U23348 ( .A1(n20279), .A2(n20332), .B1(n20331), .B2(n20278), .ZN(
        n20269) );
  AOI22_X1 U23349 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20333), .ZN(n20268) );
  OAI211_X1 U23350 ( .C1(n20336), .C2(n20284), .A(n20269), .B(n20268), .ZN(
        P2_U3154) );
  AOI22_X1 U23351 ( .A1(n20279), .A2(n20338), .B1(n20337), .B2(n20278), .ZN(
        n20271) );
  AOI22_X1 U23352 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20339), .ZN(n20270) );
  OAI211_X1 U23353 ( .C1(n20342), .C2(n20284), .A(n20271), .B(n20270), .ZN(
        P2_U3155) );
  AOI22_X1 U23354 ( .A1(n20279), .A2(n20344), .B1(n20343), .B2(n20278), .ZN(
        n20273) );
  AOI22_X1 U23355 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20345), .ZN(n20272) );
  OAI211_X1 U23356 ( .C1(n20348), .C2(n20284), .A(n20273), .B(n20272), .ZN(
        P2_U3156) );
  AOI22_X1 U23357 ( .A1(n20279), .A2(n20350), .B1(n20349), .B2(n20278), .ZN(
        n20275) );
  AOI22_X1 U23358 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20351), .ZN(n20274) );
  OAI211_X1 U23359 ( .C1(n20354), .C2(n20284), .A(n20275), .B(n20274), .ZN(
        P2_U3157) );
  AOI22_X1 U23360 ( .A1(n20279), .A2(n20356), .B1(n20355), .B2(n20278), .ZN(
        n20277) );
  AOI22_X1 U23361 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20357), .ZN(n20276) );
  OAI211_X1 U23362 ( .C1(n20360), .C2(n20284), .A(n20277), .B(n20276), .ZN(
        P2_U3158) );
  AOI22_X1 U23363 ( .A1(n20279), .A2(n20363), .B1(n20362), .B2(n20278), .ZN(
        n20283) );
  AOI22_X1 U23364 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20365), .ZN(n20282) );
  OAI211_X1 U23365 ( .C1(n20371), .C2(n20284), .A(n20283), .B(n20282), .ZN(
        P2_U3159) );
  AOI22_X1 U23366 ( .A1(n20366), .A2(n20285), .B1(n20303), .B2(n20326), .ZN(
        n20287) );
  AOI22_X1 U23367 ( .A1(n14253), .A2(n20306), .B1(n20305), .B2(n20327), .ZN(
        n20286) );
  OAI211_X1 U23368 ( .C1(n20309), .C2(n11217), .A(n20287), .B(n20286), .ZN(
        P2_U3161) );
  AOI22_X1 U23369 ( .A1(n20288), .A2(n20366), .B1(n20303), .B2(n20331), .ZN(
        n20290) );
  AOI22_X1 U23370 ( .A1(n20332), .A2(n20306), .B1(n20305), .B2(n20333), .ZN(
        n20289) );
  OAI211_X1 U23371 ( .C1(n20309), .C2(n11237), .A(n20290), .B(n20289), .ZN(
        P2_U3162) );
  AOI22_X1 U23372 ( .A1(n20366), .A2(n20291), .B1(n20303), .B2(n20337), .ZN(
        n20293) );
  AOI22_X1 U23373 ( .A1(n20338), .A2(n20306), .B1(n20305), .B2(n20339), .ZN(
        n20292) );
  OAI211_X1 U23374 ( .C1(n20309), .C2(n11271), .A(n20293), .B(n20292), .ZN(
        P2_U3163) );
  AOI22_X1 U23375 ( .A1(n20345), .A2(n20305), .B1(n20303), .B2(n20343), .ZN(
        n20296) );
  AOI22_X1 U23376 ( .A1(n20344), .A2(n20306), .B1(n20366), .B2(n20294), .ZN(
        n20295) );
  OAI211_X1 U23377 ( .C1(n20309), .C2(n11287), .A(n20296), .B(n20295), .ZN(
        P2_U3164) );
  AOI22_X1 U23378 ( .A1(n20305), .A2(n20351), .B1(n20303), .B2(n20349), .ZN(
        n20299) );
  AOI22_X1 U23379 ( .A1(n20350), .A2(n20306), .B1(n20366), .B2(n20297), .ZN(
        n20298) );
  OAI211_X1 U23380 ( .C1(n20309), .C2(n11309), .A(n20299), .B(n20298), .ZN(
        P2_U3165) );
  AOI22_X1 U23381 ( .A1(n20300), .A2(n20366), .B1(n20303), .B2(n20355), .ZN(
        n20302) );
  AOI22_X1 U23382 ( .A1(n20356), .A2(n20306), .B1(n20305), .B2(n20357), .ZN(
        n20301) );
  OAI211_X1 U23383 ( .C1(n20309), .C2(n11329), .A(n20302), .B(n20301), .ZN(
        P2_U3166) );
  AOI22_X1 U23384 ( .A1(n20366), .A2(n20304), .B1(n20303), .B2(n20362), .ZN(
        n20308) );
  AOI22_X1 U23385 ( .A1(n20363), .A2(n20306), .B1(n20305), .B2(n20365), .ZN(
        n20307) );
  OAI211_X1 U23386 ( .C1(n20309), .C2(n11353), .A(n20308), .B(n20307), .ZN(
        P2_U3167) );
  NOR2_X1 U23387 ( .A1(n20361), .A2(n20312), .ZN(n20310) );
  NAND2_X1 U23388 ( .A1(n10772), .A2(n20310), .ZN(n20318) );
  NAND2_X1 U23389 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20311), .ZN(
        n20315) );
  OAI21_X1 U23390 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20315), .A(n20312), 
        .ZN(n20313) );
  AND2_X1 U23391 ( .A1(n20318), .A2(n20313), .ZN(n20364) );
  AOI22_X1 U23392 ( .A1(n20364), .A2(n13231), .B1(n20314), .B2(n20361), .ZN(
        n20324) );
  OAI21_X1 U23393 ( .B1(n20317), .B2(n20316), .A(n20315), .ZN(n20319) );
  AND2_X1 U23394 ( .A1(n20319), .A2(n20318), .ZN(n20321) );
  OAI211_X1 U23395 ( .C1(n20361), .C2(n20101), .A(n20321), .B(n20320), .ZN(
        n20367) );
  AOI22_X1 U23396 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20322), .ZN(n20323) );
  OAI211_X1 U23397 ( .C1(n20325), .C2(n20370), .A(n20324), .B(n20323), .ZN(
        P2_U3168) );
  AOI22_X1 U23398 ( .A1(n20364), .A2(n14253), .B1(n20326), .B2(n20361), .ZN(
        n20329) );
  AOI22_X1 U23399 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20327), .ZN(n20328) );
  OAI211_X1 U23400 ( .C1(n20330), .C2(n20370), .A(n20329), .B(n20328), .ZN(
        P2_U3169) );
  AOI22_X1 U23401 ( .A1(n20364), .A2(n20332), .B1(n20331), .B2(n20361), .ZN(
        n20335) );
  AOI22_X1 U23402 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20333), .ZN(n20334) );
  OAI211_X1 U23403 ( .C1(n20336), .C2(n20370), .A(n20335), .B(n20334), .ZN(
        P2_U3170) );
  AOI22_X1 U23404 ( .A1(n20364), .A2(n20338), .B1(n20337), .B2(n20361), .ZN(
        n20341) );
  AOI22_X1 U23405 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20339), .ZN(n20340) );
  OAI211_X1 U23406 ( .C1(n20342), .C2(n20370), .A(n20341), .B(n20340), .ZN(
        P2_U3171) );
  AOI22_X1 U23407 ( .A1(n20364), .A2(n20344), .B1(n20343), .B2(n20361), .ZN(
        n20347) );
  AOI22_X1 U23408 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20345), .ZN(n20346) );
  OAI211_X1 U23409 ( .C1(n20348), .C2(n20370), .A(n20347), .B(n20346), .ZN(
        P2_U3172) );
  AOI22_X1 U23410 ( .A1(n20364), .A2(n20350), .B1(n20349), .B2(n20361), .ZN(
        n20353) );
  AOI22_X1 U23411 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20351), .ZN(n20352) );
  OAI211_X1 U23412 ( .C1(n20354), .C2(n20370), .A(n20353), .B(n20352), .ZN(
        P2_U3173) );
  AOI22_X1 U23413 ( .A1(n20364), .A2(n20356), .B1(n20355), .B2(n20361), .ZN(
        n20359) );
  AOI22_X1 U23414 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20357), .ZN(n20358) );
  OAI211_X1 U23415 ( .C1(n20360), .C2(n20370), .A(n20359), .B(n20358), .ZN(
        P2_U3174) );
  AOI22_X1 U23416 ( .A1(n20364), .A2(n20363), .B1(n20362), .B2(n20361), .ZN(
        n20369) );
  AOI22_X1 U23417 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20365), .ZN(n20368) );
  OAI211_X1 U23418 ( .C1(n20371), .C2(n20370), .A(n20369), .B(n20368), .ZN(
        P2_U3175) );
  INV_X1 U23419 ( .A(n20453), .ZN(n20372) );
  AND2_X1 U23420 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20372), .ZN(
        P2_U3179) );
  AND2_X1 U23421 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20372), .ZN(
        P2_U3180) );
  AND2_X1 U23422 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20372), .ZN(
        P2_U3181) );
  AND2_X1 U23423 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20372), .ZN(
        P2_U3182) );
  AND2_X1 U23424 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20372), .ZN(
        P2_U3183) );
  AND2_X1 U23425 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20372), .ZN(
        P2_U3184) );
  AND2_X1 U23426 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20372), .ZN(
        P2_U3185) );
  AND2_X1 U23427 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20372), .ZN(
        P2_U3186) );
  AND2_X1 U23428 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20372), .ZN(
        P2_U3187) );
  AND2_X1 U23429 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20372), .ZN(
        P2_U3188) );
  AND2_X1 U23430 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20372), .ZN(
        P2_U3189) );
  AND2_X1 U23431 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20372), .ZN(
        P2_U3190) );
  AND2_X1 U23432 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20372), .ZN(
        P2_U3191) );
  AND2_X1 U23433 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20372), .ZN(
        P2_U3192) );
  AND2_X1 U23434 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20372), .ZN(
        P2_U3193) );
  AND2_X1 U23435 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20372), .ZN(
        P2_U3194) );
  AND2_X1 U23436 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20372), .ZN(
        P2_U3195) );
  AND2_X1 U23437 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20372), .ZN(
        P2_U3196) );
  AND2_X1 U23438 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20372), .ZN(
        P2_U3197) );
  AND2_X1 U23439 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20372), .ZN(
        P2_U3198) );
  AND2_X1 U23440 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20372), .ZN(
        P2_U3199) );
  AND2_X1 U23441 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20372), .ZN(
        P2_U3200) );
  AND2_X1 U23442 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20372), .ZN(P2_U3201) );
  AND2_X1 U23443 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20372), .ZN(P2_U3202) );
  AND2_X1 U23444 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20372), .ZN(P2_U3203) );
  AND2_X1 U23445 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20372), .ZN(P2_U3204) );
  AND2_X1 U23446 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20372), .ZN(P2_U3205) );
  AND2_X1 U23447 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20372), .ZN(P2_U3206) );
  AND2_X1 U23448 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20372), .ZN(P2_U3207) );
  AND2_X1 U23449 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20372), .ZN(P2_U3208) );
  NOR2_X1 U23450 ( .A1(n20374), .A2(n20373), .ZN(n20386) );
  INV_X1 U23451 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20390) );
  OR3_X1 U23452 ( .A1(n20386), .A2(n20390), .A3(n20389), .ZN(n20376) );
  INV_X1 U23453 ( .A(n20505), .ZN(n20423) );
  AOI211_X1 U23454 ( .C1(n20938), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n20387), .B(n20423), .ZN(n20375) );
  INV_X1 U23455 ( .A(NA), .ZN(n20946) );
  NOR2_X1 U23456 ( .A1(n20946), .A2(n20378), .ZN(n20394) );
  AOI211_X1 U23457 ( .C1(n20395), .C2(n20376), .A(n20375), .B(n20394), .ZN(
        n20377) );
  INV_X1 U23458 ( .A(n20377), .ZN(P2_U3209) );
  AOI21_X1 U23459 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20938), .A(n20395), 
        .ZN(n20383) );
  NOR2_X1 U23460 ( .A1(n20390), .A2(n20383), .ZN(n20379) );
  AOI21_X1 U23461 ( .B1(n20379), .B2(n20378), .A(n20386), .ZN(n20381) );
  OAI211_X1 U23462 ( .C1(n20938), .C2(n20382), .A(n20381), .B(n20380), .ZN(
        P2_U3210) );
  AOI21_X1 U23463 ( .B1(n20385), .B2(n20384), .A(n20383), .ZN(n20393) );
  AOI22_X1 U23464 ( .A1(n20390), .A2(n20387), .B1(n20946), .B2(n20386), .ZN(
        n20388) );
  AOI211_X1 U23465 ( .C1(n20390), .C2(n20938), .A(n20389), .B(n20388), .ZN(
        n20391) );
  INV_X1 U23466 ( .A(n20391), .ZN(n20392) );
  OAI21_X1 U23467 ( .B1(n20394), .B2(n20393), .A(n20392), .ZN(P2_U3211) );
  OAI222_X1 U23468 ( .A1(n20444), .A2(n19857), .B1(n20397), .B2(n20494), .C1(
        n20396), .C2(n20445), .ZN(P2_U3212) );
  OAI222_X1 U23469 ( .A1(n20444), .A2(n13356), .B1(n20398), .B2(n20494), .C1(
        n19857), .C2(n20445), .ZN(P2_U3213) );
  OAI222_X1 U23470 ( .A1(n20444), .A2(n20400), .B1(n20399), .B2(n20494), .C1(
        n13356), .C2(n20445), .ZN(P2_U3214) );
  OAI222_X1 U23471 ( .A1(n20444), .A2(n21260), .B1(n20401), .B2(n20494), .C1(
        n20400), .C2(n20445), .ZN(P2_U3215) );
  OAI222_X1 U23472 ( .A1(n20444), .A2(n20403), .B1(n20402), .B2(n20423), .C1(
        n21260), .C2(n20445), .ZN(P2_U3216) );
  OAI222_X1 U23473 ( .A1(n20444), .A2(n20405), .B1(n20404), .B2(n20494), .C1(
        n20403), .C2(n20445), .ZN(P2_U3217) );
  INV_X1 U23474 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20407) );
  OAI222_X1 U23475 ( .A1(n20444), .A2(n20407), .B1(n20406), .B2(n20494), .C1(
        n20405), .C2(n20445), .ZN(P2_U3218) );
  OAI222_X1 U23476 ( .A1(n20444), .A2(n20409), .B1(n20408), .B2(n20423), .C1(
        n20407), .C2(n20445), .ZN(P2_U3219) );
  OAI222_X1 U23477 ( .A1(n20444), .A2(n20411), .B1(n20410), .B2(n20423), .C1(
        n20409), .C2(n20445), .ZN(P2_U3220) );
  OAI222_X1 U23478 ( .A1(n20444), .A2(n20412), .B1(n21224), .B2(n20423), .C1(
        n20411), .C2(n20445), .ZN(P2_U3221) );
  OAI222_X1 U23479 ( .A1(n20444), .A2(n20414), .B1(n20413), .B2(n20423), .C1(
        n20412), .C2(n20445), .ZN(P2_U3222) );
  OAI222_X1 U23480 ( .A1(n20444), .A2(n14496), .B1(n20415), .B2(n20423), .C1(
        n20414), .C2(n20445), .ZN(P2_U3223) );
  OAI222_X1 U23481 ( .A1(n20444), .A2(n20417), .B1(n20416), .B2(n20423), .C1(
        n14496), .C2(n20445), .ZN(P2_U3224) );
  OAI222_X1 U23482 ( .A1(n20444), .A2(n16306), .B1(n20418), .B2(n20423), .C1(
        n20417), .C2(n20445), .ZN(P2_U3225) );
  OAI222_X1 U23483 ( .A1(n20444), .A2(n21255), .B1(n21122), .B2(n20423), .C1(
        n16306), .C2(n20445), .ZN(P2_U3226) );
  OAI222_X1 U23484 ( .A1(n20444), .A2(n20420), .B1(n20419), .B2(n20423), .C1(
        n21255), .C2(n20445), .ZN(P2_U3227) );
  INV_X1 U23485 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20422) );
  OAI222_X1 U23486 ( .A1(n20444), .A2(n20422), .B1(n20421), .B2(n20423), .C1(
        n20420), .C2(n20445), .ZN(P2_U3228) );
  OAI222_X1 U23487 ( .A1(n20444), .A2(n20425), .B1(n20424), .B2(n20423), .C1(
        n20422), .C2(n20445), .ZN(P2_U3229) );
  OAI222_X1 U23488 ( .A1(n20444), .A2(n20427), .B1(n20426), .B2(n20494), .C1(
        n20425), .C2(n20445), .ZN(P2_U3230) );
  OAI222_X1 U23489 ( .A1(n20444), .A2(n20429), .B1(n20428), .B2(n20494), .C1(
        n20427), .C2(n20445), .ZN(P2_U3231) );
  OAI222_X1 U23490 ( .A1(n20444), .A2(n16220), .B1(n20430), .B2(n20494), .C1(
        n20429), .C2(n20445), .ZN(P2_U3232) );
  OAI222_X1 U23491 ( .A1(n20444), .A2(n20432), .B1(n20431), .B2(n20494), .C1(
        n16220), .C2(n20445), .ZN(P2_U3233) );
  OAI222_X1 U23492 ( .A1(n20444), .A2(n15954), .B1(n20433), .B2(n20494), .C1(
        n20432), .C2(n20445), .ZN(P2_U3234) );
  OAI222_X1 U23493 ( .A1(n20444), .A2(n21294), .B1(n20434), .B2(n20494), .C1(
        n15954), .C2(n20445), .ZN(P2_U3235) );
  OAI222_X1 U23494 ( .A1(n20444), .A2(n20436), .B1(n20435), .B2(n20494), .C1(
        n21294), .C2(n20445), .ZN(P2_U3236) );
  INV_X1 U23495 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20439) );
  OAI222_X1 U23496 ( .A1(n20444), .A2(n20439), .B1(n20437), .B2(n20494), .C1(
        n20436), .C2(n20445), .ZN(P2_U3237) );
  INV_X1 U23497 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20440) );
  OAI222_X1 U23498 ( .A1(n20445), .A2(n20439), .B1(n20438), .B2(n20494), .C1(
        n20440), .C2(n20444), .ZN(P2_U3238) );
  OAI222_X1 U23499 ( .A1(n20444), .A2(n20442), .B1(n20441), .B2(n20494), .C1(
        n20440), .C2(n20445), .ZN(P2_U3239) );
  OAI222_X1 U23500 ( .A1(n20444), .A2(n11406), .B1(n20443), .B2(n20494), .C1(
        n20442), .C2(n20445), .ZN(P2_U3240) );
  OAI222_X1 U23501 ( .A1(n20444), .A2(n16888), .B1(n20446), .B2(n20494), .C1(
        n11406), .C2(n20445), .ZN(P2_U3241) );
  OAI22_X1 U23502 ( .A1(n20505), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20494), .ZN(n20447) );
  INV_X1 U23503 ( .A(n20447), .ZN(P2_U3585) );
  AOI22_X1 U23504 ( .A1(n20494), .A2(n20448), .B1(n21240), .B2(n20505), .ZN(
        P2_U3586) );
  OAI22_X1 U23505 ( .A1(n20505), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20494), .ZN(n20449) );
  INV_X1 U23506 ( .A(n20449), .ZN(P2_U3587) );
  OAI22_X1 U23507 ( .A1(n20505), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20494), .ZN(n20450) );
  INV_X1 U23508 ( .A(n20450), .ZN(P2_U3588) );
  OAI21_X1 U23509 ( .B1(n20453), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20452), 
        .ZN(n20451) );
  INV_X1 U23510 ( .A(n20451), .ZN(P2_U3591) );
  OAI21_X1 U23511 ( .B1(n20453), .B2(n21188), .A(n20452), .ZN(P2_U3592) );
  INV_X1 U23512 ( .A(n20491), .ZN(n20490) );
  NAND2_X1 U23513 ( .A1(n20454), .A2(n20471), .ZN(n20464) );
  NAND3_X1 U23514 ( .A1(n20478), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20455), 
        .ZN(n20456) );
  NAND2_X1 U23515 ( .A1(n20456), .A2(n20482), .ZN(n20465) );
  NAND2_X1 U23516 ( .A1(n20464), .A2(n20465), .ZN(n20461) );
  AOI222_X1 U23517 ( .A1(n20461), .A2(n20460), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20459), .C1(n20458), .C2(n20457), .ZN(n20462) );
  AOI22_X1 U23518 ( .A1(n20490), .A2(n20463), .B1(n20462), .B2(n20491), .ZN(
        P2_U3602) );
  OAI21_X1 U23519 ( .B1(n20466), .B2(n20465), .A(n20464), .ZN(n20467) );
  AOI21_X1 U23520 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20468), .A(n20467), 
        .ZN(n20469) );
  AOI22_X1 U23521 ( .A1(n20490), .A2(n20470), .B1(n20469), .B2(n20491), .ZN(
        P2_U3603) );
  INV_X1 U23522 ( .A(n20471), .ZN(n20477) );
  INV_X1 U23523 ( .A(n20472), .ZN(n20473) );
  NAND3_X1 U23524 ( .A1(n20478), .A2(n20482), .A3(n20473), .ZN(n20476) );
  NAND2_X1 U23525 ( .A1(n20474), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20475) );
  OAI211_X1 U23526 ( .C1(n20478), .C2(n20477), .A(n20476), .B(n20475), .ZN(
        n20479) );
  INV_X1 U23527 ( .A(n20479), .ZN(n20480) );
  AOI22_X1 U23528 ( .A1(n20490), .A2(n20481), .B1(n20480), .B2(n20491), .ZN(
        P2_U3604) );
  INV_X1 U23529 ( .A(n20482), .ZN(n20486) );
  INV_X1 U23530 ( .A(n20483), .ZN(n20485) );
  OAI22_X1 U23531 ( .A1(n20487), .A2(n20486), .B1(n20485), .B2(n20484), .ZN(
        n20488) );
  AOI21_X1 U23532 ( .B1(n20492), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20488), 
        .ZN(n20489) );
  OAI22_X1 U23533 ( .A1(n20492), .A2(n20491), .B1(n20490), .B2(n20489), .ZN(
        P2_U3605) );
  AOI22_X1 U23534 ( .A1(n20494), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20493), 
        .B2(n20505), .ZN(P2_U3608) );
  INV_X1 U23535 ( .A(n20495), .ZN(n20501) );
  INV_X1 U23536 ( .A(n20496), .ZN(n20497) );
  OR2_X1 U23537 ( .A1(n20498), .A2(n20497), .ZN(n20499) );
  OAI211_X1 U23538 ( .C1(n20502), .C2(n20501), .A(n20500), .B(n20499), .ZN(
        n20504) );
  MUX2_X1 U23539 ( .A(P2_MORE_REG_SCAN_IN), .B(n20504), .S(n20503), .Z(
        P2_U3609) );
  MUX2_X1 U23540 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .B(P2_M_IO_N_REG_SCAN_IN), 
        .S(n20505), .Z(P2_U3611) );
  AND2_X1 U23541 ( .A1(n20942), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n20507) );
  INV_X1 U23542 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20506) );
  INV_X1 U23543 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20944) );
  NAND2_X1 U23544 ( .A1(n20944), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21024) );
  INV_X1 U23545 ( .A(n21024), .ZN(n21025) );
  AOI21_X1 U23546 ( .B1(n20507), .B2(n20506), .A(n21025), .ZN(P1_U2802) );
  OAI21_X1 U23547 ( .B1(n20509), .B2(n20508), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20510) );
  OAI21_X1 U23548 ( .B1(n20511), .B2(n9922), .A(n20510), .ZN(P1_U2803) );
  NOR2_X1 U23549 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20513) );
  INV_X1 U23550 ( .A(n21025), .ZN(n21038) );
  OAI21_X1 U23551 ( .B1(n20513), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21038), .ZN(
        n20512) );
  OAI21_X1 U23552 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21024), .A(n20512), 
        .ZN(P1_U2804) );
  AOI21_X1 U23553 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20942), .A(n21025), 
        .ZN(n21002) );
  OAI21_X1 U23554 ( .B1(BS16), .B2(n20513), .A(n21002), .ZN(n21000) );
  OAI21_X1 U23555 ( .B1(n21002), .B2(n20514), .A(n21000), .ZN(P1_U2805) );
  INV_X1 U23556 ( .A(n20515), .ZN(n20518) );
  OAI21_X1 U23557 ( .B1(n20518), .B2(n20517), .A(n20516), .ZN(P1_U2806) );
  NOR2_X1 U23558 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n21289) );
  AOI211_X1 U23559 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_3__SCAN_IN), .B(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20519) );
  INV_X1 U23560 ( .A(P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20937) );
  INV_X1 U23561 ( .A(P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n21119) );
  NAND4_X1 U23562 ( .A1(n21289), .A2(n20519), .A3(n20937), .A4(n21119), .ZN(
        n20527) );
  OR4_X1 U23563 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20526) );
  OR4_X1 U23564 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20525) );
  NOR4_X1 U23565 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20523) );
  NOR4_X1 U23566 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_14__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20522) );
  NOR4_X1 U23567 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20521) );
  NOR4_X1 U23568 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20520) );
  NAND4_X1 U23569 ( .A1(n20523), .A2(n20522), .A3(n20521), .A4(n20520), .ZN(
        n20524) );
  INV_X1 U23570 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20529) );
  NOR3_X1 U23571 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20530) );
  OAI21_X1 U23572 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20530), .A(n21020), .ZN(
        n20528) );
  OAI21_X1 U23573 ( .B1(n21020), .B2(n20529), .A(n20528), .ZN(P1_U2807) );
  INV_X1 U23574 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21001) );
  AOI21_X1 U23575 ( .B1(n21016), .B2(n21001), .A(n20530), .ZN(n20532) );
  INV_X1 U23576 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20531) );
  INV_X1 U23577 ( .A(n21020), .ZN(n21022) );
  AOI22_X1 U23578 ( .A1(n21020), .A2(n20532), .B1(n20531), .B2(n21022), .ZN(
        P1_U2808) );
  INV_X1 U23579 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20534) );
  AOI22_X1 U23580 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n20602), .B1(n20595), .B2(
        n21039), .ZN(n20533) );
  OAI211_X1 U23581 ( .C1(n20581), .C2(n20534), .A(n20533), .B(n16808), .ZN(
        n20535) );
  AOI21_X1 U23582 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n20536), .A(n20535), .ZN(
        n20539) );
  AOI22_X1 U23583 ( .A1(n21043), .A2(n20554), .B1(n20604), .B2(n20537), .ZN(
        n20538) );
  OAI211_X1 U23584 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n20540), .A(n20539), .B(
        n20538), .ZN(P1_U2831) );
  NOR3_X1 U23585 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20578), .A3(n20544), .ZN(
        n20543) );
  AOI21_X1 U23586 ( .B1(n20593), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n13116), .ZN(n20541) );
  INV_X1 U23587 ( .A(n20541), .ZN(n20542) );
  AOI211_X1 U23588 ( .C1(n20602), .C2(P1_EBX_REG_7__SCAN_IN), .A(n20543), .B(
        n20542), .ZN(n20549) );
  AOI21_X1 U23589 ( .B1(n20596), .B2(n20544), .A(n20565), .ZN(n20552) );
  OAI22_X1 U23590 ( .A1(n20552), .A2(n20962), .B1(n20545), .B2(n20583), .ZN(
        n20546) );
  AOI21_X1 U23591 ( .B1(n20547), .B2(n20554), .A(n20546), .ZN(n20548) );
  OAI211_X1 U23592 ( .C1(n20580), .C2(n20550), .A(n20549), .B(n20548), .ZN(
        P1_U2833) );
  AOI21_X1 U23593 ( .B1(n20593), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13116), .ZN(n20558) );
  AOI22_X1 U23594 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n20602), .B1(n20595), .B2(
        n9813), .ZN(n20557) );
  INV_X1 U23595 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20959) );
  OAI22_X1 U23596 ( .A1(n20552), .A2(n20959), .B1(n20551), .B2(n20583), .ZN(
        n20553) );
  AOI21_X1 U23597 ( .B1(n20611), .B2(n20554), .A(n20553), .ZN(n20556) );
  NAND4_X1 U23598 ( .A1(n20596), .A2(P1_REIP_REG_5__SCAN_IN), .A3(n20564), 
        .A4(n20959), .ZN(n20555) );
  NAND4_X1 U23599 ( .A1(n20558), .A2(n20557), .A3(n20556), .A4(n20555), .ZN(
        P1_U2834) );
  OAI21_X1 U23600 ( .B1(n20581), .B2(n20559), .A(n16808), .ZN(n20563) );
  NAND2_X1 U23601 ( .A1(n20596), .A2(n20564), .ZN(n20561) );
  OAI22_X1 U23602 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20561), .B1(n20580), 
        .B2(n20560), .ZN(n20562) );
  AOI211_X1 U23603 ( .C1(P1_EBX_REG_5__SCAN_IN), .C2(n20602), .A(n20563), .B(
        n20562), .ZN(n20571) );
  INV_X1 U23604 ( .A(n20564), .ZN(n20566) );
  AOI21_X1 U23605 ( .B1(n20596), .B2(n20566), .A(n20565), .ZN(n20573) );
  INV_X1 U23606 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20567) );
  OAI22_X1 U23607 ( .A1(n20568), .A2(n20585), .B1(n20573), .B2(n20567), .ZN(
        n20569) );
  INV_X1 U23608 ( .A(n20569), .ZN(n20570) );
  OAI211_X1 U23609 ( .C1(n20572), .C2(n20583), .A(n20571), .B(n20570), .ZN(
        P1_U2835) );
  INV_X1 U23610 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21095) );
  INV_X1 U23611 ( .A(n20573), .ZN(n20576) );
  AOI22_X1 U23612 ( .A1(n20576), .A2(P1_REIP_REG_4__SCAN_IN), .B1(n20575), 
        .B2(n20574), .ZN(n20591) );
  NOR3_X1 U23613 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20578), .A3(n20577), .ZN(
        n20589) );
  OAI22_X1 U23614 ( .A1(n20582), .A2(n20581), .B1(n20580), .B2(n20579), .ZN(
        n20588) );
  OAI22_X1 U23615 ( .A1(n20586), .A2(n20585), .B1(n20584), .B2(n20583), .ZN(
        n20587) );
  NOR4_X1 U23616 ( .A1(n13116), .A2(n20589), .A3(n20588), .A4(n20587), .ZN(
        n20590) );
  OAI211_X1 U23617 ( .C1(n21095), .C2(n20592), .A(n20591), .B(n20590), .ZN(
        P1_U2836) );
  AOI22_X1 U23618 ( .A1(n20595), .A2(n20594), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20593), .ZN(n20598) );
  NAND4_X1 U23619 ( .A1(n20596), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .A4(n20955), .ZN(n20597) );
  OAI211_X1 U23620 ( .C1(n20600), .C2(n20599), .A(n20598), .B(n20597), .ZN(
        n20601) );
  AOI21_X1 U23621 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(n20602), .A(n20601), .ZN(
        n20609) );
  INV_X1 U23622 ( .A(n20603), .ZN(n20605) );
  AOI22_X1 U23623 ( .A1(n20607), .A2(n20606), .B1(n20605), .B2(n20604), .ZN(
        n20608) );
  OAI211_X1 U23624 ( .C1(n20610), .C2(n20955), .A(n20609), .B(n20608), .ZN(
        P1_U2837) );
  AOI22_X1 U23625 ( .A1(n20611), .A2(n21042), .B1(n21040), .B2(n9813), .ZN(
        n20612) );
  OAI21_X1 U23626 ( .B1(n20618), .B2(n21295), .A(n20612), .ZN(P1_U2866) );
  INV_X1 U23627 ( .A(n20613), .ZN(n20615) );
  AOI22_X1 U23628 ( .A1(n20615), .A2(n21042), .B1(n21040), .B2(n20614), .ZN(
        n20616) );
  OAI21_X1 U23629 ( .B1(n20618), .B2(n20617), .A(n20616), .ZN(P1_U2871) );
  AOI22_X1 U23630 ( .A1(n21029), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20620) );
  OAI21_X1 U23631 ( .B1(n20621), .B2(n20649), .A(n20620), .ZN(P1_U2921) );
  AOI22_X1 U23632 ( .A1(n21029), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20622) );
  OAI21_X1 U23633 ( .B1(n21179), .B2(n20649), .A(n20622), .ZN(P1_U2922) );
  AOI22_X1 U23634 ( .A1(n21029), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20623) );
  OAI21_X1 U23635 ( .B1(n20624), .B2(n20649), .A(n20623), .ZN(P1_U2923) );
  AOI22_X1 U23636 ( .A1(n21029), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20644), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20625) );
  OAI21_X1 U23637 ( .B1(n20626), .B2(n20649), .A(n20625), .ZN(P1_U2924) );
  AOI22_X1 U23638 ( .A1(n21029), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20627) );
  OAI21_X1 U23639 ( .B1(n20628), .B2(n20649), .A(n20627), .ZN(P1_U2925) );
  AOI22_X1 U23640 ( .A1(n21029), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20629) );
  OAI21_X1 U23641 ( .B1(n20630), .B2(n20649), .A(n20629), .ZN(P1_U2926) );
  AOI22_X1 U23642 ( .A1(n21029), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20631) );
  OAI21_X1 U23643 ( .B1(n20632), .B2(n20649), .A(n20631), .ZN(P1_U2927) );
  AOI22_X1 U23644 ( .A1(n21029), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20633) );
  OAI21_X1 U23645 ( .B1(n20634), .B2(n20649), .A(n20633), .ZN(P1_U2928) );
  AOI22_X1 U23646 ( .A1(n21029), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20635) );
  OAI21_X1 U23647 ( .B1(n14122), .B2(n20649), .A(n20635), .ZN(P1_U2929) );
  AOI22_X1 U23648 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20644), .B1(n20647), 
        .B2(P1_LWORD_REG_6__SCAN_IN), .ZN(n20636) );
  OAI21_X1 U23649 ( .B1(n13977), .B2(n20649), .A(n20636), .ZN(P1_U2930) );
  INV_X1 U23650 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20638) );
  AOI22_X1 U23651 ( .A1(n21029), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20637) );
  OAI21_X1 U23652 ( .B1(n20638), .B2(n20649), .A(n20637), .ZN(P1_U2931) );
  AOI22_X1 U23653 ( .A1(n21029), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20639) );
  OAI21_X1 U23654 ( .B1(n21197), .B2(n20649), .A(n20639), .ZN(P1_U2932) );
  AOI22_X1 U23655 ( .A1(n21029), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20646), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20640) );
  OAI21_X1 U23656 ( .B1(n20641), .B2(n20649), .A(n20640), .ZN(P1_U2933) );
  AOI22_X1 U23657 ( .A1(n21029), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20644), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20642) );
  OAI21_X1 U23658 ( .B1(n20643), .B2(n20649), .A(n20642), .ZN(P1_U2934) );
  AOI22_X1 U23659 ( .A1(n21029), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20644), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20645) );
  OAI21_X1 U23660 ( .B1(n21256), .B2(n20649), .A(n20645), .ZN(P1_U2935) );
  AOI22_X1 U23661 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20647), .B1(n20646), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20648) );
  OAI21_X1 U23662 ( .B1(n20650), .B2(n20649), .A(n20648), .ZN(P1_U2936) );
  OAI22_X1 U23663 ( .A1(n20654), .A2(n20653), .B1(n20652), .B2(n20651), .ZN(
        n20655) );
  INV_X1 U23664 ( .A(n20655), .ZN(n20662) );
  OAI22_X1 U23665 ( .A1(n20658), .A2(n20657), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20656), .ZN(n20659) );
  NAND4_X1 U23666 ( .A1(n20662), .A2(n20661), .A3(n20660), .A4(n20659), .ZN(
        P1_U3031) );
  AND2_X1 U23667 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20663), .ZN(
        P1_U3032) );
  NOR3_X1 U23668 ( .A1(n20689), .A2(n20688), .A3(n20807), .ZN(n20664) );
  NOR2_X1 U23669 ( .A1(n20807), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20808) );
  NOR2_X1 U23670 ( .A1(n20664), .A2(n20808), .ZN(n20672) );
  INV_X1 U23671 ( .A(n20672), .ZN(n20666) );
  NOR2_X1 U23672 ( .A1(n20736), .A2(n20868), .ZN(n20671) );
  NAND2_X1 U23673 ( .A1(n20779), .A2(n20667), .ZN(n20668) );
  INV_X1 U23674 ( .A(n20668), .ZN(n20687) );
  AOI22_X1 U23675 ( .A1(n20688), .A2(n20882), .B1(n20874), .B2(n20687), .ZN(
        n20674) );
  AOI22_X1 U23676 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20669), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20668), .ZN(n20670) );
  OAI211_X1 U23677 ( .C1(n20672), .C2(n20671), .A(n20700), .B(n20670), .ZN(
        n20690) );
  AOI22_X1 U23678 ( .A1(n20690), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n20875), .B2(n20689), .ZN(n20673) );
  OAI211_X1 U23679 ( .C1(n20693), .C2(n20885), .A(n20674), .B(n20673), .ZN(
        P1_U3033) );
  AOI22_X1 U23680 ( .A1(n20688), .A2(n20888), .B1(n20886), .B2(n20687), .ZN(
        n20676) );
  AOI22_X1 U23681 ( .A1(n20690), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n20887), .B2(n20689), .ZN(n20675) );
  OAI211_X1 U23682 ( .C1(n20693), .C2(n20891), .A(n20676), .B(n20675), .ZN(
        P1_U3034) );
  AOI22_X1 U23683 ( .A1(n20688), .A2(n20894), .B1(n20892), .B2(n20687), .ZN(
        n20678) );
  AOI22_X1 U23684 ( .A1(n20690), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n20893), .B2(n20689), .ZN(n20677) );
  OAI211_X1 U23685 ( .C1(n20693), .C2(n20897), .A(n20678), .B(n20677), .ZN(
        P1_U3035) );
  AOI22_X1 U23686 ( .A1(n20688), .A2(n20900), .B1(n20898), .B2(n20687), .ZN(
        n20680) );
  AOI22_X1 U23687 ( .A1(n20690), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n20899), .B2(n20689), .ZN(n20679) );
  OAI211_X1 U23688 ( .C1(n20693), .C2(n20903), .A(n20680), .B(n20679), .ZN(
        P1_U3036) );
  AOI22_X1 U23689 ( .A1(n20688), .A2(n20906), .B1(n20904), .B2(n20687), .ZN(
        n20682) );
  AOI22_X1 U23690 ( .A1(n20690), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n20905), .B2(n20689), .ZN(n20681) );
  OAI211_X1 U23691 ( .C1(n20693), .C2(n20909), .A(n20682), .B(n20681), .ZN(
        P1_U3037) );
  AOI22_X1 U23692 ( .A1(n20688), .A2(n20912), .B1(n20910), .B2(n20687), .ZN(
        n20684) );
  AOI22_X1 U23693 ( .A1(n20690), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n20911), .B2(n20689), .ZN(n20683) );
  OAI211_X1 U23694 ( .C1(n20693), .C2(n20915), .A(n20684), .B(n20683), .ZN(
        P1_U3038) );
  AOI22_X1 U23695 ( .A1(n20688), .A2(n20918), .B1(n20916), .B2(n20687), .ZN(
        n20686) );
  AOI22_X1 U23696 ( .A1(n20690), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n20917), .B2(n20689), .ZN(n20685) );
  OAI211_X1 U23697 ( .C1(n20693), .C2(n20921), .A(n20686), .B(n20685), .ZN(
        P1_U3039) );
  AOI22_X1 U23698 ( .A1(n20688), .A2(n20927), .B1(n20923), .B2(n20687), .ZN(
        n20692) );
  AOI22_X1 U23699 ( .A1(n20690), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n20924), .B2(n20689), .ZN(n20691) );
  OAI211_X1 U23700 ( .C1(n20693), .C2(n20931), .A(n20692), .B(n20691), .ZN(
        P1_U3040) );
  NOR2_X1 U23701 ( .A1(n20770), .A2(n20807), .ZN(n20696) );
  AOI21_X1 U23702 ( .B1(n20696), .B2(n20727), .A(n20808), .ZN(n20705) );
  INV_X1 U23703 ( .A(n20705), .ZN(n20697) );
  NOR2_X1 U23704 ( .A1(n20736), .A2(n13840), .ZN(n20704) );
  NOR2_X1 U23705 ( .A1(n20701), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20777) );
  NOR3_X1 U23706 ( .A1(n20698), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20742) );
  NAND2_X1 U23707 ( .A1(n20779), .A2(n20742), .ZN(n20726) );
  OAI22_X1 U23708 ( .A1(n20727), .A2(n20816), .B1(n20815), .B2(n20726), .ZN(
        n20699) );
  INV_X1 U23709 ( .A(n20699), .ZN(n20707) );
  INV_X1 U23710 ( .A(n20700), .ZN(n20819) );
  OAI21_X1 U23711 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20701), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20702) );
  INV_X1 U23712 ( .A(n20702), .ZN(n20780) );
  AOI211_X1 U23713 ( .C1(n20726), .C2(P1_STATE2_REG_3__SCAN_IN), .A(n20819), 
        .B(n20780), .ZN(n20703) );
  AOI22_X1 U23714 ( .A1(n20729), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n20875), .B2(n20770), .ZN(n20706) );
  OAI211_X1 U23715 ( .C1(n20732), .C2(n20885), .A(n20707), .B(n20706), .ZN(
        P1_U3049) );
  OAI22_X1 U23716 ( .A1(n20727), .A2(n20827), .B1(n20826), .B2(n20726), .ZN(
        n20708) );
  INV_X1 U23717 ( .A(n20708), .ZN(n20710) );
  AOI22_X1 U23718 ( .A1(n20729), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n20887), .B2(n20770), .ZN(n20709) );
  OAI211_X1 U23719 ( .C1(n20732), .C2(n20891), .A(n20710), .B(n20709), .ZN(
        P1_U3050) );
  OAI22_X1 U23720 ( .A1(n20727), .A2(n20832), .B1(n20831), .B2(n20726), .ZN(
        n20711) );
  INV_X1 U23721 ( .A(n20711), .ZN(n20713) );
  AOI22_X1 U23722 ( .A1(n20729), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n20893), .B2(n20770), .ZN(n20712) );
  OAI211_X1 U23723 ( .C1(n20732), .C2(n20897), .A(n20713), .B(n20712), .ZN(
        P1_U3051) );
  OAI22_X1 U23724 ( .A1(n20727), .A2(n20837), .B1(n20836), .B2(n20726), .ZN(
        n20714) );
  INV_X1 U23725 ( .A(n20714), .ZN(n20716) );
  AOI22_X1 U23726 ( .A1(n20729), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n20899), .B2(n20770), .ZN(n20715) );
  OAI211_X1 U23727 ( .C1(n20732), .C2(n20903), .A(n20716), .B(n20715), .ZN(
        P1_U3052) );
  OAI22_X1 U23728 ( .A1(n20727), .A2(n20842), .B1(n20841), .B2(n20726), .ZN(
        n20717) );
  INV_X1 U23729 ( .A(n20717), .ZN(n20719) );
  AOI22_X1 U23730 ( .A1(n20729), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n20905), .B2(n20770), .ZN(n20718) );
  OAI211_X1 U23731 ( .C1(n20732), .C2(n20909), .A(n20719), .B(n20718), .ZN(
        P1_U3053) );
  OAI22_X1 U23732 ( .A1(n20727), .A2(n20847), .B1(n20846), .B2(n20726), .ZN(
        n20720) );
  INV_X1 U23733 ( .A(n20720), .ZN(n20722) );
  AOI22_X1 U23734 ( .A1(n20729), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n20911), .B2(n20770), .ZN(n20721) );
  OAI211_X1 U23735 ( .C1(n20732), .C2(n20915), .A(n20722), .B(n20721), .ZN(
        P1_U3054) );
  OAI22_X1 U23736 ( .A1(n20727), .A2(n20852), .B1(n20851), .B2(n20726), .ZN(
        n20723) );
  INV_X1 U23737 ( .A(n20723), .ZN(n20725) );
  AOI22_X1 U23738 ( .A1(n20729), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n20917), .B2(n20770), .ZN(n20724) );
  OAI211_X1 U23739 ( .C1(n20732), .C2(n20921), .A(n20725), .B(n20724), .ZN(
        P1_U3055) );
  OAI22_X1 U23740 ( .A1(n20727), .A2(n20858), .B1(n20857), .B2(n20726), .ZN(
        n20728) );
  INV_X1 U23741 ( .A(n20728), .ZN(n20731) );
  AOI22_X1 U23742 ( .A1(n20729), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n20924), .B2(n20770), .ZN(n20730) );
  OAI211_X1 U23743 ( .C1(n20732), .C2(n20931), .A(n20731), .B(n20730), .ZN(
        P1_U3056) );
  AOI21_X1 U23744 ( .B1(n20734), .B2(n20733), .A(n20807), .ZN(n20741) );
  OR2_X1 U23745 ( .A1(n20736), .A2(n20735), .ZN(n20739) );
  NAND2_X1 U23746 ( .A1(n20738), .A2(n20737), .ZN(n20767) );
  NAND2_X1 U23747 ( .A1(n20739), .A2(n20767), .ZN(n20745) );
  NOR2_X1 U23748 ( .A1(n20815), .A2(n20767), .ZN(n20740) );
  AOI21_X1 U23749 ( .B1(n20769), .B2(n20875), .A(n20740), .ZN(n20748) );
  INV_X1 U23750 ( .A(n20741), .ZN(n20746) );
  OR2_X1 U23751 ( .A1(n20866), .A2(n20742), .ZN(n20743) );
  OAI211_X1 U23752 ( .C1(n20746), .C2(n20745), .A(n20744), .B(n20743), .ZN(
        n20771) );
  AOI22_X1 U23753 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n20882), .B2(n20770), .ZN(n20747) );
  OAI211_X1 U23754 ( .C1(n20774), .C2(n20885), .A(n20748), .B(n20747), .ZN(
        P1_U3057) );
  NOR2_X1 U23755 ( .A1(n20826), .A2(n20767), .ZN(n20749) );
  AOI21_X1 U23756 ( .B1(n20769), .B2(n20887), .A(n20749), .ZN(n20751) );
  AOI22_X1 U23757 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n20888), .B2(n20770), .ZN(n20750) );
  OAI211_X1 U23758 ( .C1(n20774), .C2(n20891), .A(n20751), .B(n20750), .ZN(
        P1_U3058) );
  NOR2_X1 U23759 ( .A1(n20831), .A2(n20767), .ZN(n20752) );
  AOI21_X1 U23760 ( .B1(n20769), .B2(n20893), .A(n20752), .ZN(n20754) );
  AOI22_X1 U23761 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n20894), .B2(n20770), .ZN(n20753) );
  OAI211_X1 U23762 ( .C1(n20774), .C2(n20897), .A(n20754), .B(n20753), .ZN(
        P1_U3059) );
  NOR2_X1 U23763 ( .A1(n20836), .A2(n20767), .ZN(n20755) );
  AOI21_X1 U23764 ( .B1(n20770), .B2(n20900), .A(n20755), .ZN(n20757) );
  AOI22_X1 U23765 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n20769), .B2(n20899), .ZN(n20756) );
  OAI211_X1 U23766 ( .C1(n20774), .C2(n20903), .A(n20757), .B(n20756), .ZN(
        P1_U3060) );
  NOR2_X1 U23767 ( .A1(n20841), .A2(n20767), .ZN(n20758) );
  AOI21_X1 U23768 ( .B1(n20770), .B2(n20906), .A(n20758), .ZN(n20760) );
  AOI22_X1 U23769 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n20769), .B2(n20905), .ZN(n20759) );
  OAI211_X1 U23770 ( .C1(n20774), .C2(n20909), .A(n20760), .B(n20759), .ZN(
        P1_U3061) );
  NOR2_X1 U23771 ( .A1(n20846), .A2(n20767), .ZN(n20761) );
  AOI21_X1 U23772 ( .B1(n20770), .B2(n20912), .A(n20761), .ZN(n20763) );
  AOI22_X1 U23773 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n20769), .B2(n20911), .ZN(n20762) );
  OAI211_X1 U23774 ( .C1(n20774), .C2(n20915), .A(n20763), .B(n20762), .ZN(
        P1_U3062) );
  NOR2_X1 U23775 ( .A1(n20851), .A2(n20767), .ZN(n20764) );
  AOI21_X1 U23776 ( .B1(n20769), .B2(n20917), .A(n20764), .ZN(n20766) );
  AOI22_X1 U23777 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n20918), .B2(n20770), .ZN(n20765) );
  OAI211_X1 U23778 ( .C1(n20774), .C2(n20921), .A(n20766), .B(n20765), .ZN(
        P1_U3063) );
  NOR2_X1 U23779 ( .A1(n20857), .A2(n20767), .ZN(n20768) );
  AOI21_X1 U23780 ( .B1(n20769), .B2(n20924), .A(n20768), .ZN(n20773) );
  AOI22_X1 U23781 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n20927), .B2(n20770), .ZN(n20772) );
  OAI211_X1 U23782 ( .C1(n20774), .C2(n20931), .A(n20773), .B(n20772), .ZN(
        P1_U3064) );
  NOR3_X1 U23783 ( .A1(n20801), .A2(n20802), .A3(n20807), .ZN(n20775) );
  NOR2_X1 U23784 ( .A1(n20775), .A2(n20808), .ZN(n20785) );
  INV_X1 U23785 ( .A(n20785), .ZN(n20778) );
  AND2_X1 U23786 ( .A1(n20776), .A2(n20868), .ZN(n20784) );
  NAND2_X1 U23787 ( .A1(n20779), .A2(n10340), .ZN(n20782) );
  INV_X1 U23788 ( .A(n20782), .ZN(n20800) );
  AOI22_X1 U23789 ( .A1(n20801), .A2(n20882), .B1(n20874), .B2(n20800), .ZN(
        n20787) );
  INV_X1 U23790 ( .A(n20876), .ZN(n20781) );
  AOI211_X1 U23791 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20782), .A(n20781), 
        .B(n20780), .ZN(n20783) );
  AOI22_X1 U23792 ( .A1(n20803), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n20875), .B2(n20802), .ZN(n20786) );
  OAI211_X1 U23793 ( .C1(n20806), .C2(n20885), .A(n20787), .B(n20786), .ZN(
        P1_U3081) );
  AOI22_X1 U23794 ( .A1(n20801), .A2(n20888), .B1(n20886), .B2(n20800), .ZN(
        n20789) );
  AOI22_X1 U23795 ( .A1(n20803), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n20887), .B2(n20802), .ZN(n20788) );
  OAI211_X1 U23796 ( .C1(n20806), .C2(n20891), .A(n20789), .B(n20788), .ZN(
        P1_U3082) );
  AOI22_X1 U23797 ( .A1(n20801), .A2(n20894), .B1(n20892), .B2(n20800), .ZN(
        n20791) );
  AOI22_X1 U23798 ( .A1(n20803), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n20893), .B2(n20802), .ZN(n20790) );
  OAI211_X1 U23799 ( .C1(n20806), .C2(n20897), .A(n20791), .B(n20790), .ZN(
        P1_U3083) );
  AOI22_X1 U23800 ( .A1(n20801), .A2(n20900), .B1(n20898), .B2(n20800), .ZN(
        n20793) );
  AOI22_X1 U23801 ( .A1(n20803), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n20899), .B2(n20802), .ZN(n20792) );
  OAI211_X1 U23802 ( .C1(n20806), .C2(n20903), .A(n20793), .B(n20792), .ZN(
        P1_U3084) );
  AOI22_X1 U23803 ( .A1(n20801), .A2(n20906), .B1(n20904), .B2(n20800), .ZN(
        n20795) );
  AOI22_X1 U23804 ( .A1(n20803), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n20905), .B2(n20802), .ZN(n20794) );
  OAI211_X1 U23805 ( .C1(n20806), .C2(n20909), .A(n20795), .B(n20794), .ZN(
        P1_U3085) );
  AOI22_X1 U23806 ( .A1(n20801), .A2(n20912), .B1(n20910), .B2(n20800), .ZN(
        n20797) );
  AOI22_X1 U23807 ( .A1(n20803), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n20911), .B2(n20802), .ZN(n20796) );
  OAI211_X1 U23808 ( .C1(n20806), .C2(n20915), .A(n20797), .B(n20796), .ZN(
        P1_U3086) );
  AOI22_X1 U23809 ( .A1(n20801), .A2(n20918), .B1(n20916), .B2(n20800), .ZN(
        n20799) );
  AOI22_X1 U23810 ( .A1(n20803), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n20917), .B2(n20802), .ZN(n20798) );
  OAI211_X1 U23811 ( .C1(n20806), .C2(n20921), .A(n20799), .B(n20798), .ZN(
        P1_U3087) );
  AOI22_X1 U23812 ( .A1(n20801), .A2(n20927), .B1(n20923), .B2(n20800), .ZN(
        n20805) );
  AOI22_X1 U23813 ( .A1(n20803), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n20924), .B2(n20802), .ZN(n20804) );
  OAI211_X1 U23814 ( .C1(n20806), .C2(n20931), .A(n20805), .B(n20804), .ZN(
        P1_U3088) );
  NOR2_X1 U23815 ( .A1(n20861), .A2(n20807), .ZN(n20809) );
  AOI21_X1 U23816 ( .B1(n20809), .B2(n20859), .A(n20808), .ZN(n20823) );
  INV_X1 U23817 ( .A(n20823), .ZN(n20813) );
  AND2_X1 U23818 ( .A1(n20810), .A2(n20868), .ZN(n20822) );
  OR2_X1 U23819 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20814), .ZN(
        n20856) );
  OAI22_X1 U23820 ( .A1(n20859), .A2(n20816), .B1(n20815), .B2(n20856), .ZN(
        n20817) );
  INV_X1 U23821 ( .A(n20817), .ZN(n20825) );
  INV_X1 U23822 ( .A(n20818), .ZN(n20820) );
  AOI211_X1 U23823 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20856), .A(n20820), 
        .B(n20819), .ZN(n20821) );
  AOI22_X1 U23824 ( .A1(n20862), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n20875), .B2(n20861), .ZN(n20824) );
  OAI211_X1 U23825 ( .C1(n20865), .C2(n20885), .A(n20825), .B(n20824), .ZN(
        P1_U3113) );
  OAI22_X1 U23826 ( .A1(n20859), .A2(n20827), .B1(n20826), .B2(n20856), .ZN(
        n20828) );
  INV_X1 U23827 ( .A(n20828), .ZN(n20830) );
  AOI22_X1 U23828 ( .A1(n20862), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n20887), .B2(n20861), .ZN(n20829) );
  OAI211_X1 U23829 ( .C1(n20865), .C2(n20891), .A(n20830), .B(n20829), .ZN(
        P1_U3114) );
  OAI22_X1 U23830 ( .A1(n20859), .A2(n20832), .B1(n20831), .B2(n20856), .ZN(
        n20833) );
  INV_X1 U23831 ( .A(n20833), .ZN(n20835) );
  AOI22_X1 U23832 ( .A1(n20862), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n20893), .B2(n20861), .ZN(n20834) );
  OAI211_X1 U23833 ( .C1(n20865), .C2(n20897), .A(n20835), .B(n20834), .ZN(
        P1_U3115) );
  OAI22_X1 U23834 ( .A1(n20859), .A2(n20837), .B1(n20836), .B2(n20856), .ZN(
        n20838) );
  INV_X1 U23835 ( .A(n20838), .ZN(n20840) );
  AOI22_X1 U23836 ( .A1(n20862), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n20899), .B2(n20861), .ZN(n20839) );
  OAI211_X1 U23837 ( .C1(n20865), .C2(n20903), .A(n20840), .B(n20839), .ZN(
        P1_U3116) );
  OAI22_X1 U23838 ( .A1(n20859), .A2(n20842), .B1(n20841), .B2(n20856), .ZN(
        n20843) );
  INV_X1 U23839 ( .A(n20843), .ZN(n20845) );
  AOI22_X1 U23840 ( .A1(n20862), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n20905), .B2(n20861), .ZN(n20844) );
  OAI211_X1 U23841 ( .C1(n20865), .C2(n20909), .A(n20845), .B(n20844), .ZN(
        P1_U3117) );
  OAI22_X1 U23842 ( .A1(n20859), .A2(n20847), .B1(n20846), .B2(n20856), .ZN(
        n20848) );
  INV_X1 U23843 ( .A(n20848), .ZN(n20850) );
  AOI22_X1 U23844 ( .A1(n20862), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n20911), .B2(n20861), .ZN(n20849) );
  OAI211_X1 U23845 ( .C1(n20865), .C2(n20915), .A(n20850), .B(n20849), .ZN(
        P1_U3118) );
  OAI22_X1 U23846 ( .A1(n20859), .A2(n20852), .B1(n20851), .B2(n20856), .ZN(
        n20853) );
  INV_X1 U23847 ( .A(n20853), .ZN(n20855) );
  AOI22_X1 U23848 ( .A1(n20862), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n20917), .B2(n20861), .ZN(n20854) );
  OAI211_X1 U23849 ( .C1(n20865), .C2(n20921), .A(n20855), .B(n20854), .ZN(
        P1_U3119) );
  OAI22_X1 U23850 ( .A1(n20859), .A2(n20858), .B1(n20857), .B2(n20856), .ZN(
        n20860) );
  INV_X1 U23851 ( .A(n20860), .ZN(n20864) );
  AOI22_X1 U23852 ( .A1(n20862), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n20924), .B2(n20861), .ZN(n20863) );
  OAI211_X1 U23853 ( .C1(n20865), .C2(n20931), .A(n20864), .B(n20863), .ZN(
        P1_U3120) );
  OAI21_X1 U23854 ( .B1(n20926), .B2(n20925), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20867) );
  NAND2_X1 U23855 ( .A1(n20867), .A2(n20866), .ZN(n20881) );
  INV_X1 U23856 ( .A(n20881), .ZN(n20872) );
  NOR2_X1 U23857 ( .A1(n20869), .A2(n20868), .ZN(n20880) );
  NOR2_X1 U23858 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20873), .ZN(
        n20922) );
  AOI22_X1 U23859 ( .A1(n20925), .A2(n20875), .B1(n20874), .B2(n20922), .ZN(
        n20884) );
  OAI21_X1 U23860 ( .B1(n12826), .B2(n20922), .A(n20876), .ZN(n20877) );
  AOI21_X1 U23861 ( .B1(n20878), .B2(P1_STATE2_REG_2__SCAN_IN), .A(n20877), 
        .ZN(n20879) );
  AOI22_X1 U23862 ( .A1(n20928), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n20882), .B2(n20926), .ZN(n20883) );
  OAI211_X1 U23863 ( .C1(n20932), .C2(n20885), .A(n20884), .B(n20883), .ZN(
        P1_U3129) );
  AOI22_X1 U23864 ( .A1(n20925), .A2(n20887), .B1(n20886), .B2(n20922), .ZN(
        n20890) );
  AOI22_X1 U23865 ( .A1(n20928), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n20888), .B2(n20926), .ZN(n20889) );
  OAI211_X1 U23866 ( .C1(n20932), .C2(n20891), .A(n20890), .B(n20889), .ZN(
        P1_U3130) );
  AOI22_X1 U23867 ( .A1(n20925), .A2(n20893), .B1(n20892), .B2(n20922), .ZN(
        n20896) );
  AOI22_X1 U23868 ( .A1(n20928), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n20894), .B2(n20926), .ZN(n20895) );
  OAI211_X1 U23869 ( .C1(n20932), .C2(n20897), .A(n20896), .B(n20895), .ZN(
        P1_U3131) );
  AOI22_X1 U23870 ( .A1(n20925), .A2(n20899), .B1(n20898), .B2(n20922), .ZN(
        n20902) );
  AOI22_X1 U23871 ( .A1(n20928), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n20900), .B2(n20926), .ZN(n20901) );
  OAI211_X1 U23872 ( .C1(n20932), .C2(n20903), .A(n20902), .B(n20901), .ZN(
        P1_U3132) );
  AOI22_X1 U23873 ( .A1(n20925), .A2(n20905), .B1(n20904), .B2(n20922), .ZN(
        n20908) );
  AOI22_X1 U23874 ( .A1(n20928), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n20906), .B2(n20926), .ZN(n20907) );
  OAI211_X1 U23875 ( .C1(n20932), .C2(n20909), .A(n20908), .B(n20907), .ZN(
        P1_U3133) );
  AOI22_X1 U23876 ( .A1(n20925), .A2(n20911), .B1(n20910), .B2(n20922), .ZN(
        n20914) );
  AOI22_X1 U23877 ( .A1(n20928), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n20912), .B2(n20926), .ZN(n20913) );
  OAI211_X1 U23878 ( .C1(n20932), .C2(n20915), .A(n20914), .B(n20913), .ZN(
        P1_U3134) );
  AOI22_X1 U23879 ( .A1(n20925), .A2(n20917), .B1(n20916), .B2(n20922), .ZN(
        n20920) );
  AOI22_X1 U23880 ( .A1(n20928), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n20918), .B2(n20926), .ZN(n20919) );
  OAI211_X1 U23881 ( .C1(n20932), .C2(n20921), .A(n20920), .B(n20919), .ZN(
        P1_U3135) );
  AOI22_X1 U23882 ( .A1(n20925), .A2(n20924), .B1(n20923), .B2(n20922), .ZN(
        n20930) );
  AOI22_X1 U23883 ( .A1(n20928), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n20927), .B2(n20926), .ZN(n20929) );
  OAI211_X1 U23884 ( .C1(n20932), .C2(n20931), .A(n20930), .B(n20929), .ZN(
        P1_U3136) );
  NOR2_X1 U23885 ( .A1(n9922), .A2(n21133), .ZN(n20935) );
  OAI21_X1 U23886 ( .B1(n20935), .B2(n14046), .A(n20934), .ZN(P1_U3163) );
  INV_X1 U23887 ( .A(n21002), .ZN(n20936) );
  AND2_X1 U23888 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20936), .ZN(
        P1_U3164) );
  AND2_X1 U23889 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20936), .ZN(
        P1_U3165) );
  AND2_X1 U23890 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20936), .ZN(
        P1_U3166) );
  AND2_X1 U23891 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20936), .ZN(
        P1_U3167) );
  AND2_X1 U23892 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20936), .ZN(
        P1_U3168) );
  AND2_X1 U23893 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20936), .ZN(
        P1_U3169) );
  AND2_X1 U23894 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20936), .ZN(
        P1_U3170) );
  AND2_X1 U23895 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20936), .ZN(
        P1_U3171) );
  AND2_X1 U23896 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20936), .ZN(
        P1_U3172) );
  NOR2_X1 U23897 ( .A1(n21002), .A2(n21119), .ZN(P1_U3173) );
  AND2_X1 U23898 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20936), .ZN(
        P1_U3174) );
  AND2_X1 U23899 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20936), .ZN(
        P1_U3175) );
  AND2_X1 U23900 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20936), .ZN(
        P1_U3176) );
  INV_X1 U23901 ( .A(P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n21253) );
  NOR2_X1 U23902 ( .A1(n21002), .A2(n21253), .ZN(P1_U3177) );
  AND2_X1 U23903 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20936), .ZN(
        P1_U3178) );
  AND2_X1 U23904 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20936), .ZN(
        P1_U3179) );
  AND2_X1 U23905 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20936), .ZN(
        P1_U3180) );
  AND2_X1 U23906 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20936), .ZN(
        P1_U3181) );
  AND2_X1 U23907 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20936), .ZN(
        P1_U3182) );
  INV_X1 U23908 ( .A(P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21205) );
  NOR2_X1 U23909 ( .A1(n21002), .A2(n21205), .ZN(P1_U3183) );
  AND2_X1 U23910 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20936), .ZN(
        P1_U3184) );
  AND2_X1 U23911 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20936), .ZN(
        P1_U3185) );
  AND2_X1 U23912 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20936), .ZN(P1_U3186) );
  AND2_X1 U23913 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20936), .ZN(P1_U3187) );
  AND2_X1 U23914 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20936), .ZN(P1_U3188) );
  AND2_X1 U23915 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20936), .ZN(P1_U3189) );
  AND2_X1 U23916 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20936), .ZN(P1_U3190) );
  AND2_X1 U23917 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20936), .ZN(P1_U3191) );
  AND2_X1 U23918 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20936), .ZN(P1_U3192) );
  NOR2_X1 U23919 ( .A1(n21002), .A2(n20937), .ZN(P1_U3193) );
  AOI21_X1 U23920 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20943), .A(n20944), 
        .ZN(n20948) );
  INV_X1 U23921 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21037) );
  OAI22_X1 U23922 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20946), .B1(n12593), 
        .B2(n20938), .ZN(n20939) );
  NOR3_X1 U23923 ( .A1(n20940), .A2(n21037), .A3(n20939), .ZN(n20941) );
  OAI22_X1 U23924 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20948), .B1(n21025), 
        .B2(n20941), .ZN(P1_U3194) );
  AOI21_X1 U23925 ( .B1(n20943), .B2(n20946), .A(n20942), .ZN(n20950) );
  OAI211_X1 U23926 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21037), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20949) );
  NOR3_X1 U23927 ( .A1(n21037), .A2(NA), .A3(n20944), .ZN(n20945) );
  OAI22_X1 U23928 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20946), .B1(
        P1_STATE_REG_2__SCAN_IN), .B2(n20945), .ZN(n20947) );
  OAI22_X1 U23929 ( .A1(n20950), .A2(n20949), .B1(n20948), .B2(n20947), .ZN(
        P1_U3196) );
  OR2_X1 U23930 ( .A1(n21024), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20984) );
  INV_X1 U23931 ( .A(n20984), .ZN(n20992) );
  OR2_X1 U23932 ( .A1(n20951), .A2(n21038), .ZN(n20981) );
  INV_X1 U23933 ( .A(n20981), .ZN(n20993) );
  AOI222_X1 U23934 ( .A1(n20992), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20993), .ZN(n20952) );
  INV_X1 U23935 ( .A(n20952), .ZN(P1_U3197) );
  AOI222_X1 U23936 ( .A1(n20993), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21038), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20992), .ZN(n20953) );
  INV_X1 U23937 ( .A(n20953), .ZN(P1_U3198) );
  OAI222_X1 U23938 ( .A1(n20981), .A2(n20955), .B1(n20954), .B2(n21025), .C1(
        n20957), .C2(n20984), .ZN(P1_U3199) );
  AOI22_X1 U23939 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n21038), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20992), .ZN(n20956) );
  OAI21_X1 U23940 ( .B1(n20957), .B2(n20981), .A(n20956), .ZN(P1_U3200) );
  AOI22_X1 U23941 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n21038), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20993), .ZN(n20958) );
  OAI21_X1 U23942 ( .B1(n20959), .B2(n20984), .A(n20958), .ZN(P1_U3201) );
  AOI222_X1 U23943 ( .A1(n20993), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20992), .ZN(n20960) );
  INV_X1 U23944 ( .A(n20960), .ZN(P1_U3202) );
  AOI22_X1 U23945 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21038), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20992), .ZN(n20961) );
  OAI21_X1 U23946 ( .B1(n20962), .B2(n20981), .A(n20961), .ZN(P1_U3203) );
  AOI22_X1 U23947 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n21038), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20993), .ZN(n20963) );
  OAI21_X1 U23948 ( .B1(n20964), .B2(n20984), .A(n20963), .ZN(P1_U3204) );
  AOI222_X1 U23949 ( .A1(n20993), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21038), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20992), .ZN(n20965) );
  INV_X1 U23950 ( .A(n20965), .ZN(P1_U3205) );
  AOI222_X1 U23951 ( .A1(n20992), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20993), .ZN(n20966) );
  INV_X1 U23952 ( .A(n20966), .ZN(P1_U3206) );
  AOI222_X1 U23953 ( .A1(n20993), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20992), .ZN(n20967) );
  INV_X1 U23954 ( .A(n20967), .ZN(P1_U3207) );
  AOI222_X1 U23955 ( .A1(n20992), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20993), .ZN(n20968) );
  INV_X1 U23956 ( .A(n20968), .ZN(P1_U3208) );
  AOI22_X1 U23957 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n21038), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20992), .ZN(n20969) );
  OAI21_X1 U23958 ( .B1(n20970), .B2(n20981), .A(n20969), .ZN(P1_U3209) );
  AOI22_X1 U23959 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n21038), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20993), .ZN(n20971) );
  OAI21_X1 U23960 ( .B1(n20972), .B2(n20984), .A(n20971), .ZN(P1_U3210) );
  AOI222_X1 U23961 ( .A1(n20993), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20992), .ZN(n20973) );
  INV_X1 U23962 ( .A(n20973), .ZN(P1_U3211) );
  AOI222_X1 U23963 ( .A1(n20993), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20992), .ZN(n20974) );
  INV_X1 U23964 ( .A(n20974), .ZN(P1_U3212) );
  AOI222_X1 U23965 ( .A1(n20993), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20992), .ZN(n20975) );
  INV_X1 U23966 ( .A(n20975), .ZN(P1_U3213) );
  AOI222_X1 U23967 ( .A1(n20993), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20992), .ZN(n20976) );
  INV_X1 U23968 ( .A(n20976), .ZN(P1_U3214) );
  AOI222_X1 U23969 ( .A1(n20993), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20992), .ZN(n20977) );
  INV_X1 U23970 ( .A(n20977), .ZN(P1_U3215) );
  AOI222_X1 U23971 ( .A1(n20992), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20993), .ZN(n20978) );
  INV_X1 U23972 ( .A(n20978), .ZN(P1_U3216) );
  AOI222_X1 U23973 ( .A1(n20993), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20992), .ZN(n20979) );
  INV_X1 U23974 ( .A(n20979), .ZN(P1_U3217) );
  AOI22_X1 U23975 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21038), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20992), .ZN(n20980) );
  OAI21_X1 U23976 ( .B1(n20982), .B2(n20981), .A(n20980), .ZN(P1_U3218) );
  AOI22_X1 U23977 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21038), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20993), .ZN(n20983) );
  OAI21_X1 U23978 ( .B1(n20985), .B2(n20984), .A(n20983), .ZN(P1_U3219) );
  AOI222_X1 U23979 ( .A1(n20993), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20992), .ZN(n20986) );
  INV_X1 U23980 ( .A(n20986), .ZN(P1_U3220) );
  AOI222_X1 U23981 ( .A1(n20993), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20992), .ZN(n20987) );
  INV_X1 U23982 ( .A(n20987), .ZN(P1_U3221) );
  AOI222_X1 U23983 ( .A1(n20993), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20992), .ZN(n20988) );
  INV_X1 U23984 ( .A(n20988), .ZN(P1_U3222) );
  AOI222_X1 U23985 ( .A1(n20993), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20992), .ZN(n20989) );
  INV_X1 U23986 ( .A(n20989), .ZN(P1_U3223) );
  AOI222_X1 U23987 ( .A1(n20992), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20993), .ZN(n20990) );
  INV_X1 U23988 ( .A(n20990), .ZN(P1_U3224) );
  AOI222_X1 U23989 ( .A1(n20993), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20992), .ZN(n20991) );
  INV_X1 U23990 ( .A(n20991), .ZN(P1_U3225) );
  AOI222_X1 U23991 ( .A1(n20993), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21024), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20992), .ZN(n20994) );
  INV_X1 U23992 ( .A(n20994), .ZN(P1_U3226) );
  OAI22_X1 U23993 ( .A1(n21024), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21025), .ZN(n20995) );
  INV_X1 U23994 ( .A(n20995), .ZN(P1_U3458) );
  OAI22_X1 U23995 ( .A1(n21038), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21025), .ZN(n20996) );
  INV_X1 U23996 ( .A(n20996), .ZN(P1_U3459) );
  OAI22_X1 U23997 ( .A1(n21038), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21025), .ZN(n20997) );
  INV_X1 U23998 ( .A(n20997), .ZN(P1_U3460) );
  OAI22_X1 U23999 ( .A1(n21038), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21025), .ZN(n20998) );
  INV_X1 U24000 ( .A(n20998), .ZN(P1_U3461) );
  OAI21_X1 U24001 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21002), .A(n21000), 
        .ZN(n20999) );
  INV_X1 U24002 ( .A(n20999), .ZN(P1_U3464) );
  OAI21_X1 U24003 ( .B1(n21002), .B2(n21001), .A(n21000), .ZN(P1_U3465) );
  INV_X1 U24004 ( .A(n21003), .ZN(n21009) );
  INV_X1 U24005 ( .A(n21004), .ZN(n21008) );
  INV_X1 U24006 ( .A(n21005), .ZN(n21006) );
  OAI222_X1 U24007 ( .A1(n21011), .A2(n21010), .B1(n21009), .B2(n21008), .C1(
        n21007), .C2(n21006), .ZN(n21013) );
  OAI22_X1 U24008 ( .A1(n21014), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21013), .B2(n21012), .ZN(n21015) );
  INV_X1 U24009 ( .A(n21015), .ZN(P1_U3472) );
  AOI21_X1 U24010 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21017) );
  AOI22_X1 U24011 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21017), .B2(n21016), .ZN(n21019) );
  INV_X1 U24012 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21018) );
  AOI22_X1 U24013 ( .A1(n21020), .A2(n21019), .B1(n21018), .B2(n21022), .ZN(
        P1_U3481) );
  INV_X1 U24014 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21023) );
  NOR2_X1 U24015 ( .A1(n21022), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21021) );
  AOI22_X1 U24016 ( .A1(n21023), .A2(n21022), .B1(n12980), .B2(n21021), .ZN(
        P1_U3482) );
  AOI22_X1 U24017 ( .A1(n21025), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21064), 
        .B2(n21024), .ZN(P1_U3483) );
  AOI211_X1 U24018 ( .C1(n21029), .C2(n21028), .A(n21027), .B(n21026), .ZN(
        n21036) );
  NAND2_X1 U24019 ( .A1(n21030), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21031) );
  OAI21_X1 U24020 ( .B1(n21032), .B2(n21031), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n21035) );
  NOR2_X1 U24021 ( .A1(n21036), .A2(n21033), .ZN(n21034) );
  AOI22_X1 U24022 ( .A1(n21037), .A2(n21036), .B1(n21035), .B2(n21034), .ZN(
        P1_U3485) );
  MUX2_X1 U24023 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21038), .Z(P1_U3486) );
  AOI222_X1 U24024 ( .A1(n21043), .A2(n21042), .B1(P1_EBX_REG_9__SCAN_IN), 
        .B2(n21041), .C1(n21040), .C2(n21039), .ZN(n21287) );
  INV_X1 U24025 ( .A(DATAI_13_), .ZN(n21046) );
  AOI22_X1 U24026 ( .A1(n21046), .A2(keyinput101), .B1(n21045), .B2(keyinput77), .ZN(n21044) );
  OAI221_X1 U24027 ( .B1(n21046), .B2(keyinput101), .C1(n21045), .C2(
        keyinput77), .A(n21044), .ZN(n21049) );
  XNOR2_X1 U24028 ( .A(n21047), .B(keyinput51), .ZN(n21048) );
  NOR2_X1 U24029 ( .A1(n21049), .A2(n21048), .ZN(n21059) );
  AOI22_X1 U24030 ( .A1(n21051), .A2(keyinput3), .B1(keyinput25), .B2(n21323), 
        .ZN(n21050) );
  OAI221_X1 U24031 ( .B1(n21051), .B2(keyinput3), .C1(n21323), .C2(keyinput25), 
        .A(n21050), .ZN(n21052) );
  INV_X1 U24032 ( .A(n21052), .ZN(n21058) );
  AOI22_X1 U24033 ( .A1(n21054), .A2(keyinput74), .B1(n11626), .B2(keyinput45), 
        .ZN(n21053) );
  OAI221_X1 U24034 ( .B1(n21054), .B2(keyinput74), .C1(n11626), .C2(keyinput45), .A(n21053), .ZN(n21055) );
  INV_X1 U24035 ( .A(n21055), .ZN(n21057) );
  XNOR2_X1 U24036 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B(keyinput71), .ZN(
        n21056) );
  AND4_X1 U24037 ( .A1(n21059), .A2(n21058), .A3(n21057), .A4(n21056), .ZN(
        n21104) );
  INV_X1 U24038 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n21061) );
  AOI22_X1 U24039 ( .A1(n21319), .A2(keyinput62), .B1(keyinput15), .B2(n21061), 
        .ZN(n21060) );
  OAI221_X1 U24040 ( .B1(n21319), .B2(keyinput62), .C1(n21061), .C2(keyinput15), .A(n21060), .ZN(n21073) );
  AOI22_X1 U24041 ( .A1(n21064), .A2(keyinput43), .B1(n21063), .B2(keyinput85), 
        .ZN(n21062) );
  OAI221_X1 U24042 ( .B1(n21064), .B2(keyinput43), .C1(n21063), .C2(keyinput85), .A(n21062), .ZN(n21072) );
  AOI22_X1 U24043 ( .A1(n21067), .A2(keyinput22), .B1(n21066), .B2(keyinput9), 
        .ZN(n21065) );
  OAI221_X1 U24044 ( .B1(n21067), .B2(keyinput22), .C1(n21066), .C2(keyinput9), 
        .A(n21065), .ZN(n21071) );
  XOR2_X1 U24045 ( .A(n11644), .B(keyinput88), .Z(n21069) );
  XNOR2_X1 U24046 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput87), .ZN(
        n21068) );
  NAND2_X1 U24047 ( .A1(n21069), .A2(n21068), .ZN(n21070) );
  NOR4_X1 U24048 ( .A1(n21073), .A2(n21072), .A3(n21071), .A4(n21070), .ZN(
        n21103) );
  AOI22_X1 U24049 ( .A1(n21076), .A2(keyinput123), .B1(keyinput90), .B2(n21075), .ZN(n21074) );
  OAI221_X1 U24050 ( .B1(n21076), .B2(keyinput123), .C1(n21075), .C2(
        keyinput90), .A(n21074), .ZN(n21086) );
  AOI22_X1 U24051 ( .A1(n21078), .A2(keyinput7), .B1(n11236), .B2(keyinput95), 
        .ZN(n21077) );
  OAI221_X1 U24052 ( .B1(n21078), .B2(keyinput7), .C1(n11236), .C2(keyinput95), 
        .A(n21077), .ZN(n21085) );
  INV_X1 U24053 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n21080) );
  AOI22_X1 U24054 ( .A1(n21081), .A2(keyinput125), .B1(n21080), .B2(keyinput44), .ZN(n21079) );
  OAI221_X1 U24055 ( .B1(n21081), .B2(keyinput125), .C1(n21080), .C2(
        keyinput44), .A(n21079), .ZN(n21084) );
  AOI22_X1 U24056 ( .A1(n21294), .A2(keyinput99), .B1(keyinput81), .B2(n21324), 
        .ZN(n21082) );
  OAI221_X1 U24057 ( .B1(n21294), .B2(keyinput99), .C1(n21324), .C2(keyinput81), .A(n21082), .ZN(n21083) );
  NOR4_X1 U24058 ( .A1(n21086), .A2(n21085), .A3(n21084), .A4(n21083), .ZN(
        n21102) );
  INV_X1 U24059 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n21088) );
  AOI22_X1 U24060 ( .A1(n21088), .A2(keyinput97), .B1(n21321), .B2(keyinput13), 
        .ZN(n21087) );
  OAI221_X1 U24061 ( .B1(n21088), .B2(keyinput97), .C1(n21321), .C2(keyinput13), .A(n21087), .ZN(n21092) );
  XNOR2_X1 U24062 ( .A(n21089), .B(keyinput50), .ZN(n21091) );
  XOR2_X1 U24063 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B(keyinput55), .Z(
        n21090) );
  OR3_X1 U24064 ( .A1(n21092), .A2(n21091), .A3(n21090), .ZN(n21100) );
  AOI22_X1 U24065 ( .A1(n21095), .A2(keyinput121), .B1(keyinput86), .B2(n21094), .ZN(n21093) );
  OAI221_X1 U24066 ( .B1(n21095), .B2(keyinput121), .C1(n21094), .C2(
        keyinput86), .A(n21093), .ZN(n21099) );
  AOI22_X1 U24067 ( .A1(n21097), .A2(keyinput92), .B1(n14046), .B2(keyinput53), 
        .ZN(n21096) );
  OAI221_X1 U24068 ( .B1(n21097), .B2(keyinput92), .C1(n14046), .C2(keyinput53), .A(n21096), .ZN(n21098) );
  NOR3_X1 U24069 ( .A1(n21100), .A2(n21099), .A3(n21098), .ZN(n21101) );
  NAND4_X1 U24070 ( .A1(n21104), .A2(n21103), .A3(n21102), .A4(n21101), .ZN(
        n21285) );
  AOI22_X1 U24071 ( .A1(n21106), .A2(keyinput33), .B1(n21296), .B2(keyinput12), 
        .ZN(n21105) );
  OAI221_X1 U24072 ( .B1(n21106), .B2(keyinput33), .C1(n21296), .C2(keyinput12), .A(n21105), .ZN(n21117) );
  AOI22_X1 U24073 ( .A1(n21109), .A2(keyinput35), .B1(n21108), .B2(keyinput67), 
        .ZN(n21107) );
  OAI221_X1 U24074 ( .B1(n21109), .B2(keyinput35), .C1(n21108), .C2(keyinput67), .A(n21107), .ZN(n21116) );
  AOI22_X1 U24075 ( .A1(n11733), .A2(keyinput61), .B1(keyinput11), .B2(n21111), 
        .ZN(n21110) );
  OAI221_X1 U24076 ( .B1(n11733), .B2(keyinput61), .C1(n21111), .C2(keyinput11), .A(n21110), .ZN(n21115) );
  AOI22_X1 U24077 ( .A1(n13996), .A2(keyinput109), .B1(keyinput23), .B2(n21113), .ZN(n21112) );
  OAI221_X1 U24078 ( .B1(n13996), .B2(keyinput109), .C1(n21113), .C2(
        keyinput23), .A(n21112), .ZN(n21114) );
  NOR4_X1 U24079 ( .A1(n21117), .A2(n21116), .A3(n21115), .A4(n21114), .ZN(
        n21160) );
  AOI22_X1 U24080 ( .A1(n21120), .A2(keyinput49), .B1(keyinput111), .B2(n21119), .ZN(n21118) );
  OAI221_X1 U24081 ( .B1(n21120), .B2(keyinput49), .C1(n21119), .C2(
        keyinput111), .A(n21118), .ZN(n21130) );
  AOI22_X1 U24082 ( .A1(n21123), .A2(keyinput70), .B1(n21122), .B2(keyinput1), 
        .ZN(n21121) );
  OAI221_X1 U24083 ( .B1(n21123), .B2(keyinput70), .C1(n21122), .C2(keyinput1), 
        .A(n21121), .ZN(n21129) );
  AOI22_X1 U24084 ( .A1(n11243), .A2(keyinput2), .B1(keyinput28), .B2(n11069), 
        .ZN(n21124) );
  OAI221_X1 U24085 ( .B1(n11243), .B2(keyinput2), .C1(n11069), .C2(keyinput28), 
        .A(n21124), .ZN(n21128) );
  INV_X1 U24086 ( .A(P3_CODEFETCH_REG_SCAN_IN), .ZN(n21292) );
  AOI22_X1 U24087 ( .A1(n21126), .A2(keyinput79), .B1(keyinput116), .B2(n21292), .ZN(n21125) );
  OAI221_X1 U24088 ( .B1(n21126), .B2(keyinput79), .C1(n21292), .C2(
        keyinput116), .A(n21125), .ZN(n21127) );
  NOR4_X1 U24089 ( .A1(n21130), .A2(n21129), .A3(n21128), .A4(n21127), .ZN(
        n21159) );
  AOI22_X1 U24090 ( .A1(n21133), .A2(keyinput8), .B1(n21132), .B2(keyinput107), 
        .ZN(n21131) );
  OAI221_X1 U24091 ( .B1(n21133), .B2(keyinput8), .C1(n21132), .C2(keyinput107), .A(n21131), .ZN(n21143) );
  AOI22_X1 U24092 ( .A1(n16166), .A2(keyinput112), .B1(keyinput37), .B2(n21135), .ZN(n21134) );
  OAI221_X1 U24093 ( .B1(n16166), .B2(keyinput112), .C1(n21135), .C2(
        keyinput37), .A(n21134), .ZN(n21142) );
  AOI22_X1 U24094 ( .A1(n21137), .A2(keyinput21), .B1(keyinput105), .B2(n21325), .ZN(n21136) );
  OAI221_X1 U24095 ( .B1(n21137), .B2(keyinput21), .C1(n21325), .C2(
        keyinput105), .A(n21136), .ZN(n21141) );
  AOI22_X1 U24096 ( .A1(n21139), .A2(keyinput27), .B1(n21320), .B2(keyinput117), .ZN(n21138) );
  OAI221_X1 U24097 ( .B1(n21139), .B2(keyinput27), .C1(n21320), .C2(
        keyinput117), .A(n21138), .ZN(n21140) );
  NOR4_X1 U24098 ( .A1(n21143), .A2(n21142), .A3(n21141), .A4(n21140), .ZN(
        n21158) );
  AOI22_X1 U24099 ( .A1(n21145), .A2(keyinput64), .B1(n10145), .B2(keyinput84), 
        .ZN(n21144) );
  OAI221_X1 U24100 ( .B1(n21145), .B2(keyinput64), .C1(n10145), .C2(keyinput84), .A(n21144), .ZN(n21156) );
  AOI22_X1 U24101 ( .A1(n10104), .A2(keyinput42), .B1(keyinput16), .B2(n21147), 
        .ZN(n21146) );
  OAI221_X1 U24102 ( .B1(n10104), .B2(keyinput42), .C1(n21147), .C2(keyinput16), .A(n21146), .ZN(n21155) );
  AOI22_X1 U24103 ( .A1(n21150), .A2(keyinput34), .B1(keyinput124), .B2(n21149), .ZN(n21148) );
  OAI221_X1 U24104 ( .B1(n21150), .B2(keyinput34), .C1(n21149), .C2(
        keyinput124), .A(n21148), .ZN(n21154) );
  AOI22_X1 U24105 ( .A1(n12705), .A2(keyinput66), .B1(n21152), .B2(keyinput104), .ZN(n21151) );
  OAI221_X1 U24106 ( .B1(n12705), .B2(keyinput66), .C1(n21152), .C2(
        keyinput104), .A(n21151), .ZN(n21153) );
  NOR4_X1 U24107 ( .A1(n21156), .A2(n21155), .A3(n21154), .A4(n21153), .ZN(
        n21157) );
  NAND4_X1 U24108 ( .A1(n21160), .A2(n21159), .A3(n21158), .A4(n21157), .ZN(
        n21284) );
  AOI22_X1 U24109 ( .A1(n10876), .A2(keyinput32), .B1(n11867), .B2(keyinput127), .ZN(n21161) );
  OAI221_X1 U24110 ( .B1(n10876), .B2(keyinput32), .C1(n11867), .C2(
        keyinput127), .A(n21161), .ZN(n21171) );
  AOI22_X1 U24111 ( .A1(n21163), .A2(keyinput93), .B1(keyinput57), .B2(n14122), 
        .ZN(n21162) );
  OAI221_X1 U24112 ( .B1(n21163), .B2(keyinput93), .C1(n14122), .C2(keyinput57), .A(n21162), .ZN(n21170) );
  AOI22_X1 U24113 ( .A1(n21166), .A2(keyinput76), .B1(n21165), .B2(keyinput46), 
        .ZN(n21164) );
  OAI221_X1 U24114 ( .B1(n21166), .B2(keyinput76), .C1(n21165), .C2(keyinput46), .A(n21164), .ZN(n21169) );
  AOI22_X1 U24115 ( .A1(n16220), .A2(keyinput56), .B1(n11309), .B2(keyinput82), 
        .ZN(n21167) );
  OAI221_X1 U24116 ( .B1(n16220), .B2(keyinput56), .C1(n11309), .C2(keyinput82), .A(n21167), .ZN(n21168) );
  NOR4_X1 U24117 ( .A1(n21171), .A2(n21170), .A3(n21169), .A4(n21168), .ZN(
        n21219) );
  AOI22_X1 U24118 ( .A1(n21174), .A2(keyinput98), .B1(keyinput113), .B2(n21173), .ZN(n21172) );
  OAI221_X1 U24119 ( .B1(n21174), .B2(keyinput98), .C1(n21173), .C2(
        keyinput113), .A(n21172), .ZN(n21185) );
  AOI22_X1 U24120 ( .A1(n21295), .A2(keyinput89), .B1(keyinput80), .B2(n21176), 
        .ZN(n21175) );
  OAI221_X1 U24121 ( .B1(n21295), .B2(keyinput89), .C1(n21176), .C2(keyinput80), .A(n21175), .ZN(n21184) );
  INV_X1 U24122 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n21178) );
  AOI22_X1 U24123 ( .A1(n21179), .A2(keyinput91), .B1(n21178), .B2(keyinput17), 
        .ZN(n21177) );
  OAI221_X1 U24124 ( .B1(n21179), .B2(keyinput91), .C1(n21178), .C2(keyinput17), .A(n21177), .ZN(n21183) );
  AOI22_X1 U24125 ( .A1(n11289), .A2(keyinput14), .B1(keyinput58), .B2(n21181), 
        .ZN(n21180) );
  OAI221_X1 U24126 ( .B1(n11289), .B2(keyinput14), .C1(n21181), .C2(keyinput58), .A(n21180), .ZN(n21182) );
  NOR4_X1 U24127 ( .A1(n21185), .A2(n21184), .A3(n21183), .A4(n21182), .ZN(
        n21218) );
  AOI22_X1 U24128 ( .A1(n21187), .A2(keyinput102), .B1(n11664), .B2(keyinput5), 
        .ZN(n21186) );
  OAI221_X1 U24129 ( .B1(n21187), .B2(keyinput102), .C1(n11664), .C2(keyinput5), .A(n21186), .ZN(n21191) );
  XOR2_X1 U24130 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B(keyinput36), .Z(
        n21190) );
  XNOR2_X1 U24131 ( .A(n21188), .B(keyinput59), .ZN(n21189) );
  OR3_X1 U24132 ( .A1(n21191), .A2(n21190), .A3(n21189), .ZN(n21200) );
  AOI22_X1 U24133 ( .A1(n21194), .A2(keyinput120), .B1(keyinput106), .B2(
        n21193), .ZN(n21192) );
  OAI221_X1 U24134 ( .B1(n21194), .B2(keyinput120), .C1(n21193), .C2(
        keyinput106), .A(n21192), .ZN(n21199) );
  AOI22_X1 U24135 ( .A1(n21197), .A2(keyinput20), .B1(keyinput18), .B2(n21196), 
        .ZN(n21195) );
  OAI221_X1 U24136 ( .B1(n21197), .B2(keyinput20), .C1(n21196), .C2(keyinput18), .A(n21195), .ZN(n21198) );
  NOR3_X1 U24137 ( .A1(n21200), .A2(n21199), .A3(n21198), .ZN(n21217) );
  AOI22_X1 U24138 ( .A1(n21203), .A2(keyinput126), .B1(n21202), .B2(
        keyinput119), .ZN(n21201) );
  OAI221_X1 U24139 ( .B1(n21203), .B2(keyinput126), .C1(n21202), .C2(
        keyinput119), .A(n21201), .ZN(n21215) );
  AOI22_X1 U24140 ( .A1(n21206), .A2(keyinput54), .B1(keyinput83), .B2(n21205), 
        .ZN(n21204) );
  OAI221_X1 U24141 ( .B1(n21206), .B2(keyinput54), .C1(n21205), .C2(keyinput83), .A(n21204), .ZN(n21214) );
  AOI22_X1 U24142 ( .A1(n21293), .A2(keyinput29), .B1(n21208), .B2(keyinput47), 
        .ZN(n21207) );
  OAI221_X1 U24143 ( .B1(n21293), .B2(keyinput29), .C1(n21208), .C2(keyinput47), .A(n21207), .ZN(n21213) );
  AOI22_X1 U24144 ( .A1(n21211), .A2(keyinput39), .B1(n21210), .B2(keyinput69), 
        .ZN(n21209) );
  OAI221_X1 U24145 ( .B1(n21211), .B2(keyinput39), .C1(n21210), .C2(keyinput69), .A(n21209), .ZN(n21212) );
  NOR4_X1 U24146 ( .A1(n21215), .A2(n21214), .A3(n21213), .A4(n21212), .ZN(
        n21216) );
  NAND4_X1 U24147 ( .A1(n21219), .A2(n21218), .A3(n21217), .A4(n21216), .ZN(
        n21283) );
  AOI22_X1 U24148 ( .A1(n21222), .A2(keyinput4), .B1(n21221), .B2(keyinput60), 
        .ZN(n21220) );
  OAI221_X1 U24149 ( .B1(n21222), .B2(keyinput4), .C1(n21221), .C2(keyinput60), 
        .A(n21220), .ZN(n21235) );
  AOI22_X1 U24150 ( .A1(n21225), .A2(keyinput10), .B1(n21224), .B2(keyinput94), 
        .ZN(n21223) );
  OAI221_X1 U24151 ( .B1(n21225), .B2(keyinput10), .C1(n21224), .C2(keyinput94), .A(n21223), .ZN(n21234) );
  AOI22_X1 U24152 ( .A1(n21228), .A2(keyinput114), .B1(n21227), .B2(keyinput0), 
        .ZN(n21226) );
  OAI221_X1 U24153 ( .B1(n21228), .B2(keyinput114), .C1(n21227), .C2(keyinput0), .A(n21226), .ZN(n21233) );
  INV_X1 U24154 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n21231) );
  AOI22_X1 U24155 ( .A1(n21231), .A2(keyinput65), .B1(n21230), .B2(keyinput38), 
        .ZN(n21229) );
  OAI221_X1 U24156 ( .B1(n21231), .B2(keyinput65), .C1(n21230), .C2(keyinput38), .A(n21229), .ZN(n21232) );
  NOR4_X1 U24157 ( .A1(n21235), .A2(n21234), .A3(n21233), .A4(n21232), .ZN(
        n21281) );
  AOI22_X1 U24158 ( .A1(n21238), .A2(keyinput103), .B1(keyinput19), .B2(n21237), .ZN(n21236) );
  OAI221_X1 U24159 ( .B1(n21238), .B2(keyinput103), .C1(n21237), .C2(
        keyinput19), .A(n21236), .ZN(n21251) );
  AOI22_X1 U24160 ( .A1(n21241), .A2(keyinput75), .B1(keyinput96), .B2(n21240), 
        .ZN(n21239) );
  OAI221_X1 U24161 ( .B1(n21241), .B2(keyinput75), .C1(n21240), .C2(keyinput96), .A(n21239), .ZN(n21250) );
  AOI22_X1 U24162 ( .A1(n21244), .A2(keyinput78), .B1(keyinput24), .B2(n21243), 
        .ZN(n21242) );
  OAI221_X1 U24163 ( .B1(n21244), .B2(keyinput78), .C1(n21243), .C2(keyinput24), .A(n21242), .ZN(n21249) );
  AOI22_X1 U24164 ( .A1(n21247), .A2(keyinput63), .B1(keyinput108), .B2(n21246), .ZN(n21245) );
  OAI221_X1 U24165 ( .B1(n21247), .B2(keyinput63), .C1(n21246), .C2(
        keyinput108), .A(n21245), .ZN(n21248) );
  NOR4_X1 U24166 ( .A1(n21251), .A2(n21250), .A3(n21249), .A4(n21248), .ZN(
        n21280) );
  AOI22_X1 U24167 ( .A1(n21326), .A2(keyinput110), .B1(keyinput73), .B2(n21253), .ZN(n21252) );
  OAI221_X1 U24168 ( .B1(n21326), .B2(keyinput110), .C1(n21253), .C2(
        keyinput73), .A(n21252), .ZN(n21264) );
  AOI22_X1 U24169 ( .A1(n21256), .A2(keyinput48), .B1(n21255), .B2(keyinput40), 
        .ZN(n21254) );
  OAI221_X1 U24170 ( .B1(n21256), .B2(keyinput48), .C1(n21255), .C2(keyinput40), .A(n21254), .ZN(n21263) );
  AOI22_X1 U24171 ( .A1(n11274), .A2(keyinput26), .B1(keyinput52), .B2(n11356), 
        .ZN(n21257) );
  OAI221_X1 U24172 ( .B1(n11274), .B2(keyinput26), .C1(n11356), .C2(keyinput52), .A(n21257), .ZN(n21262) );
  AOI22_X1 U24173 ( .A1(n21260), .A2(keyinput100), .B1(keyinput122), .B2(
        n21259), .ZN(n21258) );
  OAI221_X1 U24174 ( .B1(n21260), .B2(keyinput100), .C1(n21259), .C2(
        keyinput122), .A(n21258), .ZN(n21261) );
  NOR4_X1 U24175 ( .A1(n21264), .A2(n21263), .A3(n21262), .A4(n21261), .ZN(
        n21279) );
  AOI22_X1 U24176 ( .A1(n21322), .A2(keyinput68), .B1(keyinput30), .B2(n21266), 
        .ZN(n21265) );
  OAI221_X1 U24177 ( .B1(n21322), .B2(keyinput68), .C1(n21266), .C2(keyinput30), .A(n21265), .ZN(n21277) );
  AOI22_X1 U24178 ( .A1(n21327), .A2(keyinput115), .B1(n14849), .B2(keyinput6), 
        .ZN(n21267) );
  OAI221_X1 U24179 ( .B1(n21327), .B2(keyinput115), .C1(n14849), .C2(keyinput6), .A(n21267), .ZN(n21276) );
  INV_X1 U24180 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n21270) );
  AOI22_X1 U24181 ( .A1(n21270), .A2(keyinput41), .B1(n21269), .B2(keyinput31), 
        .ZN(n21268) );
  OAI221_X1 U24182 ( .B1(n21270), .B2(keyinput41), .C1(n21269), .C2(keyinput31), .A(n21268), .ZN(n21275) );
  INV_X1 U24183 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n21271) );
  XOR2_X1 U24184 ( .A(n21271), .B(keyinput72), .Z(n21273) );
  XNOR2_X1 U24185 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B(keyinput118), .ZN(
        n21272) );
  NAND2_X1 U24186 ( .A1(n21273), .A2(n21272), .ZN(n21274) );
  NOR4_X1 U24187 ( .A1(n21277), .A2(n21276), .A3(n21275), .A4(n21274), .ZN(
        n21278) );
  NAND4_X1 U24188 ( .A1(n21281), .A2(n21280), .A3(n21279), .A4(n21278), .ZN(
        n21282) );
  NOR4_X1 U24189 ( .A1(n21285), .A2(n21284), .A3(n21283), .A4(n21282), .ZN(
        n21286) );
  XNOR2_X1 U24190 ( .A(n21287), .B(n21286), .ZN(n21349) );
  NAND4_X1 U24191 ( .A1(n21291), .A2(n21290), .A3(n21289), .A4(n21288), .ZN(
        n21306) );
  NAND4_X1 U24192 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_5__0__SCAN_IN), .A3(P2_INSTQUEUE_REG_5__4__SCAN_IN), 
        .A4(BUF2_REG_28__SCAN_IN), .ZN(n21305) );
  NAND4_X1 U24193 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(P2_EAX_REG_18__SCAN_IN), .A4(
        BUF1_REG_20__SCAN_IN), .ZN(n21304) );
  NOR4_X1 U24194 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(n21294), .A3(n21293), .A4(
        n21292), .ZN(n21302) );
  INV_X1 U24195 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n21300) );
  NOR4_X1 U24196 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_EAX_REG_4__SCAN_IN), .A3(P1_EAX_REG_1__SCAN_IN), .A4(n21295), .ZN(
        n21298) );
  NOR4_X1 U24197 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_8__6__SCAN_IN), .A3(P1_INSTQUEUE_REG_13__6__SCAN_IN), 
        .A4(n21296), .ZN(n21297) );
  NAND3_X1 U24198 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21298), .A3(
        n21297), .ZN(n21299) );
  NOR4_X1 U24199 ( .A1(n21300), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A3(
        P1_EAX_REG_7__SCAN_IN), .A4(n21299), .ZN(n21301) );
  NAND2_X1 U24200 ( .A1(n21302), .A2(n21301), .ZN(n21303) );
  NOR4_X1 U24201 ( .A1(n21306), .A2(n21305), .A3(n21304), .A4(n21303), .ZN(
        n21347) );
  NAND4_X1 U24202 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(P2_REIP_REG_16__SCAN_IN), 
        .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(P2_DATAWIDTH_REG_1__SCAN_IN), 
        .ZN(n21310) );
  NAND4_X1 U24203 ( .A1(P2_EAX_REG_27__SCAN_IN), .A2(BUF1_REG_10__SCAN_IN), 
        .A3(BUF1_REG_16__SCAN_IN), .A4(P1_UWORD_REG_4__SCAN_IN), .ZN(n21309)
         );
  NAND4_X1 U24204 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(
        P3_REIP_REG_8__SCAN_IN), .A3(P3_EAX_REG_10__SCAN_IN), .A4(
        P3_EAX_REG_25__SCAN_IN), .ZN(n21308) );
  NAND4_X1 U24205 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAO_REG_17__SCAN_IN), .A4(
        P3_LWORD_REG_11__SCAN_IN), .ZN(n21307) );
  NOR4_X1 U24206 ( .A1(n21310), .A2(n21309), .A3(n21308), .A4(n21307), .ZN(
        n21346) );
  NAND4_X1 U24207 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        DATAI_13_), .ZN(n21314) );
  NAND4_X1 U24208 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_12__6__SCAN_IN), .A3(P2_INSTQUEUE_REG_14__5__SCAN_IN), 
        .A4(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21313) );
  NAND4_X1 U24209 ( .A1(BUF1_REG_6__SCAN_IN), .A2(BUF1_REG_4__SCAN_IN), .A3(
        P1_DATAWIDTH_REG_22__SCAN_IN), .A4(P1_LWORD_REG_0__SCAN_IN), .ZN(
        n21312) );
  NAND4_X1 U24210 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(
        P3_ADDRESS_REG_11__SCAN_IN), .A3(P1_W_R_N_REG_SCAN_IN), .A4(
        P3_BE_N_REG_1__SCAN_IN), .ZN(n21311) );
  NOR4_X1 U24211 ( .A1(n21314), .A2(n21313), .A3(n21312), .A4(n21311), .ZN(
        n21345) );
  NOR4_X1 U24212 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21318) );
  NOR4_X1 U24213 ( .A1(P2_EBX_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(P2_BE_N_REG_2__SCAN_IN), .A4(
        P2_LWORD_REG_13__SCAN_IN), .ZN(n21317) );
  NOR4_X1 U24214 ( .A1(BUF2_REG_13__SCAN_IN), .A2(P3_DATAO_REG_24__SCAN_IN), 
        .A3(P3_DATAO_REG_26__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n21316)
         );
  NOR4_X1 U24215 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_DATAO_REG_9__SCAN_IN), .A3(P3_LWORD_REG_14__SCAN_IN), .A4(
        P3_LWORD_REG_15__SCAN_IN), .ZN(n21315) );
  NAND4_X1 U24216 ( .A1(n21318), .A2(n21317), .A3(n21316), .A4(n21315), .ZN(
        n21343) );
  NOR4_X1 U24217 ( .A1(n21322), .A2(n21321), .A3(n21320), .A4(n21319), .ZN(
        n21331) );
  NOR4_X1 U24218 ( .A1(n16220), .A2(n21325), .A3(n21324), .A4(n21323), .ZN(
        n21330) );
  NOR4_X1 U24219 ( .A1(P1_EBX_REG_22__SCAN_IN), .A2(P1_EBX_REG_16__SCAN_IN), 
        .A3(BUF1_REG_5__SCAN_IN), .A4(P1_DATAO_REG_6__SCAN_IN), .ZN(n21329) );
  NOR4_X1 U24220 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n21327), .A3(n14849), 
        .A4(n21326), .ZN(n21328) );
  NAND4_X1 U24221 ( .A1(n21331), .A2(n21330), .A3(n21329), .A4(n21328), .ZN(
        n21342) );
  NOR4_X1 U24222 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_10__3__SCAN_IN), .A3(P2_INSTQUEUE_REG_9__7__SCAN_IN), 
        .A4(BUF2_REG_27__SCAN_IN), .ZN(n21335) );
  NOR4_X1 U24223 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_10__2__SCAN_IN), .A3(P2_INSTQUEUE_REG_6__2__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n21334) );
  NOR4_X1 U24224 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(DATAI_25_), .A4(DATAI_16_), 
        .ZN(n21333) );
  NOR4_X1 U24225 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(P1_EAX_REG_14__SCAN_IN), .ZN(
        n21332) );
  NAND4_X1 U24226 ( .A1(n21335), .A2(n21334), .A3(n21333), .A4(n21332), .ZN(
        n21341) );
  NOR4_X1 U24227 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_9__3__SCAN_IN), .A3(P3_INSTQUEUE_REG_8__5__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n21339) );
  NOR4_X1 U24228 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_3__2__SCAN_IN), .A3(P3_INSTQUEUE_REG_10__4__SCAN_IN), 
        .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n21338) );
  NOR4_X1 U24229 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .A3(P2_REIP_REG_5__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21337) );
  NOR4_X1 U24230 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A4(P3_REIP_REG_11__SCAN_IN), .ZN(
        n21336) );
  NAND4_X1 U24231 ( .A1(n21339), .A2(n21338), .A3(n21337), .A4(n21336), .ZN(
        n21340) );
  NOR4_X1 U24232 ( .A1(n21343), .A2(n21342), .A3(n21341), .A4(n21340), .ZN(
        n21344) );
  NAND4_X1 U24233 ( .A1(n21347), .A2(n21346), .A3(n21345), .A4(n21344), .ZN(
        n21348) );
  XNOR2_X1 U24234 ( .A(n21349), .B(n21348), .ZN(P1_U2863) );
  NOR2_X2 U12719 ( .A1(n17111), .A2(n18548), .ZN(n12371) );
  NOR2_X2 U13118 ( .A1(n17319), .A2(n18217), .ZN(n17318) );
  NOR2_X2 U12183 ( .A1(n18227), .A2(n17327), .ZN(n17326) );
  NOR2_X2 U12187 ( .A1(n17340), .A2(n18240), .ZN(n17339) );
  AND2_X2 U11204 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12868) );
  INV_X2 U11255 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13387) );
  AND2_X1 U15695 ( .A1(n12440), .A2(n12870), .ZN(n13960) );
  BUF_X2 U12477 ( .A(n15059), .Z(n15083) );
  CLKBUF_X1 U11387 ( .A(n12590), .Z(n13564) );
  NOR2_X1 U12197 ( .A1(n18295), .A2(n21230), .ZN(n18269) );
  NOR2_X1 U15517 ( .A1(n18289), .A2(n17366), .ZN(n17365) );
  BUF_X2 U11139 ( .A(n13271), .Z(n15149) );
  CLKBUF_X1 U11160 ( .A(n12560), .Z(n14992) );
  INV_X1 U11167 ( .A(n19880), .ZN(n11026) );
  CLKBUF_X3 U11185 ( .A(n12560), .Z(n15085) );
  CLKBUF_X1 U11191 ( .A(n12792), .Z(n12793) );
  NAND2_X1 U11192 ( .A1(n9755), .A2(n12552), .ZN(n12590) );
  NOR2_X1 U11203 ( .A1(n18336), .A2(n18337), .ZN(n12357) );
  CLKBUF_X2 U11727 ( .A(n15265), .Z(n9693) );
  OR2_X1 U11920 ( .A1(n17301), .A2(n18194), .ZN(n10184) );
  NOR2_X1 U12186 ( .A1(n17309), .A2(n18203), .ZN(n17308) );
  NOR2_X1 U12294 ( .A1(n18273), .A2(n17358), .ZN(n17357) );
  NOR2_X1 U12420 ( .A1(n17402), .A2(n17403), .ZN(n17401) );
  NOR2_X1 U12510 ( .A1(n18481), .A2(n18492), .ZN(n17511) );
  INV_X1 U12730 ( .A(n12362), .ZN(n10186) );
  NOR2_X1 U12898 ( .A1(n18191), .A2(n18184), .ZN(n17149) );
  AND2_X1 U13396 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n9836) );
  AND2_X1 U15162 ( .A1(n18423), .A2(n18729), .ZN(n18462) );
  CLKBUF_X1 U15513 ( .A(n10159), .Z(n9712) );
endmodule

