

module b20_C_AntiSAT_k_256_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, ADD_1068_U4, ADD_1068_U55, 
        ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, 
        ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, 
        ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, 
        ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, 
        P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, 
        P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, 
        P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, 
        P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, 
        P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, 
        P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, 
        P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, 
        P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, 
        P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, 
        P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, 
        P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, 
        P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598;

  OAI21_X1 U5023 ( .B1(n9689), .B2(n9540), .A(n9541), .ZN(n9673) );
  AOI21_X1 U5024 ( .B1(n5785), .B2(n4522), .A(n5119), .ZN(n8063) );
  NAND2_X1 U5025 ( .A1(n7588), .A2(n9371), .ZN(n7589) );
  OAI22_X1 U5026 ( .A1(n7410), .A2(n7409), .B1(n7408), .B2(n7443), .ZN(n7411)
         );
  XNOR2_X1 U5027 ( .A(n5344), .B(n5343), .ZN(n6622) );
  XNOR2_X1 U5028 ( .A(n5330), .B(n5329), .ZN(n6534) );
  NAND4_X1 U5029 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n9482)
         );
  BUF_X2 U5030 ( .A(n5955), .Z(n6490) );
  AND2_X1 U5031 ( .A1(n9967), .A2(n9962), .ZN(n5955) );
  CLKBUF_X3 U5032 ( .A(n5935), .Z(n6210) );
  OR2_X1 U5033 ( .A1(n5791), .A2(n4868), .ZN(n4866) );
  INV_X1 U5034 ( .A(n8338), .ZN(n8344) );
  INV_X1 U5036 ( .A(n7012), .ZN(n7142) );
  INV_X4 U5037 ( .A(n7142), .ZN(n8124) );
  INV_X1 U5038 ( .A(n5218), .ZN(n5548) );
  INV_X1 U5039 ( .A(n9798), .ZN(n9549) );
  NAND2_X1 U5040 ( .A1(n6382), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6448) );
  INV_X1 U5041 ( .A(n5975), .ZN(n6401) );
  CLKBUF_X2 U5042 ( .A(n5953), .Z(n6269) );
  INV_X1 U5043 ( .A(n9789), .ZN(n9774) );
  INV_X1 U5044 ( .A(n9806), .ZN(n9616) );
  OAI21_X1 U5045 ( .B1(n7797), .B2(n4833), .A(n4563), .ZN(n9271) );
  NAND2_X1 U5046 ( .A1(n7623), .A2(n7622), .ZN(n7762) );
  OAI21_X1 U5047 ( .B1(n9957), .B2(n5853), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5854) );
  NAND2_X1 U5048 ( .A1(n4940), .A2(n5328), .ZN(n5344) );
  NAND2_X1 U5049 ( .A1(n5762), .A2(n6785), .ZN(n6507) );
  AND2_X1 U5050 ( .A1(n4715), .A2(n4714), .ZN(n7410) );
  NAND2_X1 U5051 ( .A1(n5400), .A2(n5399), .ZN(n7882) );
  NAND2_X1 U5052 ( .A1(n9967), .A2(n5857), .ZN(n9224) );
  NAND4_X2 U5053 ( .A1(n5915), .A2(n5914), .A3(n5913), .A4(n5912), .ZN(n6672)
         );
  NAND2_X1 U5054 ( .A1(n6028), .A2(n6027), .ZN(n7355) );
  AOI21_X1 U5055 ( .B1(n8730), .B2(n8862), .A(n8729), .ZN(n8894) );
  INV_X1 U5056 ( .A(n10128), .ZN(n10126) );
  NAND2_X2 U5057 ( .A1(n5308), .A2(n5307), .ZN(n5310) );
  NAND2_X2 U5058 ( .A1(n5291), .A2(n5290), .ZN(n5308) );
  XNOR2_X2 U5059 ( .A(n5871), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6416) );
  NOR2_X2 U5060 ( .A1(n5242), .A2(n4744), .ZN(n5009) );
  AOI21_X2 U5061 ( .B1(n6230), .B2(n5881), .A(n5872), .ZN(n6248) );
  INV_X2 U5062 ( .A(n9967), .ZN(n5858) );
  XNOR2_X2 U5063 ( .A(n4774), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5145) );
  OAI21_X2 U5064 ( .B1(n8543), .B2(n4927), .A(n4926), .ZN(n8590) );
  XNOR2_X2 U5065 ( .A(n4929), .B(n4820), .ZN(n8543) );
  XNOR2_X2 U5066 ( .A(n5692), .B(n5691), .ZN(n7939) );
  INV_X2 U5067 ( .A(n6264), .ZN(n6736) );
  XNOR2_X1 U5068 ( .A(n8230), .B(n7649), .ZN(n8228) );
  OAI21_X2 U5069 ( .B1(n6830), .B2(n6847), .A(n6976), .ZN(n6831) );
  OAI211_X2 U5070 ( .C1(n4916), .C2(n4915), .A(n4914), .B(n6847), .ZN(n6976)
         );
  AND2_X1 U5071 ( .A1(n5048), .A2(n6363), .ZN(n9093) );
  OAI21_X1 U5072 ( .B1(n8458), .B2(n4535), .A(n8503), .ZN(n8462) );
  AOI21_X1 U5073 ( .B1(n9786), .B2(n10100), .A(n9785), .ZN(n9904) );
  AND2_X1 U5074 ( .A1(n5083), .A2(n5084), .ZN(n9570) );
  AOI21_X1 U5075 ( .B1(n9552), .B2(n4687), .A(n4690), .ZN(n4689) );
  NAND2_X1 U5076 ( .A1(n9598), .A2(n9551), .ZN(n5085) );
  AOI21_X1 U5077 ( .B1(n5082), .B2(n5081), .A(n4567), .ZN(n5078) );
  OR2_X1 U5078 ( .A1(n9438), .A2(n9232), .ZN(n9236) );
  NAND2_X1 U5079 ( .A1(n9524), .A2(n9521), .ZN(n9438) );
  AOI21_X1 U5080 ( .B1(n9012), .B2(n5331), .A(n5735), .ZN(n8719) );
  NAND2_X1 U5081 ( .A1(n5092), .A2(n9538), .ZN(n9689) );
  OR2_X1 U5082 ( .A1(n4838), .A2(n4836), .ZN(n4835) );
  NAND2_X1 U5083 ( .A1(n6400), .A2(n6399), .ZN(n9591) );
  OR2_X1 U5084 ( .A1(n8635), .A2(n4925), .ZN(n4924) );
  OAI21_X1 U5085 ( .B1(n9714), .B2(n9533), .A(n9535), .ZN(n9701) );
  OAI21_X1 U5086 ( .B1(n8827), .B2(n8151), .A(n8283), .ZN(n8079) );
  XNOR2_X1 U5087 ( .A(n5656), .B(n5669), .ZN(n7920) );
  NAND2_X1 U5088 ( .A1(n6323), .A2(n6322), .ZN(n9831) );
  NAND2_X1 U5089 ( .A1(n6195), .A2(n6194), .ZN(n9527) );
  NAND2_X1 U5090 ( .A1(n6169), .A2(n6168), .ZN(n9892) );
  NAND2_X1 U5091 ( .A1(n5416), .A2(n5415), .ZN(n7966) );
  NAND2_X1 U5092 ( .A1(n5438), .A2(n5437), .ZN(n5455) );
  NAND2_X1 U5093 ( .A1(n6083), .A2(n6082), .ZN(n7489) );
  NAND2_X1 U5094 ( .A1(n5382), .A2(n5381), .ZN(n8246) );
  NAND2_X1 U5095 ( .A1(n6622), .A2(n6024), .ZN(n6065) );
  AND2_X1 U5096 ( .A1(n4922), .A2(n4921), .ZN(n7817) );
  NAND2_X1 U5097 ( .A1(n6007), .A2(n6006), .ZN(n7274) );
  OAI21_X1 U5098 ( .B1(n7185), .B2(n7247), .A(n7251), .ZN(n7186) );
  INV_X1 U5099 ( .A(n6853), .ZN(n7204) );
  INV_X2 U5100 ( .A(n5918), .ZN(n6408) );
  AND2_X1 U5102 ( .A1(n4557), .A2(n4701), .ZN(n9242) );
  INV_X2 U5103 ( .A(n7467), .ZN(n8862) );
  INV_X1 U5104 ( .A(n6529), .ZN(n7022) );
  NAND4_X1 U5105 ( .A1(n5928), .A2(n5927), .A3(n5926), .A4(n5925), .ZN(n9483)
         );
  BUF_X1 U5106 ( .A(n5891), .Z(n9465) );
  AND2_X1 U5107 ( .A1(n6432), .A2(n5888), .ZN(n5891) );
  AND2_X2 U5108 ( .A1(n8357), .A2(n8191), .ZN(n8338) );
  XNOR2_X1 U5109 ( .A(n5750), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8357) );
  CLKBUF_X1 U5110 ( .A(n6284), .Z(n8017) );
  OR2_X1 U5111 ( .A1(n5887), .A2(n5886), .ZN(n5888) );
  OR2_X1 U5112 ( .A1(n5975), .A2(n5911), .ZN(n5913) );
  INV_X4 U5113 ( .A(n5736), .ZN(n5184) );
  OAI21_X1 U5114 ( .B1(n5885), .B2(n5870), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5871) );
  NAND2_X4 U5115 ( .A1(n9962), .A2(n5858), .ZN(n5975) );
  INV_X2 U5116 ( .A(n8698), .ZN(n8670) );
  NAND2_X1 U5117 ( .A1(n9008), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5144) );
  OR2_X1 U5118 ( .A1(n5878), .A2(n5872), .ZN(n5879) );
  XNOR2_X1 U5119 ( .A(n5854), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5857) );
  XNOR2_X1 U5120 ( .A(n5154), .B(n5153), .ZN(n6785) );
  INV_X2 U5121 ( .A(n9959), .ZN(n9964) );
  NOR2_X1 U5122 ( .A1(n5173), .A2(n5893), .ZN(n5175) );
  BUF_X4 U5123 ( .A(n8004), .Z(n7998) );
  OAI21_X1 U5124 ( .B1(n5910), .B2(n5167), .A(n5166), .ZN(n5168) );
  CLKBUF_X1 U5125 ( .A(n5910), .Z(n6511) );
  NAND2_X2 U5126 ( .A1(n4911), .A2(n4909), .ZN(n6789) );
  INV_X2 U5127 ( .A(n5910), .ZN(n8004) );
  NAND2_X2 U5128 ( .A1(n4825), .A2(n4824), .ZN(n5910) );
  NOR2_X1 U5129 ( .A1(n4910), .A2(n4661), .ZN(n4909) );
  NAND2_X1 U5130 ( .A1(n4826), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4825) );
  AND2_X1 U5131 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  AND3_X1 U5132 ( .A1(n5847), .A2(n5867), .A3(n5846), .ZN(n5851) );
  XNOR2_X1 U5133 ( .A(n5165), .B(n5164), .ZN(n8062) );
  AND2_X1 U5134 ( .A1(n4717), .A2(n5165), .ZN(n5188) );
  INV_X1 U5135 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5151) );
  INV_X4 U5136 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U5137 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5138 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5841) );
  NOR2_X1 U5139 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5842) );
  INV_X1 U5140 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5830) );
  INV_X2 U5141 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8388) );
  OAI22_X2 U5142 ( .A1(n5310), .A2(n4939), .B1(n4543), .B2(n4941), .ZN(n5350)
         );
  NAND4_X2 U5143 ( .A1(n6389), .A2(n6388), .A3(n6387), .A4(n6386), .ZN(n9806)
         );
  BUF_X4 U5144 ( .A(n5939), .Z(n4517) );
  INV_X1 U5145 ( .A(n5981), .ZN(n5939) );
  NAND2_X4 U5146 ( .A1(n6065), .A2(n6064), .ZN(n7347) );
  NAND4_X2 U5147 ( .A1(n6405), .A2(n6404), .A3(n6403), .A4(n6402), .ZN(n9797)
         );
  AOI21_X2 U5148 ( .B1(n9040), .B2(n9037), .A(n9036), .ZN(n9126) );
  OAI21_X2 U5149 ( .B1(n9158), .B2(n9161), .A(n9159), .ZN(n9040) );
  AOI21_X4 U5150 ( .B1(n9711), .B2(n9710), .A(n9274), .ZN(n9512) );
  NAND2_X1 U5151 ( .A1(n4805), .A2(n4809), .ZN(n4811) );
  AND2_X1 U5152 ( .A1(n4806), .A2(n4584), .ZN(n4805) );
  NOR2_X1 U5153 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4716) );
  AND2_X1 U5154 ( .A1(n9465), .A2(n9453), .ZN(n9282) );
  NOR2_X1 U5155 ( .A1(n4679), .A2(n4678), .ZN(n4677) );
  NAND2_X1 U5156 ( .A1(n9373), .A2(n9372), .ZN(n4679) );
  NOR2_X1 U5157 ( .A1(n4680), .A2(n9368), .ZN(n4678) );
  OAI21_X1 U5158 ( .B1(n8290), .B2(n4769), .A(n4768), .ZN(n8292) );
  NAND2_X1 U5159 ( .A1(n8283), .A2(n8344), .ZN(n4768) );
  NAND2_X1 U5160 ( .A1(n9242), .A2(n6672), .ZN(n9243) );
  NOR2_X1 U5161 ( .A1(n8580), .A2(n4819), .ZN(n4659) );
  NAND2_X1 U5162 ( .A1(n5814), .A2(n5813), .ZN(n5110) );
  OR2_X1 U5163 ( .A1(n6224), .A2(n6247), .ZN(n5032) );
  INV_X1 U5164 ( .A(n5473), .ZN(n5477) );
  INV_X1 U5165 ( .A(n7861), .ZN(n5107) );
  OR2_X1 U5166 ( .A1(n7860), .A2(n7886), .ZN(n7861) );
  INV_X1 U5167 ( .A(n4918), .ZN(n4915) );
  NAND2_X1 U5168 ( .A1(n4917), .A2(n4918), .ZN(n4914) );
  NAND2_X1 U5169 ( .A1(n4815), .A2(n4813), .ZN(n6834) );
  NOR2_X1 U5170 ( .A1(n4814), .A2(n4816), .ZN(n4813) );
  NOR2_X1 U5171 ( .A1(n6842), .A2(n6833), .ZN(n4816) );
  OR2_X1 U5172 ( .A1(n8599), .A2(n8598), .ZN(n4818) );
  INV_X1 U5173 ( .A(n5739), .ZN(n7419) );
  NAND2_X1 U5174 ( .A1(n5810), .A2(n5809), .ZN(n6462) );
  OAI21_X1 U5175 ( .B1(n8757), .B2(n4984), .A(n5688), .ZN(n4983) );
  OAI21_X1 U5176 ( .B1(n8769), .B2(n5647), .A(n5646), .ZN(n5648) );
  AND2_X1 U5177 ( .A1(n8303), .A2(n4578), .ZN(n4880) );
  OR2_X1 U5178 ( .A1(n8978), .A2(n8116), .ZN(n8299) );
  OR2_X1 U5179 ( .A1(n8393), .A2(n8492), .ZN(n8293) );
  OR2_X1 U5180 ( .A1(n8441), .A2(n8101), .ZN(n8288) );
  NOR2_X1 U5181 ( .A1(n4858), .A2(n5782), .ZN(n4857) );
  INV_X1 U5182 ( .A(n8257), .ZN(n4858) );
  NOR2_X1 U5183 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5135) );
  NOR2_X1 U5184 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5134) );
  XNOR2_X1 U5185 ( .A(n4619), .B(n5918), .ZN(n5919) );
  INV_X1 U5186 ( .A(n4538), .ZN(n5088) );
  INV_X1 U5187 ( .A(n9513), .ZN(n4841) );
  AND2_X1 U5188 ( .A1(n5062), .A2(n4579), .ZN(n5057) );
  XNOR2_X1 U5189 ( .A(n7993), .B(n7994), .ZN(n7992) );
  AND2_X1 U5190 ( .A1(n5693), .A2(n5678), .ZN(n5691) );
  AOI21_X1 U5191 ( .B1(n4963), .B2(n5516), .A(n4593), .ZN(n4962) );
  NAND2_X1 U5192 ( .A1(n4948), .A2(n4946), .ZN(n5500) );
  NOR2_X1 U5193 ( .A1(n4589), .A2(n4947), .ZN(n4946) );
  OR2_X1 U5194 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  NOR2_X1 U5195 ( .A1(n5329), .A2(n4945), .ZN(n4944) );
  INV_X1 U5196 ( .A(n5309), .ZN(n4945) );
  AOI21_X1 U5197 ( .B1(n4723), .B2(n8419), .A(n4721), .ZN(n4720) );
  INV_X1 U5198 ( .A(n8420), .ZN(n4721) );
  INV_X1 U5199 ( .A(n8529), .ZN(n8447) );
  OAI21_X1 U5200 ( .B1(n8182), .B2(n4887), .A(n4886), .ZN(n4885) );
  NOR2_X1 U5201 ( .A1(n8183), .A2(n7636), .ZN(n4886) );
  NAND2_X1 U5202 ( .A1(n8348), .A2(n4560), .ZN(n4887) );
  NOR2_X1 U5203 ( .A1(n8177), .A2(n8350), .ZN(n4765) );
  NAND2_X1 U5204 ( .A1(n6983), .A2(n4665), .ZN(n6835) );
  OR2_X1 U5205 ( .A1(n6834), .A2(n6847), .ZN(n4665) );
  NOR2_X1 U5206 ( .A1(n7256), .A2(n7191), .ZN(n7192) );
  AND2_X1 U5207 ( .A1(n7190), .A2(n7197), .ZN(n7191) );
  INV_X1 U5208 ( .A(n7258), .ZN(n7256) );
  NAND2_X1 U5209 ( .A1(n4811), .A2(n7247), .ZN(n7258) );
  NAND2_X1 U5210 ( .A1(n4629), .A2(n4628), .ZN(n7819) );
  AND2_X1 U5211 ( .A1(n4650), .A2(n4649), .ZN(n7907) );
  AND2_X1 U5212 ( .A1(n4651), .A2(n4583), .ZN(n4649) );
  NAND2_X1 U5213 ( .A1(n4667), .A2(n4666), .ZN(n4823) );
  INV_X1 U5214 ( .A(n7912), .ZN(n4666) );
  INV_X1 U5215 ( .A(n7913), .ZN(n4667) );
  NOR2_X1 U5216 ( .A1(n8632), .A2(n8847), .ZN(n4925) );
  OAI21_X1 U5217 ( .B1(n8739), .B2(n4969), .A(n4967), .ZN(n4970) );
  INV_X1 U5218 ( .A(n4968), .ZN(n4967) );
  OAI21_X1 U5219 ( .B1(n4969), .B2(n8738), .A(n5720), .ZN(n4968) );
  NAND2_X1 U5220 ( .A1(n4544), .A2(n5000), .ZN(n4999) );
  AND2_X1 U5221 ( .A1(n4998), .A2(n5370), .ZN(n4997) );
  NAND2_X1 U5222 ( .A1(n4862), .A2(n4861), .ZN(n4860) );
  NOR2_X1 U5223 ( .A1(n8152), .A2(n4757), .ZN(n4861) );
  NAND2_X1 U5224 ( .A1(n6507), .A2(n6511), .ZN(n5354) );
  AND2_X1 U5225 ( .A1(n5755), .A2(n5754), .ZN(n7467) );
  NOR2_X1 U5226 ( .A1(n8150), .A2(n4878), .ZN(n4877) );
  INV_X1 U5227 ( .A(n8308), .ZN(n4878) );
  NAND2_X1 U5228 ( .A1(n4985), .A2(n4552), .ZN(n8818) );
  NAND2_X1 U5229 ( .A1(n4988), .A2(n4989), .ZN(n4987) );
  INV_X1 U5230 ( .A(n6507), .ZN(n5547) );
  NAND2_X1 U5231 ( .A1(n4775), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4774) );
  NAND2_X1 U5232 ( .A1(n5007), .A2(n4747), .ZN(n5805) );
  NOR2_X1 U5233 ( .A1(n5242), .A2(n4742), .ZN(n4747) );
  NAND2_X1 U5234 ( .A1(n4743), .A2(n4883), .ZN(n4742) );
  INV_X1 U5235 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U5236 ( .A1(n4611), .A2(n4555), .ZN(n5045) );
  NAND2_X1 U5237 ( .A1(n6002), .A2(n5987), .ZN(n5024) );
  NAND2_X1 U5238 ( .A1(n5906), .A2(n5902), .ZN(n6647) );
  AOI21_X1 U5239 ( .B1(n4695), .B2(n6736), .A(n6437), .ZN(n4694) );
  AOI21_X1 U5240 ( .B1(n9399), .B2(n9272), .A(n4830), .ZN(n4829) );
  INV_X1 U5241 ( .A(n9400), .ZN(n4830) );
  NAND2_X1 U5242 ( .A1(n9739), .A2(n6264), .ZN(n6756) );
  NAND2_X1 U5243 ( .A1(n8384), .A2(n8383), .ZN(n8382) );
  OR2_X1 U5244 ( .A1(n7149), .A2(n7150), .ZN(n4715) );
  NAND2_X1 U5245 ( .A1(n9330), .A2(n9329), .ZN(n9333) );
  NOR2_X1 U5246 ( .A1(n8279), .A2(n8344), .ZN(n4772) );
  NAND2_X1 U5247 ( .A1(n9369), .A2(n4677), .ZN(n4676) );
  NAND2_X1 U5248 ( .A1(n4751), .A2(n8301), .ZN(n4750) );
  NOR2_X1 U5249 ( .A1(n5788), .A2(n4755), .ZN(n4754) );
  INV_X1 U5250 ( .A(n8295), .ZN(n4755) );
  NOR2_X1 U5251 ( .A1(n9664), .A2(n4559), .ZN(n4699) );
  OAI21_X1 U5252 ( .B1(n4779), .B2(n4539), .A(n4778), .ZN(n8333) );
  NOR2_X1 U5253 ( .A1(n8326), .A2(n8327), .ZN(n4778) );
  NAND2_X1 U5254 ( .A1(n4951), .A2(n4954), .ZN(n4949) );
  INV_X1 U5255 ( .A(n7980), .ZN(n4710) );
  NOR2_X1 U5256 ( .A1(n9181), .A2(n9087), .ZN(n5069) );
  INV_X1 U5257 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U5258 ( .A1(n4730), .A2(n7559), .ZN(n4729) );
  INV_X1 U5259 ( .A(n5101), .ZN(n4730) );
  NAND2_X1 U5260 ( .A1(n5108), .A2(n6915), .ZN(n7012) );
  AND2_X1 U5261 ( .A1(n6914), .A2(n6913), .ZN(n6915) );
  NAND2_X1 U5262 ( .A1(n5110), .A2(n4718), .ZN(n5108) );
  NOR2_X1 U5263 ( .A1(n5115), .A2(n4596), .ZN(n4718) );
  NAND2_X1 U5264 ( .A1(n6789), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4792) );
  OAI21_X1 U5265 ( .B1(n6978), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6977), .ZN(
        n4902) );
  NOR2_X1 U5266 ( .A1(n7817), .A2(n4920), .ZN(n7818) );
  AND2_X1 U5267 ( .A1(n7821), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U5268 ( .A1(n5719), .A2(n4971), .ZN(n4969) );
  NOR2_X1 U5269 ( .A1(n5218), .A2(n6518), .ZN(n4850) );
  NAND2_X1 U5270 ( .A1(n8539), .A2(n7011), .ZN(n8202) );
  OAI211_X1 U5271 ( .C1(n6507), .C2(n8062), .A(n5180), .B(n5179), .ZN(n5181)
         );
  OR2_X1 U5272 ( .A1(n5354), .A2(n6514), .ZN(n5180) );
  AND2_X1 U5273 ( .A1(n8310), .A2(n8311), .ZN(n8302) );
  AND2_X1 U5274 ( .A1(n8842), .A2(n4975), .ZN(n4974) );
  NAND2_X1 U5275 ( .A1(n4976), .A2(n8857), .ZN(n4975) );
  INV_X1 U5276 ( .A(n5472), .ZN(n4976) );
  NAND2_X1 U5277 ( .A1(n8996), .A2(n5495), .ZN(n8276) );
  NAND2_X1 U5278 ( .A1(n5452), .A2(n5451), .ZN(n8858) );
  NOR2_X1 U5279 ( .A1(n4856), .A2(n4853), .ZN(n4852) );
  INV_X1 U5280 ( .A(n8239), .ZN(n4853) );
  INV_X1 U5281 ( .A(n4857), .ZN(n4856) );
  INV_X1 U5282 ( .A(n8256), .ZN(n4855) );
  OR2_X1 U5283 ( .A1(n8246), .A2(n7877), .ZN(n8239) );
  AND2_X1 U5284 ( .A1(n4605), .A2(n6463), .ZN(n7096) );
  INV_X1 U5285 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U5286 ( .A1(n5133), .A2(n4745), .ZN(n4744) );
  INV_X1 U5287 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5133) );
  INV_X1 U5288 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4745) );
  AND2_X1 U5289 ( .A1(n5112), .A2(n5747), .ZN(n5111) );
  NAND2_X1 U5290 ( .A1(n5040), .A2(n5042), .ZN(n5037) );
  INV_X1 U5291 ( .A(n5041), .ZN(n5040) );
  NAND2_X1 U5292 ( .A1(n4564), .A2(n4698), .ZN(n4697) );
  NOR2_X1 U5293 ( .A1(n9318), .A2(n9525), .ZN(n4698) );
  OAI21_X1 U5294 ( .B1(n5090), .B2(n5088), .A(n4551), .ZN(n5087) );
  NOR2_X1 U5295 ( .A1(n9629), .A2(n5091), .ZN(n5090) );
  INV_X1 U5296 ( .A(n9547), .ZN(n5091) );
  OR2_X1 U5297 ( .A1(n9831), .A2(n9680), .ZN(n9515) );
  INV_X1 U5298 ( .A(n9269), .ZN(n4833) );
  OR2_X1 U5299 ( .A1(n9872), .A2(n9880), .ZN(n9390) );
  AND2_X1 U5300 ( .A1(n7798), .A2(n9380), .ZN(n4834) );
  NOR2_X1 U5301 ( .A1(n5069), .A2(n9300), .ZN(n5068) );
  INV_X1 U5302 ( .A(n5069), .ZN(n5066) );
  OR2_X1 U5303 ( .A1(n9702), .A2(n9842), .ZN(n9693) );
  NAND2_X1 U5304 ( .A1(n4831), .A2(n9273), .ZN(n9720) );
  INV_X1 U5305 ( .A(n9732), .ZN(n4831) );
  OAI21_X1 U5306 ( .B1(n7992), .B2(n10488), .A(n7997), .ZN(n8012) );
  NAND2_X1 U5307 ( .A1(n5594), .A2(n5593), .ZN(n4935) );
  NOR2_X1 U5308 ( .A1(n5609), .A2(n4938), .ZN(n4937) );
  INV_X1 U5309 ( .A(n5593), .ZN(n4938) );
  AOI21_X1 U5310 ( .B1(n4958), .B2(n4957), .A(n4956), .ZN(n4955) );
  INV_X1 U5311 ( .A(n5559), .ZN(n4956) );
  INV_X1 U5312 ( .A(n4963), .ZN(n4957) );
  OR2_X1 U5313 ( .A1(n5475), .A2(n5474), .ZN(n4948) );
  NAND2_X1 U5314 ( .A1(n5397), .A2(n5396), .ZN(n5431) );
  OAI21_X1 U5315 ( .B1(n7998), .B2(n5236), .A(n5235), .ZN(n5237) );
  NAND2_X1 U5316 ( .A1(n5910), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4965) );
  AND2_X1 U5317 ( .A1(n7557), .A2(n8536), .ZN(n5101) );
  NAND2_X1 U5318 ( .A1(n7981), .A2(n7980), .ZN(n4713) );
  OR2_X1 U5319 ( .A1(n7650), .A2(n7649), .ZN(n5100) );
  OR2_X1 U5320 ( .A1(n7556), .A2(n4729), .ZN(n7648) );
  OR2_X1 U5321 ( .A1(n5225), .A2(n6790), .ZN(n5149) );
  NAND2_X1 U5322 ( .A1(n4708), .A2(n4706), .ZN(n8429) );
  AND2_X1 U5323 ( .A1(n8099), .A2(n4707), .ZN(n4706) );
  NAND2_X1 U5324 ( .A1(n4519), .A2(n4712), .ZN(n4707) );
  INV_X1 U5325 ( .A(n8535), .ZN(n7735) );
  INV_X1 U5326 ( .A(n4729), .ZN(n4728) );
  INV_X1 U5327 ( .A(n5100), .ZN(n4726) );
  NAND2_X1 U5328 ( .A1(n5096), .A2(n5099), .ZN(n5094) );
  NAND2_X1 U5329 ( .A1(n8120), .A2(n8413), .ZN(n8473) );
  OR2_X1 U5330 ( .A1(n7981), .A2(n4712), .ZN(n4705) );
  NAND2_X1 U5331 ( .A1(n4713), .A2(n4711), .ZN(n8094) );
  AND2_X1 U5332 ( .A1(n8174), .A2(n4612), .ZN(n8175) );
  OAI21_X1 U5333 ( .B1(n8337), .B2(n8336), .A(n5121), .ZN(n4767) );
  AND2_X1 U5334 ( .A1(n7425), .A2(n7424), .ZN(n8147) );
  AND3_X1 U5335 ( .A1(n5588), .A2(n5587), .A3(n5586), .ZN(n8116) );
  AND3_X1 U5336 ( .A1(n5573), .A2(n5572), .A3(n5571), .ZN(n8412) );
  AND4_X1 U5337 ( .A1(n5406), .A2(n5405), .A3(n5404), .A4(n5403), .ZN(n7948)
         );
  INV_X1 U5338 ( .A(n5225), .ZN(n5756) );
  OR2_X1 U5339 ( .A1(n5225), .A2(n7230), .ZN(n5187) );
  XNOR2_X1 U5340 ( .A(n6803), .B(n8062), .ZN(n8051) );
  OR2_X1 U5341 ( .A1(n8062), .A2(n6778), .ZN(n4907) );
  NOR2_X1 U5342 ( .A1(n10439), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U5343 ( .A1(n4907), .A2(n4905), .ZN(n8056) );
  NOR2_X1 U5344 ( .A1(n4906), .A2(n7110), .ZN(n4905) );
  INV_X1 U5345 ( .A(n6779), .ZN(n4906) );
  NAND2_X1 U5346 ( .A1(n5188), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6779) );
  OAI21_X1 U5347 ( .B1(n6789), .B2(n6780), .A(n4908), .ZN(n10132) );
  NAND2_X1 U5348 ( .A1(n6789), .A2(n6780), .ZN(n4908) );
  NAND2_X1 U5349 ( .A1(n6789), .A2(n7230), .ZN(n6788) );
  NAND2_X1 U5350 ( .A1(n4808), .A2(n4807), .ZN(n4806) );
  INV_X1 U5351 ( .A(n6983), .ZN(n4808) );
  OR2_X1 U5352 ( .A1(n6835), .A2(n4530), .ZN(n4809) );
  NAND2_X1 U5353 ( .A1(n6834), .A2(n6847), .ZN(n6983) );
  INV_X1 U5354 ( .A(n4794), .ZN(n4793) );
  NAND2_X1 U5355 ( .A1(n7535), .A2(n4801), .ZN(n4795) );
  NOR2_X1 U5356 ( .A1(n7391), .A2(n7381), .ZN(n7520) );
  OAI21_X1 U5357 ( .B1(n7538), .B2(n7537), .A(n4781), .ZN(n7541) );
  OR2_X1 U5358 ( .A1(n7536), .A2(n7535), .ZN(n4781) );
  NAND2_X1 U5359 ( .A1(n7541), .A2(n7540), .ZN(n7820) );
  OR2_X1 U5360 ( .A1(n7520), .A2(n4923), .ZN(n4922) );
  AND2_X1 U5361 ( .A1(n7521), .A2(n7535), .ZN(n4923) );
  AND2_X1 U5362 ( .A1(n4669), .A2(n4668), .ZN(n7913) );
  NAND2_X1 U5363 ( .A1(n7909), .A2(n7910), .ZN(n4668) );
  XNOR2_X1 U5364 ( .A(n4821), .B(n4820), .ZN(n8553) );
  INV_X1 U5365 ( .A(n4821), .ZN(n8577) );
  NOR2_X1 U5366 ( .A1(n8553), .A2(n8552), .ZN(n8579) );
  AND2_X1 U5367 ( .A1(n4627), .A2(n4626), .ZN(n8608) );
  NAND2_X1 U5368 ( .A1(n8597), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4626) );
  INV_X1 U5369 ( .A(n8590), .ZN(n4627) );
  NAND2_X1 U5370 ( .A1(n4818), .A2(n4541), .ZN(n4664) );
  AND2_X1 U5371 ( .A1(n4664), .A2(n4663), .ZN(n8637) );
  INV_X1 U5372 ( .A(n8627), .ZN(n4663) );
  NAND2_X1 U5373 ( .A1(n5808), .A2(n5828), .ZN(n6926) );
  NOR2_X1 U5374 ( .A1(n5812), .A2(n7943), .ZN(n5828) );
  AOI21_X1 U5375 ( .B1(n4787), .B2(n10136), .A(n4785), .ZN(n8705) );
  NAND2_X1 U5376 ( .A1(n4786), .A2(n8702), .ZN(n4785) );
  XNOR2_X1 U5377 ( .A(n4789), .B(n4788), .ZN(n4787) );
  NOR2_X1 U5378 ( .A1(n8666), .A2(n4639), .ZN(n4637) );
  NAND2_X1 U5379 ( .A1(n8700), .A2(n8690), .ZN(n4639) );
  AOI21_X1 U5380 ( .B1(n4867), .B2(n8324), .A(n4526), .ZN(n4865) );
  NAND2_X1 U5381 ( .A1(n4860), .A2(n4523), .ZN(n7774) );
  AND2_X1 U5382 ( .A1(n8244), .A2(n8250), .ZN(n8164) );
  NAND2_X1 U5383 ( .A1(n5776), .A2(n4863), .ZN(n4862) );
  NOR2_X1 U5384 ( .A1(n7465), .A2(n4864), .ZN(n4863) );
  AND4_X1 U5385 ( .A1(n5340), .A2(n5339), .A3(n5338), .A4(n5337), .ZN(n7886)
         );
  NAND2_X1 U5386 ( .A1(n7430), .A2(n5305), .ZN(n7466) );
  AND3_X1 U5387 ( .A1(n5267), .A2(n5266), .A3(n5265), .ZN(n7309) );
  OR2_X1 U5388 ( .A1(n5218), .A2(n6515), .ZN(n5266) );
  OR2_X1 U5389 ( .A1(n5218), .A2(n6510), .ZN(n5219) );
  OR2_X1 U5390 ( .A1(n5354), .A2(n6513), .ZN(n4845) );
  INV_X1 U5391 ( .A(n4983), .ZN(n4982) );
  AND2_X1 U5392 ( .A1(n8149), .A2(n8186), .ZN(n8748) );
  INV_X1 U5393 ( .A(n4875), .ZN(n4874) );
  OAI21_X1 U5394 ( .B1(n4877), .B2(n4876), .A(n8764), .ZN(n4875) );
  INV_X1 U5395 ( .A(n8302), .ZN(n8775) );
  NOR2_X1 U5396 ( .A1(n4991), .A2(n5535), .ZN(n4990) );
  INV_X1 U5397 ( .A(n5558), .ZN(n4991) );
  INV_X1 U5398 ( .A(n5534), .ZN(n4992) );
  NAND2_X1 U5399 ( .A1(n5515), .A2(n5514), .ZN(n8828) );
  OAI21_X1 U5400 ( .B1(n8063), .B2(n5786), .A(n8288), .ZN(n8827) );
  NAND2_X1 U5401 ( .A1(n8858), .A2(n5472), .ZN(n8863) );
  NAND2_X1 U5402 ( .A1(n7955), .A2(n8266), .ZN(n5006) );
  OR2_X1 U5403 ( .A1(n7882), .A2(n7948), .ZN(n8257) );
  AND2_X1 U5404 ( .A1(n6935), .A2(n8338), .ZN(n8865) );
  INV_X1 U5405 ( .A(n8727), .ZN(n8866) );
  NAND2_X1 U5406 ( .A1(n7096), .A2(n6467), .ZN(n6938) );
  INV_X1 U5407 ( .A(n7483), .ZN(n7840) );
  OR2_X1 U5408 ( .A1(n8357), .A2(n8191), .ZN(n8476) );
  INV_X1 U5409 ( .A(n5805), .ZN(n5155) );
  AND2_X1 U5410 ( .A1(n5156), .A2(n5153), .ZN(n5012) );
  NOR2_X1 U5411 ( .A1(n4741), .A2(n4739), .ZN(n5007) );
  INV_X1 U5412 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5797) );
  OAI21_X1 U5413 ( .B1(n5796), .B2(n5113), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5798) );
  NAND2_X1 U5414 ( .A1(n5830), .A2(n5114), .ZN(n5113) );
  NAND2_X1 U5415 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n5114) );
  NAND2_X1 U5416 ( .A1(n4736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U5417 ( .A1(n5521), .A2(n5112), .ZN(n4736) );
  XNOR2_X1 U5418 ( .A(n5546), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8693) );
  NOR2_X1 U5419 ( .A1(n5380), .A2(n5379), .ZN(n7823) );
  XNOR2_X1 U5420 ( .A(n5243), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6842) );
  AND2_X1 U5421 ( .A1(n5188), .A2(n5189), .ZN(n4661) );
  AND2_X1 U5422 ( .A1(n9007), .A2(n5189), .ZN(n4910) );
  NAND2_X1 U5423 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  XNOR2_X1 U5424 ( .A(n5999), .B(n6481), .ZN(n6001) );
  NAND2_X1 U5425 ( .A1(n6907), .A2(n5987), .ZN(n5025) );
  NAND2_X1 U5426 ( .A1(n5034), .A2(n9105), .ZN(n5033) );
  NAND2_X1 U5427 ( .A1(n6224), .A2(n6225), .ZN(n5034) );
  CLKBUF_X1 U5428 ( .A(n6906), .Z(n6907) );
  XNOR2_X1 U5429 ( .A(n5938), .B(n6408), .ZN(n5944) );
  NOR2_X1 U5430 ( .A1(n5044), .A2(n5047), .ZN(n5043) );
  OR2_X1 U5431 ( .A1(n9194), .A2(n9195), .ZN(n5047) );
  INV_X1 U5432 ( .A(n5046), .ZN(n5044) );
  NAND2_X1 U5433 ( .A1(n4693), .A2(n6739), .ZN(n4692) );
  INV_X1 U5434 ( .A(n9458), .ZN(n4693) );
  AND2_X1 U5435 ( .A1(n7938), .A2(n6430), .ZN(n5875) );
  OR2_X1 U5436 ( .A1(n9635), .A2(n4891), .ZN(n4534) );
  NAND2_X1 U5437 ( .A1(n4892), .A2(n9907), .ZN(n4891) );
  NAND2_X1 U5438 ( .A1(n9911), .A2(n9602), .ZN(n5084) );
  NAND2_X1 U5439 ( .A1(n5085), .A2(n5080), .ZN(n5083) );
  AND2_X1 U5440 ( .A1(n9569), .A2(n5084), .ZN(n5082) );
  AND2_X1 U5441 ( .A1(n9518), .A2(n9422), .ZN(n9629) );
  NAND2_X1 U5442 ( .A1(n9548), .A2(n5090), .ZN(n5089) );
  NOR2_X1 U5443 ( .A1(n9664), .A2(n4839), .ZN(n4838) );
  NAND2_X1 U5444 ( .A1(n4842), .A2(n4841), .ZN(n4840) );
  NAND2_X1 U5445 ( .A1(n4840), .A2(n9514), .ZN(n9665) );
  NAND2_X1 U5446 ( .A1(n9515), .A2(n9286), .ZN(n9664) );
  INV_X1 U5447 ( .A(n5063), .ZN(n5062) );
  OAI21_X1 U5448 ( .B1(n9304), .B2(n5064), .A(n7786), .ZN(n5063) );
  NAND2_X1 U5449 ( .A1(n7797), .A2(n4834), .ZN(n9270) );
  NAND2_X1 U5450 ( .A1(n9379), .A2(n9384), .ZN(n9304) );
  AND2_X1 U5451 ( .A1(n9371), .A2(n9372), .ZN(n7493) );
  NAND2_X1 U5452 ( .A1(n7352), .A2(n7351), .ZN(n7491) );
  NAND2_X1 U5453 ( .A1(n9292), .A2(n6997), .ZN(n5074) );
  NOR2_X1 U5454 ( .A1(n5075), .A2(n5073), .ZN(n5072) );
  NAND2_X1 U5455 ( .A1(n7159), .A2(n7165), .ZN(n7158) );
  AND2_X1 U5456 ( .A1(n9242), .A2(n6963), .ZN(n6965) );
  NAND2_X1 U5457 ( .A1(n6511), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4703) );
  NAND2_X1 U5458 ( .A1(n8019), .A2(n8018), .ZN(n9777) );
  NAND2_X1 U5459 ( .A1(n6252), .A2(n6251), .ZN(n9534) );
  AND3_X1 U5460 ( .A1(n5934), .A2(n5933), .A3(n5932), .ZN(n6853) );
  NAND2_X1 U5461 ( .A1(n7083), .A2(n10077), .ZN(n10100) );
  AND2_X1 U5462 ( .A1(n6434), .A2(n9459), .ZN(n10082) );
  AND3_X1 U5463 ( .A1(n6757), .A2(n6756), .A3(n6755), .ZN(n6764) );
  OR2_X1 U5464 ( .A1(n8012), .A2(n8011), .ZN(n8014) );
  XNOR2_X1 U5465 ( .A(n5708), .B(n5723), .ZN(n9016) );
  XNOR2_X1 U5466 ( .A(n5899), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U5467 ( .A1(n5898), .A2(n5897), .ZN(n5899) );
  XNOR2_X1 U5468 ( .A(n5636), .B(n5635), .ZN(n7857) );
  NAND2_X1 U5469 ( .A1(n5876), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U5470 ( .A1(n4961), .A2(n4962), .ZN(n5561) );
  NAND2_X1 U5471 ( .A1(n5517), .A2(n4963), .ZN(n4961) );
  OR2_X1 U5472 ( .A1(n4943), .A2(n4543), .ZN(n4939) );
  INV_X1 U5473 ( .A(n4942), .ZN(n4941) );
  AND4_X1 U5474 ( .A1(n5424), .A2(n5423), .A3(n5422), .A4(n5421), .ZN(n8261)
         );
  AND2_X1 U5475 ( .A1(n5104), .A2(n7873), .ZN(n5103) );
  OR2_X1 U5476 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  AND4_X1 U5477 ( .A1(n5471), .A2(n5470), .A3(n5469), .A4(n5468), .ZN(n8436)
         );
  NAND2_X1 U5478 ( .A1(n7312), .A2(n7323), .ZN(n4714) );
  NAND2_X1 U5479 ( .A1(n8382), .A2(n4556), .ZN(n7149) );
  INV_X1 U5480 ( .A(n8795), .ZN(n8480) );
  AND2_X1 U5481 ( .A1(n5526), .A2(n5525), .ZN(n8497) );
  AND4_X1 U5482 ( .A1(n5556), .A2(n5555), .A3(n5554), .A4(n5553), .ZN(n8492)
         );
  NAND2_X1 U5483 ( .A1(n5667), .A2(n5666), .ZN(n8770) );
  INV_X1 U5484 ( .A(n8116), .ZN(n8821) );
  INV_X1 U5485 ( .A(n8412), .ZN(n8810) );
  INV_X1 U5486 ( .A(n8492), .ZN(n8830) );
  INV_X1 U5487 ( .A(n8101), .ZN(n8845) );
  INV_X1 U5488 ( .A(n8436), .ZN(n8844) );
  INV_X1 U5489 ( .A(n8261), .ZN(n8530) );
  INV_X1 U5490 ( .A(n7323), .ZN(n8537) );
  NAND2_X1 U5491 ( .A1(n8030), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n8050) );
  NOR2_X1 U5492 ( .A1(n6790), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6791) );
  NOR2_X1 U5493 ( .A1(n6814), .A2(n4784), .ZN(n6811) );
  AND2_X1 U5494 ( .A1(n6809), .A2(n4671), .ZN(n4784) );
  NAND2_X1 U5495 ( .A1(n6811), .A2(n6810), .ZN(n6840) );
  OR2_X1 U5496 ( .A1(n7816), .A2(n5383), .ZN(n4669) );
  XNOR2_X1 U5497 ( .A(n7907), .B(n7823), .ZN(n7816) );
  XNOR2_X1 U5498 ( .A(n8608), .B(n8625), .ZN(n8591) );
  NOR2_X1 U5499 ( .A1(n8657), .A2(n8656), .ZN(n8659) );
  INV_X1 U5500 ( .A(n4924), .ZN(n8655) );
  OAI21_X1 U5501 ( .B1(n5768), .B2(n7467), .A(n5767), .ZN(n8716) );
  NOR2_X1 U5502 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  XNOR2_X1 U5503 ( .A(n4970), .B(n8326), .ZN(n5768) );
  NOR2_X1 U5504 ( .A1(n8368), .A2(n8727), .ZN(n5765) );
  AND2_X1 U5505 ( .A1(n8736), .A2(n8323), .ZN(n8731) );
  AND2_X1 U5506 ( .A1(n8753), .A2(n4617), .ZN(n4616) );
  OR2_X1 U5507 ( .A1(n10161), .A2(n8751), .ZN(n4617) );
  NAND2_X1 U5508 ( .A1(n5600), .A2(n5599), .ZN(n8801) );
  OR2_X1 U5509 ( .A1(n5218), .A2(n7744), .ZN(n5599) );
  INV_X1 U5510 ( .A(n10160), .ZN(n8854) );
  AND2_X1 U5511 ( .A1(n8146), .A2(n8145), .ZN(n8886) );
  OR2_X1 U5512 ( .A1(n5218), .A2(n10472), .ZN(n8145) );
  NAND2_X1 U5513 ( .A1(n5658), .A2(n5657), .ZN(n8959) );
  OR2_X1 U5514 ( .A1(n5218), .A2(n7921), .ZN(n5657) );
  INV_X1 U5515 ( .A(n7943), .ZN(n6725) );
  INV_X1 U5516 ( .A(n9058), .ZN(n5052) );
  NAND2_X1 U5517 ( .A1(n5955), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U5518 ( .A1(n9186), .A2(n9482), .ZN(n5054) );
  NAND2_X1 U5519 ( .A1(n9215), .A2(n6672), .ZN(n5053) );
  XNOR2_X1 U5520 ( .A(n5944), .B(n5942), .ZN(n6678) );
  CLKBUF_X1 U5521 ( .A(n6676), .Z(n6677) );
  NAND2_X1 U5522 ( .A1(n9282), .A2(n6651), .ZN(n9877) );
  AND2_X1 U5523 ( .A1(n8010), .A2(n8009), .ZN(n9898) );
  NAND2_X1 U5524 ( .A1(n4762), .A2(n4759), .ZN(n8238) );
  NAND2_X1 U5525 ( .A1(n4760), .A2(n8338), .ZN(n4759) );
  NAND2_X1 U5526 ( .A1(n4763), .A2(n8344), .ZN(n4762) );
  NAND2_X1 U5527 ( .A1(n8238), .A2(n4756), .ZN(n8241) );
  NOR2_X1 U5528 ( .A1(n4758), .A2(n4757), .ZN(n4756) );
  INV_X1 U5529 ( .A(n8236), .ZN(n4758) );
  NAND2_X1 U5530 ( .A1(n8243), .A2(n7747), .ZN(n8249) );
  NAND2_X1 U5531 ( .A1(n4771), .A2(n4770), .ZN(n8290) );
  NAND2_X1 U5532 ( .A1(n8282), .A2(n8344), .ZN(n4770) );
  NAND2_X1 U5533 ( .A1(n4773), .A2(n4772), .ZN(n4771) );
  NAND2_X1 U5534 ( .A1(n4570), .A2(n8338), .ZN(n4769) );
  NAND2_X1 U5535 ( .A1(n4676), .A2(n4675), .ZN(n9375) );
  AOI21_X1 U5536 ( .B1(n4677), .B2(n4680), .A(n7621), .ZN(n4675) );
  OAI211_X1 U5537 ( .C1(n4752), .C2(n8338), .A(n4749), .B(n8802), .ZN(n4748)
         );
  AOI21_X1 U5538 ( .B1(n8294), .B2(n4754), .A(n4753), .ZN(n4752) );
  INV_X1 U5539 ( .A(n8299), .ZN(n4753) );
  NAND2_X1 U5540 ( .A1(n8321), .A2(n8748), .ZN(n4780) );
  AND2_X1 U5541 ( .A1(n4700), .A2(n4527), .ZN(n9419) );
  NAND2_X1 U5542 ( .A1(n4688), .A2(n9440), .ZN(n4687) );
  INV_X1 U5543 ( .A(n9443), .ZN(n4690) );
  OR2_X1 U5544 ( .A1(n5428), .A2(n5427), .ZN(n5432) );
  AOI21_X1 U5545 ( .B1(n8328), .B2(n8331), .A(n8330), .ZN(n8343) );
  OR2_X1 U5546 ( .A1(n8887), .A2(n8339), .ZN(n4930) );
  NOR2_X1 U5547 ( .A1(n6793), .A2(n4817), .ZN(n4814) );
  AND2_X1 U5548 ( .A1(n8667), .A2(n4790), .ZN(n8672) );
  NAND2_X1 U5549 ( .A1(n8669), .A2(n8668), .ZN(n4790) );
  INV_X1 U5550 ( .A(n5831), .ZN(n6914) );
  OAI21_X1 U5551 ( .B1(n6022), .B2(n5042), .A(n7133), .ZN(n5041) );
  NAND2_X1 U5552 ( .A1(n5041), .A2(n5039), .ZN(n5038) );
  NAND2_X1 U5553 ( .A1(n6022), .A2(n5042), .ZN(n5039) );
  OR2_X1 U5554 ( .A1(n9655), .A2(n9666), .ZN(n9417) );
  NAND2_X1 U5555 ( .A1(n9366), .A2(n9355), .ZN(n9340) );
  NAND2_X1 U5556 ( .A1(n4950), .A2(n4600), .ZN(n5734) );
  INV_X1 U5557 ( .A(n5691), .ZN(n4954) );
  AOI21_X1 U5558 ( .B1(n5691), .B2(n4953), .A(n4952), .ZN(n4951) );
  INV_X1 U5559 ( .A(n5673), .ZN(n4953) );
  INV_X1 U5560 ( .A(n5693), .ZN(n4952) );
  INV_X1 U5561 ( .A(n5591), .ZN(n5592) );
  INV_X1 U5562 ( .A(n5560), .ZN(n4960) );
  INV_X1 U5563 ( .A(SI_19_), .ZN(n5541) );
  INV_X1 U5564 ( .A(n5497), .ZN(n5498) );
  INV_X1 U5565 ( .A(n5478), .ZN(n4947) );
  INV_X1 U5566 ( .A(SI_15_), .ZN(n5476) );
  INV_X1 U5567 ( .A(n8123), .ZN(n4723) );
  AND2_X1 U5568 ( .A1(n8431), .A2(n8432), .ZN(n8099) );
  INV_X1 U5569 ( .A(n8465), .ZN(n5099) );
  AOI21_X1 U5570 ( .B1(n8465), .B2(n5098), .A(n5097), .ZN(n5096) );
  NAND2_X1 U5571 ( .A1(n4711), .A2(n4710), .ZN(n4709) );
  NAND2_X1 U5572 ( .A1(n8886), .A2(n8887), .ZN(n8181) );
  OR3_X1 U5573 ( .A1(n8172), .A2(n8819), .A3(n8807), .ZN(n8173) );
  OR4_X1 U5574 ( .A1(n8842), .A2(n8268), .A3(n8852), .A4(n8169), .ZN(n8170) );
  NOR2_X1 U5575 ( .A1(n8738), .A2(n4613), .ZN(n4612) );
  NAND2_X1 U5576 ( .A1(n8748), .A2(n4547), .ZN(n4613) );
  INV_X1 U5577 ( .A(n4930), .ZN(n8335) );
  OR2_X1 U5578 ( .A1(n8345), .A2(n5131), .ZN(n8336) );
  NAND2_X1 U5579 ( .A1(n4930), .A2(n5745), .ZN(n5131) );
  OAI21_X1 U5580 ( .B1(n6783), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6784), .ZN(
        n4917) );
  NAND2_X1 U5581 ( .A1(n4919), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U5582 ( .A1(n4904), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4903) );
  OAI211_X1 U5583 ( .C1(n4900), .C2(n4899), .A(n4898), .B(n7247), .ZN(n7251)
         );
  INV_X1 U5584 ( .A(n4903), .ZN(n4899) );
  NAND2_X1 U5585 ( .A1(n4902), .A2(n4903), .ZN(n4898) );
  NAND2_X1 U5586 ( .A1(n4823), .A2(n4822), .ZN(n4821) );
  NAND2_X1 U5587 ( .A1(n8551), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U5588 ( .A1(n4656), .A2(n4657), .ZN(n8624) );
  NAND2_X1 U5589 ( .A1(n4660), .A2(n8582), .ZN(n4657) );
  NAND2_X1 U5590 ( .A1(n4658), .A2(n4659), .ZN(n4656) );
  NAND2_X1 U5591 ( .A1(n8687), .A2(n8658), .ZN(n4643) );
  AOI21_X1 U5592 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n4789) );
  INV_X1 U5593 ( .A(n8701), .ZN(n4788) );
  NAND2_X1 U5594 ( .A1(n8704), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4786) );
  NOR2_X1 U5595 ( .A1(n8637), .A2(n4662), .ZN(n8660) );
  NOR2_X1 U5596 ( .A1(n8632), .A2(n10489), .ZN(n4662) );
  NAND2_X1 U5597 ( .A1(n4870), .A2(n8323), .ZN(n4869) );
  INV_X1 U5598 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10330) );
  INV_X1 U5599 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7525) );
  AOI21_X1 U5600 ( .B1(n5001), .B2(n5324), .A(n4521), .ZN(n5000) );
  NAND2_X1 U5601 ( .A1(n5201), .A2(n7218), .ZN(n4978) );
  INV_X1 U5602 ( .A(n5201), .ZN(n4979) );
  NAND2_X1 U5603 ( .A1(n5183), .A2(n6916), .ZN(n8199) );
  NAND2_X1 U5604 ( .A1(n5182), .A2(n5181), .ZN(n8198) );
  INV_X1 U5605 ( .A(n5115), .ZN(n5109) );
  NAND2_X1 U5606 ( .A1(n8737), .A2(n8186), .ZN(n4870) );
  AND2_X1 U5607 ( .A1(n8310), .A2(n4880), .ZN(n4872) );
  INV_X1 U5608 ( .A(n4990), .ZN(n4988) );
  OR2_X1 U5609 ( .A1(n5811), .A2(n5827), .ZN(n6467) );
  INV_X1 U5610 ( .A(n4744), .ZN(n4743) );
  INV_X1 U5611 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5143) );
  INV_X1 U5612 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5747) );
  NOR2_X1 U5613 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4740) );
  NOR2_X1 U5614 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(n5125), .ZN(n5112) );
  OR2_X1 U5615 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5125) );
  INV_X1 U5616 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U5617 ( .A1(n5521), .A2(n5520), .ZN(n5746) );
  NAND2_X1 U5618 ( .A1(n5008), .A2(n5009), .ZN(n5519) );
  AND2_X1 U5619 ( .A1(n5140), .A2(n5139), .ZN(n5008) );
  NOR2_X1 U5620 ( .A1(n6298), .A2(n5031), .ZN(n5027) );
  NAND2_X1 U5621 ( .A1(n5028), .A2(n5030), .ZN(n9046) );
  NAND2_X1 U5622 ( .A1(n5987), .A2(n7020), .ZN(n5020) );
  NAND2_X1 U5623 ( .A1(n5885), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5887) );
  INV_X1 U5624 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5881) );
  INV_X1 U5625 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5882) );
  NOR2_X1 U5626 ( .A1(n4894), .A2(n4895), .ZN(n4892) );
  OR2_X1 U5627 ( .A1(n9591), .A2(n9622), .ZN(n4894) );
  NOR2_X1 U5628 ( .A1(n9738), .A2(n9534), .ZN(n4897) );
  OAI21_X1 U5629 ( .B1(n9340), .B2(n9337), .A(n9361), .ZN(n7360) );
  INV_X1 U5630 ( .A(n7360), .ZN(n9299) );
  OR2_X1 U5631 ( .A1(n7347), .A2(n7489), .ZN(n4889) );
  INV_X1 U5632 ( .A(n6997), .ZN(n5075) );
  INV_X1 U5633 ( .A(n6995), .ZN(n5073) );
  AND2_X1 U5634 ( .A1(n9347), .A2(n9343), .ZN(n9292) );
  NOR2_X1 U5635 ( .A1(n9635), .A2(n4890), .ZN(n9587) );
  INV_X1 U5636 ( .A(n4892), .ZN(n4890) );
  AND2_X1 U5637 ( .A1(n5730), .A2(n5697), .ZN(n5725) );
  AND2_X1 U5638 ( .A1(n5673), .A2(n5655), .ZN(n5669) );
  NOR2_X1 U5639 ( .A1(n5539), .A2(n4964), .ZN(n4963) );
  INV_X1 U5640 ( .A(n5518), .ZN(n4964) );
  OR2_X1 U5641 ( .A1(n6147), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6166) );
  OAI21_X1 U5642 ( .B1(n4944), .B2(n4943), .A(n5343), .ZN(n4942) );
  INV_X1 U5643 ( .A(n5328), .ZN(n4943) );
  OR2_X1 U5644 ( .A1(n6042), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6081) );
  CLKBUF_X1 U5645 ( .A(n5970), .Z(n5988) );
  NAND2_X1 U5646 ( .A1(n5910), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5166) );
  INV_X1 U5647 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4827) );
  XNOR2_X1 U5648 ( .A(n5157), .B(n5156), .ZN(n5762) );
  NAND2_X1 U5649 ( .A1(n5805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5157) );
  AND2_X1 U5650 ( .A1(n7864), .A2(n5106), .ZN(n5105) );
  OR2_X1 U5651 ( .A1(n7730), .A2(n5107), .ZN(n5106) );
  NAND2_X1 U5652 ( .A1(n5105), .A2(n5107), .ZN(n5104) );
  AND2_X1 U5653 ( .A1(n8498), .A2(n8127), .ZN(n8420) );
  NAND2_X1 U5654 ( .A1(n7862), .A2(n7861), .ZN(n7926) );
  NAND2_X1 U5655 ( .A1(n8128), .A2(n8499), .ZN(n8502) );
  INV_X1 U5656 ( .A(n5762), .ZN(n8698) );
  AND4_X1 U5657 ( .A1(n5389), .A2(n5388), .A3(n5387), .A4(n5386), .ZN(n7877)
         );
  NAND2_X1 U5658 ( .A1(n8050), .A2(n8051), .ZN(n8049) );
  NAND2_X1 U5659 ( .A1(n5188), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6792) );
  NAND2_X1 U5660 ( .A1(n8056), .A2(n6779), .ZN(n10131) );
  NAND2_X1 U5661 ( .A1(n10147), .A2(n10146), .ZN(n10145) );
  NAND2_X1 U5662 ( .A1(n4913), .A2(n4916), .ZN(n6828) );
  INV_X1 U5663 ( .A(n4917), .ZN(n4913) );
  NOR2_X1 U5664 ( .A1(n6818), .A2(n5202), .ZN(n6817) );
  INV_X1 U5665 ( .A(n4902), .ZN(n4901) );
  NOR2_X1 U5666 ( .A1(n6831), .A2(n7328), .ZN(n6979) );
  OR2_X1 U5667 ( .A1(n5481), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5332) );
  AOI21_X1 U5668 ( .B1(n4798), .B2(n4802), .A(n4797), .ZN(n4803) );
  NAND2_X1 U5669 ( .A1(n4800), .A2(n7387), .ZN(n4797) );
  INV_X1 U5670 ( .A(n4672), .ZN(n4800) );
  OAI21_X1 U5671 ( .B1(n7258), .B2(n7259), .A(n4804), .ZN(n4672) );
  NAND2_X1 U5672 ( .A1(n7527), .A2(n4654), .ZN(n4651) );
  OR2_X1 U5673 ( .A1(n4647), .A2(n4803), .ZN(n4650) );
  NAND2_X1 U5674 ( .A1(n4653), .A2(n4648), .ZN(n4647) );
  NOR2_X1 U5675 ( .A1(n7529), .A2(n4655), .ZN(n4648) );
  NAND2_X1 U5676 ( .A1(n7820), .A2(n4586), .ZN(n7825) );
  XNOR2_X1 U5677 ( .A(n8624), .B(n8625), .ZN(n8599) );
  INV_X1 U5678 ( .A(n4818), .ZN(n8626) );
  NAND2_X1 U5679 ( .A1(n8643), .A2(n8644), .ZN(n8645) );
  NAND2_X1 U5680 ( .A1(n8645), .A2(n8646), .ZN(n8667) );
  XNOR2_X1 U5681 ( .A(n8660), .B(n8668), .ZN(n8638) );
  NAND2_X1 U5682 ( .A1(n4642), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U5683 ( .A1(n8699), .A2(n8687), .ZN(n4641) );
  NAND2_X1 U5684 ( .A1(n4644), .A2(n4643), .ZN(n4642) );
  INV_X1 U5685 ( .A(n8699), .ZN(n4644) );
  AOI21_X1 U5686 ( .B1(n8732), .B2(n5184), .A(n5718), .ZN(n8368) );
  OR2_X1 U5687 ( .A1(n5701), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U5688 ( .A1(n5660), .A2(n5659), .ZN(n5681) );
  OR2_X1 U5689 ( .A1(n5551), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U5690 ( .A1(n5527), .A2(n10330), .ZN(n5551) );
  INV_X1 U5691 ( .A(n5528), .ZN(n5527) );
  OR2_X1 U5692 ( .A1(n5508), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U5693 ( .A1(n5488), .A2(n5487), .ZN(n5508) );
  INV_X1 U5694 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5487) );
  INV_X1 U5695 ( .A(n5489), .ZN(n5488) );
  OR2_X1 U5696 ( .A1(n5466), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5489) );
  INV_X1 U5697 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5417) );
  OR2_X1 U5698 ( .A1(n5401), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5419) );
  OR2_X1 U5699 ( .A1(n5384), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U5700 ( .A1(n4996), .A2(n5000), .ZN(n7749) );
  NAND2_X1 U5701 ( .A1(n7466), .A2(n5001), .ZN(n4996) );
  AND2_X1 U5702 ( .A1(n5361), .A2(n5360), .ZN(n7865) );
  OR2_X1 U5703 ( .A1(n5335), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U5704 ( .A1(n5003), .A2(n5323), .ZN(n7638) );
  NAND2_X1 U5705 ( .A1(n5005), .A2(n5004), .ZN(n5003) );
  INV_X1 U5706 ( .A(n7466), .ZN(n5005) );
  NAND2_X1 U5707 ( .A1(n5289), .A2(n4849), .ZN(n7413) );
  NOR2_X1 U5708 ( .A1(n4548), .A2(n4850), .ZN(n4849) );
  AND4_X1 U5709 ( .A1(n5232), .A2(n5231), .A3(n5230), .A4(n5229), .ZN(n7323)
         );
  AND2_X1 U5710 ( .A1(n8219), .A2(n8211), .ZN(n8153) );
  NAND2_X1 U5711 ( .A1(n7220), .A2(n7218), .ZN(n7219) );
  NAND2_X1 U5712 ( .A1(n4602), .A2(n7104), .ZN(n7222) );
  NAND2_X1 U5713 ( .A1(n6934), .A2(n8338), .ZN(n8727) );
  OR2_X1 U5714 ( .A1(n8038), .A2(n5794), .ZN(n7753) );
  AND2_X1 U5715 ( .A1(n8352), .A2(n8185), .ZN(n5831) );
  INV_X1 U5716 ( .A(n8737), .ZN(n8738) );
  AND2_X1 U5717 ( .A1(n8323), .A2(n8322), .ZN(n8737) );
  OR2_X1 U5718 ( .A1(n5791), .A2(n4870), .ZN(n8736) );
  NAND2_X1 U5719 ( .A1(n8756), .A2(n8757), .ZN(n8755) );
  NAND2_X1 U5720 ( .A1(n4973), .A2(n4972), .ZN(n8064) );
  AOI21_X1 U5721 ( .B1(n4974), .B2(n4977), .A(n4525), .ZN(n4972) );
  AOI21_X1 U5722 ( .B1(n4855), .B2(n4857), .A(n4571), .ZN(n4854) );
  INV_X1 U5723 ( .A(SI_22_), .ZN(n10408) );
  XNOR2_X1 U5724 ( .A(n5829), .B(n5830), .ZN(n6923) );
  NAND2_X1 U5725 ( .A1(n4881), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5154) );
  NOR2_X1 U5726 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4882) );
  OR2_X1 U5727 ( .A1(n5286), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5481) );
  OR2_X1 U5728 ( .A1(n5413), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5414) );
  NOR2_X1 U5729 ( .A1(n5242), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U5730 ( .A1(n7069), .A2(n7071), .ZN(n6023) );
  CLKBUF_X1 U5731 ( .A(n5981), .Z(n5982) );
  INV_X1 U5732 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6170) );
  INV_X1 U5733 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10357) );
  OR2_X1 U5734 ( .A1(n6363), .A2(n9092), .ZN(n5046) );
  CLKBUF_X1 U5735 ( .A(n9099), .Z(n9100) );
  OR2_X1 U5736 ( .A1(n6211), .A2(n7582), .ZN(n6235) );
  INV_X1 U5737 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6234) );
  OR2_X1 U5738 ( .A1(n9126), .A2(n9125), .ZN(n5048) );
  AND2_X1 U5739 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5992) );
  INV_X1 U5740 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6638) );
  NOR2_X1 U5741 ( .A1(n6066), .A2(n6638), .ZN(n6084) );
  OR2_X1 U5742 ( .A1(n6151), .A2(n6880), .ZN(n6171) );
  OR2_X1 U5743 ( .A1(n6129), .A2(n6128), .ZN(n6151) );
  INV_X1 U5744 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9164) );
  AND2_X1 U5745 ( .A1(n6205), .A2(n6204), .ZN(n9205) );
  NAND2_X1 U5746 ( .A1(n9220), .A2(n9448), .ZN(n9462) );
  NOR2_X1 U5747 ( .A1(n5079), .A2(n9597), .ZN(n5077) );
  INV_X1 U5748 ( .A(n5082), .ZN(n5079) );
  OR2_X1 U5749 ( .A1(n9919), .A2(n9549), .ZN(n5117) );
  INV_X1 U5750 ( .A(n5087), .ZN(n5086) );
  AND2_X1 U5751 ( .A1(n6369), .A2(n6384), .ZN(n9613) );
  INV_X1 U5752 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9127) );
  NOR2_X1 U5753 ( .A1(n6351), .A2(n9127), .ZN(n6368) );
  NAND2_X1 U5754 ( .A1(n4841), .A2(n9515), .ZN(n4837) );
  INV_X1 U5755 ( .A(n9515), .ZN(n4836) );
  NOR2_X1 U5756 ( .A1(n10357), .A2(n6268), .ZN(n6287) );
  NAND2_X1 U5757 ( .A1(n4897), .A2(n4896), .ZN(n9702) );
  NAND2_X1 U5758 ( .A1(n9749), .A2(n9944), .ZN(n9738) );
  INV_X1 U5759 ( .A(n4897), .ZN(n9715) );
  OR2_X1 U5760 ( .A1(n4834), .A2(n4833), .ZN(n4832) );
  AOI21_X1 U5761 ( .B1(n5057), .B2(n5064), .A(n4561), .ZN(n5056) );
  NAND2_X1 U5762 ( .A1(n6127), .A2(n6126), .ZN(n7616) );
  AND2_X1 U5763 ( .A1(n9374), .A2(n9373), .ZN(n7590) );
  NAND2_X1 U5764 ( .A1(n5067), .A2(n5065), .ZN(n7615) );
  NAND2_X1 U5765 ( .A1(n5070), .A2(n5066), .ZN(n5065) );
  INV_X1 U5766 ( .A(n7590), .ZN(n9303) );
  NAND2_X1 U5767 ( .A1(n6996), .A2(n6995), .ZN(n7159) );
  INV_X1 U5768 ( .A(n9292), .ZN(n7165) );
  NAND2_X1 U5769 ( .A1(n4673), .A2(n6856), .ZN(n9331) );
  NAND2_X1 U5770 ( .A1(n6854), .A2(n9244), .ZN(n4673) );
  NAND2_X1 U5771 ( .A1(n9342), .A2(n9328), .ZN(n6857) );
  AND2_X1 U5772 ( .A1(n6434), .A2(n6437), .ZN(n9739) );
  NAND2_X1 U5773 ( .A1(n6965), .A2(n6853), .ZN(n6851) );
  AND2_X1 U5774 ( .A1(n9453), .A2(n6437), .ZN(n5889) );
  NAND2_X1 U5775 ( .A1(n8016), .A2(n8015), .ZN(n9507) );
  AND2_X1 U5776 ( .A1(n9556), .A2(n9280), .ZN(n9768) );
  AND3_X1 U5777 ( .A1(n6178), .A2(n6177), .A3(n6176), .ZN(n9878) );
  INV_X1 U5778 ( .A(n9879), .ZN(n10105) );
  INV_X1 U5779 ( .A(n10100), .ZN(n10111) );
  NAND2_X1 U5780 ( .A1(n6418), .A2(n7938), .ZN(n9951) );
  INV_X1 U5781 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5019) );
  INV_X1 U5782 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U5783 ( .A1(n4674), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U5784 ( .A1(n5852), .A2(n5018), .ZN(n4674) );
  XNOR2_X1 U5785 ( .A(n5874), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U5786 ( .A1(n4936), .A2(n4933), .ZN(n5618) );
  INV_X1 U5787 ( .A(n4934), .ZN(n4933) );
  OAI21_X1 U5788 ( .B1(n5609), .B2(n4935), .A(n5610), .ZN(n4934) );
  XNOR2_X1 U5789 ( .A(n6433), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U5790 ( .A1(n6432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6433) );
  OAI21_X1 U5791 ( .B1(n5517), .B2(n5516), .A(n5518), .ZN(n5540) );
  NAND2_X1 U5792 ( .A1(n4948), .A2(n5478), .ZN(n5496) );
  NAND2_X1 U5793 ( .A1(n5350), .A2(n5349), .ZN(n5372) );
  OR2_X1 U5794 ( .A1(n5237), .A2(SI_4_), .ZN(n5238) );
  AND4_X1 U5795 ( .A1(n5275), .A2(n5274), .A3(n5273), .A4(n5272), .ZN(n7564)
         );
  NOR2_X1 U5796 ( .A1(n7556), .A2(n5101), .ZN(n7560) );
  AOI21_X1 U5797 ( .B1(n4735), .B2(n8364), .A(n8522), .ZN(n8366) );
  NAND2_X1 U5798 ( .A1(n8502), .A2(n8131), .ZN(n4735) );
  AND2_X1 U5799 ( .A1(n4713), .A2(n4542), .ZN(n7984) );
  NAND2_X1 U5800 ( .A1(n5711), .A2(n5710), .ZN(n8329) );
  OR2_X1 U5801 ( .A1(n5218), .A2(n5709), .ZN(n5710) );
  NAND2_X1 U5802 ( .A1(n7648), .A2(n5100), .ZN(n7729) );
  AND4_X1 U5803 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n7106)
         );
  AND2_X1 U5804 ( .A1(n5645), .A2(n5644), .ZN(n8425) );
  NAND2_X1 U5805 ( .A1(n8473), .A2(n4520), .ZN(n4722) );
  INV_X1 U5806 ( .A(n4724), .ZN(n7731) );
  AOI21_X1 U5807 ( .B1(n7728), .B2(n4726), .A(n4568), .ZN(n4725) );
  NAND2_X1 U5808 ( .A1(n4728), .A2(n7728), .ZN(n4727) );
  NAND2_X1 U5809 ( .A1(n7731), .A2(n7730), .ZN(n7862) );
  AND2_X1 U5810 ( .A1(n6936), .A2(n6935), .ZN(n8518) );
  NAND2_X1 U5811 ( .A1(n8398), .A2(n8464), .ZN(n5095) );
  OR2_X1 U5812 ( .A1(n7944), .A2(n7948), .ZN(n7945) );
  NOR2_X1 U5813 ( .A1(n8118), .A2(n4733), .ZN(n4732) );
  INV_X1 U5814 ( .A(n4734), .ZN(n4733) );
  AND2_X1 U5815 ( .A1(n6939), .A2(n7102), .ZN(n8482) );
  INV_X1 U5816 ( .A(n8522), .ZN(n8503) );
  NAND2_X1 U5817 ( .A1(n8094), .A2(n8093), .ZN(n8523) );
  NAND2_X1 U5818 ( .A1(n4766), .A2(n4765), .ZN(n4623) );
  NAND2_X1 U5819 ( .A1(n4885), .A2(n4884), .ZN(n8351) );
  INV_X1 U5820 ( .A(n8147), .ZN(n8710) );
  INV_X1 U5821 ( .A(n8425), .ZN(n8783) );
  NAND2_X1 U5822 ( .A1(n5628), .A2(n5627), .ZN(n8795) );
  INV_X1 U5823 ( .A(n7948), .ZN(n8531) );
  INV_X1 U5824 ( .A(n7877), .ZN(n8532) );
  NAND4_X1 U5825 ( .A1(n5303), .A2(n5302), .A3(n5301), .A4(n5300), .ZN(n7649)
         );
  INV_X1 U5826 ( .A(n7564), .ZN(n8536) );
  AND3_X1 U5827 ( .A1(n5185), .A2(n5186), .A3(n5187), .ZN(n4777) );
  NAND2_X1 U5828 ( .A1(n5184), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4776) );
  CLKBUF_X1 U5829 ( .A(n6916), .Z(n8540) );
  OR2_X2 U5830 ( .A1(n6926), .A2(n6726), .ZN(n8679) );
  NAND2_X1 U5831 ( .A1(n4907), .A2(n6779), .ZN(n8054) );
  INV_X1 U5832 ( .A(n4812), .ZN(n6798) );
  OAI21_X1 U5833 ( .B1(n6820), .B2(n6794), .A(n6795), .ZN(n4812) );
  NAND2_X1 U5834 ( .A1(n6840), .A2(n4783), .ZN(n6844) );
  OR2_X1 U5835 ( .A1(n6841), .A2(n6842), .ZN(n4783) );
  NAND2_X1 U5836 ( .A1(n6844), .A2(n6843), .ZN(n6971) );
  NAND2_X1 U5837 ( .A1(n4809), .A2(n4806), .ZN(n7189) );
  NAND2_X1 U5838 ( .A1(n7260), .A2(n7258), .ZN(n4799) );
  AOI21_X1 U5839 ( .B1(n7385), .B2(n7384), .A(n4782), .ZN(n7538) );
  AND2_X1 U5840 ( .A1(n7383), .A2(n7390), .ZN(n4782) );
  OR2_X1 U5841 ( .A1(n4652), .A2(n4803), .ZN(n7530) );
  NAND2_X1 U5842 ( .A1(n4653), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4652) );
  INV_X1 U5843 ( .A(n7523), .ZN(n4921) );
  INV_X1 U5844 ( .A(n4922), .ZN(n7524) );
  INV_X1 U5845 ( .A(n4823), .ZN(n8550) );
  NOR2_X1 U5846 ( .A1(n8543), .A2(n8544), .ZN(n8563) );
  NOR2_X1 U5847 ( .A1(n8579), .A2(n8580), .ZN(n8583) );
  NAND2_X1 U5848 ( .A1(n4928), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4927) );
  NAND2_X1 U5849 ( .A1(n8564), .A2(n4928), .ZN(n4926) );
  NOR2_X1 U5850 ( .A1(n8610), .A2(n8609), .ZN(n8613) );
  INV_X1 U5851 ( .A(n4664), .ZN(n8628) );
  XNOR2_X1 U5852 ( .A(n4924), .B(n8640), .ZN(n8636) );
  NAND2_X1 U5853 ( .A1(n4640), .A2(n4645), .ZN(n4634) );
  NAND2_X1 U5854 ( .A1(n8699), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U5855 ( .A1(n10149), .A2(n4533), .ZN(n4638) );
  NOR2_X1 U5856 ( .A1(n8707), .A2(n4637), .ZN(n4636) );
  AND2_X1 U5857 ( .A1(n5621), .A2(n5620), .ZN(n8788) );
  OR2_X1 U5858 ( .A1(n5218), .A2(n10354), .ZN(n5620) );
  OR2_X1 U5859 ( .A1(n8476), .A2(n10155), .ZN(n8876) );
  NAND2_X1 U5860 ( .A1(n4860), .A2(n8240), .ZN(n7748) );
  NAND2_X1 U5861 ( .A1(n4862), .A2(n8237), .ZN(n7637) );
  AND2_X1 U5862 ( .A1(n5313), .A2(n5312), .ZN(n7647) );
  AND3_X1 U5863 ( .A1(n5246), .A2(n5245), .A3(n5244), .ZN(n8220) );
  OR2_X1 U5864 ( .A1(n5218), .A2(n5236), .ZN(n5245) );
  INV_X1 U5865 ( .A(n5770), .ZN(n7477) );
  OAI21_X1 U5866 ( .B1(n7218), .B2(n7220), .A(n7219), .ZN(n10153) );
  AND2_X1 U5867 ( .A1(n8185), .A2(n8693), .ZN(n10155) );
  OR2_X1 U5868 ( .A1(n7111), .A2(n8876), .ZN(n8856) );
  INV_X1 U5869 ( .A(n8476), .ZN(n8037) );
  AND2_X1 U5870 ( .A1(n8338), .A2(n5831), .ZN(n8038) );
  AND2_X1 U5871 ( .A1(n7102), .A2(n7101), .ZN(n10160) );
  INV_X1 U5872 ( .A(n8856), .ZN(n8849) );
  NAND2_X1 U5873 ( .A1(n4931), .A2(n8148), .ZN(n8887) );
  OR2_X1 U5874 ( .A1(n5218), .A2(n8362), .ZN(n8148) );
  NAND2_X1 U5875 ( .A1(n8361), .A2(n5331), .ZN(n4931) );
  NAND2_X1 U5876 ( .A1(n8928), .A2(n8037), .ZN(n8929) );
  INV_X2 U5877 ( .A(n8884), .ZN(n8928) );
  INV_X1 U5878 ( .A(n8887), .ZN(n8940) );
  NOR2_X1 U5879 ( .A1(n5218), .A2(n9014), .ZN(n5735) );
  AND2_X1 U5880 ( .A1(n8721), .A2(n8909), .ZN(n5793) );
  INV_X1 U5881 ( .A(n8329), .ZN(n8944) );
  OR2_X1 U5882 ( .A1(n5218), .A2(n5698), .ZN(n5699) );
  NAND2_X1 U5883 ( .A1(n5680), .A2(n5679), .ZN(n8953) );
  OR2_X1 U5884 ( .A1(n5218), .A2(n7941), .ZN(n5679) );
  INV_X1 U5885 ( .A(n4873), .ZN(n8765) );
  AOI21_X1 U5886 ( .B1(n4879), .B2(n4877), .A(n4876), .ZN(n4873) );
  NAND2_X1 U5887 ( .A1(n5638), .A2(n5637), .ZN(n8965) );
  OR2_X1 U5888 ( .A1(n5218), .A2(n8076), .ZN(n5637) );
  NAND2_X1 U5889 ( .A1(n4879), .A2(n8308), .ZN(n8776) );
  INV_X1 U5890 ( .A(n8788), .ZN(n8971) );
  NAND2_X1 U5891 ( .A1(n8910), .A2(n8303), .ZN(n8780) );
  NAND2_X1 U5892 ( .A1(n5583), .A2(n5582), .ZN(n8978) );
  OR2_X1 U5893 ( .A1(n5218), .A2(n10369), .ZN(n5582) );
  NAND2_X1 U5894 ( .A1(n5565), .A2(n5564), .ZN(n8984) );
  OR2_X1 U5895 ( .A1(n5218), .A2(n5563), .ZN(n5564) );
  NAND2_X1 U5896 ( .A1(n4986), .A2(n4989), .ZN(n8820) );
  NAND2_X1 U5897 ( .A1(n4995), .A2(n4990), .ZN(n4986) );
  NAND2_X1 U5898 ( .A1(n5550), .A2(n5549), .ZN(n8393) );
  NAND2_X1 U5899 ( .A1(n4993), .A2(n5534), .ZN(n8080) );
  NAND2_X1 U5900 ( .A1(n4995), .A2(n4994), .ZN(n4993) );
  INV_X1 U5901 ( .A(n8497), .ZN(n8989) );
  NAND2_X1 U5902 ( .A1(n5507), .A2(n5506), .ZN(n8441) );
  INV_X1 U5903 ( .A(n8440), .ZN(n8996) );
  NAND2_X1 U5904 ( .A1(n8863), .A2(n8857), .ZN(n8843) );
  NAND2_X1 U5905 ( .A1(n10580), .A2(n8037), .ZN(n9001) );
  NAND2_X1 U5906 ( .A1(n5443), .A2(n5442), .ZN(n7982) );
  NAND2_X1 U5907 ( .A1(n5006), .A2(n8263), .ZN(n7971) );
  NAND2_X1 U5908 ( .A1(n4859), .A2(n8257), .ZN(n7954) );
  NAND2_X1 U5909 ( .A1(n7843), .A2(n8256), .ZN(n4859) );
  INV_X1 U5910 ( .A(n9001), .ZN(n8995) );
  INV_X2 U5911 ( .A(n10578), .ZN(n10580) );
  INV_X1 U5912 ( .A(n6733), .ZN(n6726) );
  AND2_X1 U5913 ( .A1(n5012), .A2(n5011), .ZN(n5010) );
  INV_X1 U5914 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5011) );
  INV_X1 U5915 ( .A(n5158), .ZN(n8363) );
  INV_X1 U5916 ( .A(n5145), .ZN(n9015) );
  NAND2_X1 U5917 ( .A1(n5805), .A2(n5806), .ZN(n7943) );
  NAND2_X1 U5918 ( .A1(n5801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5802) );
  OR2_X1 U5919 ( .A1(n5798), .A2(n5797), .ZN(n5799) );
  INV_X1 U5920 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10354) );
  INV_X1 U5921 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7744) );
  INV_X1 U5922 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10369) );
  INV_X1 U5923 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7335) );
  INV_X1 U5924 ( .A(n8693), .ZN(n8352) );
  INV_X1 U5925 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7079) );
  INV_X1 U5926 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6945) );
  NOR2_X1 U5927 ( .A1(n6511), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9021) );
  INV_X1 U5928 ( .A(n7917), .ZN(n8551) );
  INV_X1 U5929 ( .A(n6973), .ZN(n6847) );
  INV_X1 U5930 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5132) );
  OR2_X1 U5931 ( .A1(n4912), .A2(n5188), .ZN(n4911) );
  NAND2_X1 U5932 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4912) );
  NAND2_X1 U5933 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5164) );
  INV_X1 U5934 ( .A(n6182), .ZN(n4620) );
  INV_X1 U5935 ( .A(n9822), .ZN(n9680) );
  CLKBUF_X1 U5936 ( .A(n6716), .Z(n6717) );
  OR2_X1 U5937 ( .A1(n6413), .A2(n6414), .ZN(n4625) );
  INV_X1 U5938 ( .A(n5014), .ZN(n5013) );
  CLKBUF_X1 U5939 ( .A(n9066), .Z(n9067) );
  CLKBUF_X1 U5940 ( .A(n9081), .Z(n9082) );
  NAND2_X1 U5941 ( .A1(n5045), .A2(n5046), .ZN(n9196) );
  NAND2_X1 U5942 ( .A1(n6907), .A2(n5022), .ZN(n7019) );
  INV_X1 U5943 ( .A(n5024), .ZN(n5022) );
  INV_X1 U5944 ( .A(n5029), .ZN(n9118) );
  AOI21_X1 U5945 ( .B1(n9100), .B2(n6224), .A(n5033), .ZN(n5029) );
  CLKBUF_X1 U5946 ( .A(n6904), .Z(n6905) );
  CLKBUF_X1 U5947 ( .A(n7601), .Z(n7602) );
  CLKBUF_X1 U5948 ( .A(n7603), .Z(n7604) );
  NAND2_X1 U5949 ( .A1(n6286), .A2(n6285), .ZN(n9842) );
  CLKBUF_X1 U5950 ( .A(n9147), .Z(n9148) );
  AOI21_X1 U5951 ( .B1(n5123), .B2(n6269), .A(n6239), .ZN(n9869) );
  OR2_X1 U5952 ( .A1(n6458), .A2(n6454), .ZN(n9189) );
  CLKBUF_X1 U5953 ( .A(n7069), .Z(n7070) );
  OR2_X1 U5954 ( .A1(n6519), .A2(n5948), .ZN(n6007) );
  AND2_X1 U5955 ( .A1(n6448), .A2(n6385), .ZN(n9599) );
  OR2_X1 U5956 ( .A1(n6458), .A2(n6444), .ZN(n9209) );
  AND2_X1 U5957 ( .A1(n6459), .A2(n9557), .ZN(n9218) );
  AND2_X1 U5958 ( .A1(n6442), .A2(n6435), .ZN(n9206) );
  NAND3_X1 U5959 ( .A1(n6504), .A2(P1_STATE_REG_SCAN_IN), .A3(n6523), .ZN(
        n9219) );
  AND2_X1 U5960 ( .A1(n9457), .A2(n4692), .ZN(n4691) );
  INV_X1 U5961 ( .A(n9878), .ZN(n10106) );
  INV_X1 U5962 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5236) );
  INV_X1 U5963 ( .A(n6672), .ZN(n6752) );
  OR2_X1 U5964 ( .A1(n10033), .A2(n10032), .ZN(n10035) );
  NAND2_X1 U5965 ( .A1(n5083), .A2(n5082), .ZN(n9568) );
  INV_X1 U5966 ( .A(n9797), .ZN(n9602) );
  INV_X1 U5967 ( .A(n5089), .ZN(n9627) );
  NAND2_X1 U5968 ( .A1(n9548), .A2(n9547), .ZN(n9625) );
  NAND2_X1 U5969 ( .A1(n4838), .A2(n4840), .ZN(n9668) );
  NAND2_X1 U5970 ( .A1(n6232), .A2(n6231), .ZN(n9743) );
  NAND2_X1 U5971 ( .A1(n9270), .A2(n9269), .ZN(n9763) );
  NAND2_X1 U5972 ( .A1(n5060), .A2(n5059), .ZN(n5058) );
  NAND2_X1 U5973 ( .A1(n5061), .A2(n7761), .ZN(n7787) );
  NAND2_X1 U5974 ( .A1(n7759), .A2(n9304), .ZN(n5061) );
  NAND2_X1 U5975 ( .A1(n6150), .A2(n6149), .ZN(n7760) );
  NAND2_X1 U5976 ( .A1(n7491), .A2(n7490), .ZN(n7587) );
  OR2_X1 U5977 ( .A1(n6962), .A2(n6264), .ZN(n9740) );
  NAND2_X1 U5978 ( .A1(n7158), .A2(n6997), .ZN(n6998) );
  INV_X1 U5979 ( .A(n9740), .ZN(n10053) );
  INV_X1 U5980 ( .A(n9767), .ZN(n10059) );
  INV_X1 U5981 ( .A(n9752), .ZN(n10050) );
  NAND2_X1 U5982 ( .A1(n4702), .A2(n5949), .ZN(n4701) );
  OAI21_X1 U5983 ( .B1(n6514), .B2(n5910), .A(n4703), .ZN(n4702) );
  OR2_X1 U5984 ( .A1(n10063), .A2(n4606), .ZN(n9752) );
  INV_X2 U5985 ( .A(n10056), .ZN(n10063) );
  OR2_X1 U5986 ( .A1(n6756), .A2(n9219), .ZN(n9557) );
  NAND2_X1 U5987 ( .A1(n10105), .A2(n6672), .ZN(n10069) );
  INV_X1 U5988 ( .A(n9889), .ZN(n9819) );
  AND2_X2 U5989 ( .A1(n6764), .A2(n6759), .ZN(n10128) );
  INV_X1 U5990 ( .A(n9507), .ZN(n9902) );
  OAI211_X1 U5991 ( .C1(n9778), .C2(n10068), .A(n9779), .B(n9780), .ZN(n9903)
         );
  INV_X1 U5992 ( .A(n9578), .ZN(n9907) );
  INV_X1 U5993 ( .A(n9591), .ZN(n9911) );
  INV_X1 U5994 ( .A(n9233), .ZN(n9915) );
  INV_X1 U5995 ( .A(n9622), .ZN(n9919) );
  INV_X1 U5996 ( .A(n9743), .ZN(n9944) );
  NAND2_X1 U5997 ( .A1(n10119), .A2(n10082), .ZN(n9948) );
  XNOR2_X1 U5998 ( .A(n8008), .B(n8007), .ZN(n9960) );
  NAND2_X1 U5999 ( .A1(n8014), .A2(n8003), .ZN(n8008) );
  INV_X1 U6000 ( .A(n5857), .ZN(n9962) );
  CLKBUF_X1 U6001 ( .A(n6540), .Z(n6541) );
  XNOR2_X1 U6002 ( .A(n5898), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7938) );
  INV_X1 U6003 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10438) );
  NOR2_X1 U6004 ( .A1(n6511), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9959) );
  INV_X1 U6005 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7646) );
  INV_X1 U6006 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7334) );
  INV_X1 U6007 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10338) );
  INV_X1 U6008 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10453) );
  INV_X1 U6009 ( .A(n7036), .ZN(n7374) );
  INV_X1 U6010 ( .A(n5197), .ZN(n5194) );
  INV_X1 U6011 ( .A(n4715), .ZN(n7311) );
  NAND2_X1 U6012 ( .A1(n10143), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U6013 ( .A1(n8050), .A2(n4609), .ZN(n8031) );
  INV_X1 U6014 ( .A(n4669), .ZN(n7908) );
  XNOR2_X1 U6015 ( .A(n8659), .B(n4646), .ZN(n8686) );
  INV_X1 U6016 ( .A(n4615), .ZN(n4614) );
  OAI21_X1 U6017 ( .B1(n8956), .B2(n8882), .A(n4616), .ZN(n4615) );
  AOI21_X1 U6018 ( .B1(n9186), .B2(n6672), .A(n5050), .ZN(n6674) );
  NOR2_X1 U6019 ( .A1(n5052), .A2(n5051), .ZN(n5050) );
  AND2_X1 U6020 ( .A1(n5054), .A2(n5053), .ZN(n6680) );
  OAI21_X1 U6021 ( .B1(n9484), .B2(n6752), .A(n5049), .ZN(P1_U3555) );
  NAND2_X1 U6022 ( .A1(n9484), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U6023 ( .A1(n4844), .A2(n4843), .ZN(P1_U3519) );
  NAND2_X1 U6024 ( .A1(n10117), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4843) );
  NAND2_X1 U6025 ( .A1(n9903), .A2(n10119), .ZN(n4844) );
  XNOR2_X1 U6026 ( .A(n5879), .B(P1_IR_REG_20__SCAN_IN), .ZN(n5890) );
  INV_X1 U6027 ( .A(n5890), .ZN(n6437) );
  INV_X1 U6028 ( .A(n7527), .ZN(n4653) );
  AND2_X1 U6029 ( .A1(n5055), .A2(n5056), .ZN(n4518) );
  INV_X1 U6030 ( .A(n6984), .ZN(n4807) );
  AND2_X1 U6031 ( .A1(n4572), .A2(n4709), .ZN(n4519) );
  INV_X1 U6032 ( .A(n7259), .ZN(n4802) );
  AND2_X1 U6033 ( .A1(n8121), .A2(n4587), .ZN(n4520) );
  AND2_X1 U6034 ( .A1(n7732), .A2(n8534), .ZN(n4521) );
  NOR2_X1 U6035 ( .A1(n8838), .A2(n8189), .ZN(n4522) );
  INV_X1 U6036 ( .A(n7020), .ZN(n5026) );
  INV_X1 U6037 ( .A(n7529), .ZN(n4654) );
  NAND2_X1 U6038 ( .A1(n5852), .A2(n5116), .ZN(n5873) );
  AND2_X1 U6039 ( .A1(n8244), .A2(n8240), .ZN(n4523) );
  INV_X1 U6040 ( .A(n5064), .ZN(n5059) );
  NAND2_X1 U6041 ( .A1(n4565), .A2(n7761), .ZN(n5064) );
  INV_X1 U6042 ( .A(n5081), .ZN(n5080) );
  NAND2_X1 U6043 ( .A1(n9582), .A2(n4546), .ZN(n5081) );
  NOR2_X1 U6044 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n4524) );
  NAND2_X1 U6045 ( .A1(n4562), .A2(n5323), .ZN(n5002) );
  NOR2_X1 U6046 ( .A1(n8440), .A2(n5495), .ZN(n4525) );
  INV_X1 U6047 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4746) );
  NOR2_X1 U6048 ( .A1(n8329), .A2(n8368), .ZN(n4526) );
  AND2_X1 U6049 ( .A1(n5288), .A2(n5481), .ZN(n7184) );
  INV_X1 U6050 ( .A(n7184), .ZN(n4904) );
  AND3_X1 U6051 ( .A1(n9416), .A2(n4699), .A3(n4582), .ZN(n4527) );
  AND2_X1 U6052 ( .A1(n5094), .A2(n8407), .ZN(n4528) );
  NOR2_X1 U6053 ( .A1(n7497), .A2(n4889), .ZN(n4529) );
  NAND2_X1 U6054 ( .A1(n4807), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4530) );
  OR2_X1 U6055 ( .A1(n5016), .A2(n5015), .ZN(n7802) );
  INV_X1 U6056 ( .A(n8464), .ZN(n5098) );
  OR2_X1 U6057 ( .A1(n7290), .A2(n4889), .ZN(n4531) );
  NAND2_X1 U6058 ( .A1(n5013), .A2(n6062), .ZN(n7510) );
  OR2_X1 U6059 ( .A1(n10129), .A2(n4608), .ZN(n4532) );
  AND2_X1 U6060 ( .A1(n8689), .A2(n8697), .ZN(n4533) );
  NAND2_X1 U6061 ( .A1(n8910), .A2(n4880), .ZN(n4879) );
  NAND2_X1 U6062 ( .A1(n8199), .A2(n8198), .ZN(n7095) );
  INV_X1 U6063 ( .A(n8828), .ZN(n4995) );
  AND2_X1 U6064 ( .A1(n4722), .A2(n8123), .ZN(n4535) );
  INV_X1 U6065 ( .A(n7134), .ZN(n5042) );
  INV_X1 U6066 ( .A(n5009), .ZN(n5286) );
  AND2_X1 U6067 ( .A1(n8473), .A2(n8121), .ZN(n4536) );
  AND2_X1 U6068 ( .A1(n5095), .A2(n8465), .ZN(n4537) );
  INV_X1 U6069 ( .A(n8539), .ZN(n5200) );
  NAND2_X1 U6070 ( .A1(n9922), .A2(n9821), .ZN(n4538) );
  NAND2_X1 U6071 ( .A1(n4791), .A2(n6807), .ZN(n6793) );
  OR2_X1 U6072 ( .A1(n8738), .A2(n8188), .ZN(n4539) );
  INV_X1 U6073 ( .A(n9224), .ZN(n5923) );
  XOR2_X1 U6074 ( .A(n8329), .B(n8368), .Z(n4540) );
  OR2_X1 U6075 ( .A1(n8625), .A2(n8624), .ZN(n4541) );
  AND2_X1 U6076 ( .A1(n5486), .A2(n5485), .ZN(n8440) );
  NAND2_X1 U6077 ( .A1(n7979), .A2(n8530), .ZN(n4542) );
  INV_X1 U6078 ( .A(n4712), .ZN(n4711) );
  NAND2_X1 U6079 ( .A1(n7983), .A2(n4542), .ZN(n4712) );
  INV_X1 U6080 ( .A(n8237), .ZN(n4757) );
  NOR2_X1 U6081 ( .A1(n5342), .A2(SI_9_), .ZN(n4543) );
  OR2_X1 U6082 ( .A1(n7865), .A2(n7868), .ZN(n4544) );
  AND2_X1 U6083 ( .A1(n5089), .A2(n4538), .ZN(n4545) );
  NAND2_X1 U6084 ( .A1(n9233), .A2(n9806), .ZN(n4546) );
  AND2_X1 U6085 ( .A1(n8302), .A2(n8764), .ZN(n4547) );
  AND2_X1 U6086 ( .A1(n5547), .A2(n7184), .ZN(n4548) );
  NOR2_X1 U6087 ( .A1(n5791), .A2(n5790), .ZN(n4549) );
  NAND2_X1 U6088 ( .A1(n5188), .A2(n4716), .ZN(n5242) );
  AND4_X1 U6089 ( .A1(n5142), .A2(n5141), .A3(n5797), .A4(n5830), .ZN(n4550)
         );
  OR2_X1 U6090 ( .A1(n9622), .A2(n9798), .ZN(n4551) );
  INV_X1 U6091 ( .A(n5324), .ZN(n5004) );
  NAND2_X1 U6092 ( .A1(n5007), .A2(n5009), .ZN(n5803) );
  NAND2_X1 U6093 ( .A1(n5188), .A2(n5189), .ZN(n5207) );
  AND2_X1 U6094 ( .A1(n8819), .A2(n4987), .ZN(n4552) );
  NOR2_X1 U6095 ( .A1(n5159), .A2(n5158), .ZN(n4553) );
  OR2_X1 U6096 ( .A1(n9317), .A2(n4697), .ZN(n4554) );
  INV_X1 U6097 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5886) );
  NOR2_X1 U6098 ( .A1(n9092), .A2(n9125), .ZN(n4555) );
  AND2_X1 U6099 ( .A1(n9390), .A2(n9392), .ZN(n9762) );
  AND2_X1 U6100 ( .A1(n5294), .A2(n5332), .ZN(n7197) );
  OR2_X1 U6101 ( .A1(n7148), .A2(n7244), .ZN(n4556) );
  OR2_X1 U6102 ( .A1(n5949), .A2(n6544), .ZN(n4557) );
  NAND2_X1 U6103 ( .A1(n9935), .A2(n9537), .ZN(n4558) );
  AND2_X1 U6104 ( .A1(n9415), .A2(n9414), .ZN(n4559) );
  AND2_X1 U6105 ( .A1(n5130), .A2(n8181), .ZN(n4560) );
  INV_X1 U6106 ( .A(n5535), .ZN(n4994) );
  INV_X1 U6107 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5189) );
  AND2_X1 U6108 ( .A1(n9370), .A2(n9368), .ZN(n9300) );
  OR2_X1 U6109 ( .A1(n7616), .A2(n9176), .ZN(n9374) );
  NOR2_X1 U6110 ( .A1(n9527), .A2(n9754), .ZN(n4561) );
  INV_X1 U6111 ( .A(n5031), .ZN(n5030) );
  OAI21_X1 U6112 ( .B1(n5033), .B2(n5032), .A(n6246), .ZN(n5031) );
  OR2_X1 U6113 ( .A1(n7732), .A2(n8534), .ZN(n4562) );
  OAI21_X1 U6114 ( .B1(n7497), .B2(n9475), .A(n7490), .ZN(n5070) );
  INV_X1 U6115 ( .A(n5706), .ZN(n4971) );
  OAI21_X1 U6116 ( .B1(n7260), .B2(n4796), .A(n4793), .ZN(n7527) );
  AND2_X1 U6117 ( .A1(n9762), .A2(n4832), .ZN(n4563) );
  AND2_X1 U6118 ( .A1(n9462), .A2(n9225), .ZN(n4564) );
  OR2_X1 U6119 ( .A1(n9892), .A2(n10106), .ZN(n4565) );
  INV_X1 U6120 ( .A(n9514), .ZN(n4839) );
  OR2_X1 U6121 ( .A1(n7259), .A2(n7387), .ZN(n4796) );
  INV_X1 U6122 ( .A(n4893), .ZN(n9603) );
  NOR3_X1 U6123 ( .A1(n9635), .A2(n4895), .A3(n9622), .ZN(n4893) );
  INV_X1 U6124 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5139) );
  INV_X1 U6125 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4883) );
  INV_X1 U6126 ( .A(n4804), .ZN(n4801) );
  NAND2_X1 U6127 ( .A1(n7386), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4804) );
  AND4_X1 U6128 ( .A1(n5747), .A2(n5520), .A3(n5522), .A4(n5143), .ZN(n4566)
         );
  NOR2_X1 U6129 ( .A1(n9907), .A2(n9774), .ZN(n4567) );
  AND2_X1 U6130 ( .A1(n7727), .A2(n7735), .ZN(n4568) );
  OR2_X1 U6131 ( .A1(n5557), .A2(n4992), .ZN(n4569) );
  AND2_X1 U6132 ( .A1(n8293), .A2(n8287), .ZN(n4570) );
  NOR2_X1 U6133 ( .A1(n8260), .A2(n8530), .ZN(n4571) );
  AND2_X1 U6134 ( .A1(n8095), .A2(n8093), .ZN(n4572) );
  INV_X1 U6135 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9007) );
  INV_X1 U6136 ( .A(n7387), .ZN(n7535) );
  INV_X1 U6137 ( .A(n7497), .ZN(n9181) );
  INV_X1 U6138 ( .A(n8193), .ZN(n4847) );
  OR2_X1 U6139 ( .A1(n8947), .A2(n8728), .ZN(n8323) );
  AND2_X1 U6140 ( .A1(n8268), .A2(n8263), .ZN(n4573) );
  AND2_X1 U6141 ( .A1(n6297), .A2(n9134), .ZN(n4574) );
  AND2_X1 U6142 ( .A1(n8209), .A2(n7218), .ZN(n4575) );
  OR2_X1 U6143 ( .A1(n5026), .A2(n6001), .ZN(n4576) );
  NOR2_X1 U6144 ( .A1(n5033), .A2(n6247), .ZN(n4577) );
  NAND2_X1 U6145 ( .A1(n8788), .A2(n8795), .ZN(n4578) );
  NAND2_X1 U6146 ( .A1(n9527), .A2(n9754), .ZN(n4579) );
  AND2_X1 U6147 ( .A1(n8299), .A2(n8298), .ZN(n4580) );
  INV_X1 U6148 ( .A(n8310), .ZN(n4876) );
  OR2_X1 U6149 ( .A1(n8965), .A2(n8425), .ZN(n8310) );
  AND2_X1 U6150 ( .A1(n8132), .A2(n8131), .ZN(n4581) );
  NAND2_X1 U6151 ( .A1(n4839), .A2(n9444), .ZN(n4582) );
  NAND2_X1 U6152 ( .A1(n7821), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4583) );
  NAND2_X1 U6153 ( .A1(n4904), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4584) );
  INV_X1 U6154 ( .A(n5668), .ZN(n4984) );
  INV_X1 U6155 ( .A(n9284), .ZN(n9436) );
  OR2_X1 U6156 ( .A1(n8886), .A2(n8710), .ZN(n4585) );
  NAND2_X1 U6157 ( .A1(n4569), .A2(n5558), .ZN(n4989) );
  INV_X1 U6158 ( .A(n4868), .ZN(n4867) );
  NAND2_X1 U6159 ( .A1(n4869), .A2(n4540), .ZN(n4868) );
  INV_X1 U6160 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5520) );
  NAND2_X2 U6161 ( .A1(n6504), .A2(n5889), .ZN(n6377) );
  INV_X1 U6162 ( .A(n6377), .ZN(n6394) );
  INV_X2 U6163 ( .A(n6377), .ZN(n6360) );
  NAND2_X2 U6164 ( .A1(n5158), .A2(n5145), .ZN(n5736) );
  INV_X1 U6165 ( .A(n8578), .ZN(n4820) );
  NAND2_X1 U6166 ( .A1(n4705), .A2(n4519), .ZN(n8430) );
  NAND2_X1 U6167 ( .A1(n4704), .A2(n8396), .ZN(n8398) );
  NAND2_X1 U6168 ( .A1(n8109), .A2(n8486), .ZN(n8394) );
  INV_X1 U6169 ( .A(n8587), .ZN(n8597) );
  OR2_X1 U6170 ( .A1(n7822), .A2(n7821), .ZN(n4586) );
  INV_X1 U6171 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4966) );
  NAND2_X1 U6172 ( .A1(n5058), .A2(n5062), .ZN(n9528) );
  INV_X1 U6173 ( .A(n8406), .ZN(n5097) );
  OR2_X1 U6174 ( .A1(n8374), .A2(n8795), .ZN(n4587) );
  OR2_X1 U6175 ( .A1(n9911), .A2(n9218), .ZN(n4588) );
  NOR2_X1 U6176 ( .A1(n5498), .A2(SI_16_), .ZN(n4589) );
  NOR2_X1 U6177 ( .A1(n8563), .A2(n8564), .ZN(n4590) );
  NOR2_X1 U6178 ( .A1(n8583), .A2(n8582), .ZN(n4591) );
  INV_X1 U6179 ( .A(n4819), .ZN(n4660) );
  NOR2_X1 U6180 ( .A1(n8587), .A2(n8581), .ZN(n4819) );
  OR2_X1 U6181 ( .A1(n9907), .A2(n9889), .ZN(n4592) );
  AND2_X1 U6182 ( .A1(n5538), .A2(SI_18_), .ZN(n4593) );
  INV_X1 U6183 ( .A(n4959), .ZN(n4958) );
  NAND2_X1 U6184 ( .A1(n4962), .A2(n4960), .ZN(n4959) );
  OR2_X1 U6185 ( .A1(n9907), .A2(n9948), .ZN(n4594) );
  AND2_X1 U6186 ( .A1(n7797), .A2(n9380), .ZN(n4595) );
  XNOR2_X1 U6187 ( .A(n5802), .B(P2_IR_REG_25__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U6188 ( .A1(n6267), .A2(n6266), .ZN(n9935) );
  INV_X1 U6189 ( .A(n9935), .ZN(n4896) );
  OAI21_X1 U6190 ( .B1(n5807), .B2(n5808), .A(n6725), .ZN(n5811) );
  OAI21_X1 U6191 ( .B1(n5796), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5829) );
  INV_X1 U6192 ( .A(n7218), .ZN(n5769) );
  INV_X1 U6193 ( .A(n8857), .ZN(n4977) );
  NAND2_X1 U6194 ( .A1(n5781), .A2(n8239), .ZN(n7843) );
  NAND2_X1 U6195 ( .A1(n6023), .A2(n6022), .ZN(n7132) );
  OR2_X1 U6196 ( .A1(n8185), .A2(n8191), .ZN(n4596) );
  NAND2_X1 U6197 ( .A1(n5025), .A2(n6001), .ZN(n7018) );
  NAND2_X1 U6198 ( .A1(n6098), .A2(n6097), .ZN(n9169) );
  INV_X1 U6199 ( .A(n9169), .ZN(n5015) );
  NAND2_X1 U6200 ( .A1(n7192), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7260) );
  NOR2_X1 U6201 ( .A1(n4803), .A2(n7527), .ZN(n4597) );
  AND2_X1 U6202 ( .A1(n6060), .A2(n6062), .ZN(n4598) );
  AND2_X1 U6203 ( .A1(n4650), .A2(n4651), .ZN(n4599) );
  AND2_X1 U6204 ( .A1(n5726), .A2(n4949), .ZN(n4600) );
  INV_X1 U6205 ( .A(n5002), .ZN(n5001) );
  NOR2_X1 U6206 ( .A1(n7290), .A2(n7347), .ZN(n4601) );
  AND2_X1 U6207 ( .A1(n7218), .A2(n7221), .ZN(n4602) );
  INV_X1 U6208 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n4655) );
  AND2_X1 U6209 ( .A1(n4799), .A2(n4802), .ZN(n4603) );
  AND2_X1 U6210 ( .A1(n10134), .A2(n4634), .ZN(n4604) );
  AND2_X1 U6211 ( .A1(n5110), .A2(n5109), .ZN(n4605) );
  XNOR2_X1 U6212 ( .A(n5752), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8191) );
  AND2_X2 U6213 ( .A1(n6764), .A2(n6763), .ZN(n10119) );
  NAND2_X1 U6214 ( .A1(n6434), .A2(n5890), .ZN(n4606) );
  OR2_X1 U6215 ( .A1(n8699), .A2(n8688), .ZN(n4607) );
  INV_X1 U6216 ( .A(n4810), .ZN(n6985) );
  NOR2_X1 U6217 ( .A1(n6835), .A2(n5248), .ZN(n4810) );
  AND2_X1 U6218 ( .A1(n4640), .A2(n4607), .ZN(n4608) );
  INV_X1 U6219 ( .A(n8658), .ZN(n4646) );
  OR2_X1 U6220 ( .A1(n8030), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4609) );
  INV_X1 U6221 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U6222 ( .A1(n4610), .A2(n4691), .ZN(n9471) );
  NAND2_X1 U6223 ( .A1(n4694), .A2(n4696), .ZN(n4610) );
  OR3_X2 U6224 ( .A1(n7360), .A2(n7359), .A3(n7358), .ZN(n9252) );
  NAND2_X1 U6225 ( .A1(n9788), .A2(n4592), .ZN(P1_U3550) );
  NAND2_X1 U6226 ( .A1(n9906), .A2(n4594), .ZN(P1_U3518) );
  OAI211_X2 U6227 ( .C1(n9268), .C2(n9240), .A(n9239), .B(n9441), .ZN(n9275)
         );
  AOI211_X1 U6228 ( .C1(n9898), .C2(n9507), .A(n9278), .B(n9277), .ZN(n9279)
         );
  NAND2_X2 U6229 ( .A1(n9610), .A2(n9609), .ZN(n9608) );
  NAND2_X1 U6230 ( .A1(n9594), .A2(n9520), .ZN(n9581) );
  OAI21_X1 U6231 ( .B1(n9512), .B2(n4837), .A(n4835), .ZN(n9643) );
  NOR2_X2 U6232 ( .A1(n6333), .A2(n6332), .ZN(n9158) );
  NAND2_X1 U6233 ( .A1(n7603), .A2(n6080), .ZN(n6098) );
  NAND2_X1 U6234 ( .A1(n4622), .A2(n4577), .ZN(n5028) );
  NOR2_X1 U6235 ( .A1(n9193), .A2(n4625), .ZN(n6487) );
  NAND2_X1 U6236 ( .A1(n9149), .A2(n6165), .ZN(n6183) );
  NAND2_X1 U6237 ( .A1(n9081), .A2(n6146), .ZN(n9147) );
  INV_X1 U6238 ( .A(n9126), .ZN(n4611) );
  NAND2_X1 U6239 ( .A1(n6145), .A2(n9079), .ZN(n9081) );
  XNOR2_X1 U6240 ( .A(n5967), .B(n5965), .ZN(n6718) );
  NAND2_X1 U6241 ( .A1(n5023), .A2(n4576), .ZN(n7069) );
  NAND2_X1 U6242 ( .A1(n5191), .A2(n5190), .ZN(n5197) );
  NAND2_X1 U6243 ( .A1(n5258), .A2(n5257), .ZN(n5276) );
  AOI21_X1 U6244 ( .B1(n8184), .B2(n7636), .A(n8185), .ZN(n4884) );
  NAND2_X1 U6245 ( .A1(n4621), .A2(n4620), .ZN(n6184) );
  INV_X1 U6246 ( .A(n6183), .ZN(n4621) );
  NAND3_X1 U6247 ( .A1(n4550), .A2(n4740), .A3(n5137), .ZN(n4739) );
  NAND2_X1 U6248 ( .A1(n4618), .A2(n4614), .ZN(P2_U3207) );
  OR2_X1 U6249 ( .A1(n8951), .A2(n10163), .ZN(n4618) );
  NAND2_X1 U6250 ( .A1(n8755), .A2(n5668), .ZN(n8747) );
  NAND2_X1 U6251 ( .A1(n5155), .A2(n5012), .ZN(n4775) );
  OAI21_X1 U6252 ( .B1(n7844), .B2(n5408), .A(n5407), .ZN(n7955) );
  NAND2_X1 U6253 ( .A1(n5916), .A2(n5917), .ZN(n4619) );
  AND2_X1 U6254 ( .A1(n6645), .A2(n5907), .ZN(n9061) );
  NAND2_X1 U6255 ( .A1(n6646), .A2(n6647), .ZN(n6645) );
  NAND2_X1 U6256 ( .A1(n5028), .A2(n5027), .ZN(n5035) );
  INV_X1 U6257 ( .A(n9099), .ZN(n4622) );
  NAND2_X1 U6258 ( .A1(n5984), .A2(n5983), .ZN(n6906) );
  NAND2_X1 U6259 ( .A1(n9068), .A2(n6321), .ZN(n6333) );
  INV_X1 U6260 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U6261 ( .A1(n6250), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U6262 ( .A1(n5017), .A2(n7803), .ZN(n5016) );
  OAI21_X2 U6263 ( .B1(n5517), .B2(n4959), .A(n4955), .ZN(n5578) );
  OAI21_X1 U6264 ( .B1(n5595), .B2(n5594), .A(n5593), .ZN(n5608) );
  OAI21_X1 U6265 ( .B1(n6436), .B2(n6487), .A(n9206), .ZN(n6461) );
  NAND2_X1 U6266 ( .A1(n4750), .A2(n8338), .ZN(n4749) );
  NAND3_X1 U6267 ( .A1(n4623), .A2(n8351), .A3(n4585), .ZN(n8353) );
  NAND2_X1 U6268 ( .A1(n4748), .A2(n8307), .ZN(n8316) );
  NAND2_X1 U6269 ( .A1(n8300), .A2(n4580), .ZN(n4751) );
  NAND2_X1 U6270 ( .A1(n8281), .A2(n8280), .ZN(n4773) );
  NAND2_X1 U6271 ( .A1(n4737), .A2(n8259), .ZN(n8264) );
  AOI21_X1 U6272 ( .B1(n8317), .B2(n8764), .A(n4780), .ZN(n4779) );
  NAND2_X1 U6273 ( .A1(n4624), .A2(n5190), .ZN(n5177) );
  NAND2_X1 U6274 ( .A1(n5170), .A2(n5169), .ZN(n4624) );
  OR2_X2 U6275 ( .A1(n9645), .A2(n9546), .ZN(n9548) );
  NAND2_X1 U6276 ( .A1(n9598), .A2(n5077), .ZN(n5076) );
  NAND2_X1 U6277 ( .A1(n9536), .A2(n4558), .ZN(n5092) );
  OAI21_X2 U6278 ( .B1(n9734), .B2(n9530), .A(n9532), .ZN(n9714) );
  NAND2_X1 U6279 ( .A1(n5285), .A2(n5291), .ZN(n6519) );
  INV_X1 U6280 ( .A(n5168), .ZN(n5170) );
  AND2_X2 U6281 ( .A1(n5045), .A2(n5043), .ZN(n9193) );
  NAND2_X1 U6282 ( .A1(n5014), .A2(n6062), .ZN(n7601) );
  NOR2_X1 U6283 ( .A1(n7819), .A2(n7777), .ZN(n7894) );
  NAND2_X1 U6284 ( .A1(n7818), .A2(n7823), .ZN(n4628) );
  INV_X1 U6285 ( .A(n7895), .ZN(n4629) );
  INV_X1 U6286 ( .A(n8562), .ZN(n4929) );
  NOR2_X1 U6287 ( .A1(n8636), .A2(n8639), .ZN(n8656) );
  NOR2_X1 U6288 ( .A1(n8613), .A2(n8612), .ZN(n8635) );
  OAI21_X2 U6289 ( .B1(P1_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n5151), .ZN(n4824) );
  OR2_X2 U6290 ( .A1(n9236), .A2(n9285), .ZN(n9268) );
  NAND2_X1 U6291 ( .A1(n5372), .A2(n5371), .ZN(n5394) );
  INV_X1 U6292 ( .A(n8333), .ZN(n8330) );
  XNOR2_X1 U6293 ( .A(n5727), .B(n5725), .ZN(n9019) );
  NAND2_X1 U6294 ( .A1(n9319), .A2(n4554), .ZN(n4695) );
  INV_X1 U6295 ( .A(n8349), .ZN(n4932) );
  NAND2_X1 U6296 ( .A1(n4767), .A2(n4932), .ZN(n4766) );
  MUX2_X1 U6297 ( .A(n5171), .B(n5172), .S(n5910), .Z(n5173) );
  AOI21_X2 U6298 ( .B1(n9581), .B2(n9523), .A(n9522), .ZN(n9567) );
  NAND2_X2 U6299 ( .A1(n5500), .A2(n5499), .ZN(n5517) );
  NAND2_X1 U6300 ( .A1(n8659), .A2(n4532), .ZN(n4631) );
  INV_X1 U6301 ( .A(n4630), .ZN(n4633) );
  OAI21_X1 U6302 ( .B1(n8691), .B2(n4638), .A(n4636), .ZN(n4630) );
  OAI21_X1 U6303 ( .B1(n8659), .B2(n4604), .A(n4631), .ZN(n4632) );
  NAND3_X1 U6304 ( .A1(n4635), .A2(n4633), .A3(n4632), .ZN(P2_U3201) );
  NAND3_X1 U6305 ( .A1(n8691), .A2(n10149), .A3(n8700), .ZN(n4635) );
  INV_X1 U6306 ( .A(n8579), .ZN(n4658) );
  NAND2_X1 U6307 ( .A1(n4792), .A2(n10145), .ZN(n4791) );
  NAND2_X1 U6308 ( .A1(n6793), .A2(n4670), .ZN(n6821) );
  NAND3_X1 U6309 ( .A1(n4792), .A2(n10145), .A3(n4671), .ZN(n4670) );
  INV_X1 U6310 ( .A(n6807), .ZN(n4671) );
  OR2_X1 U6311 ( .A1(n9331), .A2(n7000), .ZN(n9330) );
  INV_X2 U6312 ( .A(n6206), .ZN(n5852) );
  AND2_X2 U6313 ( .A1(n5116), .A2(n5019), .ZN(n5018) );
  NAND2_X1 U6314 ( .A1(n9371), .A2(n9370), .ZN(n4680) );
  NAND2_X1 U6315 ( .A1(n9413), .A2(n9399), .ZN(n9401) );
  NAND2_X1 U6316 ( .A1(n4681), .A2(n9733), .ZN(n9413) );
  NAND2_X1 U6317 ( .A1(n4683), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U6318 ( .A1(n9388), .A2(n9463), .ZN(n4682) );
  NOR2_X1 U6319 ( .A1(n4684), .A2(n9398), .ZN(n4683) );
  AND2_X1 U6320 ( .A1(n9387), .A2(n9444), .ZN(n4684) );
  NAND2_X1 U6321 ( .A1(n4685), .A2(n4689), .ZN(n9446) );
  NAND3_X1 U6322 ( .A1(n9435), .A2(n4686), .A3(n9552), .ZN(n4685) );
  NAND3_X1 U6323 ( .A1(n4688), .A2(n9284), .A3(n9440), .ZN(n4686) );
  NAND2_X1 U6324 ( .A1(n9434), .A2(n9436), .ZN(n4688) );
  NAND3_X1 U6325 ( .A1(n9455), .A2(n6264), .A3(n4554), .ZN(n4696) );
  NAND4_X1 U6326 ( .A1(n9402), .A2(n9404), .A3(n9674), .A4(n9403), .ZN(n4700)
         );
  NAND2_X2 U6327 ( .A1(n6443), .A2(n6540), .ZN(n5949) );
  NAND2_X1 U6328 ( .A1(n5949), .A2(n7998), .ZN(n5948) );
  NAND2_X1 U6329 ( .A1(n5949), .A2(n5910), .ZN(n6284) );
  NAND2_X1 U6330 ( .A1(n8398), .A2(n5096), .ZN(n5093) );
  NAND2_X1 U6331 ( .A1(n8394), .A2(n8395), .ZN(n4704) );
  NAND2_X1 U6332 ( .A1(n7981), .A2(n4519), .ZN(n4708) );
  NAND3_X1 U6333 ( .A1(n8473), .A2(n4520), .A3(n8419), .ZN(n4719) );
  NAND2_X1 U6334 ( .A1(n4719), .A2(n4720), .ZN(n8422) );
  OAI21_X1 U6335 ( .B1(n7556), .B2(n4727), .A(n4725), .ZN(n4724) );
  NAND2_X1 U6336 ( .A1(n8408), .A2(n4734), .ZN(n8119) );
  NAND2_X1 U6337 ( .A1(n8408), .A2(n4732), .ZN(n4731) );
  NAND2_X1 U6338 ( .A1(n8121), .A2(n4731), .ZN(n8475) );
  OR2_X1 U6339 ( .A1(n8117), .A2(n8821), .ZN(n4734) );
  INV_X1 U6340 ( .A(n8264), .ZN(n8267) );
  NAND2_X1 U6341 ( .A1(n4738), .A2(n8256), .ZN(n4737) );
  NAND3_X1 U6342 ( .A1(n8254), .A2(n8255), .A3(n8253), .ZN(n4738) );
  NAND3_X1 U6343 ( .A1(n8201), .A2(n7218), .A3(n8200), .ZN(n8208) );
  NAND3_X1 U6344 ( .A1(n4566), .A2(n5136), .A3(n5138), .ZN(n4741) );
  AND4_X1 U6345 ( .A1(n5136), .A2(n5138), .A3(n5137), .A4(n4746), .ZN(n5140)
         );
  NAND3_X1 U6346 ( .A1(n5136), .A2(n5138), .A3(n5137), .ZN(n5480) );
  NAND3_X1 U6347 ( .A1(n4761), .A2(n8237), .A3(n8232), .ZN(n4760) );
  NAND3_X1 U6348 ( .A1(n8229), .A2(n8228), .A3(n8227), .ZN(n4761) );
  NAND3_X1 U6349 ( .A1(n4764), .A2(n8218), .A3(n8233), .ZN(n4763) );
  NAND3_X1 U6350 ( .A1(n8217), .A2(n8216), .A3(n8228), .ZN(n4764) );
  NAND2_X2 U6351 ( .A1(n4777), .A2(n4776), .ZN(n8539) );
  MUX2_X1 U6352 ( .A(n6802), .B(n7110), .S(n8698), .Z(n6803) );
  OAI21_X1 U6353 ( .B1(n7258), .B2(n4796), .A(n4795), .ZN(n4794) );
  INV_X1 U6354 ( .A(n7260), .ZN(n4798) );
  INV_X1 U6355 ( .A(n4811), .ZN(n7190) );
  NAND2_X1 U6356 ( .A1(n6820), .A2(n6795), .ZN(n4815) );
  INV_X1 U6357 ( .A(n6795), .ZN(n4817) );
  MUX2_X1 U6358 ( .A(n9024), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6359 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9024), .S(n6507), .Z(n8035) );
  NAND2_X1 U6360 ( .A1(n4827), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4826) );
  NAND2_X1 U6361 ( .A1(n9732), .A2(n9399), .ZN(n4828) );
  NAND2_X1 U6362 ( .A1(n4828), .A2(n4829), .ZN(n9711) );
  AND2_X2 U6363 ( .A1(n7762), .A2(n9384), .ZN(n5129) );
  NAND2_X2 U6364 ( .A1(n7589), .A2(n7590), .ZN(n7623) );
  INV_X1 U6365 ( .A(n9512), .ZN(n4842) );
  NAND3_X1 U6366 ( .A1(n5199), .A2(n4846), .A3(n4845), .ZN(n7013) );
  OR2_X1 U6367 ( .A1(n6507), .A2(n6789), .ZN(n4846) );
  NAND2_X1 U6368 ( .A1(n8199), .A2(n4847), .ZN(n4848) );
  AND2_X2 U6369 ( .A1(n8202), .A2(n8203), .ZN(n7218) );
  NAND2_X1 U6370 ( .A1(n4848), .A2(n8198), .ZN(n7220) );
  NAND2_X1 U6371 ( .A1(n5781), .A2(n4852), .ZN(n4851) );
  NAND2_X1 U6372 ( .A1(n4851), .A2(n4854), .ZN(n7970) );
  NAND2_X1 U6373 ( .A1(n5776), .A2(n8218), .ZN(n7470) );
  INV_X1 U6374 ( .A(n8218), .ZN(n4864) );
  NAND2_X2 U6375 ( .A1(n4866), .A2(n4865), .ZN(n8178) );
  NAND2_X1 U6376 ( .A1(n8910), .A2(n4872), .ZN(n4871) );
  NAND2_X1 U6377 ( .A1(n4871), .A2(n4874), .ZN(n8763) );
  NAND3_X1 U6378 ( .A1(n5007), .A2(n5009), .A3(n4882), .ZN(n4881) );
  OR2_X1 U6379 ( .A1(n8806), .A2(n5788), .ZN(n5789) );
  OAI21_X1 U6380 ( .B1(n8079), .B2(n8078), .A(n8293), .ZN(n8817) );
  NAND2_X1 U6381 ( .A1(n8803), .A2(n8802), .ZN(n8910) );
  NAND2_X1 U6382 ( .A1(n7239), .A2(n8212), .ZN(n7320) );
  OAI21_X1 U6383 ( .B1(n8817), .B2(n5787), .A(n8295), .ZN(n8806) );
  AND2_X2 U6384 ( .A1(n9628), .A2(n9518), .ZN(n9610) );
  NAND2_X2 U6385 ( .A1(n6045), .A2(n6044), .ZN(n7285) );
  NAND2_X1 U6386 ( .A1(n5771), .A2(n8219), .ZN(n7240) );
  NAND2_X1 U6387 ( .A1(n7240), .A2(n8209), .ZN(n7239) );
  AND2_X1 U6388 ( .A1(n5135), .A2(n5134), .ZN(n5136) );
  INV_X1 U6389 ( .A(n8837), .ZN(n5785) );
  NOR3_X2 U6390 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .A3(
        P2_IR_REG_14__SCAN_IN), .ZN(n5138) );
  NAND2_X2 U6391 ( .A1(n9957), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5896) );
  NAND3_X2 U6392 ( .A1(n5018), .A2(n5852), .A3(n4524), .ZN(n9957) );
  INV_X1 U6393 ( .A(n7290), .ZN(n4888) );
  NAND2_X1 U6394 ( .A1(n4888), .A2(n4529), .ZN(n7593) );
  INV_X1 U6395 ( .A(n9242), .ZN(n10074) );
  NOR2_X1 U6396 ( .A1(n9635), .A2(n9622), .ZN(n9617) );
  INV_X1 U6397 ( .A(n9915), .ZN(n4895) );
  NOR2_X2 U6398 ( .A1(n9751), .A2(n9872), .ZN(n9749) );
  NAND2_X1 U6399 ( .A1(n6976), .A2(n6831), .ZN(n4900) );
  NAND2_X1 U6400 ( .A1(n7182), .A2(n4903), .ZN(n7185) );
  NAND2_X1 U6401 ( .A1(n4900), .A2(n4901), .ZN(n7182) );
  NAND2_X1 U6402 ( .A1(n10131), .A2(n10132), .ZN(n10130) );
  NAND2_X1 U6403 ( .A1(n6828), .A2(n4918), .ZN(n6830) );
  NAND2_X1 U6404 ( .A1(n6782), .A2(n6818), .ZN(n4916) );
  INV_X1 U6405 ( .A(n6842), .ZN(n4919) );
  INV_X1 U6406 ( .A(n8566), .ZN(n4928) );
  NAND2_X1 U6407 ( .A1(n5595), .A2(n4937), .ZN(n4936) );
  INV_X1 U6408 ( .A(n5618), .ZN(n5615) );
  NAND2_X1 U6409 ( .A1(n5310), .A2(n4944), .ZN(n4940) );
  NAND2_X1 U6410 ( .A1(n5310), .A2(n5309), .ZN(n5330) );
  OAI21_X1 U6411 ( .B1(n5674), .B2(n4954), .A(n4951), .ZN(n5727) );
  NAND2_X1 U6412 ( .A1(n5674), .A2(n4951), .ZN(n4950) );
  NAND2_X1 U6413 ( .A1(n5674), .A2(n5673), .ZN(n5692) );
  OAI21_X1 U6414 ( .B1(n5910), .B2(n4966), .A(n4965), .ZN(n5193) );
  AOI21_X1 U6415 ( .B1(n8739), .B2(n8738), .A(n5706), .ZN(n8724) );
  NAND2_X1 U6416 ( .A1(n8858), .A2(n4974), .ZN(n4973) );
  OAI211_X1 U6417 ( .C1(n4980), .C2(n4979), .A(n5221), .B(n4978), .ZN(n5223)
         );
  NAND2_X1 U6418 ( .A1(n7104), .A2(n7221), .ZN(n4980) );
  NAND2_X1 U6419 ( .A1(n7223), .A2(n5201), .ZN(n7232) );
  NAND2_X1 U6420 ( .A1(n4980), .A2(n5769), .ZN(n7223) );
  INV_X1 U6421 ( .A(n5648), .ZN(n8756) );
  NAND2_X1 U6422 ( .A1(n4981), .A2(n4982), .ZN(n5690) );
  NAND2_X1 U6423 ( .A1(n5648), .A2(n5668), .ZN(n4981) );
  NAND2_X1 U6424 ( .A1(n8828), .A2(n4989), .ZN(n4985) );
  OAI21_X1 U6425 ( .B1(n7466), .B2(n4999), .A(n4997), .ZN(n7772) );
  NAND3_X1 U6426 ( .A1(n5000), .A2(n4544), .A3(n5002), .ZN(n4998) );
  NAND2_X1 U6427 ( .A1(n5006), .A2(n4573), .ZN(n5452) );
  NAND2_X1 U6428 ( .A1(n5155), .A2(n5010), .ZN(n9008) );
  NAND2_X1 U6429 ( .A1(n6060), .A2(n7511), .ZN(n5014) );
  NAND2_X1 U6430 ( .A1(n7601), .A2(n7605), .ZN(n7603) );
  NAND2_X1 U6431 ( .A1(n5016), .A2(n9169), .ZN(n6122) );
  NAND2_X1 U6432 ( .A1(n6096), .A2(n6095), .ZN(n5017) );
  AND2_X1 U6433 ( .A1(n5017), .A2(n9169), .ZN(n7801) );
  NAND2_X1 U6434 ( .A1(n5020), .A2(n5024), .ZN(n5021) );
  NAND2_X1 U6435 ( .A1(n6906), .A2(n5021), .ZN(n5023) );
  NAND2_X1 U6436 ( .A1(n5035), .A2(n4574), .ZN(n6303) );
  NAND2_X1 U6437 ( .A1(n6023), .A2(n5038), .ZN(n5036) );
  NAND2_X1 U6438 ( .A1(n5036), .A2(n5037), .ZN(n6059) );
  INV_X1 U6439 ( .A(n5048), .ZN(n9124) );
  XNOR2_X1 U6440 ( .A(n6672), .B(n10074), .ZN(n6748) );
  INV_X1 U6441 ( .A(n7759), .ZN(n5060) );
  NAND2_X1 U6442 ( .A1(n7759), .A2(n5057), .ZN(n5055) );
  NAND2_X1 U6443 ( .A1(n7352), .A2(n5068), .ZN(n5067) );
  NAND2_X1 U6444 ( .A1(n6996), .A2(n5072), .ZN(n5071) );
  NAND3_X1 U6445 ( .A1(n5074), .A2(n9294), .A3(n5071), .ZN(n7050) );
  NAND2_X1 U6446 ( .A1(n5076), .A2(n5078), .ZN(n9553) );
  AND2_X1 U6447 ( .A1(n4546), .A2(n5085), .ZN(n9583) );
  OAI21_X1 U6448 ( .B1(n9548), .B2(n5088), .A(n5086), .ZN(n9550) );
  NAND2_X1 U6449 ( .A1(n5093), .A2(n4528), .ZN(n8408) );
  NOR2_X2 U6450 ( .A1(n7411), .A2(n7412), .ZN(n7556) );
  NAND2_X1 U6451 ( .A1(n7731), .A2(n5105), .ZN(n5102) );
  NAND2_X1 U6452 ( .A1(n5102), .A2(n5103), .ZN(n7875) );
  NAND2_X1 U6453 ( .A1(n5521), .A2(n5111), .ZN(n5751) );
  INV_X1 U6454 ( .A(n5751), .ZN(n5749) );
  NAND2_X1 U6455 ( .A1(n8502), .A2(n4581), .ZN(n8365) );
  NOR2_X2 U6456 ( .A1(n7593), .A2(n7616), .ZN(n7625) );
  MUX2_X2 U6457 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8941), .S(n10580), .Z(n8942) );
  MUX2_X2 U6458 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8941), .S(n8928), .Z(n8895)
         );
  AND2_X2 U6459 ( .A1(n8363), .A2(n9015), .ZN(n5224) );
  OR2_X1 U6460 ( .A1(n8711), .A2(n5736), .ZN(n7425) );
  NAND2_X1 U6461 ( .A1(n5798), .A2(n5797), .ZN(n5801) );
  INV_X1 U6462 ( .A(n10149), .ZN(n8666) );
  AND2_X1 U6463 ( .A1(n6796), .A2(n8670), .ZN(n10149) );
  AND2_X1 U6464 ( .A1(n5812), .A2(n7943), .ZN(n5115) );
  AND4_X2 U6465 ( .A1(n5851), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(n5116)
         );
  AND2_X1 U6466 ( .A1(n9101), .A2(n6222), .ZN(n5118) );
  NOR2_X1 U6467 ( .A1(n8189), .A2(n5784), .ZN(n5119) );
  AND2_X1 U6468 ( .A1(n5128), .A2(n5834), .ZN(n5120) );
  NOR2_X1 U6469 ( .A1(n8342), .A2(n8341), .ZN(n5121) );
  NOR2_X1 U6470 ( .A1(n6106), .A2(n6085), .ZN(n5122) );
  NOR2_X1 U6471 ( .A1(n6236), .A2(n6253), .ZN(n5123) );
  AND2_X1 U6472 ( .A1(n5277), .A2(n5262), .ZN(n5124) );
  INV_X1 U6473 ( .A(n8865), .ZN(n7469) );
  INV_X1 U6474 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5813) );
  INV_X1 U6475 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5192) );
  INV_X1 U6476 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5167) );
  AND4_X1 U6477 ( .A1(n5450), .A2(n5449), .A3(n5448), .A4(n5447), .ZN(n8515)
         );
  XNOR2_X1 U6478 ( .A(n5753), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8350) );
  AND2_X1 U6479 ( .A1(n7425), .A2(n5761), .ZN(n8339) );
  NAND2_X1 U6480 ( .A1(n8440), .A2(n8864), .ZN(n5126) );
  INV_X1 U6481 ( .A(n8186), .ZN(n5790) );
  OR2_X1 U6482 ( .A1(n8719), .A2(n9001), .ZN(n5127) );
  OR2_X1 U6483 ( .A1(n8719), .A2(n8929), .ZN(n5128) );
  AND2_X1 U6484 ( .A1(n8180), .A2(n8179), .ZN(n5130) );
  AND2_X1 U6485 ( .A1(n7102), .A2(n5811), .ZN(n6724) );
  NAND2_X2 U6486 ( .A1(n7111), .A2(n8854), .ZN(n10161) );
  INV_X1 U6487 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5864) );
  INV_X1 U6488 ( .A(n5935), .ZN(n6233) );
  INV_X1 U6489 ( .A(n8339), .ZN(n8340) );
  NOR2_X1 U6490 ( .A1(n8338), .A2(n8340), .ZN(n8341) );
  INV_X1 U6491 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5141) );
  INV_X1 U6492 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5748) );
  INV_X1 U6493 ( .A(n6058), .ZN(n6056) );
  OR2_X1 U6494 ( .A1(n5724), .A2(n5723), .ZN(n5728) );
  INV_X1 U6496 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5869) );
  INV_X1 U6497 ( .A(n9272), .ZN(n9273) );
  OR2_X1 U6498 ( .A1(n7927), .A2(n8533), .ZN(n7863) );
  INV_X1 U6499 ( .A(n5603), .ZN(n5602) );
  NAND2_X1 U6500 ( .A1(n8329), .A2(n8740), .ZN(n5720) );
  INV_X1 U6501 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7987) );
  INV_X1 U6502 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10411) );
  OR2_X1 U6503 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  AND2_X1 U6504 ( .A1(n5670), .A2(n5669), .ZN(n5671) );
  INV_X1 U6505 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5866) );
  INV_X1 U6506 ( .A(SI_17_), .ZN(n5501) );
  NAND2_X1 U6507 ( .A1(n7998), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5235) );
  INV_X1 U6508 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5156) );
  INV_X1 U6509 ( .A(n8364), .ZN(n8132) );
  INV_X1 U6510 ( .A(n8350), .ZN(n8185) );
  NAND2_X1 U6511 ( .A1(n5602), .A2(n5601), .ZN(n5622) );
  NOR2_X1 U6512 ( .A1(n5228), .A2(n7110), .ZN(n5160) );
  NOR2_X1 U6513 ( .A1(n6821), .A2(n7235), .ZN(n6820) );
  NOR2_X1 U6514 ( .A1(n8662), .A2(n8661), .ZN(n8664) );
  INV_X1 U6515 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10456) );
  INV_X1 U6516 ( .A(n5569), .ZN(n5568) );
  OAI22_X1 U6517 ( .A1(n7772), .A2(n5390), .B1(n7776), .B2(n7877), .ZN(n7844)
         );
  AND2_X1 U6518 ( .A1(n5763), .A2(n6507), .ZN(n6934) );
  INV_X1 U6519 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6046) );
  INV_X1 U6520 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6128) );
  NOR2_X1 U6521 ( .A1(n6223), .A2(n5118), .ZN(n6224) );
  INV_X1 U6522 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6880) );
  AND2_X1 U6523 ( .A1(n6084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6106) );
  INV_X1 U6524 ( .A(n6490), .ZN(n6086) );
  INV_X1 U6525 ( .A(n9312), .ZN(n9519) );
  INV_X1 U6526 ( .A(n9527), .ZN(n7788) );
  OR2_X1 U6527 ( .A1(n9951), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6419) );
  INV_X1 U6528 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9954) );
  INV_X1 U6529 ( .A(SI_20_), .ZN(n5577) );
  OR2_X1 U6530 ( .A1(n6166), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6167) );
  OR2_X1 U6531 ( .A1(n6469), .A2(n6468), .ZN(n6933) );
  OR2_X1 U6532 ( .A1(n5639), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U6533 ( .A1(n8119), .A2(n8118), .ZN(n8121) );
  NAND2_X1 U6534 ( .A1(n6936), .A2(n6934), .ZN(n8516) );
  AND2_X1 U6535 ( .A1(n7102), .A2(n8038), .ZN(n8355) );
  NAND2_X1 U6536 ( .A1(n8680), .A2(n8696), .ZN(n8681) );
  OR2_X1 U6537 ( .A1(n5584), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U6538 ( .A1(n5568), .A2(n10456), .ZN(n5584) );
  OR2_X1 U6539 ( .A1(n7732), .A2(n7886), .ZN(n8240) );
  AND3_X1 U6540 ( .A1(n6467), .A2(n7102), .A3(n6924), .ZN(n7098) );
  OR2_X1 U6541 ( .A1(n6047), .A2(n6046), .ZN(n6066) );
  NOR2_X1 U6542 ( .A1(n6324), .A2(n9164), .ZN(n6336) );
  AND2_X1 U6543 ( .A1(n6439), .A2(n9950), .ZN(n6442) );
  AND2_X1 U6544 ( .A1(n9558), .A2(n6449), .ZN(n9572) );
  INV_X1 U6545 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7582) );
  INV_X1 U6546 ( .A(n9542), .ZN(n9692) );
  NAND2_X1 U6547 ( .A1(n7789), .A2(n7788), .ZN(n9751) );
  INV_X1 U6548 ( .A(n7789), .ZN(n7791) );
  INV_X1 U6549 ( .A(n9475), .ZN(n9087) );
  NAND4_X1 U6550 ( .A1(n5979), .A2(n5978), .A3(n5977), .A4(n5976), .ZN(n6529)
         );
  NAND2_X1 U6551 ( .A1(n6381), .A2(n6380), .ZN(n9233) );
  INV_X1 U6552 ( .A(n9739), .ZN(n9750) );
  INV_X1 U6553 ( .A(n9478), .ZN(n7609) );
  NAND2_X1 U6554 ( .A1(n6419), .A2(n9953), .ZN(n6762) );
  AOI22_X1 U6555 ( .A1(n7146), .A2(n7145), .B1(n5200), .B2(n7144), .ZN(n8384)
         );
  AOI21_X1 U6556 ( .B1(n7142), .B2(n8047), .A(n4847), .ZN(n7009) );
  INV_X1 U6557 ( .A(n8520), .ZN(n8510) );
  AND2_X1 U6558 ( .A1(n8482), .A2(n8037), .ZN(n8527) );
  AND2_X1 U6559 ( .A1(n5687), .A2(n5686), .ZN(n8367) );
  AND4_X1 U6560 ( .A1(n5513), .A2(n5512), .A3(n5511), .A4(n5510), .ZN(n8101)
         );
  INV_X1 U6561 ( .A(n8703), .ZN(n10136) );
  INV_X1 U6562 ( .A(n8706), .ZN(n10143) );
  INV_X1 U6563 ( .A(n8665), .ZN(n8684) );
  AND2_X1 U6564 ( .A1(n10161), .A2(n7452), .ZN(n8872) );
  INV_X1 U6565 ( .A(n8929), .ZN(n8925) );
  OAI21_X1 U6566 ( .B1(n5816), .B2(n6462), .A(n5815), .ZN(n7097) );
  AND2_X1 U6567 ( .A1(n8257), .A2(n8258), .ZN(n8256) );
  OR3_X1 U6568 ( .A1(n7548), .A2(n7449), .A3(n7448), .ZN(n10174) );
  NAND2_X1 U6569 ( .A1(n7753), .A2(n7483), .ZN(n8909) );
  OR2_X1 U6570 ( .A1(n6938), .A2(n6466), .ZN(n6473) );
  AND2_X1 U6571 ( .A1(n6926), .A2(n6733), .ZN(n7102) );
  INV_X1 U6572 ( .A(n9209), .ZN(n9186) );
  INV_X1 U6573 ( .A(n9218), .ZN(n9142) );
  AND2_X1 U6574 ( .A1(n6259), .A2(n6258), .ZN(n9860) );
  AND3_X1 U6575 ( .A1(n6215), .A2(n6214), .A3(n6213), .ZN(n9880) );
  NAND2_X1 U6576 ( .A1(n5955), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5926) );
  INV_X1 U6577 ( .A(n9494), .ZN(n10039) );
  XNOR2_X1 U6578 ( .A(n9553), .B(n9552), .ZN(n9772) );
  AND2_X1 U6579 ( .A1(n9327), .A2(n9406), .ZN(n9710) );
  AND2_X1 U6580 ( .A1(n9288), .A2(n9400), .ZN(n9721) );
  AND2_X1 U6581 ( .A1(n6747), .A2(n6746), .ZN(n10068) );
  INV_X1 U6582 ( .A(n9877), .ZN(n10104) );
  INV_X1 U6583 ( .A(n10068), .ZN(n10116) );
  AND2_X1 U6584 ( .A1(n6762), .A2(n6761), .ZN(n6763) );
  AND2_X1 U6585 ( .A1(n6043), .A2(n6081), .ZN(n6630) );
  INV_X1 U6586 ( .A(n9971), .ZN(n6768) );
  INV_X1 U6587 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10293) );
  INV_X1 U6588 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10305) );
  AND2_X1 U6589 ( .A1(n6931), .A2(n6930), .ZN(n8520) );
  NAND2_X1 U6590 ( .A1(n6921), .A2(n6920), .ZN(n8522) );
  INV_X1 U6591 ( .A(n8367), .ZN(n8758) );
  OAI211_X1 U6592 ( .C1(n5739), .C2(n8799), .A(n5606), .B(n5605), .ZN(n8809)
         );
  INV_X1 U6593 ( .A(n8515), .ZN(n8867) );
  OR2_X1 U6594 ( .A1(P2_U3150), .A2(n6777), .ZN(n10141) );
  OR2_X1 U6595 ( .A1(n8679), .A2(n8354), .ZN(n8703) );
  AOI21_X1 U6596 ( .B1(n8684), .B2(n10149), .A(n8683), .ZN(n8685) );
  OR2_X1 U6597 ( .A1(n8029), .A2(n8670), .ZN(n10129) );
  INV_X1 U6598 ( .A(n8872), .ZN(n8882) );
  INV_X1 U6599 ( .A(n10161), .ZN(n10163) );
  NAND2_X1 U6600 ( .A1(n8928), .A2(n8909), .ZN(n8930) );
  OR2_X1 U6601 ( .A1(n7097), .A2(n5833), .ZN(n8884) );
  NAND2_X1 U6602 ( .A1(n10580), .A2(n8909), .ZN(n9003) );
  AND2_X1 U6603 ( .A1(n6473), .A2(n6472), .ZN(n10578) );
  INV_X1 U6604 ( .A(n6724), .ZN(n6698) );
  AND2_X1 U6605 ( .A1(n6923), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6733) );
  INV_X1 U6606 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7921) );
  INV_X1 U6607 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7237) );
  INV_X1 U6608 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10469) );
  INV_X1 U6609 ( .A(n9831), .ZN(n9663) );
  INV_X1 U6610 ( .A(n9206), .ZN(n9145) );
  INV_X1 U6611 ( .A(n9860), .ZN(n9704) );
  INV_X1 U6612 ( .A(n9880), .ZN(n9735) );
  OR2_X1 U6613 ( .A1(n9996), .A2(n6651), .ZN(n10027) );
  INV_X1 U6614 ( .A(n10030), .ZN(n10048) );
  OR2_X1 U6615 ( .A1(n10063), .A2(n10068), .ZN(n9746) );
  OR2_X1 U6616 ( .A1(n10063), .A2(n7084), .ZN(n9767) );
  NAND2_X1 U6617 ( .A1(n6962), .A2(n9557), .ZN(n10056) );
  NAND2_X1 U6618 ( .A1(n10128), .A2(n10082), .ZN(n9889) );
  INV_X1 U6619 ( .A(n9534), .ZN(n9940) );
  INV_X1 U6620 ( .A(n10119), .ZN(n10117) );
  INV_X1 U6621 ( .A(n10065), .ZN(n10066) );
  AND2_X1 U6622 ( .A1(n9951), .A2(n9950), .ZN(n10065) );
  INV_X1 U6623 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7743) );
  INV_X1 U6624 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10319) );
  INV_X1 U6625 ( .A(n6709), .ZN(n6874) );
  INV_X1 U6626 ( .A(n8679), .ZN(P2_U3893) );
  INV_X1 U6627 ( .A(n9484), .ZN(P1_U3973) );
  NOR2_X1 U6628 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5137) );
  NOR2_X1 U6629 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5142) );
  XNOR2_X2 U6630 ( .A(n5144), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6631 ( .A1(n5224), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5150) );
  NAND2_X4 U6632 ( .A1(n8363), .A2(n5145), .ZN(n5225) );
  INV_X1 U6633 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6790) );
  INV_X1 U6634 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5146) );
  OR2_X1 U6635 ( .A1(n5736), .A2(n5146), .ZN(n5148) );
  NAND2_X1 U6636 ( .A1(n5158), .A2(n9015), .ZN(n5228) );
  INV_X1 U6637 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10439) );
  OR2_X1 U6638 ( .A1(n5228), .A2(n10439), .ZN(n5147) );
  NAND2_X1 U6639 ( .A1(n6511), .A2(SI_0_), .ZN(n5152) );
  XNOR2_X1 U6640 ( .A(n5152), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9024) );
  INV_X1 U6641 ( .A(n8035), .ZN(n8047) );
  OR2_X1 U6642 ( .A1(n7106), .A2(n8047), .ZN(n7105) );
  NAND2_X1 U6643 ( .A1(n5184), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5163) );
  INV_X1 U6644 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7110) );
  INV_X1 U6645 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6802) );
  OR2_X1 U6646 ( .A1(n6802), .A2(n9015), .ZN(n5159) );
  NOR2_X1 U6647 ( .A1(n5160), .A2(n4553), .ZN(n5162) );
  NAND2_X1 U6648 ( .A1(n5224), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5161) );
  NAND3_X1 U6649 ( .A1(n5163), .A2(n5162), .A3(n5161), .ZN(n6916) );
  INV_X1 U6650 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6651 ( .A1(n5168), .A2(SI_1_), .ZN(n5190) );
  INV_X1 U6652 ( .A(SI_1_), .ZN(n5169) );
  INV_X1 U6653 ( .A(n5177), .ZN(n5174) );
  INV_X1 U6654 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5172) );
  INV_X1 U6655 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5171) );
  INV_X1 U6656 ( .A(SI_0_), .ZN(n5893) );
  NAND2_X1 U6657 ( .A1(n5174), .A2(n5175), .ZN(n5191) );
  INV_X1 U6658 ( .A(n5175), .ZN(n5176) );
  NAND2_X1 U6659 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  NAND2_X1 U6660 ( .A1(n5191), .A2(n5178), .ZN(n6514) );
  NAND2_X2 U6661 ( .A1(n6507), .A2(n7998), .ZN(n5218) );
  INV_X1 U6662 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6509) );
  OR2_X1 U6663 ( .A1(n5218), .A2(n6509), .ZN(n5179) );
  INV_X1 U6664 ( .A(n5181), .ZN(n5183) );
  INV_X1 U6665 ( .A(n6916), .ZN(n5182) );
  NAND2_X1 U6666 ( .A1(n7105), .A2(n7095), .ZN(n7104) );
  NAND2_X1 U6667 ( .A1(n5182), .A2(n5183), .ZN(n7221) );
  NAND2_X1 U6668 ( .A1(n5224), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5186) );
  INV_X1 U6669 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6780) );
  OR2_X1 U6670 ( .A1(n5228), .A2(n6780), .ZN(n5185) );
  NAND2_X1 U6671 ( .A1(n5193), .A2(SI_2_), .ZN(n5209) );
  OAI21_X1 U6672 ( .B1(n5193), .B2(SI_2_), .A(n5209), .ZN(n5195) );
  NAND2_X1 U6673 ( .A1(n5194), .A2(n5195), .ZN(n5198) );
  INV_X1 U6674 ( .A(n5195), .ZN(n5196) );
  NAND2_X1 U6675 ( .A1(n5197), .A2(n5196), .ZN(n5210) );
  NAND2_X1 U6676 ( .A1(n5198), .A2(n5210), .ZN(n6513) );
  OR2_X1 U6677 ( .A1(n5218), .A2(n5192), .ZN(n5199) );
  INV_X1 U6678 ( .A(n7013), .ZN(n7011) );
  NAND2_X1 U6679 ( .A1(n5200), .A2(n7013), .ZN(n8203) );
  NAND2_X1 U6680 ( .A1(n5200), .A2(n7011), .ZN(n5201) );
  NAND2_X1 U6681 ( .A1(n5224), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5206) );
  OR2_X1 U6682 ( .A1(n5225), .A2(n7235), .ZN(n5205) );
  OR2_X1 U6683 ( .A1(n5736), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5204) );
  INV_X1 U6684 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5202) );
  OR2_X1 U6685 ( .A1(n5228), .A2(n5202), .ZN(n5203) );
  AND4_X2 U6686 ( .A1(n5206), .A2(n5205), .A3(n5204), .A4(n5203), .ZN(n7244)
         );
  NAND2_X1 U6687 ( .A1(n5207), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5208) );
  XNOR2_X1 U6688 ( .A(n5208), .B(n5132), .ZN(n6807) );
  NAND2_X1 U6689 ( .A1(n5210), .A2(n5209), .ZN(n5216) );
  MUX2_X1 U6690 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n8004), .Z(n5211) );
  NAND2_X1 U6691 ( .A1(n5211), .A2(SI_3_), .ZN(n5233) );
  INV_X1 U6692 ( .A(n5211), .ZN(n5213) );
  INV_X1 U6693 ( .A(SI_3_), .ZN(n5212) );
  NAND2_X1 U6694 ( .A1(n5213), .A2(n5212), .ZN(n5214) );
  AND2_X1 U6695 ( .A1(n5233), .A2(n5214), .ZN(n5215) );
  NAND2_X1 U6696 ( .A1(n5216), .A2(n5215), .ZN(n5234) );
  OR2_X1 U6697 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  NAND2_X1 U6698 ( .A1(n5234), .A2(n5217), .ZN(n6512) );
  OR2_X1 U6699 ( .A1(n5354), .A2(n6512), .ZN(n5220) );
  INV_X1 U6700 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6510) );
  OAI211_X1 U6701 ( .C1(n6507), .C2(n6807), .A(n5220), .B(n5219), .ZN(n5770)
         );
  OR2_X1 U6702 ( .A1(n7244), .A2(n7477), .ZN(n5221) );
  NAND2_X1 U6703 ( .A1(n7244), .A2(n7477), .ZN(n5222) );
  NAND2_X1 U6704 ( .A1(n5223), .A2(n5222), .ZN(n7241) );
  BUF_X4 U6705 ( .A(n5224), .Z(n7420) );
  NAND2_X1 U6706 ( .A1(n7420), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5232) );
  INV_X1 U6707 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6833) );
  OR2_X1 U6708 ( .A1(n5225), .A2(n6833), .ZN(n5231) );
  INV_X1 U6709 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6710 ( .A1(n8388), .A2(n5226), .ZN(n5251) );
  NAND2_X1 U6711 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5227) );
  AND2_X1 U6712 ( .A1(n5251), .A2(n5227), .ZN(n7453) );
  OR2_X1 U6713 ( .A1(n5736), .A2(n7453), .ZN(n5230) );
  CLKBUF_X3 U6714 ( .A(n5228), .Z(n5739) );
  INV_X1 U6715 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6829) );
  OR2_X1 U6716 ( .A1(n5739), .A2(n6829), .ZN(n5229) );
  NAND2_X1 U6717 ( .A1(n5234), .A2(n5233), .ZN(n5240) );
  NAND2_X1 U6718 ( .A1(n5237), .A2(SI_4_), .ZN(n5257) );
  AND2_X1 U6719 ( .A1(n5238), .A2(n5257), .ZN(n5239) );
  NAND2_X1 U6720 ( .A1(n5240), .A2(n5239), .ZN(n5258) );
  OR2_X1 U6721 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  NAND2_X1 U6722 ( .A1(n5258), .A2(n5241), .ZN(n6516) );
  OR2_X1 U6723 ( .A1(n5354), .A2(n6516), .ZN(n5246) );
  NAND2_X1 U6724 ( .A1(n5242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6725 ( .A1(n5547), .A2(n6842), .ZN(n5244) );
  INV_X1 U6726 ( .A(n8220), .ZN(n5774) );
  NAND2_X1 U6727 ( .A1(n8537), .A2(n5774), .ZN(n5772) );
  NAND2_X1 U6728 ( .A1(n7241), .A2(n5772), .ZN(n5247) );
  NAND2_X1 U6729 ( .A1(n7323), .A2(n8220), .ZN(n5773) );
  NAND2_X1 U6730 ( .A1(n5247), .A2(n5773), .ZN(n7322) );
  NAND2_X1 U6731 ( .A1(n7420), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5256) );
  INV_X1 U6732 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5248) );
  OR2_X1 U6733 ( .A1(n5225), .A2(n5248), .ZN(n5255) );
  INV_X1 U6734 ( .A(n5251), .ZN(n5250) );
  INV_X1 U6735 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6736 ( .A1(n5250), .A2(n5249), .ZN(n5270) );
  NAND2_X1 U6737 ( .A1(n5251), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5252) );
  AND2_X1 U6738 ( .A1(n5270), .A2(n5252), .ZN(n7313) );
  OR2_X1 U6739 ( .A1(n5736), .A2(n7313), .ZN(n5254) );
  INV_X1 U6740 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7328) );
  OR2_X1 U6741 ( .A1(n5739), .A2(n7328), .ZN(n5253) );
  NAND4_X1 U6742 ( .A1(n5256), .A2(n5255), .A3(n5254), .A4(n5253), .ZN(n7443)
         );
  INV_X1 U6743 ( .A(n7443), .ZN(n7243) );
  MUX2_X1 U6744 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7998), .Z(n5259) );
  NAND2_X1 U6745 ( .A1(n5259), .A2(SI_5_), .ZN(n5277) );
  INV_X1 U6746 ( .A(n5259), .ZN(n5261) );
  INV_X1 U6747 ( .A(SI_5_), .ZN(n5260) );
  NAND2_X1 U6748 ( .A1(n5261), .A2(n5260), .ZN(n5262) );
  XNOR2_X1 U6749 ( .A(n5276), .B(n5124), .ZN(n6521) );
  OR2_X1 U6750 ( .A1(n5354), .A2(n6521), .ZN(n5267) );
  INV_X1 U6751 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6515) );
  OR2_X1 U6752 ( .A1(n5263), .A2(n9007), .ZN(n5264) );
  XNOR2_X1 U6753 ( .A(n5264), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6973) );
  NAND2_X1 U6754 ( .A1(n5547), .A2(n6973), .ZN(n5265) );
  INV_X1 U6755 ( .A(n7309), .ZN(n7330) );
  NAND2_X1 U6756 ( .A1(n7243), .A2(n7330), .ZN(n8213) );
  NAND2_X1 U6757 ( .A1(n7443), .A2(n7309), .ZN(n8221) );
  NAND2_X1 U6758 ( .A1(n8213), .A2(n8221), .ZN(n8158) );
  NAND2_X1 U6759 ( .A1(n7322), .A2(n8158), .ZN(n7321) );
  NAND2_X1 U6760 ( .A1(n7243), .A2(n7309), .ZN(n5268) );
  NAND2_X1 U6761 ( .A1(n7321), .A2(n5268), .ZN(n7439) );
  NAND2_X1 U6762 ( .A1(n5756), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5275) );
  INV_X2 U6763 ( .A(n7420), .ZN(n5759) );
  INV_X1 U6764 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5269) );
  OR2_X1 U6765 ( .A1(n5759), .A2(n5269), .ZN(n5274) );
  OR2_X2 U6766 ( .A1(n5270), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6767 ( .A1(n5270), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5271) );
  AND2_X1 U6768 ( .A1(n5317), .A2(n5271), .ZN(n7546) );
  OR2_X1 U6769 ( .A1(n5736), .A2(n7546), .ZN(n5273) );
  INV_X1 U6770 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7183) );
  OR2_X1 U6771 ( .A1(n5739), .A2(n7183), .ZN(n5272) );
  INV_X1 U6772 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U6773 ( .A1(n5276), .A2(n5124), .ZN(n5278) );
  NAND2_X1 U6774 ( .A1(n5278), .A2(n5277), .ZN(n5284) );
  MUX2_X1 U6775 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7998), .Z(n5279) );
  NAND2_X1 U6776 ( .A1(n5279), .A2(SI_6_), .ZN(n5290) );
  INV_X1 U6777 ( .A(n5279), .ZN(n5281) );
  INV_X1 U6778 ( .A(SI_6_), .ZN(n5280) );
  NAND2_X1 U6779 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  AND2_X1 U6780 ( .A1(n5290), .A2(n5282), .ZN(n5283) );
  NAND2_X1 U6781 ( .A1(n5284), .A2(n5283), .ZN(n5291) );
  OR2_X1 U6782 ( .A1(n5284), .A2(n5283), .ZN(n5285) );
  OR2_X1 U6783 ( .A1(n6519), .A2(n5354), .ZN(n5289) );
  NAND2_X1 U6784 ( .A1(n5286), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5287) );
  MUX2_X1 U6785 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5287), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5288) );
  NAND2_X1 U6786 ( .A1(n8536), .A2(n7413), .ZN(n7437) );
  NAND2_X1 U6787 ( .A1(n7439), .A2(n7437), .ZN(n7428) );
  MUX2_X1 U6788 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7998), .Z(n5292) );
  NAND2_X1 U6789 ( .A1(n5292), .A2(SI_7_), .ZN(n5309) );
  OAI21_X1 U6790 ( .B1(n5292), .B2(SI_7_), .A(n5309), .ZN(n5306) );
  XNOR2_X1 U6791 ( .A(n5308), .B(n5306), .ZN(n6531) );
  INV_X2 U6792 ( .A(n5354), .ZN(n5331) );
  NAND2_X1 U6793 ( .A1(n6531), .A2(n5331), .ZN(n5296) );
  NAND2_X1 U6794 ( .A1(n5481), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5293) );
  MUX2_X1 U6795 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5293), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5294) );
  AOI22_X1 U6796 ( .A1(n5548), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5547), .B2(
        n7197), .ZN(n5295) );
  NAND2_X1 U6797 ( .A1(n5296), .A2(n5295), .ZN(n8230) );
  NAND2_X1 U6798 ( .A1(n5756), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5303) );
  INV_X1 U6799 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5297) );
  OR2_X1 U6800 ( .A1(n5759), .A2(n5297), .ZN(n5302) );
  INV_X1 U6801 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5298) );
  XNOR2_X1 U6802 ( .A(n5317), .B(n5298), .ZN(n7568) );
  OR2_X1 U6803 ( .A1(n5736), .A2(n7568), .ZN(n5301) );
  INV_X1 U6804 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5299) );
  OR2_X1 U6805 ( .A1(n5739), .A2(n5299), .ZN(n5300) );
  INV_X1 U6806 ( .A(n7413), .ZN(n7547) );
  NAND2_X1 U6807 ( .A1(n7564), .A2(n7547), .ZN(n7438) );
  INV_X1 U6808 ( .A(n7438), .ZN(n7441) );
  NOR2_X1 U6809 ( .A1(n8228), .A2(n7441), .ZN(n5304) );
  NAND2_X1 U6810 ( .A1(n7428), .A2(n5304), .ZN(n7430) );
  NAND2_X1 U6811 ( .A1(n8230), .A2(n7649), .ZN(n5305) );
  INV_X1 U6812 ( .A(n5306), .ZN(n5307) );
  MUX2_X1 U6813 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n7998), .Z(n5325) );
  XNOR2_X1 U6814 ( .A(n5325), .B(SI_8_), .ZN(n5329) );
  NAND2_X1 U6815 ( .A1(n6534), .A2(n5331), .ZN(n5313) );
  NAND2_X1 U6816 ( .A1(n5332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5311) );
  XNOR2_X1 U6817 ( .A(n5311), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7390) );
  AOI22_X1 U6818 ( .A1(n5548), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5547), .B2(
        n7390), .ZN(n5312) );
  NAND2_X1 U6819 ( .A1(n5756), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5322) );
  INV_X1 U6820 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5314) );
  OR2_X1 U6821 ( .A1(n5759), .A2(n5314), .ZN(n5321) );
  INV_X1 U6822 ( .A(n5317), .ZN(n5316) );
  NOR2_X1 U6823 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n5315) );
  NAND2_X1 U6824 ( .A1(n5316), .A2(n5315), .ZN(n5335) );
  OAI21_X1 U6825 ( .B1(n5317), .B2(P2_REG3_REG_7__SCAN_IN), .A(
        P2_REG3_REG_8__SCAN_IN), .ZN(n5318) );
  AND2_X1 U6826 ( .A1(n5335), .A2(n5318), .ZN(n7471) );
  OR2_X1 U6827 ( .A1(n5736), .A2(n7471), .ZN(n5320) );
  INV_X1 U6828 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7389) );
  OR2_X1 U6829 ( .A1(n5739), .A2(n7389), .ZN(n5319) );
  NAND4_X1 U6830 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .ZN(n8535)
         );
  NOR2_X1 U6831 ( .A1(n7647), .A2(n7735), .ZN(n5324) );
  NAND2_X1 U6832 ( .A1(n7647), .A2(n7735), .ZN(n5323) );
  INV_X1 U6833 ( .A(n5325), .ZN(n5327) );
  INV_X1 U6834 ( .A(SI_8_), .ZN(n5326) );
  NAND2_X1 U6835 ( .A1(n5327), .A2(n5326), .ZN(n5328) );
  INV_X1 U6836 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6624) );
  MUX2_X1 U6837 ( .A(n10469), .B(n6624), .S(n8004), .Z(n5341) );
  XNOR2_X1 U6838 ( .A(n5341), .B(SI_9_), .ZN(n5343) );
  NAND2_X1 U6839 ( .A1(n6622), .A2(n5331), .ZN(n5334) );
  NOR2_X1 U6840 ( .A1(n5332), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5375) );
  OR2_X1 U6841 ( .A1(n5375), .A2(n9007), .ZN(n5356) );
  XNOR2_X1 U6842 ( .A(n5356), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7387) );
  AOI22_X1 U6843 ( .A1(n5548), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5547), .B2(
        n7387), .ZN(n5333) );
  NAND2_X1 U6844 ( .A1(n5334), .A2(n5333), .ZN(n7732) );
  NAND2_X1 U6845 ( .A1(n7420), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5340) );
  OR2_X1 U6846 ( .A1(n5225), .A2(n4655), .ZN(n5339) );
  NAND2_X1 U6847 ( .A1(n5335), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5336) );
  AND2_X1 U6848 ( .A1(n5364), .A2(n5336), .ZN(n7738) );
  OR2_X1 U6849 ( .A1(n5736), .A2(n7738), .ZN(n5338) );
  INV_X1 U6850 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7381) );
  OR2_X1 U6851 ( .A1(n5739), .A2(n7381), .ZN(n5337) );
  INV_X1 U6852 ( .A(n7886), .ZN(n8534) );
  INV_X1 U6853 ( .A(n5341), .ZN(n5342) );
  MUX2_X1 U6854 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n8004), .Z(n5345) );
  NAND2_X1 U6855 ( .A1(n5345), .A2(SI_10_), .ZN(n5371) );
  INV_X1 U6856 ( .A(n5345), .ZN(n5347) );
  INV_X1 U6857 ( .A(SI_10_), .ZN(n5346) );
  NAND2_X1 U6858 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  NAND2_X1 U6859 ( .A1(n5371), .A2(n5348), .ZN(n5351) );
  INV_X1 U6860 ( .A(n5351), .ZN(n5349) );
  INV_X1 U6861 ( .A(n5350), .ZN(n5352) );
  NAND2_X1 U6862 ( .A1(n5352), .A2(n5351), .ZN(n5353) );
  NAND2_X1 U6863 ( .A1(n5372), .A2(n5353), .ZN(n6621) );
  OR2_X1 U6864 ( .A1(n6621), .A2(n5354), .ZN(n5361) );
  INV_X1 U6865 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6866 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U6867 ( .A1(n5357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5359) );
  INV_X1 U6868 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5358) );
  XNOR2_X1 U6869 ( .A(n5359), .B(n5358), .ZN(n7821) );
  INV_X1 U6870 ( .A(n7821), .ZN(n7539) );
  AOI22_X1 U6871 ( .A1(n5548), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5547), .B2(
        n7539), .ZN(n5360) );
  NAND2_X1 U6872 ( .A1(n5756), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5369) );
  INV_X1 U6873 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5362) );
  OR2_X1 U6874 ( .A1(n5759), .A2(n5362), .ZN(n5368) );
  INV_X1 U6875 ( .A(n5364), .ZN(n5363) );
  NAND2_X1 U6876 ( .A1(n5363), .A2(n7525), .ZN(n5384) );
  NAND2_X1 U6877 ( .A1(n5364), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5365) );
  AND2_X1 U6878 ( .A1(n5384), .A2(n5365), .ZN(n7889) );
  OR2_X1 U6879 ( .A1(n5736), .A2(n7889), .ZN(n5367) );
  INV_X1 U6880 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7754) );
  OR2_X1 U6881 ( .A1(n5739), .A2(n7754), .ZN(n5366) );
  NAND4_X1 U6882 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n8533)
         );
  INV_X1 U6883 ( .A(n8533), .ZN(n7868) );
  NAND2_X1 U6884 ( .A1(n7865), .A2(n7868), .ZN(n5370) );
  MUX2_X1 U6885 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n8004), .Z(n5395) );
  XNOR2_X1 U6886 ( .A(n5395), .B(SI_11_), .ZN(n5373) );
  XNOR2_X1 U6887 ( .A(n5394), .B(n5373), .ZN(n6682) );
  NAND2_X1 U6888 ( .A1(n6682), .A2(n5331), .ZN(n5382) );
  NOR2_X1 U6889 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5374) );
  AND2_X1 U6890 ( .A1(n5375), .A2(n5374), .ZN(n5378) );
  NOR2_X1 U6891 ( .A1(n5378), .A2(n9007), .ZN(n5376) );
  MUX2_X1 U6892 ( .A(n9007), .B(n5376), .S(P2_IR_REG_11__SCAN_IN), .Z(n5380)
         );
  INV_X1 U6893 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6894 ( .A1(n5378), .A2(n5377), .ZN(n5413) );
  INV_X1 U6895 ( .A(n5413), .ZN(n5379) );
  AOI22_X1 U6896 ( .A1(n5548), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5547), .B2(
        n7823), .ZN(n5381) );
  NAND2_X1 U6897 ( .A1(n7420), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5389) );
  INV_X1 U6898 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5383) );
  OR2_X1 U6899 ( .A1(n5225), .A2(n5383), .ZN(n5388) );
  INV_X1 U6900 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7777) );
  OR2_X1 U6901 ( .A1(n5739), .A2(n7777), .ZN(n5387) );
  NAND2_X1 U6902 ( .A1(n5384), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5385) );
  AND2_X1 U6903 ( .A1(n5401), .A2(n5385), .ZN(n7934) );
  OR2_X1 U6904 ( .A1(n5736), .A2(n7934), .ZN(n5386) );
  NOR2_X1 U6905 ( .A1(n8246), .A2(n8532), .ZN(n5390) );
  INV_X1 U6906 ( .A(n8246), .ZN(n7776) );
  INV_X1 U6907 ( .A(n5395), .ZN(n5392) );
  INV_X1 U6908 ( .A(SI_11_), .ZN(n5391) );
  NAND2_X1 U6909 ( .A1(n5392), .A2(n5391), .ZN(n5393) );
  NAND2_X1 U6910 ( .A1(n5394), .A2(n5393), .ZN(n5397) );
  NAND2_X1 U6911 ( .A1(n5395), .A2(SI_11_), .ZN(n5396) );
  MUX2_X1 U6912 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n8004), .Z(n5410) );
  XNOR2_X1 U6913 ( .A(n5410), .B(SI_12_), .ZN(n5409) );
  XNOR2_X1 U6914 ( .A(n5431), .B(n5409), .ZN(n6729) );
  NAND2_X1 U6915 ( .A1(n6729), .A2(n5331), .ZN(n5400) );
  NAND2_X1 U6916 ( .A1(n5413), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5398) );
  XNOR2_X1 U6917 ( .A(n5398), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7917) );
  AOI22_X1 U6918 ( .A1(n5548), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5547), .B2(
        n7917), .ZN(n5399) );
  NAND2_X1 U6919 ( .A1(n7420), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5406) );
  INV_X1 U6920 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7911) );
  OR2_X1 U6921 ( .A1(n5225), .A2(n7911), .ZN(n5405) );
  NAND2_X1 U6922 ( .A1(n5401), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5402) );
  AND2_X1 U6923 ( .A1(n5419), .A2(n5402), .ZN(n7880) );
  OR2_X1 U6924 ( .A1(n5736), .A2(n7880), .ZN(n5404) );
  INV_X1 U6925 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7852) );
  OR2_X1 U6926 ( .A1(n5739), .A2(n7852), .ZN(n5403) );
  AND2_X1 U6927 ( .A1(n7882), .A2(n8531), .ZN(n5408) );
  OR2_X1 U6928 ( .A1(n7882), .A2(n8531), .ZN(n5407) );
  INV_X1 U6929 ( .A(n5409), .ZN(n5429) );
  NAND2_X1 U6930 ( .A1(n5431), .A2(n5429), .ZN(n5411) );
  NAND2_X1 U6931 ( .A1(n5410), .A2(SI_12_), .ZN(n5434) );
  NAND2_X1 U6932 ( .A1(n5411), .A2(n5434), .ZN(n5412) );
  MUX2_X1 U6933 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n8004), .Z(n5425) );
  XNOR2_X1 U6934 ( .A(n5425), .B(SI_13_), .ZN(n5426) );
  XNOR2_X1 U6935 ( .A(n5412), .B(n5426), .ZN(n6714) );
  NAND2_X1 U6936 ( .A1(n6714), .A2(n5331), .ZN(n5416) );
  NAND2_X1 U6937 ( .A1(n5414), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5440) );
  XNOR2_X1 U6938 ( .A(n5440), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8578) );
  AOI22_X1 U6939 ( .A1(n5548), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5547), .B2(
        n8578), .ZN(n5415) );
  NAND2_X1 U6940 ( .A1(n7420), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5424) );
  INV_X1 U6941 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8552) );
  OR2_X1 U6942 ( .A1(n5225), .A2(n8552), .ZN(n5423) );
  INV_X1 U6943 ( .A(n5419), .ZN(n5418) );
  NAND2_X1 U6944 ( .A1(n5418), .A2(n5417), .ZN(n5445) );
  NAND2_X1 U6945 ( .A1(n5419), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5420) );
  AND2_X1 U6946 ( .A1(n5445), .A2(n5420), .ZN(n7960) );
  OR2_X1 U6947 ( .A1(n5736), .A2(n7960), .ZN(n5422) );
  INV_X1 U6948 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8544) );
  OR2_X1 U6949 ( .A1(n5739), .A2(n8544), .ZN(n5421) );
  NAND2_X1 U6950 ( .A1(n7966), .A2(n8530), .ZN(n8266) );
  OR2_X1 U6951 ( .A1(n7966), .A2(n8530), .ZN(n8263) );
  NAND2_X1 U6952 ( .A1(n5425), .A2(SI_13_), .ZN(n5433) );
  INV_X1 U6953 ( .A(n5433), .ZN(n5428) );
  INV_X1 U6954 ( .A(n5426), .ZN(n5427) );
  AND2_X1 U6955 ( .A1(n5429), .A2(n5432), .ZN(n5430) );
  NAND2_X1 U6956 ( .A1(n5431), .A2(n5430), .ZN(n5438) );
  INV_X1 U6957 ( .A(n5432), .ZN(n5436) );
  AND2_X1 U6958 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  MUX2_X1 U6959 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n8004), .Z(n5456) );
  XNOR2_X1 U6960 ( .A(n5456), .B(SI_14_), .ZN(n5453) );
  XNOR2_X1 U6961 ( .A(n5455), .B(n5453), .ZN(n6770) );
  NAND2_X1 U6962 ( .A1(n6770), .A2(n5331), .ZN(n5443) );
  INV_X1 U6963 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6964 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  NAND2_X1 U6965 ( .A1(n5441), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5461) );
  XNOR2_X1 U6966 ( .A(n5461), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8587) );
  AOI22_X1 U6967 ( .A1(n5548), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8587), .B2(
        n5547), .ZN(n5442) );
  NAND2_X1 U6968 ( .A1(n7420), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5450) );
  INV_X1 U6969 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8581) );
  OR2_X1 U6970 ( .A1(n5225), .A2(n8581), .ZN(n5449) );
  INV_X1 U6971 ( .A(n5445), .ZN(n5444) );
  NAND2_X1 U6972 ( .A1(n5444), .A2(n7987), .ZN(n5466) );
  NAND2_X1 U6973 ( .A1(n5445), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5446) );
  AND2_X1 U6974 ( .A1(n5466), .A2(n5446), .ZN(n7986) );
  OR2_X1 U6975 ( .A1(n5736), .A2(n7986), .ZN(n5448) );
  INV_X1 U6976 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8565) );
  OR2_X1 U6977 ( .A1(n5739), .A2(n8565), .ZN(n5447) );
  OR2_X1 U6978 ( .A1(n7982), .A2(n8515), .ZN(n8271) );
  NAND2_X1 U6979 ( .A1(n7982), .A2(n8515), .ZN(n8272) );
  NAND2_X1 U6980 ( .A1(n8271), .A2(n8272), .ZN(n8268) );
  NAND2_X1 U6981 ( .A1(n7982), .A2(n8867), .ZN(n5451) );
  INV_X1 U6982 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U6983 ( .A1(n5455), .A2(n5454), .ZN(n5458) );
  NAND2_X1 U6984 ( .A1(n5456), .A2(SI_14_), .ZN(n5457) );
  NAND2_X1 U6985 ( .A1(n5458), .A2(n5457), .ZN(n5475) );
  MUX2_X1 U6986 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n8004), .Z(n5473) );
  XNOR2_X1 U6987 ( .A(n5473), .B(SI_15_), .ZN(n5459) );
  XNOR2_X1 U6988 ( .A(n5475), .B(n5459), .ZN(n6767) );
  NAND2_X1 U6989 ( .A1(n6767), .A2(n5331), .ZN(n5465) );
  INV_X1 U6990 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6991 ( .A1(n5461), .A2(n5460), .ZN(n5462) );
  NAND2_X1 U6992 ( .A1(n5462), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5463) );
  XNOR2_X1 U6993 ( .A(n5463), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8625) );
  AOI22_X1 U6994 ( .A1(n8625), .A2(n5547), .B1(n5548), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6995 ( .A1(n5465), .A2(n5464), .ZN(n8853) );
  NAND2_X1 U6996 ( .A1(n7420), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5471) );
  INV_X1 U6997 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8598) );
  OR2_X1 U6998 ( .A1(n5225), .A2(n8598), .ZN(n5470) );
  NAND2_X1 U6999 ( .A1(n5466), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5467) );
  AND2_X1 U7000 ( .A1(n5489), .A2(n5467), .ZN(n8855) );
  OR2_X1 U7001 ( .A1(n5736), .A2(n8855), .ZN(n5469) );
  INV_X1 U7002 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10421) );
  OR2_X1 U7003 ( .A1(n5739), .A2(n10421), .ZN(n5468) );
  OR2_X1 U7004 ( .A1(n8853), .A2(n8844), .ZN(n5472) );
  NAND2_X1 U7005 ( .A1(n8853), .A2(n8844), .ZN(n8857) );
  NOR2_X1 U7006 ( .A1(n5477), .A2(n5476), .ZN(n5474) );
  NAND2_X1 U7007 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  MUX2_X1 U7008 ( .A(n6945), .B(n10453), .S(n8004), .Z(n5497) );
  XNOR2_X1 U7009 ( .A(n5497), .B(SI_16_), .ZN(n5479) );
  XNOR2_X1 U7010 ( .A(n5496), .B(n5479), .ZN(n6944) );
  NAND2_X1 U7011 ( .A1(n6944), .A2(n5331), .ZN(n5486) );
  OR2_X1 U7012 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  NAND2_X1 U7013 ( .A1(n5482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5483) );
  MUX2_X1 U7014 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5483), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5484) );
  NAND2_X1 U7015 ( .A1(n5484), .A2(n5519), .ZN(n8641) );
  INV_X1 U7016 ( .A(n8641), .ZN(n8632) );
  AOI22_X1 U7017 ( .A1(n5548), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5547), .B2(
        n8632), .ZN(n5485) );
  NAND2_X1 U7018 ( .A1(n7420), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5494) );
  INV_X1 U7019 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10489) );
  OR2_X1 U7020 ( .A1(n5225), .A2(n10489), .ZN(n5493) );
  NAND2_X1 U7021 ( .A1(n5489), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5490) );
  AND2_X1 U7022 ( .A1(n5508), .A2(n5490), .ZN(n8434) );
  OR2_X1 U7023 ( .A1(n5736), .A2(n8434), .ZN(n5492) );
  INV_X1 U7024 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8847) );
  OR2_X1 U7025 ( .A1(n5739), .A2(n8847), .ZN(n5491) );
  NAND4_X1 U7026 ( .A1(n5494), .A2(n5493), .A3(n5492), .A4(n5491), .ZN(n8864)
         );
  INV_X1 U7027 ( .A(n8864), .ZN(n5495) );
  NAND2_X1 U7028 ( .A1(n5126), .A2(n8276), .ZN(n8842) );
  NAND2_X1 U7029 ( .A1(n5498), .A2(SI_16_), .ZN(n5499) );
  MUX2_X1 U7030 ( .A(n7079), .B(n10319), .S(n7998), .Z(n5502) );
  NAND2_X1 U7031 ( .A1(n5502), .A2(n5501), .ZN(n5518) );
  INV_X1 U7032 ( .A(n5502), .ZN(n5503) );
  NAND2_X1 U7033 ( .A1(n5503), .A2(SI_17_), .ZN(n5504) );
  NAND2_X1 U7034 ( .A1(n5518), .A2(n5504), .ZN(n5516) );
  XNOR2_X1 U7035 ( .A(n5517), .B(n5516), .ZN(n7078) );
  NAND2_X1 U7036 ( .A1(n7078), .A2(n5331), .ZN(n5507) );
  NAND2_X1 U7037 ( .A1(n5519), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5505) );
  XNOR2_X1 U7038 ( .A(n5505), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8668) );
  AOI22_X1 U7039 ( .A1(n5548), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5547), .B2(
        n8668), .ZN(n5506) );
  NAND2_X1 U7040 ( .A1(n7420), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5513) );
  INV_X1 U7041 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10346) );
  OR2_X1 U7042 ( .A1(n5225), .A2(n10346), .ZN(n5512) );
  INV_X1 U7043 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8639) );
  OR2_X1 U7044 ( .A1(n5739), .A2(n8639), .ZN(n5511) );
  NAND2_X1 U7045 ( .A1(n5508), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5509) );
  AND2_X1 U7046 ( .A1(n5528), .A2(n5509), .ZN(n8448) );
  OR2_X1 U7047 ( .A1(n5736), .A2(n8448), .ZN(n5510) );
  AND2_X1 U7048 ( .A1(n8441), .A2(n8101), .ZN(n5786) );
  INV_X1 U7049 ( .A(n5786), .ZN(n8278) );
  NAND2_X1 U7050 ( .A1(n8288), .A2(n8278), .ZN(n8190) );
  NAND2_X1 U7051 ( .A1(n8064), .A2(n8190), .ZN(n5515) );
  NAND2_X1 U7052 ( .A1(n8441), .A2(n8845), .ZN(n5514) );
  MUX2_X1 U7053 ( .A(n7237), .B(n10338), .S(n7998), .Z(n5537) );
  XNOR2_X1 U7054 ( .A(n5537), .B(SI_18_), .ZN(n5536) );
  XNOR2_X1 U7055 ( .A(n5540), .B(n5536), .ZN(n7236) );
  NAND2_X1 U7056 ( .A1(n7236), .A2(n5331), .ZN(n5526) );
  INV_X1 U7057 ( .A(n5519), .ZN(n5521) );
  NAND2_X1 U7058 ( .A1(n5746), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7059 ( .A1(n5523), .A2(n5522), .ZN(n5545) );
  OR2_X1 U7060 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  AND2_X1 U7061 ( .A1(n5545), .A2(n5524), .ZN(n8696) );
  AOI22_X1 U7062 ( .A1(n5548), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5547), .B2(
        n8696), .ZN(n5525) );
  NAND2_X1 U7063 ( .A1(n5528), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5529) );
  AND2_X1 U7064 ( .A1(n5551), .A2(n5529), .ZN(n8833) );
  OR2_X1 U7065 ( .A1(n5736), .A2(n8833), .ZN(n5533) );
  INV_X1 U7066 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8922) );
  OR2_X1 U7067 ( .A1(n5225), .A2(n8922), .ZN(n5532) );
  INV_X1 U7068 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10285) );
  OR2_X1 U7069 ( .A1(n5759), .A2(n10285), .ZN(n5531) );
  INV_X1 U7070 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8832) );
  OR2_X1 U7071 ( .A1(n5739), .A2(n8832), .ZN(n5530) );
  NAND4_X1 U7072 ( .A1(n5533), .A2(n5532), .A3(n5531), .A4(n5530), .ZN(n8529)
         );
  NOR2_X1 U7073 ( .A1(n8497), .A2(n8447), .ZN(n5535) );
  NAND2_X1 U7074 ( .A1(n8497), .A2(n8447), .ZN(n5534) );
  INV_X1 U7075 ( .A(n5536), .ZN(n5539) );
  INV_X1 U7076 ( .A(n5537), .ZN(n5538) );
  MUX2_X1 U7077 ( .A(n7335), .B(n7334), .S(n7998), .Z(n5542) );
  NAND2_X1 U7078 ( .A1(n5542), .A2(n5541), .ZN(n5559) );
  INV_X1 U7079 ( .A(n5542), .ZN(n5543) );
  NAND2_X1 U7080 ( .A1(n5543), .A2(SI_19_), .ZN(n5544) );
  NAND2_X1 U7081 ( .A1(n5559), .A2(n5544), .ZN(n5560) );
  XNOR2_X1 U7082 ( .A(n5561), .B(n5560), .ZN(n7333) );
  NAND2_X1 U7083 ( .A1(n7333), .A2(n5331), .ZN(n5550) );
  NAND2_X1 U7084 ( .A1(n5545), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5546) );
  AOI22_X1 U7085 ( .A1(n5548), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8693), .B2(
        n5547), .ZN(n5549) );
  NAND2_X1 U7086 ( .A1(n5551), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7087 ( .A1(n5569), .A2(n5552), .ZN(n8402) );
  NAND2_X1 U7088 ( .A1(n5184), .A2(n8402), .ZN(n5556) );
  INV_X1 U7089 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8082) );
  OR2_X1 U7090 ( .A1(n5759), .A2(n8082), .ZN(n5555) );
  INV_X1 U7091 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8692) );
  OR2_X1 U7092 ( .A1(n5225), .A2(n8692), .ZN(n5554) );
  INV_X1 U7093 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8088) );
  OR2_X1 U7094 ( .A1(n5739), .A2(n8088), .ZN(n5553) );
  NOR2_X1 U7095 ( .A1(n8393), .A2(n8830), .ZN(n5557) );
  NAND2_X1 U7096 ( .A1(n8393), .A2(n8830), .ZN(n5558) );
  MUX2_X1 U7097 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7998), .Z(n5575) );
  XNOR2_X1 U7098 ( .A(n5575), .B(n5577), .ZN(n5562) );
  XNOR2_X1 U7099 ( .A(n5578), .B(n5562), .ZN(n7553) );
  NAND2_X1 U7100 ( .A1(n7553), .A2(n5331), .ZN(n5565) );
  INV_X1 U7101 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7102 ( .A1(n7420), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7103 ( .A1(n5756), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5566) );
  AND2_X1 U7104 ( .A1(n5567), .A2(n5566), .ZN(n5573) );
  NAND2_X1 U7105 ( .A1(n5569), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7106 ( .A1(n5584), .A2(n5570), .ZN(n8824) );
  NAND2_X1 U7107 ( .A1(n8824), .A2(n5184), .ZN(n5572) );
  NAND2_X1 U7108 ( .A1(n7419), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5571) );
  NOR2_X1 U7109 ( .A1(n8984), .A2(n8412), .ZN(n5787) );
  INV_X1 U7110 ( .A(n5787), .ZN(n8298) );
  NAND2_X1 U7111 ( .A1(n8984), .A2(n8412), .ZN(n8295) );
  NAND2_X1 U7112 ( .A1(n8298), .A2(n8295), .ZN(n8819) );
  OR2_X1 U7113 ( .A1(n8984), .A2(n8810), .ZN(n5574) );
  NAND2_X1 U7114 ( .A1(n8818), .A2(n5574), .ZN(n8808) );
  INV_X1 U7115 ( .A(n5575), .ZN(n5576) );
  OAI21_X1 U7116 ( .B1(n5578), .B2(n5577), .A(n5576), .ZN(n5580) );
  NAND2_X1 U7117 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  NAND2_X1 U7118 ( .A1(n5580), .A2(n5579), .ZN(n5595) );
  MUX2_X1 U7119 ( .A(n10369), .B(n7646), .S(n7998), .Z(n5591) );
  XNOR2_X1 U7120 ( .A(n5591), .B(SI_21_), .ZN(n5581) );
  XNOR2_X1 U7121 ( .A(n5595), .B(n5581), .ZN(n7635) );
  NAND2_X1 U7122 ( .A1(n7635), .A2(n5331), .ZN(n5583) );
  NAND2_X1 U7123 ( .A1(n5584), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7124 ( .A1(n5603), .A2(n5585), .ZN(n8813) );
  NAND2_X1 U7125 ( .A1(n8813), .A2(n5184), .ZN(n5588) );
  AOI22_X1 U7126 ( .A1(n7420), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n5756), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7127 ( .A1(n7419), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5586) );
  AND2_X1 U7128 ( .A1(n8978), .A2(n8116), .ZN(n5788) );
  INV_X1 U7129 ( .A(n5788), .ZN(n8301) );
  NAND2_X1 U7130 ( .A1(n8299), .A2(n8301), .ZN(n8807) );
  NAND2_X1 U7131 ( .A1(n8808), .A2(n8807), .ZN(n5590) );
  OR2_X1 U7132 ( .A1(n8978), .A2(n8821), .ZN(n5589) );
  NAND2_X1 U7133 ( .A1(n5590), .A2(n5589), .ZN(n8793) );
  NOR2_X1 U7134 ( .A1(n5592), .A2(SI_21_), .ZN(n5594) );
  NAND2_X1 U7135 ( .A1(n5592), .A2(SI_21_), .ZN(n5593) );
  MUX2_X1 U7136 ( .A(n7744), .B(n7743), .S(n7998), .Z(n5596) );
  NAND2_X1 U7137 ( .A1(n5596), .A2(n10408), .ZN(n5610) );
  INV_X1 U7138 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7139 ( .A1(n5597), .A2(SI_22_), .ZN(n5598) );
  NAND2_X1 U7140 ( .A1(n5610), .A2(n5598), .ZN(n5609) );
  XNOR2_X1 U7141 ( .A(n5608), .B(n5609), .ZN(n7742) );
  NAND2_X1 U7142 ( .A1(n7742), .A2(n5331), .ZN(n5600) );
  INV_X1 U7143 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8799) );
  INV_X1 U7144 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7145 ( .A1(n5603), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7146 ( .A1(n5622), .A2(n5604), .ZN(n8797) );
  NAND2_X1 U7147 ( .A1(n8797), .A2(n5184), .ZN(n5606) );
  AOI22_X1 U7148 ( .A1(n7420), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n5756), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n5605) );
  XNOR2_X1 U7149 ( .A(n8801), .B(n8809), .ZN(n8802) );
  INV_X1 U7150 ( .A(n8802), .ZN(n8794) );
  NAND2_X1 U7151 ( .A1(n8793), .A2(n8794), .ZN(n8792) );
  OR2_X1 U7152 ( .A1(n8801), .A2(n8809), .ZN(n5607) );
  NAND2_X1 U7153 ( .A1(n8792), .A2(n5607), .ZN(n8782) );
  MUX2_X1 U7154 ( .A(n10354), .B(n10438), .S(n7998), .Z(n5612) );
  INV_X1 U7155 ( .A(SI_23_), .ZN(n5611) );
  NAND2_X1 U7156 ( .A1(n5612), .A2(n5611), .ZN(n5650) );
  INV_X1 U7157 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7158 ( .A1(n5613), .A2(SI_23_), .ZN(n5614) );
  NAND2_X1 U7159 ( .A1(n5650), .A2(n5614), .ZN(n5616) );
  NAND2_X1 U7160 ( .A1(n5615), .A2(n5616), .ZN(n5619) );
  INV_X1 U7161 ( .A(n5616), .ZN(n5617) );
  NAND2_X1 U7162 ( .A1(n5618), .A2(n5617), .ZN(n5652) );
  NAND2_X1 U7163 ( .A1(n5619), .A2(n5652), .ZN(n7814) );
  NAND2_X1 U7164 ( .A1(n7814), .A2(n5331), .ZN(n5621) );
  OR2_X2 U7165 ( .A1(n5622), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7166 ( .A1(n5622), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7167 ( .A1(n5639), .A2(n5623), .ZN(n8786) );
  NAND2_X1 U7168 ( .A1(n8786), .A2(n5184), .ZN(n5628) );
  INV_X1 U7169 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U7170 ( .A1(n7420), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7171 ( .A1(n5756), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5624) );
  OAI211_X1 U7172 ( .C1(n8785), .C2(n5739), .A(n5625), .B(n5624), .ZN(n5626)
         );
  INV_X1 U7173 ( .A(n5626), .ZN(n5627) );
  OR2_X1 U7174 ( .A1(n8788), .A2(n8480), .ZN(n5629) );
  NAND2_X1 U7175 ( .A1(n8782), .A2(n5629), .ZN(n5631) );
  NAND2_X1 U7176 ( .A1(n8788), .A2(n8480), .ZN(n5630) );
  NAND2_X1 U7177 ( .A1(n5631), .A2(n5630), .ZN(n8769) );
  NAND2_X1 U7178 ( .A1(n5652), .A2(n5650), .ZN(n5636) );
  INV_X1 U7179 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8076) );
  INV_X1 U7180 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7858) );
  MUX2_X1 U7181 ( .A(n8076), .B(n7858), .S(n7998), .Z(n5633) );
  INV_X1 U7182 ( .A(SI_24_), .ZN(n5632) );
  NAND2_X1 U7183 ( .A1(n5633), .A2(n5632), .ZN(n5649) );
  INV_X1 U7184 ( .A(n5633), .ZN(n5634) );
  NAND2_X1 U7185 ( .A1(n5634), .A2(SI_24_), .ZN(n5670) );
  AND2_X1 U7186 ( .A1(n5649), .A2(n5670), .ZN(n5635) );
  NAND2_X1 U7187 ( .A1(n7857), .A2(n5331), .ZN(n5638) );
  NAND2_X1 U7188 ( .A1(n5639), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U7189 ( .A1(n5661), .A2(n5640), .ZN(n8772) );
  NAND2_X1 U7190 ( .A1(n8772), .A2(n5184), .ZN(n5645) );
  INV_X1 U7191 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10295) );
  NAND2_X1 U7192 ( .A1(n7420), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7193 ( .A1(n7419), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5641) );
  OAI211_X1 U7194 ( .C1(n5225), .C2(n10295), .A(n5642), .B(n5641), .ZN(n5643)
         );
  INV_X1 U7195 ( .A(n5643), .ZN(n5644) );
  NOR2_X1 U7196 ( .A1(n8965), .A2(n8783), .ZN(n5647) );
  NAND2_X1 U7197 ( .A1(n8965), .A2(n8783), .ZN(n5646) );
  AND2_X1 U7198 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  NAND2_X1 U7199 ( .A1(n5652), .A2(n5651), .ZN(n5672) );
  AND2_X1 U7200 ( .A1(n5672), .A2(n5670), .ZN(n5656) );
  INV_X1 U7201 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7923) );
  MUX2_X1 U7202 ( .A(n7921), .B(n7923), .S(n7998), .Z(n5653) );
  INV_X1 U7203 ( .A(SI_25_), .ZN(n10356) );
  NAND2_X1 U7204 ( .A1(n5653), .A2(n10356), .ZN(n5673) );
  INV_X1 U7205 ( .A(n5653), .ZN(n5654) );
  NAND2_X1 U7206 ( .A1(n5654), .A2(SI_25_), .ZN(n5655) );
  NAND2_X1 U7207 ( .A1(n7920), .A2(n5331), .ZN(n5658) );
  INV_X1 U7208 ( .A(n5661), .ZN(n5660) );
  INV_X1 U7209 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7210 ( .A1(n5661), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7211 ( .A1(n5681), .A2(n5662), .ZN(n8762) );
  NAND2_X1 U7212 ( .A1(n8762), .A2(n5184), .ZN(n5667) );
  INV_X1 U7213 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10400) );
  NAND2_X1 U7214 ( .A1(n7420), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7215 ( .A1(n7419), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5663) );
  OAI211_X1 U7216 ( .C1(n5225), .C2(n10400), .A(n5664), .B(n5663), .ZN(n5665)
         );
  INV_X1 U7217 ( .A(n5665), .ZN(n5666) );
  XNOR2_X1 U7218 ( .A(n8959), .B(n8770), .ZN(n8764) );
  INV_X1 U7219 ( .A(n8764), .ZN(n8757) );
  OR2_X1 U7220 ( .A1(n8959), .A2(n8770), .ZN(n5668) );
  NAND2_X1 U7221 ( .A1(n5672), .A2(n5671), .ZN(n5674) );
  INV_X1 U7222 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7941) );
  INV_X1 U7223 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10451) );
  MUX2_X1 U7224 ( .A(n7941), .B(n10451), .S(n7998), .Z(n5676) );
  INV_X1 U7225 ( .A(SI_26_), .ZN(n5675) );
  NAND2_X1 U7226 ( .A1(n5676), .A2(n5675), .ZN(n5693) );
  INV_X1 U7227 ( .A(n5676), .ZN(n5677) );
  NAND2_X1 U7228 ( .A1(n5677), .A2(SI_26_), .ZN(n5678) );
  NAND2_X1 U7229 ( .A1(n7939), .A2(n5331), .ZN(n5680) );
  OR2_X2 U7230 ( .A1(n5681), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U7231 ( .A1(n5681), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7232 ( .A1(n5701), .A2(n5682), .ZN(n8752) );
  NAND2_X1 U7233 ( .A1(n8752), .A2(n5184), .ZN(n5687) );
  INV_X1 U7234 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U7235 ( .A1(n7420), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7236 ( .A1(n5756), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5683) );
  OAI211_X1 U7237 ( .C1(n8751), .C2(n5739), .A(n5684), .B(n5683), .ZN(n5685)
         );
  INV_X1 U7238 ( .A(n5685), .ZN(n5686) );
  NAND2_X1 U7239 ( .A1(n8953), .A2(n8758), .ZN(n5688) );
  OR2_X1 U7240 ( .A1(n8953), .A2(n8758), .ZN(n5689) );
  NAND2_X1 U7241 ( .A1(n5690), .A2(n5689), .ZN(n8739) );
  INV_X1 U7242 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5698) );
  INV_X1 U7243 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9973) );
  MUX2_X1 U7244 ( .A(n5698), .B(n9973), .S(n7998), .Z(n5695) );
  INV_X1 U7245 ( .A(SI_27_), .ZN(n5694) );
  NAND2_X1 U7246 ( .A1(n5695), .A2(n5694), .ZN(n5730) );
  INV_X1 U7247 ( .A(n5695), .ZN(n5696) );
  NAND2_X1 U7248 ( .A1(n5696), .A2(SI_27_), .ZN(n5697) );
  NAND2_X1 U7249 ( .A1(n9019), .A2(n5331), .ZN(n5700) );
  NAND2_X2 U7250 ( .A1(n5700), .A2(n5699), .ZN(n8947) );
  NAND2_X1 U7251 ( .A1(n5701), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U7252 ( .A1(n5713), .A2(n5702), .ZN(n8743) );
  INV_X1 U7253 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10399) );
  NAND2_X1 U7254 ( .A1(n7420), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U7255 ( .A1(n7419), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5703) );
  OAI211_X1 U7256 ( .C1(n5225), .C2(n10399), .A(n5704), .B(n5703), .ZN(n5705)
         );
  AOI21_X2 U7257 ( .B1(n8743), .B2(n5184), .A(n5705), .ZN(n8728) );
  NAND2_X1 U7258 ( .A1(n8947), .A2(n8728), .ZN(n8322) );
  INV_X1 U7259 ( .A(n8728), .ZN(n8749) );
  NOR2_X1 U7260 ( .A1(n8947), .A2(n8749), .ZN(n5706) );
  NAND2_X1 U7261 ( .A1(n5727), .A2(n5725), .ZN(n5707) );
  NAND2_X1 U7262 ( .A1(n5707), .A2(n5730), .ZN(n5708) );
  INV_X1 U7263 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5709) );
  INV_X1 U7264 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9970) );
  MUX2_X1 U7265 ( .A(n5709), .B(n9970), .S(n7998), .Z(n5722) );
  XNOR2_X1 U7266 ( .A(n5722), .B(SI_28_), .ZN(n5723) );
  NAND2_X1 U7267 ( .A1(n9016), .A2(n5331), .ZN(n5711) );
  INV_X1 U7268 ( .A(n5713), .ZN(n5712) );
  INV_X1 U7269 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U7270 ( .A1(n5712), .A2(n8138), .ZN(n8711) );
  NAND2_X1 U7271 ( .A1(n5713), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7272 ( .A1(n8711), .A2(n5714), .ZN(n8732) );
  INV_X1 U7273 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U7274 ( .A1(n7419), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7275 ( .A1(n5756), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5715) );
  OAI211_X1 U7276 ( .C1(n5759), .C2(n5717), .A(n5716), .B(n5715), .ZN(n5718)
         );
  NAND2_X1 U7277 ( .A1(n8944), .A2(n8368), .ZN(n5719) );
  INV_X1 U7278 ( .A(n8368), .ZN(n8740) );
  INV_X1 U7279 ( .A(SI_28_), .ZN(n5721) );
  NAND2_X1 U7280 ( .A1(n5722), .A2(n5721), .ZN(n5729) );
  INV_X1 U7281 ( .A(n5729), .ZN(n5724) );
  AND2_X1 U7282 ( .A1(n5725), .A2(n5728), .ZN(n5726) );
  INV_X1 U7283 ( .A(n5728), .ZN(n5732) );
  AND2_X1 U7284 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  NAND2_X1 U7285 ( .A1(n5734), .A2(n5733), .ZN(n7993) );
  INV_X1 U7286 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9014) );
  INV_X1 U7287 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9968) );
  MUX2_X1 U7288 ( .A(n9014), .B(n9968), .S(n7998), .Z(n7994) );
  XNOR2_X1 U7289 ( .A(n7992), .B(SI_29_), .ZN(n9012) );
  INV_X1 U7290 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7291 ( .A1(n7420), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7292 ( .A1(n5756), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U7293 ( .C1(n5740), .C2(n5739), .A(n5738), .B(n5737), .ZN(n5741)
         );
  INV_X1 U7294 ( .A(n5741), .ZN(n5742) );
  NAND2_X1 U7295 ( .A1(n7425), .A2(n5742), .ZN(n8725) );
  AND2_X1 U7296 ( .A1(n8719), .A2(n8725), .ZN(n8334) );
  INV_X1 U7297 ( .A(n8334), .ZN(n5745) );
  INV_X1 U7298 ( .A(n8719), .ZN(n5744) );
  INV_X1 U7299 ( .A(n8725), .ZN(n5743) );
  NAND2_X1 U7300 ( .A1(n5744), .A2(n5743), .ZN(n8179) );
  NAND2_X1 U7301 ( .A1(n5745), .A2(n8179), .ZN(n8326) );
  INV_X1 U7302 ( .A(n8326), .ZN(n8328) );
  NAND2_X1 U7303 ( .A1(n5749), .A2(n5748), .ZN(n5796) );
  NAND2_X1 U7304 ( .A1(n5796), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7305 ( .A1(n8357), .A2(n8693), .ZN(n5755) );
  NAND2_X1 U7306 ( .A1(n5751), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7307 ( .A1(n8191), .A2(n8350), .ZN(n5754) );
  INV_X1 U7308 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U7309 ( .A1(n7419), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7310 ( .A1(n5756), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5757) );
  OAI211_X1 U7311 ( .C1(n5759), .C2(n10397), .A(n5758), .B(n5757), .ZN(n5760)
         );
  INV_X1 U7312 ( .A(n5760), .ZN(n5761) );
  INV_X1 U7313 ( .A(n6785), .ZN(n8354) );
  NAND2_X1 U7314 ( .A1(n8354), .A2(n8698), .ZN(n5763) );
  INV_X1 U7315 ( .A(n6934), .ZN(n6935) );
  NAND2_X1 U7316 ( .A1(n6507), .A2(P2_B_REG_SCAN_IN), .ZN(n5764) );
  NAND2_X1 U7317 ( .A1(n8865), .A2(n5764), .ZN(n8708) );
  NOR2_X1 U7318 ( .A1(n8339), .A2(n8708), .ZN(n5766) );
  NAND2_X1 U7319 ( .A1(n7106), .A2(n8035), .ZN(n8193) );
  NAND2_X1 U7320 ( .A1(n7219), .A2(n8203), .ZN(n7231) );
  NAND2_X1 U7321 ( .A1(n7244), .A2(n5770), .ZN(n8219) );
  INV_X1 U7322 ( .A(n7244), .ZN(n8538) );
  NAND2_X1 U7323 ( .A1(n8538), .A2(n7477), .ZN(n8211) );
  NAND2_X1 U7324 ( .A1(n7231), .A2(n8153), .ZN(n5771) );
  NAND2_X1 U7325 ( .A1(n5773), .A2(n5772), .ZN(n8209) );
  NAND2_X1 U7326 ( .A1(n7323), .A2(n5774), .ZN(n8212) );
  NAND2_X1 U7327 ( .A1(n7320), .A2(n8221), .ZN(n7446) );
  NAND2_X1 U7328 ( .A1(n7564), .A2(n7413), .ZN(n8216) );
  AND2_X1 U7329 ( .A1(n8213), .A2(n8216), .ZN(n8225) );
  NAND2_X1 U7330 ( .A1(n7446), .A2(n8225), .ZN(n5775) );
  NAND2_X1 U7331 ( .A1(n8536), .A2(n7547), .ZN(n8227) );
  NAND2_X1 U7332 ( .A1(n5775), .A2(n8227), .ZN(n7427) );
  NAND2_X1 U7333 ( .A1(n7427), .A2(n8228), .ZN(n5776) );
  INV_X1 U7334 ( .A(n8230), .ZN(n7558) );
  NAND2_X1 U7335 ( .A1(n7558), .A2(n7649), .ZN(n8218) );
  AND2_X1 U7336 ( .A1(n7647), .A2(n8535), .ZN(n7465) );
  INV_X1 U7337 ( .A(n7647), .ZN(n5777) );
  NAND2_X1 U7338 ( .A1(n5777), .A2(n7735), .ZN(n8237) );
  NAND2_X1 U7339 ( .A1(n7732), .A2(n7886), .ZN(n8236) );
  NAND2_X1 U7340 ( .A1(n8240), .A2(n8236), .ZN(n8152) );
  AND2_X1 U7341 ( .A1(n7865), .A2(n8533), .ZN(n7747) );
  NAND2_X1 U7342 ( .A1(n8246), .A2(n7877), .ZN(n8234) );
  INV_X1 U7343 ( .A(n8234), .ZN(n5779) );
  INV_X1 U7344 ( .A(n7865), .ZN(n7869) );
  NAND2_X1 U7345 ( .A1(n7869), .A2(n7868), .ZN(n8250) );
  INV_X1 U7346 ( .A(n8250), .ZN(n5778) );
  NOR2_X1 U7347 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  NAND2_X1 U7348 ( .A1(n7774), .A2(n5780), .ZN(n5781) );
  NAND2_X1 U7349 ( .A1(n7882), .A2(n7948), .ZN(n8258) );
  NOR2_X1 U7350 ( .A1(n7966), .A2(n8261), .ZN(n5782) );
  INV_X1 U7351 ( .A(n7966), .ZN(n8260) );
  NAND2_X1 U7352 ( .A1(n7970), .A2(n8271), .ZN(n5783) );
  NAND2_X1 U7353 ( .A1(n5783), .A2(n8272), .ZN(n8837) );
  AND2_X1 U7354 ( .A1(n8853), .A2(n8436), .ZN(n8838) );
  INV_X1 U7355 ( .A(n8276), .ZN(n8189) );
  OR2_X1 U7356 ( .A1(n8853), .A2(n8436), .ZN(n8839) );
  AND2_X1 U7357 ( .A1(n5126), .A2(n8839), .ZN(n5784) );
  AND2_X1 U7358 ( .A1(n8497), .A2(n8529), .ZN(n8151) );
  NAND2_X1 U7359 ( .A1(n8989), .A2(n8447), .ZN(n8283) );
  AND2_X1 U7360 ( .A1(n8393), .A2(n8492), .ZN(n8078) );
  NAND2_X1 U7361 ( .A1(n5789), .A2(n8299), .ZN(n8803) );
  INV_X1 U7362 ( .A(n8809), .ZN(n8413) );
  OR2_X1 U7363 ( .A1(n8801), .A2(n8413), .ZN(n8303) );
  NAND2_X1 U7364 ( .A1(n8971), .A2(n8480), .ZN(n8308) );
  AND2_X1 U7365 ( .A1(n8965), .A2(n8425), .ZN(n8150) );
  INV_X1 U7366 ( .A(n8770), .ZN(n8318) );
  OR2_X1 U7367 ( .A1(n8959), .A2(n8318), .ZN(n8319) );
  NAND2_X1 U7368 ( .A1(n8763), .A2(n8319), .ZN(n8746) );
  NOR2_X1 U7369 ( .A1(n8953), .A2(n8367), .ZN(n8187) );
  NOR2_X1 U7370 ( .A1(n8746), .A2(n8187), .ZN(n5791) );
  NAND2_X1 U7371 ( .A1(n8953), .A2(n8367), .ZN(n8186) );
  XNOR2_X1 U7372 ( .A(n8178), .B(n8326), .ZN(n8721) );
  INV_X1 U7373 ( .A(n8357), .ZN(n7746) );
  NAND2_X1 U7374 ( .A1(n8191), .A2(n8185), .ZN(n6913) );
  NAND2_X1 U7375 ( .A1(n7746), .A2(n6913), .ZN(n5792) );
  NAND2_X1 U7376 ( .A1(n5792), .A2(n8352), .ZN(n5794) );
  INV_X1 U7377 ( .A(n10155), .ZN(n6937) );
  OR2_X1 U7378 ( .A1(n6937), .A2(n8357), .ZN(n7483) );
  NOR2_X1 U7379 ( .A1(n8716), .A2(n5793), .ZN(n6474) );
  OR2_X1 U7380 ( .A1(n5794), .A2(n8185), .ZN(n5795) );
  NAND2_X1 U7381 ( .A1(n5795), .A2(n8344), .ZN(n5816) );
  NAND2_X1 U7382 ( .A1(n5801), .A2(n5799), .ZN(n5812) );
  INV_X1 U7383 ( .A(P2_B_REG_SCAN_IN), .ZN(n5800) );
  XNOR2_X1 U7384 ( .A(n5812), .B(n5800), .ZN(n5807) );
  NAND2_X1 U7385 ( .A1(n5803), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5804) );
  MUX2_X1 U7386 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5804), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5806) );
  OR2_X1 U7387 ( .A1(n5811), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5810) );
  OR2_X1 U7388 ( .A1(n5808), .A2(n6725), .ZN(n5809) );
  INV_X1 U7389 ( .A(n5811), .ZN(n5814) );
  NAND2_X1 U7390 ( .A1(n4605), .A2(n5816), .ZN(n5815) );
  NOR2_X1 U7391 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .ZN(
        n5820) );
  NOR4_X1 U7392 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n5819) );
  NOR4_X1 U7393 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5818) );
  NOR4_X1 U7394 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5817) );
  NAND4_X1 U7395 ( .A1(n5820), .A2(n5819), .A3(n5818), .A4(n5817), .ZN(n5826)
         );
  NOR4_X1 U7396 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5824) );
  NOR4_X1 U7397 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5823) );
  NOR4_X1 U7398 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5822) );
  NOR4_X1 U7399 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n5821) );
  NAND4_X1 U7400 ( .A1(n5824), .A2(n5823), .A3(n5822), .A4(n5821), .ZN(n5825)
         );
  NOR2_X1 U7401 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  NAND2_X1 U7402 ( .A1(n8338), .A2(n6914), .ZN(n6924) );
  INV_X1 U7403 ( .A(n4605), .ZN(n5832) );
  NAND2_X1 U7404 ( .A1(n5832), .A2(n6462), .ZN(n6469) );
  INV_X1 U7405 ( .A(n8191), .ZN(n7636) );
  NAND2_X1 U7406 ( .A1(n7840), .A2(n7636), .ZN(n7100) );
  NAND3_X1 U7407 ( .A1(n7098), .A2(n6469), .A3(n7100), .ZN(n5833) );
  OR2_X1 U7408 ( .A1(n6474), .A2(n8884), .ZN(n5835) );
  NAND2_X1 U7409 ( .A1(n8884), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7410 ( .A1(n5835), .A2(n5120), .ZN(P2_U3488) );
  NOR2_X1 U7411 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5839) );
  NOR2_X2 U7412 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5838) );
  NOR2_X2 U7413 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5837) );
  NOR2_X2 U7414 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5836) );
  AND4_X2 U7415 ( .A1(n5839), .A2(n5838), .A3(n5837), .A4(n5836), .ZN(n5845)
         );
  NOR2_X2 U7416 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5929) );
  NOR2_X1 U7417 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5840) );
  NAND2_X1 U7418 ( .A1(n5929), .A2(n5840), .ZN(n5970) );
  INV_X1 U7419 ( .A(n5970), .ZN(n5844) );
  NAND3_X2 U7420 ( .A1(n5845), .A2(n5844), .A3(n5843), .ZN(n6206) );
  NOR2_X1 U7421 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5850) );
  NOR2_X1 U7422 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5849) );
  NOR2_X1 U7423 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5848) );
  NAND2_X1 U7424 ( .A1(n9954), .A2(n5895), .ZN(n5853) );
  NAND2_X1 U7425 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5855) );
  NAND2_X1 U7426 ( .A1(n5896), .A2(n5855), .ZN(n5856) );
  XNOR2_X2 U7427 ( .A(n5856), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U7428 ( .A1(n5923), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7429 ( .A1(n5857), .A2(n5858), .ZN(n6200) );
  INV_X2 U7430 ( .A(n6200), .ZN(n5953) );
  NAND2_X1 U7431 ( .A1(n5953), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7432 ( .A1(n5955), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5860) );
  INV_X1 U7433 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6545) );
  OR2_X1 U7434 ( .A1(n5975), .A2(n6545), .ZN(n5859) );
  NAND4_X1 U7435 ( .A1(n5862), .A2(n5861), .A3(n5860), .A4(n5859), .ZN(n6689)
         );
  INV_X1 U7436 ( .A(n6206), .ZN(n5863) );
  NAND2_X1 U7437 ( .A1(n5863), .A2(n5847), .ZN(n5880) );
  NAND3_X1 U7438 ( .A1(n5864), .A2(n5882), .A3(n5881), .ZN(n5865) );
  NOR2_X2 U7439 ( .A1(n5880), .A2(n5865), .ZN(n5878) );
  NAND2_X1 U7440 ( .A1(n5878), .A2(n5866), .ZN(n5876) );
  INV_X1 U7441 ( .A(n5876), .ZN(n5868) );
  INV_X1 U7442 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7443 ( .A1(n5868), .A2(n5867), .ZN(n5885) );
  NAND2_X1 U7444 ( .A1(n5886), .A2(n5869), .ZN(n5870) );
  INV_X1 U7445 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7446 ( .A1(n5873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5874) );
  NAND2_X2 U7447 ( .A1(n6416), .A2(n5875), .ZN(n6504) );
  XNOR2_X2 U7448 ( .A(n5877), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U7449 ( .A1(n6689), .A2(n6394), .ZN(n5901) );
  NAND2_X1 U7450 ( .A1(n5880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6230) );
  INV_X1 U7451 ( .A(n6248), .ZN(n5883) );
  NAND2_X1 U7452 ( .A1(n5883), .A2(n5882), .ZN(n6250) );
  XNOR2_X2 U7453 ( .A(n5884), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6264) );
  NAND2_X2 U7454 ( .A1(n6736), .A2(n6437), .ZN(n9459) );
  NAND2_X1 U7455 ( .A1(n5887), .A2(n5886), .ZN(n6432) );
  NAND2_X1 U7456 ( .A1(n5889), .A2(n6264), .ZN(n7082) );
  OAI211_X2 U7457 ( .C1(n9459), .C2(n9465), .A(n6504), .B(n7082), .ZN(n5981)
         );
  MUX2_X1 U7458 ( .A(n6264), .B(n5890), .S(n9453), .Z(n5892) );
  NOR2_X2 U7459 ( .A1(n5891), .A2(n9453), .ZN(n6434) );
  OAI21_X2 U7460 ( .B1(n5892), .B2(n6434), .A(n6504), .ZN(n5918) );
  NAND2_X2 U7461 ( .A1(n5981), .A2(n5918), .ZN(n5947) );
  INV_X1 U7462 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6547) );
  NOR2_X1 U7463 ( .A1(n5910), .A2(n5893), .ZN(n5894) );
  XNOR2_X1 U7464 ( .A(n5894), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9974) );
  XNOR2_X2 U7465 ( .A(n5896), .B(n5895), .ZN(n6443) );
  NAND2_X1 U7466 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n5897) );
  MUX2_X1 U7467 ( .A(n6547), .B(n9974), .S(n5949), .Z(n6963) );
  INV_X1 U7468 ( .A(n6963), .ZN(n6741) );
  NAND2_X1 U7469 ( .A1(n5947), .A2(n6741), .ZN(n5900) );
  AND2_X1 U7470 ( .A1(n5901), .A2(n5900), .ZN(n5906) );
  OR2_X1 U7471 ( .A1(n6504), .A2(n6545), .ZN(n5902) );
  NAND2_X1 U7472 ( .A1(n6689), .A2(n4517), .ZN(n5905) );
  OAI22_X1 U7473 ( .A1(n6963), .A2(n6377), .B1(n6547), .B2(n6504), .ZN(n5903)
         );
  INV_X1 U7474 ( .A(n5903), .ZN(n5904) );
  NAND2_X1 U7475 ( .A1(n5905), .A2(n5904), .ZN(n6646) );
  NAND2_X1 U7476 ( .A1(n5906), .A2(n6408), .ZN(n5907) );
  INV_X1 U7477 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7478 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5908) );
  XNOR2_X1 U7479 ( .A(n5909), .B(n5908), .ZN(n6544) );
  NAND2_X1 U7480 ( .A1(n5947), .A2(n10074), .ZN(n5917) );
  NAND2_X1 U7481 ( .A1(n5953), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7482 ( .A1(n5923), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5914) );
  INV_X1 U7483 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7484 ( .A1(n6672), .A2(n6394), .ZN(n5916) );
  AOI22_X1 U7485 ( .A1(n6672), .A2(n4517), .B1(n6394), .B2(n10074), .ZN(n5920)
         );
  XNOR2_X1 U7486 ( .A(n5919), .B(n5920), .ZN(n9059) );
  NAND2_X1 U7487 ( .A1(n9061), .A2(n9059), .ZN(n9060) );
  INV_X1 U7488 ( .A(n5919), .ZN(n5921) );
  NAND2_X1 U7489 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  NAND2_X1 U7490 ( .A1(n9060), .A2(n5922), .ZN(n6676) );
  NAND2_X1 U7491 ( .A1(n5923), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7492 ( .A1(n5953), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5927) );
  INV_X1 U7493 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5924) );
  OR2_X1 U7494 ( .A1(n5975), .A2(n5924), .ZN(n5925) );
  NAND2_X1 U7495 ( .A1(n9483), .A2(n6394), .ZN(n5937) );
  OR2_X1 U7496 ( .A1(n6513), .A2(n5948), .ZN(n5934) );
  OR2_X1 U7497 ( .A1(n6284), .A2(n4966), .ZN(n5933) );
  OR2_X1 U7498 ( .A1(n5929), .A2(n5872), .ZN(n5931) );
  INV_X1 U7499 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7500 ( .A1(n5931), .A2(n5930), .ZN(n5950) );
  OAI21_X1 U7501 ( .B1(n5931), .B2(n5930), .A(n5950), .ZN(n6664) );
  OR2_X1 U7502 ( .A1(n5949), .A2(n6664), .ZN(n5932) );
  NAND2_X1 U7503 ( .A1(n5947), .A2(n7204), .ZN(n5936) );
  NAND2_X1 U7504 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  NAND2_X1 U7505 ( .A1(n9483), .A2(n4517), .ZN(n5941) );
  NAND2_X1 U7506 ( .A1(n7204), .A2(n6394), .ZN(n5940) );
  NAND2_X1 U7507 ( .A1(n5941), .A2(n5940), .ZN(n5942) );
  NAND2_X1 U7508 ( .A1(n6676), .A2(n6678), .ZN(n5946) );
  INV_X1 U7509 ( .A(n5942), .ZN(n5943) );
  NAND2_X1 U7510 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  NAND2_X1 U7511 ( .A1(n5946), .A2(n5945), .ZN(n6716) );
  NAND2_X1 U7514 ( .A1(n5950), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5951) );
  XNOR2_X1 U7515 ( .A(n5951), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6559) );
  AOI22_X1 U7516 ( .A1(n6265), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n6522), .B2(
        n6559), .ZN(n5952) );
  OAI21_X1 U7517 ( .B1(n6512), .B2(n5948), .A(n5952), .ZN(n10049) );
  NAND2_X1 U7518 ( .A1(n5935), .A2(n10049), .ZN(n5961) );
  NAND2_X1 U7519 ( .A1(n6489), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5959) );
  INV_X1 U7520 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7521 ( .A1(n5953), .A2(n5954), .ZN(n5958) );
  NAND2_X1 U7522 ( .A1(n6490), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5957) );
  INV_X1 U7523 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6566) );
  OR2_X1 U7524 ( .A1(n5975), .A2(n6566), .ZN(n5956) );
  NAND2_X1 U7525 ( .A1(n9482), .A2(n6394), .ZN(n5960) );
  NAND2_X1 U7526 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  XNOR2_X1 U7527 ( .A(n5962), .B(n6408), .ZN(n5967) );
  NAND2_X1 U7528 ( .A1(n9482), .A2(n4517), .ZN(n5964) );
  NAND2_X1 U7529 ( .A1(n10049), .A2(n6360), .ZN(n5963) );
  NAND2_X1 U7530 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  NAND2_X1 U7531 ( .A1(n6716), .A2(n6718), .ZN(n5969) );
  INV_X1 U7532 ( .A(n5965), .ZN(n5966) );
  NAND2_X1 U7533 ( .A1(n5967), .A2(n5966), .ZN(n5968) );
  NAND2_X1 U7534 ( .A1(n5969), .A2(n5968), .ZN(n6904) );
  INV_X1 U7535 ( .A(n6904), .ZN(n5984) );
  OR2_X1 U7536 ( .A1(n6516), .A2(n5948), .ZN(n5973) );
  NAND2_X1 U7537 ( .A1(n5988), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5971) );
  XNOR2_X1 U7538 ( .A(n5971), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U7539 ( .A1(n6265), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6522), .B2(
        n10003), .ZN(n5972) );
  AND2_X2 U7540 ( .A1(n5973), .A2(n5972), .ZN(n10085) );
  INV_X2 U7541 ( .A(n9224), .ZN(n6489) );
  NAND2_X1 U7542 ( .A1(n6489), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5979) );
  NOR2_X1 U7543 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5974) );
  NOR2_X1 U7544 ( .A1(n5992), .A2(n5974), .ZN(n7163) );
  NAND2_X1 U7545 ( .A1(n5953), .A2(n7163), .ZN(n5978) );
  NAND2_X1 U7546 ( .A1(n6490), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7547 ( .A1(n6401), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5976) );
  OAI22_X1 U7548 ( .A1(n10085), .A2(n6233), .B1(n7022), .B2(n6377), .ZN(n5980)
         );
  XNOR2_X1 U7549 ( .A(n5980), .B(n6481), .ZN(n5986) );
  OAI22_X1 U7550 ( .A1(n10085), .A2(n6377), .B1(n7022), .B2(n5982), .ZN(n5985)
         );
  XNOR2_X1 U7551 ( .A(n5986), .B(n5985), .ZN(n6909) );
  INV_X1 U7552 ( .A(n6909), .ZN(n5983) );
  NAND2_X1 U7553 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  OR2_X1 U7554 ( .A1(n6521), .A2(n5948), .ZN(n5991) );
  OR2_X1 U7555 ( .A1(n5988), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7556 ( .A1(n6003), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5989) );
  XNOR2_X1 U7557 ( .A(n5989), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U7558 ( .A1(n6265), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6522), .B2(
        n6587), .ZN(n5990) );
  NAND2_X1 U7559 ( .A1(n5991), .A2(n5990), .ZN(n7048) );
  NAND2_X1 U7560 ( .A1(n7048), .A2(n6210), .ZN(n5998) );
  NAND2_X1 U7561 ( .A1(n6489), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7562 ( .A1(n5992), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6009) );
  OAI21_X1 U7563 ( .B1(n5992), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6009), .ZN(
        n7088) );
  INV_X1 U7564 ( .A(n7088), .ZN(n7026) );
  NAND2_X1 U7565 ( .A1(n6269), .A2(n7026), .ZN(n5995) );
  NAND2_X1 U7566 ( .A1(n6490), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7567 ( .A1(n6401), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5993) );
  NAND4_X1 U7568 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n9481)
         );
  NAND2_X1 U7569 ( .A1(n9481), .A2(n6360), .ZN(n5997) );
  NAND2_X1 U7570 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  AND2_X1 U7571 ( .A1(n9481), .A2(n4517), .ZN(n6000) );
  AOI21_X1 U7572 ( .B1(n7048), .B2(n6360), .A(n6000), .ZN(n7020) );
  INV_X1 U7573 ( .A(n6001), .ZN(n6002) );
  NOR2_X1 U7574 ( .A1(n6003), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6040) );
  OR2_X1 U7575 ( .A1(n6040), .A2(n5872), .ZN(n6005) );
  INV_X1 U7576 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7577 ( .A1(n6005), .A2(n6004), .ZN(n6025) );
  OAI21_X1 U7578 ( .B1(n6005), .B2(n6004), .A(n6025), .ZN(n6611) );
  INV_X1 U7579 ( .A(n6611), .ZN(n6597) );
  AOI22_X1 U7580 ( .A1(n6265), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6522), .B2(
        n6597), .ZN(n6006) );
  NAND2_X1 U7581 ( .A1(n7274), .A2(n6210), .ZN(n6016) );
  NAND2_X1 U7582 ( .A1(n6489), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6014) );
  INV_X1 U7583 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6008) );
  NOR2_X1 U7584 ( .A1(n6009), .A2(n6008), .ZN(n6029) );
  AND2_X1 U7585 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  NOR2_X1 U7586 ( .A1(n6029), .A2(n6010), .ZN(n7273) );
  NAND2_X1 U7587 ( .A1(n5953), .A2(n7273), .ZN(n6013) );
  NAND2_X1 U7588 ( .A1(n6490), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7589 ( .A1(n6401), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6011) );
  NAND4_X1 U7590 ( .A1(n6014), .A2(n6013), .A3(n6012), .A4(n6011), .ZN(n9480)
         );
  NAND2_X1 U7591 ( .A1(n9480), .A2(n6360), .ZN(n6015) );
  NAND2_X1 U7592 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  XNOR2_X1 U7593 ( .A(n6017), .B(n6481), .ZN(n6019) );
  AND2_X1 U7594 ( .A1(n9480), .A2(n4517), .ZN(n6018) );
  AOI21_X1 U7595 ( .B1(n7274), .B2(n6360), .A(n6018), .ZN(n6020) );
  XNOR2_X1 U7596 ( .A(n6019), .B(n6020), .ZN(n7071) );
  INV_X1 U7597 ( .A(n6019), .ZN(n6021) );
  NAND2_X1 U7598 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  INV_X2 U7599 ( .A(n5948), .ZN(n6024) );
  NAND2_X1 U7600 ( .A1(n6531), .A2(n6024), .ZN(n6028) );
  NAND2_X1 U7601 ( .A1(n6025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6026) );
  XNOR2_X1 U7602 ( .A(n6026), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6631) );
  AOI22_X1 U7603 ( .A1(n6265), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6522), .B2(
        n6631), .ZN(n6027) );
  NAND2_X1 U7604 ( .A1(n6029), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6047) );
  OR2_X1 U7605 ( .A1(n6029), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6030) );
  AND2_X1 U7606 ( .A1(n6047), .A2(n6030), .ZN(n7299) );
  NAND2_X1 U7607 ( .A1(n6269), .A2(n7299), .ZN(n6034) );
  NAND2_X1 U7608 ( .A1(n6489), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7609 ( .A1(n6490), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6032) );
  INV_X1 U7610 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6609) );
  OR2_X1 U7611 ( .A1(n5975), .A2(n6609), .ZN(n6031) );
  NAND4_X1 U7612 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(n9479)
         );
  AND2_X1 U7613 ( .A1(n9479), .A2(n4517), .ZN(n6035) );
  AOI21_X1 U7614 ( .B1(n7355), .B2(n6360), .A(n6035), .ZN(n7134) );
  NAND2_X1 U7615 ( .A1(n7355), .A2(n6210), .ZN(n6037) );
  NAND2_X1 U7616 ( .A1(n9479), .A2(n6360), .ZN(n6036) );
  NAND2_X1 U7617 ( .A1(n6037), .A2(n6036), .ZN(n6038) );
  XNOR2_X1 U7618 ( .A(n6038), .B(n6481), .ZN(n7133) );
  INV_X1 U7619 ( .A(n6059), .ZN(n6057) );
  NAND2_X1 U7620 ( .A1(n6534), .A2(n6024), .ZN(n6045) );
  NOR2_X1 U7621 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6039) );
  NAND2_X1 U7622 ( .A1(n6040), .A2(n6039), .ZN(n6042) );
  NAND2_X1 U7623 ( .A1(n6042), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6041) );
  MUX2_X1 U7624 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6041), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n6043) );
  AOI22_X1 U7625 ( .A1(n6265), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6522), .B2(
        n6630), .ZN(n6044) );
  NAND2_X1 U7626 ( .A1(n7285), .A2(n6210), .ZN(n6054) );
  NAND2_X1 U7627 ( .A1(n6489), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7628 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  AND2_X1 U7629 ( .A1(n6066), .A2(n6048), .ZN(n7516) );
  NAND2_X1 U7630 ( .A1(n6269), .A2(n7516), .ZN(n6051) );
  NAND2_X1 U7631 ( .A1(n6490), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6050) );
  INV_X1 U7632 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6625) );
  OR2_X1 U7633 ( .A1(n5975), .A2(n6625), .ZN(n6049) );
  NAND4_X1 U7634 ( .A1(n6052), .A2(n6051), .A3(n6050), .A4(n6049), .ZN(n9478)
         );
  NAND2_X1 U7635 ( .A1(n9478), .A2(n6360), .ZN(n6053) );
  NAND2_X1 U7636 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  XNOR2_X1 U7637 ( .A(n6055), .B(n6481), .ZN(n6058) );
  NAND2_X1 U7638 ( .A1(n6057), .A2(n6056), .ZN(n6062) );
  AND2_X1 U7639 ( .A1(n9478), .A2(n4517), .ZN(n6061) );
  AOI21_X1 U7640 ( .B1(n7285), .B2(n6360), .A(n6061), .ZN(n7511) );
  NAND2_X1 U7641 ( .A1(n6081), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6063) );
  XNOR2_X1 U7642 ( .A(n6063), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6699) );
  AOI22_X1 U7643 ( .A1(n6265), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6522), .B2(
        n6699), .ZN(n6064) );
  NAND2_X1 U7644 ( .A1(n7347), .A2(n6210), .ZN(n6074) );
  AND2_X1 U7645 ( .A1(n6066), .A2(n6638), .ZN(n6067) );
  NOR2_X1 U7646 ( .A1(n6084), .A2(n6067), .ZN(n7611) );
  NAND2_X1 U7647 ( .A1(n6269), .A2(n7611), .ZN(n6072) );
  NAND2_X1 U7648 ( .A1(n6489), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7649 ( .A1(n6490), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6070) );
  INV_X1 U7650 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6068) );
  OR2_X1 U7651 ( .A1(n5975), .A2(n6068), .ZN(n6069) );
  NAND4_X1 U7652 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n9477)
         );
  NAND2_X1 U7653 ( .A1(n9477), .A2(n6360), .ZN(n6073) );
  NAND2_X1 U7654 ( .A1(n6074), .A2(n6073), .ZN(n6075) );
  XNOR2_X1 U7655 ( .A(n6075), .B(n6481), .ZN(n6077) );
  AND2_X1 U7656 ( .A1(n9477), .A2(n4517), .ZN(n6076) );
  AOI21_X1 U7657 ( .B1(n7347), .B2(n6360), .A(n6076), .ZN(n6078) );
  XNOR2_X1 U7658 ( .A(n6077), .B(n6078), .ZN(n7605) );
  INV_X1 U7659 ( .A(n6077), .ZN(n6079) );
  NAND2_X1 U7660 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  INV_X1 U7661 ( .A(n6098), .ZN(n6096) );
  OR2_X1 U7662 ( .A1(n6621), .A2(n5948), .ZN(n6083) );
  NOR2_X1 U7663 ( .A1(n6081), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6124) );
  OR2_X1 U7664 ( .A1(n6124), .A2(n5872), .ZN(n6101) );
  XNOR2_X1 U7665 ( .A(n6101), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6709) );
  AOI22_X1 U7666 ( .A1(n6265), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6522), .B2(
        n6709), .ZN(n6082) );
  NAND2_X1 U7667 ( .A1(n7489), .A2(n6210), .ZN(n6093) );
  NAND2_X1 U7668 ( .A1(n6489), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6091) );
  NOR2_X1 U7669 ( .A1(n6084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7670 ( .A1(n6269), .A2(n5122), .ZN(n6090) );
  INV_X1 U7671 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6087) );
  OR2_X1 U7672 ( .A1(n6086), .A2(n6087), .ZN(n6089) );
  INV_X1 U7673 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6702) );
  OR2_X1 U7674 ( .A1(n5975), .A2(n6702), .ZN(n6088) );
  NAND4_X1 U7675 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n9476)
         );
  NAND2_X1 U7676 ( .A1(n9476), .A2(n6360), .ZN(n6092) );
  NAND2_X1 U7677 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  XNOR2_X1 U7678 ( .A(n6094), .B(n6408), .ZN(n6097) );
  INV_X1 U7679 ( .A(n6097), .ZN(n6095) );
  AND2_X1 U7680 ( .A1(n9476), .A2(n4517), .ZN(n6099) );
  AOI21_X1 U7681 ( .B1(n7489), .B2(n6360), .A(n6099), .ZN(n7803) );
  NAND2_X1 U7682 ( .A1(n6682), .A2(n6024), .ZN(n6105) );
  INV_X1 U7683 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7684 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  NAND2_X1 U7685 ( .A1(n6102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6103) );
  XNOR2_X1 U7686 ( .A(n6103), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6872) );
  AOI22_X1 U7687 ( .A1(n6872), .A2(n6522), .B1(n6265), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7688 ( .A1(n6105), .A2(n6104), .ZN(n7497) );
  NAND2_X1 U7689 ( .A1(n7497), .A2(n6210), .ZN(n6114) );
  NAND2_X1 U7690 ( .A1(n6489), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7691 ( .A1(n6106), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6129) );
  OR2_X1 U7692 ( .A1(n6106), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6107) );
  AND2_X1 U7693 ( .A1(n6129), .A2(n6107), .ZN(n9178) );
  NAND2_X1 U7694 ( .A1(n6269), .A2(n9178), .ZN(n6111) );
  INV_X1 U7695 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6108) );
  OR2_X1 U7696 ( .A1(n6086), .A2(n6108), .ZN(n6110) );
  INV_X1 U7697 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6865) );
  OR2_X1 U7698 ( .A1(n5975), .A2(n6865), .ZN(n6109) );
  NAND4_X1 U7699 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n9475)
         );
  NAND2_X1 U7700 ( .A1(n9475), .A2(n6360), .ZN(n6113) );
  NAND2_X1 U7701 ( .A1(n6114), .A2(n6113), .ZN(n6115) );
  XNOR2_X1 U7702 ( .A(n6115), .B(n6408), .ZN(n6117) );
  AND2_X1 U7703 ( .A1(n9475), .A2(n4517), .ZN(n6116) );
  AOI21_X1 U7704 ( .B1(n7497), .B2(n6360), .A(n6116), .ZN(n6118) );
  NAND2_X1 U7705 ( .A1(n6117), .A2(n6118), .ZN(n9078) );
  INV_X1 U7706 ( .A(n6117), .ZN(n6120) );
  INV_X1 U7707 ( .A(n6118), .ZN(n6119) );
  NAND2_X1 U7708 ( .A1(n6120), .A2(n6119), .ZN(n6121) );
  AND2_X1 U7709 ( .A1(n9078), .A2(n6121), .ZN(n9170) );
  NAND2_X1 U7710 ( .A1(n6122), .A2(n9170), .ZN(n9077) );
  NAND2_X1 U7711 ( .A1(n9077), .A2(n9078), .ZN(n6145) );
  NAND2_X1 U7712 ( .A1(n6729), .A2(n6024), .ZN(n6127) );
  NOR2_X1 U7713 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6123) );
  NAND2_X1 U7714 ( .A1(n6124), .A2(n6123), .ZN(n6147) );
  NAND2_X1 U7715 ( .A1(n6147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6125) );
  XNOR2_X1 U7716 ( .A(n6125), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6871) );
  AOI22_X1 U7717 ( .A1(n6265), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6871), .B2(
        n6522), .ZN(n6126) );
  NAND2_X1 U7718 ( .A1(n7616), .A2(n6210), .ZN(n6137) );
  NAND2_X1 U7719 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  AND2_X1 U7720 ( .A1(n6151), .A2(n6130), .ZN(n9089) );
  NAND2_X1 U7721 ( .A1(n6269), .A2(n9089), .ZN(n6135) );
  NAND2_X1 U7722 ( .A1(n6489), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7723 ( .A1(n6490), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6133) );
  INV_X1 U7724 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6131) );
  OR2_X1 U7725 ( .A1(n5975), .A2(n6131), .ZN(n6132) );
  NAND4_X1 U7726 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n10103)
         );
  NAND2_X1 U7727 ( .A1(n10103), .A2(n6360), .ZN(n6136) );
  NAND2_X1 U7728 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  XNOR2_X1 U7729 ( .A(n6138), .B(n6408), .ZN(n6140) );
  AND2_X1 U7730 ( .A1(n10103), .A2(n4517), .ZN(n6139) );
  AOI21_X1 U7731 ( .B1(n7616), .B2(n6360), .A(n6139), .ZN(n6141) );
  NAND2_X1 U7732 ( .A1(n6140), .A2(n6141), .ZN(n6146) );
  INV_X1 U7733 ( .A(n6140), .ZN(n6143) );
  INV_X1 U7734 ( .A(n6141), .ZN(n6142) );
  NAND2_X1 U7735 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  AND2_X1 U7736 ( .A1(n6146), .A2(n6144), .ZN(n9079) );
  NAND2_X1 U7737 ( .A1(n6714), .A2(n6024), .ZN(n6150) );
  NAND2_X1 U7738 ( .A1(n6166), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6148) );
  XNOR2_X1 U7739 ( .A(n6148), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7037) );
  AOI22_X1 U7740 ( .A1(n7037), .A2(n6522), .B1(n6265), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7741 ( .A1(n7760), .A2(n6210), .ZN(n6159) );
  NAND2_X1 U7742 ( .A1(n6489), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7743 ( .A1(n6151), .A2(n6880), .ZN(n6152) );
  AND2_X1 U7744 ( .A1(n6171), .A2(n6152), .ZN(n9155) );
  NAND2_X1 U7745 ( .A1(n6269), .A2(n9155), .ZN(n6156) );
  NAND2_X1 U7746 ( .A1(n6490), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6155) );
  INV_X1 U7747 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6153) );
  OR2_X1 U7748 ( .A1(n5975), .A2(n6153), .ZN(n6154) );
  NAND4_X1 U7749 ( .A1(n6157), .A2(n6156), .A3(n6155), .A4(n6154), .ZN(n9474)
         );
  NAND2_X1 U7750 ( .A1(n9474), .A2(n6360), .ZN(n6158) );
  NAND2_X1 U7751 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  XNOR2_X1 U7752 ( .A(n6160), .B(n6481), .ZN(n6162) );
  AND2_X1 U7753 ( .A1(n9474), .A2(n4517), .ZN(n6161) );
  AOI21_X1 U7754 ( .B1(n7760), .B2(n6360), .A(n6161), .ZN(n6163) );
  XNOR2_X1 U7755 ( .A(n6162), .B(n6163), .ZN(n9150) );
  NAND2_X1 U7756 ( .A1(n9147), .A2(n9150), .ZN(n9149) );
  INV_X1 U7757 ( .A(n6162), .ZN(n6164) );
  NAND2_X1 U7758 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7759 ( .A1(n6770), .A2(n6024), .ZN(n6169) );
  NAND2_X1 U7760 ( .A1(n6167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6191) );
  XNOR2_X1 U7761 ( .A(n6191), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7036) );
  AOI22_X1 U7762 ( .A1(n7036), .A2(n6522), .B1(n6265), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7763 ( .A1(n9892), .A2(n6210), .ZN(n6180) );
  NOR2_X2 U7764 ( .A1(n6171), .A2(n6170), .ZN(n6196) );
  AND2_X1 U7765 ( .A1(n6171), .A2(n6170), .ZN(n6172) );
  NOR2_X1 U7766 ( .A1(n6196), .A2(n6172), .ZN(n9032) );
  NAND2_X1 U7767 ( .A1(n9032), .A2(n5953), .ZN(n6178) );
  INV_X1 U7768 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6174) );
  INV_X1 U7769 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6173) );
  OAI22_X1 U7770 ( .A1(n6086), .A2(n6174), .B1(n9224), .B2(n6173), .ZN(n6175)
         );
  INV_X1 U7771 ( .A(n6175), .ZN(n6177) );
  INV_X1 U7772 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7370) );
  OR2_X1 U7773 ( .A1(n5975), .A2(n7370), .ZN(n6176) );
  OR2_X1 U7774 ( .A1(n9878), .A2(n6377), .ZN(n6179) );
  NAND2_X1 U7775 ( .A1(n6180), .A2(n6179), .ZN(n6181) );
  XNOR2_X1 U7776 ( .A(n6181), .B(n6408), .ZN(n6182) );
  NAND2_X1 U7777 ( .A1(n6183), .A2(n6182), .ZN(n6189) );
  NAND2_X1 U7778 ( .A1(n6184), .A2(n6189), .ZN(n9027) );
  INV_X1 U7779 ( .A(n9027), .ZN(n6188) );
  NAND2_X1 U7780 ( .A1(n9892), .A2(n6360), .ZN(n6186) );
  OR2_X1 U7781 ( .A1(n9878), .A2(n5982), .ZN(n6185) );
  NAND2_X1 U7782 ( .A1(n6186), .A2(n6185), .ZN(n9028) );
  INV_X1 U7783 ( .A(n9028), .ZN(n6187) );
  NAND2_X1 U7784 ( .A1(n6188), .A2(n6187), .ZN(n9025) );
  NAND2_X1 U7785 ( .A1(n9025), .A2(n6189), .ZN(n9099) );
  NAND2_X1 U7786 ( .A1(n6767), .A2(n6024), .ZN(n6195) );
  INV_X1 U7787 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7788 ( .A1(n6191), .A2(n6190), .ZN(n6192) );
  NAND2_X1 U7789 ( .A1(n6192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6193) );
  XNOR2_X1 U7790 ( .A(n6193), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7576) );
  AOI22_X1 U7791 ( .A1(n7576), .A2(n6522), .B1(n6265), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7792 ( .A1(n9527), .A2(n6210), .ZN(n6202) );
  NAND2_X1 U7793 ( .A1(n6196), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6211) );
  OR2_X1 U7794 ( .A1(n6196), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7795 ( .A1(n6211), .A2(n6197), .ZN(n9211) );
  AOI22_X1 U7796 ( .A1(n6489), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n6490), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n6199) );
  INV_X1 U7797 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9887) );
  OR2_X1 U7798 ( .A1(n5975), .A2(n9887), .ZN(n6198) );
  OAI211_X1 U7799 ( .C1(n9211), .C2(n6200), .A(n6199), .B(n6198), .ZN(n9754)
         );
  NAND2_X1 U7800 ( .A1(n9754), .A2(n6360), .ZN(n6201) );
  NAND2_X1 U7801 ( .A1(n6202), .A2(n6201), .ZN(n6203) );
  XNOR2_X1 U7802 ( .A(n6203), .B(n6408), .ZN(n6221) );
  NAND2_X1 U7803 ( .A1(n9527), .A2(n6360), .ZN(n6205) );
  NAND2_X1 U7804 ( .A1(n9754), .A2(n4517), .ZN(n6204) );
  AND2_X1 U7805 ( .A1(n6221), .A2(n9205), .ZN(n6225) );
  NAND2_X1 U7806 ( .A1(n6944), .A2(n6024), .ZN(n6209) );
  NAND2_X1 U7807 ( .A1(n6206), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6207) );
  XNOR2_X1 U7808 ( .A(n6207), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7574) );
  AOI22_X1 U7809 ( .A1(n6265), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6522), .B2(
        n7574), .ZN(n6208) );
  NAND2_X2 U7810 ( .A1(n6209), .A2(n6208), .ZN(n9872) );
  NAND2_X1 U7811 ( .A1(n9872), .A2(n6210), .ZN(n6217) );
  NAND2_X1 U7812 ( .A1(n6211), .A2(n7582), .ZN(n6212) );
  AND2_X1 U7813 ( .A1(n6235), .A2(n6212), .ZN(n9756) );
  NAND2_X1 U7814 ( .A1(n9756), .A2(n5953), .ZN(n6215) );
  AOI22_X1 U7815 ( .A1(n6489), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n6490), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n6214) );
  INV_X1 U7816 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7703) );
  OR2_X1 U7817 ( .A1(n5975), .A2(n7703), .ZN(n6213) );
  NAND2_X1 U7818 ( .A1(n9735), .A2(n6360), .ZN(n6216) );
  NAND2_X1 U7819 ( .A1(n6217), .A2(n6216), .ZN(n6218) );
  XNOR2_X1 U7820 ( .A(n6218), .B(n6481), .ZN(n6226) );
  NAND2_X1 U7821 ( .A1(n9872), .A2(n6360), .ZN(n6220) );
  OR2_X1 U7822 ( .A1(n9880), .A2(n5982), .ZN(n6219) );
  NAND2_X1 U7823 ( .A1(n6220), .A2(n6219), .ZN(n6227) );
  NAND2_X1 U7824 ( .A1(n6226), .A2(n6227), .ZN(n9106) );
  INV_X1 U7825 ( .A(n9106), .ZN(n6223) );
  INV_X1 U7826 ( .A(n6221), .ZN(n9101) );
  INV_X1 U7827 ( .A(n9205), .ZN(n6222) );
  INV_X1 U7828 ( .A(n6226), .ZN(n6229) );
  INV_X1 U7829 ( .A(n6227), .ZN(n6228) );
  NAND2_X1 U7830 ( .A1(n6229), .A2(n6228), .ZN(n9105) );
  NAND2_X1 U7831 ( .A1(n7078), .A2(n6024), .ZN(n6232) );
  XNOR2_X1 U7832 ( .A(n6230), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10042) );
  AOI22_X1 U7833 ( .A1(n6265), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6522), .B2(
        n10042), .ZN(n6231) );
  NAND2_X1 U7834 ( .A1(n9743), .A2(n6210), .ZN(n6241) );
  AND2_X1 U7835 ( .A1(n6235), .A2(n6234), .ZN(n6236) );
  NOR2_X2 U7836 ( .A1(n6235), .A2(n6234), .ZN(n6253) );
  INV_X1 U7837 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U7838 ( .A1(n6489), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7839 ( .A1(n6490), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6237) );
  OAI211_X1 U7840 ( .C1(n10307), .C2(n5975), .A(n6238), .B(n6237), .ZN(n6239)
         );
  OR2_X1 U7841 ( .A1(n9869), .A2(n6377), .ZN(n6240) );
  NAND2_X1 U7842 ( .A1(n6241), .A2(n6240), .ZN(n6242) );
  XNOR2_X1 U7843 ( .A(n6242), .B(n6408), .ZN(n9116) );
  NOR2_X1 U7844 ( .A1(n9869), .A2(n5982), .ZN(n6243) );
  AOI21_X1 U7845 ( .B1(n9743), .B2(n6360), .A(n6243), .ZN(n9115) );
  AND2_X1 U7846 ( .A1(n9116), .A2(n9115), .ZN(n6247) );
  INV_X1 U7847 ( .A(n9116), .ZN(n6245) );
  INV_X1 U7848 ( .A(n9115), .ZN(n6244) );
  NAND2_X1 U7849 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  NAND2_X1 U7850 ( .A1(n7236), .A2(n6024), .ZN(n6252) );
  NAND2_X1 U7851 ( .A1(n6248), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6249) );
  AND2_X1 U7852 ( .A1(n6250), .A2(n6249), .ZN(n9489) );
  AOI22_X1 U7853 ( .A1(n6265), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6522), .B2(
        n9489), .ZN(n6251) );
  OR2_X1 U7854 ( .A1(n6253), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7855 ( .A1(n6253), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6268) );
  AND2_X1 U7856 ( .A1(n6254), .A2(n6268), .ZN(n9717) );
  NAND2_X1 U7857 ( .A1(n9717), .A2(n5953), .ZN(n6259) );
  INV_X1 U7858 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10457) );
  NAND2_X1 U7859 ( .A1(n6489), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7860 ( .A1(n6401), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6255) );
  OAI211_X1 U7861 ( .C1(n6086), .C2(n10457), .A(n6256), .B(n6255), .ZN(n6257)
         );
  INV_X1 U7862 ( .A(n6257), .ZN(n6258) );
  NOR2_X1 U7863 ( .A1(n9860), .A2(n5982), .ZN(n6260) );
  AOI21_X1 U7864 ( .B1(n9534), .B2(n6360), .A(n6260), .ZN(n9184) );
  NAND2_X1 U7865 ( .A1(n9534), .A2(n6210), .ZN(n6262) );
  NAND2_X1 U7866 ( .A1(n9704), .A2(n6360), .ZN(n6261) );
  NAND2_X1 U7867 ( .A1(n6262), .A2(n6261), .ZN(n6263) );
  XNOR2_X1 U7868 ( .A(n6263), .B(n6408), .ZN(n9047) );
  NAND2_X1 U7869 ( .A1(n7333), .A2(n6024), .ZN(n6267) );
  AOI22_X1 U7870 ( .A1(n6265), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6522), .B2(
        n6264), .ZN(n6266) );
  NAND2_X1 U7871 ( .A1(n9935), .A2(n6210), .ZN(n6275) );
  AOI21_X1 U7872 ( .B1(n10357), .B2(n6268), .A(n6287), .ZN(n9705) );
  NAND2_X1 U7873 ( .A1(n6269), .A2(n9705), .ZN(n6273) );
  NAND2_X1 U7874 ( .A1(n6489), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7875 ( .A1(n6490), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6271) );
  INV_X1 U7876 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9852) );
  OR2_X1 U7877 ( .A1(n5975), .A2(n9852), .ZN(n6270) );
  NAND4_X1 U7878 ( .A1(n6273), .A2(n6272), .A3(n6271), .A4(n6270), .ZN(n9537)
         );
  NAND2_X1 U7879 ( .A1(n9537), .A2(n6360), .ZN(n6274) );
  NAND2_X1 U7880 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  XNOR2_X1 U7881 ( .A(n6276), .B(n6481), .ZN(n6279) );
  NAND2_X1 U7882 ( .A1(n9935), .A2(n6360), .ZN(n6278) );
  NAND2_X1 U7883 ( .A1(n9537), .A2(n4517), .ZN(n6277) );
  NAND2_X1 U7884 ( .A1(n6278), .A2(n6277), .ZN(n9049) );
  NAND2_X1 U7885 ( .A1(n6279), .A2(n9049), .ZN(n9135) );
  OAI21_X1 U7886 ( .B1(n9184), .B2(n9047), .A(n9135), .ZN(n6298) );
  INV_X1 U7887 ( .A(n6279), .ZN(n9050) );
  NAND2_X1 U7888 ( .A1(n9047), .A2(n9184), .ZN(n6280) );
  NAND2_X1 U7889 ( .A1(n6280), .A2(n9049), .ZN(n6283) );
  INV_X1 U7890 ( .A(n9184), .ZN(n6281) );
  NOR2_X1 U7891 ( .A1(n9049), .A2(n6281), .ZN(n6282) );
  AOI22_X1 U7892 ( .A1(n9050), .A2(n6283), .B1(n6282), .B2(n9047), .ZN(n6297)
         );
  NAND2_X1 U7893 ( .A1(n7553), .A2(n6024), .ZN(n6286) );
  INV_X1 U7894 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7555) );
  OR2_X1 U7895 ( .A1(n8017), .A2(n7555), .ZN(n6285) );
  NAND2_X1 U7896 ( .A1(n9842), .A2(n6210), .ZN(n6294) );
  NAND2_X1 U7897 ( .A1(n6489), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6292) );
  INV_X1 U7898 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9139) );
  INV_X1 U7899 ( .A(n6287), .ZN(n6288) );
  NAND2_X1 U7900 ( .A1(n6287), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6308) );
  INV_X1 U7901 ( .A(n6308), .ZN(n6306) );
  AOI21_X1 U7902 ( .B1(n9139), .B2(n6288), .A(n6306), .ZN(n9695) );
  NAND2_X1 U7903 ( .A1(n6269), .A2(n9695), .ZN(n6291) );
  NAND2_X1 U7904 ( .A1(n6490), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7905 ( .A1(n6401), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6289) );
  NAND4_X1 U7906 ( .A1(n6292), .A2(n6291), .A3(n6290), .A4(n6289), .ZN(n9287)
         );
  NAND2_X1 U7907 ( .A1(n9287), .A2(n6360), .ZN(n6293) );
  NAND2_X1 U7908 ( .A1(n6294), .A2(n6293), .ZN(n6295) );
  XNOR2_X1 U7909 ( .A(n6295), .B(n6408), .ZN(n6299) );
  AND2_X1 U7910 ( .A1(n9287), .A2(n4517), .ZN(n6296) );
  AOI21_X1 U7911 ( .B1(n9842), .B2(n6360), .A(n6296), .ZN(n6300) );
  NAND2_X1 U7912 ( .A1(n6299), .A2(n6300), .ZN(n9134) );
  INV_X1 U7913 ( .A(n6299), .ZN(n6302) );
  INV_X1 U7914 ( .A(n6300), .ZN(n6301) );
  NAND2_X1 U7915 ( .A1(n6302), .A2(n6301), .ZN(n9133) );
  NAND2_X1 U7916 ( .A1(n6303), .A2(n9133), .ZN(n9066) );
  INV_X1 U7917 ( .A(n9066), .ZN(n6318) );
  NAND2_X1 U7918 ( .A1(n7635), .A2(n6024), .ZN(n6305) );
  OR2_X1 U7919 ( .A1(n8017), .A2(n7646), .ZN(n6304) );
  NAND2_X2 U7920 ( .A1(n6305), .A2(n6304), .ZN(n9682) );
  NAND2_X1 U7921 ( .A1(n9682), .A2(n6210), .ZN(n6314) );
  NAND2_X1 U7922 ( .A1(n6489), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6312) );
  INV_X1 U7923 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U7924 ( .A1(n6306), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6324) );
  INV_X1 U7925 ( .A(n6324), .ZN(n6307) );
  AOI21_X1 U7926 ( .B1(n9071), .B2(n6308), .A(n6307), .ZN(n9683) );
  NAND2_X1 U7927 ( .A1(n6269), .A2(n9683), .ZN(n6311) );
  NAND2_X1 U7928 ( .A1(n6490), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7929 ( .A1(n6401), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6309) );
  NAND4_X1 U7930 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n9542)
         );
  NAND2_X1 U7931 ( .A1(n9542), .A2(n6360), .ZN(n6313) );
  NAND2_X1 U7932 ( .A1(n6314), .A2(n6313), .ZN(n6315) );
  XNOR2_X1 U7933 ( .A(n6315), .B(n6408), .ZN(n6320) );
  AND2_X1 U7934 ( .A1(n9542), .A2(n4517), .ZN(n6316) );
  AOI21_X1 U7935 ( .B1(n9682), .B2(n6360), .A(n6316), .ZN(n6319) );
  XNOR2_X1 U7936 ( .A(n6320), .B(n6319), .ZN(n9070) );
  INV_X1 U7937 ( .A(n9070), .ZN(n6317) );
  NAND2_X1 U7938 ( .A1(n6318), .A2(n6317), .ZN(n9068) );
  NAND2_X1 U7939 ( .A1(n6320), .A2(n6319), .ZN(n6321) );
  NAND2_X1 U7940 ( .A1(n7742), .A2(n6024), .ZN(n6323) );
  OR2_X1 U7941 ( .A1(n8017), .A2(n7743), .ZN(n6322) );
  NAND2_X1 U7942 ( .A1(n9831), .A2(n6210), .ZN(n6330) );
  NAND2_X1 U7943 ( .A1(n6489), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6328) );
  AOI21_X1 U7944 ( .B1(n9164), .B2(n6324), .A(n6336), .ZN(n9661) );
  NAND2_X1 U7945 ( .A1(n6269), .A2(n9661), .ZN(n6327) );
  NAND2_X1 U7946 ( .A1(n6490), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7947 ( .A1(n6401), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6325) );
  NAND4_X1 U7948 ( .A1(n6328), .A2(n6327), .A3(n6326), .A4(n6325), .ZN(n9822)
         );
  NAND2_X1 U7949 ( .A1(n9822), .A2(n6360), .ZN(n6329) );
  NAND2_X1 U7950 ( .A1(n6330), .A2(n6329), .ZN(n6331) );
  XNOR2_X1 U7951 ( .A(n6331), .B(n6408), .ZN(n6332) );
  OAI22_X1 U7952 ( .A1(n9663), .A2(n6377), .B1(n9680), .B2(n5982), .ZN(n9161)
         );
  NAND2_X1 U7953 ( .A1(n6333), .A2(n6332), .ZN(n9159) );
  NAND2_X1 U7954 ( .A1(n7814), .A2(n6024), .ZN(n6335) );
  OR2_X1 U7955 ( .A1(n8017), .A2(n10438), .ZN(n6334) );
  NAND2_X2 U7956 ( .A1(n6335), .A2(n6334), .ZN(n9655) );
  NAND2_X1 U7957 ( .A1(n9655), .A2(n6210), .ZN(n6343) );
  NAND2_X1 U7958 ( .A1(n6336), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6351) );
  OAI21_X1 U7959 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n6336), .A(n6351), .ZN(
        n6337) );
  INV_X1 U7960 ( .A(n6337), .ZN(n9647) );
  NAND2_X1 U7961 ( .A1(n5953), .A2(n9647), .ZN(n6341) );
  NAND2_X1 U7962 ( .A1(n5923), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6340) );
  INV_X1 U7963 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10409) );
  OR2_X1 U7964 ( .A1(n6086), .A2(n10409), .ZN(n6339) );
  NAND2_X1 U7965 ( .A1(n6401), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6338) );
  NAND4_X1 U7966 ( .A1(n6341), .A2(n6340), .A3(n6339), .A4(n6338), .ZN(n9631)
         );
  NAND2_X1 U7967 ( .A1(n9631), .A2(n6360), .ZN(n6342) );
  NAND2_X1 U7968 ( .A1(n6343), .A2(n6342), .ZN(n6344) );
  XNOR2_X1 U7969 ( .A(n6344), .B(n6481), .ZN(n6348) );
  NAND2_X1 U7970 ( .A1(n9655), .A2(n6360), .ZN(n6346) );
  NAND2_X1 U7971 ( .A1(n9631), .A2(n4517), .ZN(n6345) );
  NAND2_X1 U7972 ( .A1(n6346), .A2(n6345), .ZN(n6347) );
  NAND2_X1 U7973 ( .A1(n6348), .A2(n6347), .ZN(n9037) );
  NOR2_X1 U7974 ( .A1(n6348), .A2(n6347), .ZN(n9036) );
  NAND2_X1 U7975 ( .A1(n7857), .A2(n6024), .ZN(n6350) );
  OR2_X1 U7976 ( .A1(n8017), .A2(n7858), .ZN(n6349) );
  NAND2_X2 U7977 ( .A1(n6350), .A2(n6349), .ZN(n9922) );
  NAND2_X1 U7978 ( .A1(n9922), .A2(n6210), .ZN(n6357) );
  AOI21_X1 U7979 ( .B1(n6351), .B2(n9127), .A(n6368), .ZN(n9636) );
  NAND2_X1 U7980 ( .A1(n5953), .A2(n9636), .ZN(n6355) );
  NAND2_X1 U7981 ( .A1(n6489), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U7982 ( .A1(n6401), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6353) );
  INV_X1 U7983 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10467) );
  OR2_X1 U7984 ( .A1(n6086), .A2(n10467), .ZN(n6352) );
  NAND4_X1 U7985 ( .A1(n6355), .A2(n6354), .A3(n6353), .A4(n6352), .ZN(n9821)
         );
  NAND2_X1 U7986 ( .A1(n9821), .A2(n6360), .ZN(n6356) );
  NAND2_X1 U7987 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  XNOR2_X1 U7988 ( .A(n6358), .B(n6408), .ZN(n6362) );
  AND2_X1 U7989 ( .A1(n9821), .A2(n4517), .ZN(n6359) );
  AOI21_X1 U7990 ( .B1(n9922), .B2(n6360), .A(n6359), .ZN(n6361) );
  NAND2_X1 U7991 ( .A1(n6362), .A2(n6361), .ZN(n6363) );
  OAI21_X1 U7992 ( .B1(n6362), .B2(n6361), .A(n6363), .ZN(n9125) );
  NAND2_X1 U7993 ( .A1(n7920), .A2(n6024), .ZN(n6365) );
  OR2_X1 U7994 ( .A1(n8017), .A2(n7923), .ZN(n6364) );
  NAND2_X2 U7995 ( .A1(n6365), .A2(n6364), .ZN(n9622) );
  NAND2_X1 U7996 ( .A1(n9622), .A2(n6210), .ZN(n6375) );
  NAND2_X1 U7997 ( .A1(n5923), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6373) );
  INV_X1 U7998 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6367) );
  INV_X1 U7999 ( .A(n6368), .ZN(n6366) );
  NAND2_X1 U8000 ( .A1(n6367), .A2(n6366), .ZN(n6369) );
  AND2_X2 U8001 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n6368), .ZN(n6382) );
  INV_X1 U8002 ( .A(n6382), .ZN(n6384) );
  NAND2_X1 U8003 ( .A1(n5953), .A2(n9613), .ZN(n6372) );
  NAND2_X1 U8004 ( .A1(n6490), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U8005 ( .A1(n6401), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6370) );
  NAND4_X1 U8006 ( .A1(n6373), .A2(n6372), .A3(n6371), .A4(n6370), .ZN(n9798)
         );
  NAND2_X1 U8007 ( .A1(n9798), .A2(n6360), .ZN(n6374) );
  NAND2_X1 U8008 ( .A1(n6375), .A2(n6374), .ZN(n6376) );
  XNOR2_X1 U8009 ( .A(n6376), .B(n6481), .ZN(n6379) );
  OAI22_X1 U8010 ( .A1(n9919), .A2(n6377), .B1(n9549), .B2(n5982), .ZN(n6378)
         );
  XNOR2_X1 U8011 ( .A(n6379), .B(n6378), .ZN(n9092) );
  NOR2_X1 U8012 ( .A1(n6379), .A2(n6378), .ZN(n9195) );
  NAND2_X1 U8013 ( .A1(n7939), .A2(n6024), .ZN(n6381) );
  OR2_X1 U8014 ( .A1(n8017), .A2(n10451), .ZN(n6380) );
  NAND2_X1 U8015 ( .A1(n9233), .A2(n6210), .ZN(n6391) );
  INV_X1 U8016 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U8017 ( .A1(n6384), .A2(n6383), .ZN(n6385) );
  NAND2_X1 U8018 ( .A1(n5953), .A2(n9599), .ZN(n6389) );
  NAND2_X1 U8019 ( .A1(n6489), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U8020 ( .A1(n6490), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U8021 ( .A1(n6401), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8022 ( .A1(n9806), .A2(n6360), .ZN(n6390) );
  NAND2_X1 U8023 ( .A1(n6391), .A2(n6390), .ZN(n6392) );
  XNOR2_X1 U8024 ( .A(n6392), .B(n6408), .ZN(n6395) );
  AND2_X1 U8025 ( .A1(n9806), .A2(n4517), .ZN(n6393) );
  AOI21_X1 U8026 ( .B1(n9233), .B2(n6360), .A(n6393), .ZN(n6396) );
  XNOR2_X1 U8027 ( .A(n6395), .B(n6396), .ZN(n9194) );
  INV_X1 U8028 ( .A(n6395), .ZN(n6398) );
  INV_X1 U8029 ( .A(n6396), .ZN(n6397) );
  AND2_X1 U8030 ( .A1(n6398), .A2(n6397), .ZN(n6414) );
  NAND2_X1 U8031 ( .A1(n9019), .A2(n6024), .ZN(n6400) );
  OR2_X1 U8032 ( .A1(n8017), .A2(n9973), .ZN(n6399) );
  NAND2_X1 U8033 ( .A1(n9591), .A2(n6210), .ZN(n6407) );
  XNOR2_X1 U8034 ( .A(n6448), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U8035 ( .A1(n5953), .A2(n9584), .ZN(n6405) );
  NAND2_X1 U8036 ( .A1(n5923), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U8037 ( .A1(n6490), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6403) );
  NAND2_X1 U8038 ( .A1(n6401), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U8039 ( .A1(n9797), .A2(n6360), .ZN(n6406) );
  NAND2_X1 U8040 ( .A1(n6407), .A2(n6406), .ZN(n6409) );
  XNOR2_X1 U8041 ( .A(n6409), .B(n6408), .ZN(n6412) );
  AND2_X1 U8042 ( .A1(n9797), .A2(n4517), .ZN(n6410) );
  AOI21_X1 U8043 ( .B1(n9591), .B2(n6360), .A(n6410), .ZN(n6411) );
  NAND2_X1 U8044 ( .A1(n6412), .A2(n6411), .ZN(n6497) );
  OAI21_X1 U8045 ( .B1(n6412), .B2(n6411), .A(n6497), .ZN(n6413) );
  OAI21_X1 U8046 ( .B1(n9193), .B2(n6414), .A(n6413), .ZN(n6415) );
  INV_X1 U8047 ( .A(n6415), .ZN(n6436) );
  INV_X1 U8048 ( .A(n6430), .ZN(n7925) );
  NAND2_X1 U8049 ( .A1(n7925), .A2(P1_B_REG_SCAN_IN), .ZN(n6417) );
  MUX2_X1 U8050 ( .A(n6417), .B(P1_B_REG_SCAN_IN), .S(n6416), .Z(n6418) );
  OR2_X1 U8051 ( .A1(n6416), .A2(n7938), .ZN(n9953) );
  NOR4_X1 U8052 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6428) );
  NOR4_X1 U8053 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6427) );
  INV_X1 U8054 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10064) );
  INV_X1 U8055 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10316) );
  INV_X1 U8056 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10272) );
  INV_X1 U8057 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10335) );
  NAND4_X1 U8058 ( .A1(n10064), .A2(n10316), .A3(n10272), .A4(n10335), .ZN(
        n6425) );
  NOR4_X1 U8059 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6423) );
  NOR4_X1 U8060 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6422) );
  NOR4_X1 U8061 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6421) );
  NOR4_X1 U8062 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6420) );
  NAND4_X1 U8063 ( .A1(n6423), .A2(n6422), .A3(n6421), .A4(n6420), .ZN(n6424)
         );
  NOR4_X1 U8064 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n6425), .A4(n6424), .ZN(n6426) );
  NAND3_X1 U8065 ( .A1(n6428), .A2(n6427), .A3(n6426), .ZN(n6753) );
  NOR2_X1 U8066 ( .A1(n6753), .A2(n10411), .ZN(n6429) );
  OR2_X1 U8067 ( .A1(n9951), .A2(n6429), .ZN(n6431) );
  OR2_X1 U8068 ( .A1(n7938), .A2(n6430), .ZN(n9952) );
  NAND2_X1 U8069 ( .A1(n6431), .A2(n9952), .ZN(n6686) );
  NOR2_X1 U8070 ( .A1(n6762), .A2(n6686), .ZN(n6439) );
  INV_X1 U8071 ( .A(n6505), .ZN(n6523) );
  INV_X1 U8072 ( .A(n9219), .ZN(n9950) );
  NOR2_X1 U8073 ( .A1(n10082), .A2(n9282), .ZN(n6435) );
  INV_X1 U8074 ( .A(n6756), .ZN(n6438) );
  NAND2_X1 U8075 ( .A1(n9282), .A2(n9459), .ZN(n6687) );
  OAI21_X1 U8076 ( .B1(n6439), .B2(n6438), .A(n6687), .ZN(n6671) );
  INV_X1 U8077 ( .A(n6504), .ZN(n6440) );
  OAI21_X1 U8078 ( .B1(n6671), .B2(n6440), .A(P1_STATE_REG_SCAN_IN), .ZN(n6441) );
  NAND2_X1 U8079 ( .A1(n6505), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9466) );
  NAND2_X2 U8080 ( .A1(n6441), .A2(n9466), .ZN(n9210) );
  INV_X1 U8081 ( .A(n6442), .ZN(n6458) );
  NAND2_X1 U8082 ( .A1(n9282), .A2(n6443), .ZN(n9879) );
  OR2_X1 U8083 ( .A1(n9879), .A2(n9459), .ZN(n6444) );
  NAND2_X1 U8084 ( .A1(n6489), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6453) );
  INV_X1 U8085 ( .A(n6448), .ZN(n6446) );
  AND2_X1 U8086 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6445) );
  NAND2_X1 U8087 ( .A1(n6446), .A2(n6445), .ZN(n9558) );
  INV_X1 U8088 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6455) );
  INV_X1 U8089 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6447) );
  OAI21_X1 U8090 ( .B1(n6448), .B2(n6455), .A(n6447), .ZN(n6449) );
  NAND2_X1 U8091 ( .A1(n5953), .A2(n9572), .ZN(n6452) );
  NAND2_X1 U8092 ( .A1(n6490), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6451) );
  INV_X1 U8093 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9787) );
  OR2_X1 U8094 ( .A1(n5975), .A2(n9787), .ZN(n6450) );
  NAND4_X1 U8095 ( .A1(n6453), .A2(n6452), .A3(n6451), .A4(n6450), .ZN(n9789)
         );
  NOR2_X1 U8096 ( .A1(n9209), .A2(n9774), .ZN(n6457) );
  INV_X1 U8097 ( .A(n6443), .ZN(n6651) );
  OR2_X1 U8098 ( .A1(n9877), .A2(n9459), .ZN(n6454) );
  OAI22_X1 U8099 ( .A1(n9189), .A2(n9616), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6455), .ZN(n6456) );
  AOI211_X1 U8100 ( .C1(n9584), .C2(n9210), .A(n6457), .B(n6456), .ZN(n6460)
         );
  OR2_X1 U8101 ( .A1(n6458), .A2(n4606), .ZN(n6459) );
  NAND3_X1 U8102 ( .A1(n6461), .A2(n6460), .A3(n4588), .ZN(P1_U3214) );
  INV_X1 U8103 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6475) );
  INV_X1 U8104 ( .A(n6462), .ZN(n6463) );
  NOR2_X1 U8105 ( .A1(n4596), .A2(n8352), .ZN(n6464) );
  AND2_X1 U8106 ( .A1(n6464), .A2(n8357), .ZN(n6919) );
  AND2_X1 U8107 ( .A1(n7102), .A2(n6919), .ZN(n6465) );
  NOR2_X1 U8108 ( .A1(n8355), .A2(n6465), .ZN(n6466) );
  INV_X1 U8109 ( .A(n6467), .ZN(n6468) );
  INV_X1 U8110 ( .A(n6933), .ZN(n6471) );
  OR2_X1 U8111 ( .A1(n8037), .A2(n8338), .ZN(n6918) );
  OAI21_X1 U8112 ( .B1(n6918), .B2(n6919), .A(n8876), .ZN(n6922) );
  AND2_X1 U8113 ( .A1(n7102), .A2(n6922), .ZN(n6470) );
  NAND2_X1 U8114 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  MUX2_X1 U8115 ( .A(n6475), .B(n6474), .S(n10580), .Z(n6476) );
  NAND2_X1 U8116 ( .A1(n6476), .A2(n5127), .ZN(P2_U3456) );
  NAND2_X1 U8117 ( .A1(n9016), .A2(n6024), .ZN(n6478) );
  OR2_X1 U8118 ( .A1(n8017), .A2(n9970), .ZN(n6477) );
  NAND2_X2 U8119 ( .A1(n6478), .A2(n6477), .ZN(n9578) );
  NAND2_X1 U8120 ( .A1(n9578), .A2(n6210), .ZN(n6480) );
  NAND2_X1 U8121 ( .A1(n9789), .A2(n6360), .ZN(n6479) );
  NAND2_X1 U8122 ( .A1(n6480), .A2(n6479), .ZN(n6482) );
  XNOR2_X1 U8123 ( .A(n6482), .B(n6481), .ZN(n6484) );
  AOI22_X1 U8124 ( .A1(n9578), .A2(n6360), .B1(n4517), .B2(n9789), .ZN(n6483)
         );
  XNOR2_X1 U8125 ( .A(n6484), .B(n6483), .ZN(n6486) );
  INV_X1 U8126 ( .A(n6486), .ZN(n6498) );
  NAND3_X1 U8127 ( .A1(n6498), .A2(n9206), .A3(n6497), .ZN(n6485) );
  OR2_X2 U8128 ( .A1(n6487), .A2(n6485), .ZN(n6503) );
  NAND3_X1 U8129 ( .A1(n6487), .A2(n6486), .A3(n9206), .ZN(n6502) );
  INV_X1 U8130 ( .A(n9558), .ZN(n6488) );
  NAND2_X1 U8131 ( .A1(n5953), .A2(n6488), .ZN(n6494) );
  NAND2_X1 U8132 ( .A1(n6489), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U8133 ( .A1(n6490), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6492) );
  INV_X1 U8134 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10454) );
  OR2_X1 U8135 ( .A1(n5975), .A2(n10454), .ZN(n6491) );
  NAND4_X1 U8136 ( .A1(n6494), .A2(n6493), .A3(n6492), .A4(n6491), .ZN(n9781)
         );
  INV_X1 U8137 ( .A(n9781), .ZN(n9575) );
  NAND2_X1 U8138 ( .A1(n9210), .A2(n9572), .ZN(n6496) );
  INV_X1 U8139 ( .A(n9189), .ZN(n9215) );
  AOI22_X1 U8140 ( .A1(n9215), .A2(n9797), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6495) );
  OAI211_X1 U8141 ( .C1(n9575), .C2(n9209), .A(n6496), .B(n6495), .ZN(n6500)
         );
  NOR3_X1 U8142 ( .A1(n6498), .A2(n6497), .A3(n9145), .ZN(n6499) );
  AOI211_X1 U8143 ( .C1(n9578), .C2(n9142), .A(n6500), .B(n6499), .ZN(n6501)
         );
  NAND3_X1 U8144 ( .A1(n6503), .A2(n6502), .A3(n6501), .ZN(P1_U3220) );
  OR3_X2 U8145 ( .A1(n6505), .A2(n6504), .A3(P1_U3086), .ZN(n9484) );
  NAND2_X1 U8146 ( .A1(n6926), .A2(n8344), .ZN(n6506) );
  NAND2_X1 U8147 ( .A1(n6506), .A2(n6923), .ZN(n6786) );
  NAND2_X1 U8148 ( .A1(n6786), .A2(n6507), .ZN(n6508) );
  NAND2_X1 U8149 ( .A1(n6508), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  AND2_X1 U8150 ( .A1(n6511), .A2(P2_U3151), .ZN(n7811) );
  INV_X2 U8151 ( .A(n7811), .ZN(n9023) );
  INV_X2 U8152 ( .A(n9021), .ZN(n9013) );
  OAI222_X1 U8153 ( .A1(P2_U3151), .A2(n8062), .B1(n9023), .B2(n6514), .C1(
        n6509), .C2(n9013), .ZN(P2_U3294) );
  OAI222_X1 U8154 ( .A1(P2_U3151), .A2(n6807), .B1(n9023), .B2(n6512), .C1(
        n6510), .C2(n9013), .ZN(P2_U3292) );
  OAI222_X1 U8155 ( .A1(P2_U3151), .A2(n6789), .B1(n9023), .B2(n6513), .C1(
        n5192), .C2(n9013), .ZN(P2_U3293) );
  NAND2_X2 U8156 ( .A1(n6511), .A2(P1_U3086), .ZN(n9971) );
  INV_X1 U8157 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10483) );
  INV_X1 U8158 ( .A(n6559), .ZN(n6576) );
  OAI222_X1 U8159 ( .A1(n9971), .A2(n10483), .B1(n9964), .B2(n6512), .C1(n6576), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U8160 ( .A1(n9971), .A2(n4966), .B1(n9964), .B2(n6513), .C1(n6664), 
        .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U8161 ( .A1(n4919), .A2(P2_U3151), .B1(n9013), .B2(n5236), .C1(
        n6516), .C2(n9023), .ZN(P2_U3291) );
  OAI222_X1 U8162 ( .A1(n9964), .A2(n6514), .B1(n9971), .B2(n5167), .C1(
        P1_U3086), .C2(n6544), .ZN(P1_U3354) );
  OAI222_X1 U8163 ( .A1(n6847), .A2(P2_U3151), .B1(n9023), .B2(n6521), .C1(
        n6515), .C2(n9013), .ZN(P2_U3290) );
  INV_X1 U8164 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6517) );
  INV_X1 U8165 ( .A(n10003), .ZN(n10012) );
  OAI222_X1 U8166 ( .A1(n9971), .A2(n6517), .B1(n9964), .B2(n6516), .C1(n10012), .C2(P1_U3086), .ZN(P1_U3351) );
  OAI222_X1 U8167 ( .A1(P2_U3151), .A2(n4904), .B1(n9023), .B2(n6519), .C1(
        n6518), .C2(n9013), .ZN(P2_U3289) );
  INV_X1 U8168 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6520) );
  OAI222_X1 U8169 ( .A1(n9971), .A2(n6520), .B1(n9964), .B2(n6519), .C1(n6611), 
        .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U8170 ( .A(n6587), .ZN(n6596) );
  INV_X1 U8171 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6670) );
  OAI222_X1 U8172 ( .A1(P1_U3086), .A2(n6596), .B1(n9964), .B2(n6521), .C1(
        n9971), .C2(n6670), .ZN(P1_U3350) );
  AOI21_X1 U8173 ( .B1(n6523), .B2(n9282), .A(n6522), .ZN(n6539) );
  INV_X1 U8174 ( .A(n6539), .ZN(n6524) );
  NAND2_X1 U8175 ( .A1(n9219), .A2(n9466), .ZN(n6538) );
  AND2_X1 U8176 ( .A1(n6524), .A2(n6538), .ZN(n10030) );
  NOR2_X1 U8177 ( .A1(n10030), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8178 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10472) );
  INV_X1 U8179 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6527) );
  INV_X1 U8180 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8027) );
  OR2_X1 U8181 ( .A1(n5975), .A2(n8027), .ZN(n6526) );
  INV_X1 U8182 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9896) );
  OR2_X1 U8183 ( .A1(n6086), .A2(n9896), .ZN(n6525) );
  OAI211_X1 U8184 ( .C1(n9224), .C2(n6527), .A(n6526), .B(n6525), .ZN(n9280)
         );
  NAND2_X1 U8185 ( .A1(n9280), .A2(P1_U3973), .ZN(n6528) );
  OAI21_X1 U8186 ( .B1(P1_U3973), .B2(n10472), .A(n6528), .ZN(P1_U3585) );
  NAND2_X1 U8187 ( .A1(n6529), .A2(P1_U3973), .ZN(n6530) );
  OAI21_X1 U8188 ( .B1(P1_U3973), .B2(n5236), .A(n6530), .ZN(P1_U3558) );
  INV_X1 U8189 ( .A(n7197), .ZN(n7247) );
  INV_X1 U8190 ( .A(n6531), .ZN(n6533) );
  INV_X1 U8191 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6532) );
  OAI222_X1 U8192 ( .A1(n7247), .A2(P2_U3151), .B1(n9023), .B2(n6533), .C1(
        n6532), .C2(n9013), .ZN(P2_U3288) );
  INV_X1 U8193 ( .A(n6631), .ZN(n6618) );
  INV_X1 U8194 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6668) );
  OAI222_X1 U8195 ( .A1(P1_U3086), .A2(n6618), .B1(n9964), .B2(n6533), .C1(
        n9971), .C2(n6668), .ZN(P1_U3348) );
  INV_X1 U8196 ( .A(n7390), .ZN(n7386) );
  INV_X1 U8197 ( .A(n6534), .ZN(n6536) );
  INV_X1 U8198 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6535) );
  OAI222_X1 U8199 ( .A1(n7386), .A2(P2_U3151), .B1(n9023), .B2(n6536), .C1(
        n6535), .C2(n9013), .ZN(P2_U3287) );
  INV_X1 U8200 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6537) );
  INV_X1 U8201 ( .A(n6630), .ZN(n9984) );
  OAI222_X1 U8202 ( .A1(n9971), .A2(n6537), .B1(n9964), .B2(n6536), .C1(
        P1_U3086), .C2(n9984), .ZN(P1_U3347) );
  NAND2_X1 U8203 ( .A1(n6539), .A2(n6538), .ZN(n9996) );
  OR3_X1 U8204 ( .A1(n9996), .A2(n6541), .A3(n6443), .ZN(n9494) );
  XNOR2_X1 U8205 ( .A(n6544), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6554) );
  INV_X1 U8206 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6697) );
  AND2_X1 U8207 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6649) );
  XNOR2_X1 U8208 ( .A(n6554), .B(n6649), .ZN(n6551) );
  INV_X1 U8209 ( .A(n6544), .ZN(n6555) );
  INV_X1 U8210 ( .A(n10027), .ZN(n10041) );
  INV_X1 U8211 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6542) );
  INV_X1 U8212 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6966) );
  OAI22_X1 U8213 ( .A1(n10048), .A2(n6542), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6966), .ZN(n6543) );
  AOI21_X1 U8214 ( .B1(n6555), .B2(n10041), .A(n6543), .ZN(n6550) );
  INV_X1 U8215 ( .A(n6541), .ZN(n6648) );
  OR2_X1 U8216 ( .A1(n9996), .A2(n6648), .ZN(n9493) );
  INV_X1 U8217 ( .A(n9493), .ZN(n10043) );
  MUX2_X1 U8218 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n5911), .S(n6544), .Z(n6546)
         );
  OR3_X1 U8219 ( .A1(n6546), .A2(n6545), .A3(n6547), .ZN(n6657) );
  OAI21_X1 U8220 ( .B1(n6545), .B2(n6547), .A(n6546), .ZN(n6548) );
  NAND3_X1 U8221 ( .A1(n10043), .A2(n6657), .A3(n6548), .ZN(n6549) );
  OAI211_X1 U8222 ( .C1(n9494), .C2(n6551), .A(n6550), .B(n6549), .ZN(P1_U3244) );
  INV_X1 U8223 ( .A(n6664), .ZN(n6558) );
  NAND2_X1 U8224 ( .A1(n6555), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6656) );
  MUX2_X1 U8225 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n5924), .S(n6664), .Z(n6655)
         );
  AOI21_X1 U8226 ( .B1(n6657), .B2(n6656), .A(n6655), .ZN(n6659) );
  AOI21_X1 U8227 ( .B1(n6558), .B2(P1_REG1_REG_2__SCAN_IN), .A(n6659), .ZN(
        n6553) );
  MUX2_X1 U8228 ( .A(n6566), .B(P1_REG1_REG_3__SCAN_IN), .S(n6559), .Z(n6552)
         );
  NOR2_X1 U8229 ( .A1(n6553), .A2(n6552), .ZN(n10002) );
  AOI211_X1 U8230 ( .C1(n6553), .C2(n6552), .A(n10002), .B(n9493), .ZN(n6563)
         );
  XNOR2_X1 U8231 ( .A(n6664), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U8232 ( .A1(n6554), .A2(n6649), .ZN(n6557) );
  NAND2_X1 U8233 ( .A1(n6555), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U8234 ( .A1(n6557), .A2(n6556), .ZN(n6653) );
  AOI22_X1 U8235 ( .A1(n6654), .A2(n6653), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n6558), .ZN(n6561) );
  INV_X1 U8236 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10057) );
  MUX2_X1 U8237 ( .A(n10057), .B(P1_REG2_REG_3__SCAN_IN), .S(n6559), .Z(n6560)
         );
  NOR2_X1 U8238 ( .A1(n6561), .A2(n6560), .ZN(n10009) );
  AOI211_X1 U8239 ( .C1(n6561), .C2(n6560), .A(n10009), .B(n9494), .ZN(n6562)
         );
  NOR2_X1 U8240 ( .A1(n6563), .A2(n6562), .ZN(n6565) );
  NOR2_X1 U8241 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5954), .ZN(n6720) );
  AOI21_X1 U8242 ( .B1(n10030), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6720), .ZN(
        n6564) );
  OAI211_X1 U8243 ( .C1(n6576), .C2(n10027), .A(n6565), .B(n6564), .ZN(
        P1_U3246) );
  NAND2_X1 U8244 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7023) );
  NOR2_X1 U8245 ( .A1(n6576), .A2(n6566), .ZN(n9997) );
  INV_X1 U8246 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6567) );
  MUX2_X1 U8247 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6567), .S(n10003), .Z(n6568)
         );
  OAI21_X1 U8248 ( .B1(n10002), .B2(n9997), .A(n6568), .ZN(n10000) );
  INV_X1 U8249 ( .A(n10000), .ZN(n6569) );
  AOI21_X1 U8250 ( .B1(n10003), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6569), .ZN(
        n6572) );
  INV_X1 U8251 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6570) );
  MUX2_X1 U8252 ( .A(n6570), .B(P1_REG1_REG_5__SCAN_IN), .S(n6587), .Z(n6571)
         );
  NOR2_X1 U8253 ( .A1(n6572), .A2(n6571), .ZN(n6589) );
  AOI211_X1 U8254 ( .C1(n6572), .C2(n6571), .A(n6589), .B(n9493), .ZN(n6573)
         );
  INV_X1 U8255 ( .A(n6573), .ZN(n6574) );
  NAND2_X1 U8256 ( .A1(n7023), .A2(n6574), .ZN(n6575) );
  AOI21_X1 U8257 ( .B1(n10030), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6575), .ZN(
        n6586) );
  NOR2_X1 U8258 ( .A1(n6576), .A2(n10057), .ZN(n10004) );
  INV_X1 U8259 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6577) );
  MUX2_X1 U8260 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6577), .S(n10003), .Z(n6578)
         );
  OAI21_X1 U8261 ( .B1(n10009), .B2(n10004), .A(n6578), .ZN(n10007) );
  INV_X1 U8262 ( .A(n10007), .ZN(n6580) );
  NOR2_X1 U8263 ( .A1(n10012), .A2(n6577), .ZN(n6581) );
  INV_X1 U8264 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7087) );
  MUX2_X1 U8265 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7087), .S(n6587), .Z(n6579)
         );
  OAI21_X1 U8266 ( .B1(n6580), .B2(n6581), .A(n6579), .ZN(n6595) );
  INV_X1 U8267 ( .A(n6581), .ZN(n6583) );
  MUX2_X1 U8268 ( .A(n7087), .B(P1_REG2_REG_5__SCAN_IN), .S(n6587), .Z(n6582)
         );
  NAND3_X1 U8269 ( .A1(n10007), .A2(n6583), .A3(n6582), .ZN(n6584) );
  NAND3_X1 U8270 ( .A1(n10039), .A2(n6595), .A3(n6584), .ZN(n6585) );
  OAI211_X1 U8271 ( .C1(n10027), .C2(n6596), .A(n6586), .B(n6585), .ZN(
        P1_U3248) );
  AND2_X1 U8272 ( .A1(n6587), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6590) );
  MUX2_X1 U8273 ( .A(n10123), .B(P1_REG1_REG_6__SCAN_IN), .S(n6611), .Z(n6588)
         );
  OAI21_X1 U8274 ( .B1(n6589), .B2(n6590), .A(n6588), .ZN(n6610) );
  INV_X1 U8275 ( .A(n6589), .ZN(n6593) );
  INV_X1 U8276 ( .A(n6590), .ZN(n6592) );
  INV_X1 U8277 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10123) );
  MUX2_X1 U8278 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10123), .S(n6611), .Z(n6591)
         );
  NAND3_X1 U8279 ( .A1(n6593), .A2(n6592), .A3(n6591), .ZN(n6594) );
  NAND3_X1 U8280 ( .A1(n6610), .A2(n10043), .A3(n6594), .ZN(n6604) );
  NAND2_X1 U8281 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n7072) );
  OAI21_X1 U8282 ( .B1(n7087), .B2(n6596), .A(n6595), .ZN(n6600) );
  INV_X1 U8283 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6598) );
  MUX2_X1 U8284 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6598), .S(n6597), .Z(n6599)
         );
  NAND2_X1 U8285 ( .A1(n6600), .A2(n6599), .ZN(n6605) );
  OAI211_X1 U8286 ( .C1(n6600), .C2(n6599), .A(n10039), .B(n6605), .ZN(n6601)
         );
  NAND2_X1 U8287 ( .A1(n7072), .A2(n6601), .ZN(n6602) );
  AOI21_X1 U8288 ( .B1(n10030), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6602), .ZN(
        n6603) );
  OAI211_X1 U8289 ( .C1(n10027), .C2(n6611), .A(n6604), .B(n6603), .ZN(
        P1_U3249) );
  OAI21_X1 U8290 ( .B1(n6598), .B2(n6611), .A(n6605), .ZN(n6608) );
  INV_X1 U8291 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6606) );
  AOI22_X1 U8292 ( .A1(n6631), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6606), .B2(
        n6618), .ZN(n6607) );
  NAND2_X1 U8293 ( .A1(n6607), .A2(n6608), .ZN(n6632) );
  OAI211_X1 U8294 ( .C1(n6608), .C2(n6607), .A(n10039), .B(n6632), .ZN(n6617)
         );
  NAND2_X1 U8295 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7136) );
  MUX2_X1 U8296 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6609), .S(n6631), .Z(n6613)
         );
  OAI21_X1 U8297 ( .B1(n10123), .B2(n6611), .A(n6610), .ZN(n6612) );
  NAND2_X1 U8298 ( .A1(n6613), .A2(n6612), .ZN(n6626) );
  OAI211_X1 U8299 ( .C1(n6613), .C2(n6612), .A(n10043), .B(n6626), .ZN(n6614)
         );
  NAND2_X1 U8300 ( .A1(n7136), .A2(n6614), .ZN(n6615) );
  AOI21_X1 U8301 ( .B1(n10030), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6615), .ZN(
        n6616) );
  OAI211_X1 U8302 ( .C1(n10027), .C2(n6618), .A(n6617), .B(n6616), .ZN(
        P1_U3250) );
  INV_X1 U8303 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6619) );
  OAI222_X1 U8304 ( .A1(n9971), .A2(n6619), .B1(n9964), .B2(n6621), .C1(n6874), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8305 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6620) );
  OAI222_X1 U8306 ( .A1(P2_U3151), .A2(n7821), .B1(n9023), .B2(n6621), .C1(
        n6620), .C2(n9013), .ZN(P2_U3285) );
  INV_X1 U8307 ( .A(n6622), .ZN(n6623) );
  OAI222_X1 U8308 ( .A1(P2_U3151), .A2(n7535), .B1(n9023), .B2(n6623), .C1(
        n10469), .C2(n9013), .ZN(P2_U3286) );
  INV_X1 U8309 ( .A(n6699), .ZN(n6708) );
  OAI222_X1 U8310 ( .A1(n9971), .A2(n6624), .B1(n9964), .B2(n6623), .C1(n6708), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  AOI22_X1 U8311 ( .A1(n6699), .A2(n6068), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6708), .ZN(n6629) );
  MUX2_X1 U8312 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6625), .S(n6630), .Z(n9977)
         );
  NAND2_X1 U8313 ( .A1(n6631), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U8314 ( .A1(n6627), .A2(n6626), .ZN(n9978) );
  NAND2_X1 U8315 ( .A1(n9977), .A2(n9978), .ZN(n9976) );
  OAI21_X1 U8316 ( .B1(n6625), .B2(n9984), .A(n9976), .ZN(n6628) );
  NOR2_X1 U8317 ( .A1(n6629), .A2(n6628), .ZN(n6700) );
  AOI21_X1 U8318 ( .B1(n6629), .B2(n6628), .A(n6700), .ZN(n6643) );
  INV_X1 U8319 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U8320 ( .A1(n6699), .A2(n10344), .B1(P1_REG2_REG_9__SCAN_IN), .B2(
        n6708), .ZN(n6636) );
  INV_X1 U8321 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6634) );
  AOI22_X1 U8322 ( .A1(n6630), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6634), .B2(
        n9984), .ZN(n9980) );
  NAND2_X1 U8323 ( .A1(n6631), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U8324 ( .A1(n6633), .A2(n6632), .ZN(n9981) );
  NAND2_X1 U8325 ( .A1(n9980), .A2(n9981), .ZN(n9979) );
  OAI21_X1 U8326 ( .B1(n6634), .B2(n9984), .A(n9979), .ZN(n6635) );
  NOR2_X1 U8327 ( .A1(n6636), .A2(n6635), .ZN(n6707) );
  AOI21_X1 U8328 ( .B1(n6636), .B2(n6635), .A(n6707), .ZN(n6637) );
  OR2_X1 U8329 ( .A1(n6637), .A2(n9494), .ZN(n6640) );
  NOR2_X1 U8330 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6638), .ZN(n7607) );
  AOI21_X1 U8331 ( .B1(n10030), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7607), .ZN(
        n6639) );
  OAI211_X1 U8332 ( .C1(n10027), .C2(n6708), .A(n6640), .B(n6639), .ZN(n6641)
         );
  INV_X1 U8333 ( .A(n6641), .ZN(n6642) );
  OAI21_X1 U8334 ( .B1(n6643), .B2(n9493), .A(n6642), .ZN(P1_U3252) );
  INV_X1 U8335 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10372) );
  NOR2_X1 U8336 ( .A1(n6724), .A2(n10372), .ZN(P2_U3240) );
  INV_X1 U8337 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10300) );
  NOR2_X1 U8338 ( .A1(n6724), .A2(n10300), .ZN(P2_U3245) );
  INV_X1 U8339 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6644) );
  NOR2_X1 U8340 ( .A1(n6724), .A2(n6644), .ZN(P2_U3235) );
  INV_X1 U8341 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10486) );
  NOR2_X1 U8342 ( .A1(n6724), .A2(n10486), .ZN(P2_U3236) );
  INV_X1 U8343 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10396) );
  NOR2_X1 U8344 ( .A1(n6724), .A2(n10396), .ZN(P2_U3254) );
  INV_X1 U8345 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10347) );
  NOR2_X1 U8346 ( .A1(n6724), .A2(n10347), .ZN(P2_U3262) );
  OAI21_X1 U8347 ( .B1(n6647), .B2(n6646), .A(n6645), .ZN(n6675) );
  MUX2_X1 U8348 ( .A(n6675), .B(n6649), .S(n6648), .Z(n6652) );
  OR2_X1 U8349 ( .A1(n6541), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6650) );
  AND2_X1 U8350 ( .A1(n6651), .A2(n6650), .ZN(n9989) );
  NOR2_X1 U8351 ( .A1(n9989), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9988) );
  AOI211_X1 U8352 ( .C1(n6652), .C2(n6651), .A(n9988), .B(n9484), .ZN(n10014)
         );
  XOR2_X1 U8353 ( .A(n6654), .B(n6653), .Z(n6661) );
  AND3_X1 U8354 ( .A1(n6657), .A2(n6656), .A3(n6655), .ZN(n6658) );
  NOR3_X1 U8355 ( .A1(n9493), .A2(n6659), .A3(n6658), .ZN(n6660) );
  AOI21_X1 U8356 ( .B1(n10039), .B2(n6661), .A(n6660), .ZN(n6663) );
  AOI22_X1 U8357 ( .A1(n10030), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6662) );
  OAI211_X1 U8358 ( .C1(n6664), .C2(n10027), .A(n6663), .B(n6662), .ZN(n6665)
         );
  OR2_X1 U8359 ( .A1(n10014), .A2(n6665), .ZN(P1_U3245) );
  NAND2_X1 U8360 ( .A1(n9287), .A2(P1_U3973), .ZN(n6666) );
  OAI21_X1 U8361 ( .B1(n5563), .B2(P1_U3973), .A(n6666), .ZN(P1_U3574) );
  NAND2_X1 U8362 ( .A1(P2_U3893), .A2(n7649), .ZN(n6667) );
  OAI21_X1 U8363 ( .B1(P2_U3893), .B2(n6668), .A(n6667), .ZN(P2_U3498) );
  NAND2_X1 U8364 ( .A1(P2_U3893), .A2(n7443), .ZN(n6669) );
  OAI21_X1 U8365 ( .B1(P2_U3893), .B2(n6670), .A(n6669), .ZN(P2_U3496) );
  OR2_X1 U8366 ( .A1(n6671), .A2(n9219), .ZN(n9058) );
  NAND2_X1 U8367 ( .A1(n9142), .A2(n6741), .ZN(n6673) );
  OAI211_X1 U8368 ( .C1(n6675), .C2(n9145), .A(n6674), .B(n6673), .ZN(P1_U3232) );
  XOR2_X1 U8369 ( .A(n6678), .B(n6677), .Z(n6681) );
  AOI22_X1 U8370 ( .A1(n9142), .A2(n7204), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9058), .ZN(n6679) );
  OAI211_X1 U8371 ( .C1(n6681), .C2(n9145), .A(n6680), .B(n6679), .ZN(P1_U3237) );
  INV_X1 U8372 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6683) );
  INV_X1 U8373 ( .A(n6682), .ZN(n6685) );
  INV_X1 U8374 ( .A(n6872), .ZN(n10026) );
  OAI222_X1 U8375 ( .A1(n9971), .A2(n6683), .B1(n9964), .B2(n6685), .C1(
        P1_U3086), .C2(n10026), .ZN(P1_U3344) );
  INV_X1 U8376 ( .A(n7823), .ZN(n7910) );
  INV_X1 U8377 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6684) );
  OAI222_X1 U8378 ( .A1(n7910), .A2(P2_U3151), .B1(n9023), .B2(n6685), .C1(
        n6684), .C2(n9013), .ZN(P2_U3284) );
  INV_X1 U8379 ( .A(n6686), .ZN(n6688) );
  NAND2_X1 U8380 ( .A1(n9950), .A2(n6687), .ZN(n6758) );
  INV_X1 U8381 ( .A(n6758), .ZN(n6761) );
  NAND3_X1 U8382 ( .A1(n6688), .A2(n6761), .A3(n6762), .ZN(n6962) );
  NOR2_X1 U8383 ( .A1(n6689), .A2(n6963), .ZN(n6954) );
  INV_X1 U8384 ( .A(n6954), .ZN(n6690) );
  NAND2_X1 U8385 ( .A1(n6689), .A2(n6963), .ZN(n9245) );
  AND2_X1 U8386 ( .A1(n6690), .A2(n9245), .ZN(n10067) );
  INV_X1 U8387 ( .A(n9459), .ZN(n6739) );
  NAND2_X1 U8388 ( .A1(n9282), .A2(n6739), .ZN(n6738) );
  INV_X1 U8389 ( .A(n6738), .ZN(n6691) );
  NOR3_X1 U8390 ( .A1(n10067), .A2(n6434), .A3(n6691), .ZN(n6695) );
  INV_X1 U8391 ( .A(n6434), .ZN(n6737) );
  NOR2_X1 U8392 ( .A1(n6737), .A2(n6963), .ZN(n10071) );
  AND2_X1 U8393 ( .A1(n6264), .A2(n6437), .ZN(n9456) );
  INV_X1 U8394 ( .A(n9456), .ZN(n6692) );
  NAND2_X1 U8395 ( .A1(n10071), .A2(n6692), .ZN(n6693) );
  OAI211_X1 U8396 ( .C1(n9557), .C2(n5051), .A(n10069), .B(n6693), .ZN(n6694)
         );
  OAI21_X1 U8397 ( .B1(n6695), .B2(n6694), .A(n10056), .ZN(n6696) );
  OAI21_X1 U8398 ( .B1(n6697), .B2(n10056), .A(n6696), .ZN(P1_U3293) );
  AND2_X1 U8399 ( .A1(n6698), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8400 ( .A1(n6698), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8401 ( .A1(n6698), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8402 ( .A1(n6698), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8403 ( .A1(n6698), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8404 ( .A1(n6698), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8405 ( .A1(n6698), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8406 ( .A1(n6698), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8407 ( .A1(n6698), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8408 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7805) );
  INV_X1 U8409 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7677) );
  NOR2_X1 U8410 ( .A1(n6699), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6701) );
  NOR2_X1 U8411 ( .A1(n6701), .A2(n6700), .ZN(n6704) );
  MUX2_X1 U8412 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6702), .S(n6709), .Z(n6703)
         );
  NAND2_X1 U8413 ( .A1(n6703), .A2(n6704), .ZN(n6866) );
  OAI211_X1 U8414 ( .C1(n6704), .C2(n6703), .A(n6866), .B(n10043), .ZN(n6705)
         );
  OAI21_X1 U8415 ( .B1(n10048), .B2(n7677), .A(n6705), .ZN(n6706) );
  NOR2_X1 U8416 ( .A1(n7805), .A2(n6706), .ZN(n6713) );
  AOI21_X1 U8417 ( .B1(n6708), .B2(n10344), .A(n6707), .ZN(n6711) );
  INV_X1 U8418 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6875) );
  AOI22_X1 U8419 ( .A1(n6709), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n6875), .B2(
        n6874), .ZN(n6710) );
  NAND2_X1 U8420 ( .A1(n6710), .A2(n6711), .ZN(n6873) );
  OAI211_X1 U8421 ( .C1(n6711), .C2(n6710), .A(n10039), .B(n6873), .ZN(n6712)
         );
  OAI211_X1 U8422 ( .C1(n10027), .C2(n6874), .A(n6713), .B(n6712), .ZN(
        P1_U3253) );
  INV_X1 U8423 ( .A(n6714), .ZN(n6734) );
  AOI22_X1 U8424 ( .A1(n8578), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n9021), .ZN(n6715) );
  OAI21_X1 U8425 ( .B1(n6734), .B2(n9023), .A(n6715), .ZN(P2_U3282) );
  XOR2_X1 U8426 ( .A(n6718), .B(n6717), .Z(n6723) );
  INV_X1 U8427 ( .A(n10049), .ZN(n6993) );
  INV_X1 U8428 ( .A(n9483), .ZN(n6855) );
  OAI22_X1 U8429 ( .A1(n9218), .A2(n6993), .B1(n6855), .B2(n9189), .ZN(n6719)
         );
  AOI211_X1 U8430 ( .C1(n9186), .C2(n6529), .A(n6720), .B(n6719), .ZN(n6722)
         );
  NAND2_X1 U8431 ( .A1(n9210), .A2(n5954), .ZN(n6721) );
  OAI211_X1 U8432 ( .C1(n6723), .C2(n9145), .A(n6722), .B(n6721), .ZN(P1_U3218) );
  INV_X1 U8433 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6728) );
  NOR3_X1 U8434 ( .A1(n5808), .A2(n6726), .A3(n6725), .ZN(n6727) );
  AOI21_X1 U8435 ( .B1(n6698), .B2(n6728), .A(n6727), .ZN(P2_U3377) );
  INV_X1 U8436 ( .A(n6729), .ZN(n6731) );
  INV_X1 U8437 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6730) );
  OAI222_X1 U8438 ( .A1(n8551), .A2(P2_U3151), .B1(n9023), .B2(n6731), .C1(
        n6730), .C2(n9013), .ZN(P2_U3283) );
  INV_X1 U8439 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6732) );
  INV_X1 U8440 ( .A(n6871), .ZN(n6899) );
  OAI222_X1 U8441 ( .A1(n9971), .A2(n6732), .B1(n9964), .B2(n6731), .C1(
        P1_U3086), .C2(n6899), .ZN(P1_U3343) );
  AOI22_X1 U8442 ( .A1(n6698), .A2(n5813), .B1(n6733), .B2(n5115), .ZN(
        P2_U3376) );
  INV_X1 U8443 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6735) );
  INV_X1 U8444 ( .A(n7037), .ZN(n7033) );
  OAI222_X1 U8445 ( .A1(n9971), .A2(n6735), .B1(n9964), .B2(n6734), .C1(
        P1_U3086), .C2(n7033), .ZN(P1_U3342) );
  AND2_X1 U8446 ( .A1(n6698), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8447 ( .A1(n6698), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8448 ( .A1(n6698), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8449 ( .A1(n6698), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8450 ( .A1(n6698), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8451 ( .A1(n6698), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8452 ( .A1(n6698), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8453 ( .A1(n6698), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8454 ( .A1(n6698), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8455 ( .A1(n6698), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8456 ( .A1(n6698), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8457 ( .A1(n6698), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8458 ( .A1(n6698), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8459 ( .A1(n6698), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8460 ( .A1(n6698), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8461 ( .A1(n9465), .A2(n6736), .ZN(n6740) );
  OAI211_X1 U8462 ( .C1(n6740), .C2(n6739), .A(n6738), .B(n6737), .ZN(n7083)
         );
  INV_X1 U8463 ( .A(n9465), .ZN(n9454) );
  NAND2_X1 U8464 ( .A1(n9454), .A2(n6264), .ZN(n9463) );
  OR2_X1 U8465 ( .A1(n9463), .A2(n5890), .ZN(n10077) );
  INV_X1 U8466 ( .A(n6748), .ZN(n6742) );
  NAND2_X1 U8467 ( .A1(n6689), .A2(n6741), .ZN(n6947) );
  NAND2_X1 U8468 ( .A1(n6742), .A2(n6947), .ZN(n6950) );
  NAND2_X1 U8469 ( .A1(n6752), .A2(n9242), .ZN(n6743) );
  NAND2_X1 U8470 ( .A1(n6950), .A2(n6743), .ZN(n6744) );
  XNOR2_X1 U8471 ( .A(n9483), .B(n7204), .ZN(n9290) );
  INV_X1 U8472 ( .A(n9290), .ZN(n6750) );
  NAND2_X1 U8473 ( .A1(n6744), .A2(n6750), .ZN(n6849) );
  OAI21_X1 U8474 ( .B1(n6744), .B2(n6750), .A(n6849), .ZN(n7205) );
  OR2_X1 U8475 ( .A1(n6965), .A2(n6853), .ZN(n6745) );
  AND3_X1 U8476 ( .A1(n6851), .A2(n6745), .A3(n9739), .ZN(n7203) );
  INV_X1 U8477 ( .A(n9482), .ZN(n6994) );
  NAND2_X1 U8478 ( .A1(n9465), .A2(n6264), .ZN(n6747) );
  NAND2_X1 U8479 ( .A1(n9453), .A2(n5890), .ZN(n6746) );
  NAND2_X1 U8480 ( .A1(n6748), .A2(n6954), .ZN(n6953) );
  NAND2_X1 U8481 ( .A1(n6752), .A2(n10074), .ZN(n6749) );
  NAND2_X1 U8482 ( .A1(n6953), .A2(n6749), .ZN(n6854) );
  XNOR2_X1 U8483 ( .A(n6854), .B(n6750), .ZN(n6751) );
  OAI222_X1 U8484 ( .A1(n9877), .A2(n6752), .B1(n9879), .B2(n6994), .C1(n10068), .C2(n6751), .ZN(n7201) );
  AOI211_X1 U8485 ( .C1(n10100), .C2(n7205), .A(n7203), .B(n7201), .ZN(n6766)
         );
  OAI21_X1 U8486 ( .B1(n9951), .B2(P1_D_REG_1__SCAN_IN), .A(n9952), .ZN(n6757)
         );
  INV_X1 U8487 ( .A(n9951), .ZN(n6754) );
  NAND2_X1 U8488 ( .A1(n6754), .A2(n6753), .ZN(n6755) );
  NOR2_X1 U8489 ( .A1(n6762), .A2(n6758), .ZN(n6759) );
  AOI22_X1 U8490 ( .A1(n9819), .A2(n7204), .B1(n10126), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6760) );
  OAI21_X1 U8491 ( .B1(n6766), .B2(n10126), .A(n6760), .ZN(P1_U3524) );
  INV_X1 U8492 ( .A(n9948), .ZN(n9936) );
  AOI22_X1 U8493 ( .A1(n9936), .A2(n7204), .B1(n10117), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n6765) );
  OAI21_X1 U8494 ( .B1(n6766), .B2(n10117), .A(n6765), .ZN(P1_U3459) );
  INV_X1 U8495 ( .A(n6767), .ZN(n6775) );
  AOI22_X1 U8496 ( .A1(n7576), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n6768), .ZN(n6769) );
  OAI21_X1 U8497 ( .B1(n6775), .B2(n9964), .A(n6769), .ZN(P1_U3340) );
  INV_X1 U8498 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6771) );
  INV_X1 U8499 ( .A(n6770), .ZN(n6773) );
  OAI222_X1 U8500 ( .A1(n9971), .A2(n6771), .B1(n9964), .B2(n6773), .C1(
        P1_U3086), .C2(n7374), .ZN(P1_U3341) );
  INV_X1 U8501 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6772) );
  OAI222_X1 U8502 ( .A1(n8597), .A2(P2_U3151), .B1(n9023), .B2(n6773), .C1(
        n6772), .C2(n9013), .ZN(P2_U3281) );
  INV_X1 U8503 ( .A(n8625), .ZN(n8614) );
  INV_X1 U8504 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6774) );
  OAI222_X1 U8505 ( .A1(n8614), .A2(P2_U3151), .B1(n9023), .B2(n6775), .C1(
        n6774), .C2(n9013), .ZN(P2_U3280) );
  NOR2_X1 U8506 ( .A1(n8670), .A2(P2_U3151), .ZN(n9020) );
  NAND2_X1 U8507 ( .A1(n6786), .A2(n9020), .ZN(n6776) );
  MUX2_X1 U8508 ( .A(n8679), .B(n6776), .S(n6785), .Z(n8706) );
  INV_X1 U8509 ( .A(n6923), .ZN(n7812) );
  NOR2_X1 U8510 ( .A1(n6926), .A2(n7812), .ZN(n6777) );
  INV_X1 U8511 ( .A(n10141), .ZN(n8704) );
  INV_X1 U8512 ( .A(n6789), .ZN(n10144) );
  OAI21_X1 U8513 ( .B1(n10144), .B2(n6780), .A(n10130), .ZN(n6781) );
  NAND2_X1 U8514 ( .A1(n6781), .A2(n6807), .ZN(n6782) );
  OAI21_X1 U8515 ( .B1(n6781), .B2(n6807), .A(n6782), .ZN(n6818) );
  INV_X1 U8516 ( .A(n6782), .ZN(n6783) );
  MUX2_X1 U8517 ( .A(n6829), .B(P2_REG2_REG_4__SCAN_IN), .S(n6842), .Z(n6784)
         );
  OR3_X1 U8518 ( .A1(n6817), .A2(n6784), .A3(n6783), .ZN(n6787) );
  NOR2_X1 U8519 ( .A1(n6785), .A2(P2_U3151), .ZN(n9017) );
  AND2_X1 U8520 ( .A1(n6786), .A2(n9017), .ZN(n6796) );
  INV_X1 U8521 ( .A(n6796), .ZN(n8029) );
  AOI21_X1 U8522 ( .B1(n6828), .B2(n6787), .A(n10129), .ZN(n6801) );
  INV_X1 U8523 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7230) );
  OAI21_X1 U8524 ( .B1(n6789), .B2(n7230), .A(n6788), .ZN(n10147) );
  OAI21_X1 U8525 ( .B1(n8062), .B2(n6791), .A(n6792), .ZN(n8048) );
  OAI21_X1 U8526 ( .B1(n8048), .B2(n6802), .A(n6792), .ZN(n10146) );
  INV_X1 U8527 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7235) );
  INV_X1 U8528 ( .A(n6793), .ZN(n6794) );
  MUX2_X1 U8529 ( .A(n6833), .B(P2_REG1_REG_4__SCAN_IN), .S(n6842), .Z(n6795)
         );
  NOR3_X1 U8530 ( .A1(n6820), .A2(n6795), .A3(n6794), .ZN(n6797) );
  OAI21_X1 U8531 ( .B1(n6798), .B2(n6797), .A(n10149), .ZN(n6799) );
  NAND2_X1 U8532 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U8533 ( .A1(n6799), .A2(n7151), .ZN(n6800) );
  AOI211_X1 U8534 ( .C1(n8704), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6801), .B(
        n6800), .ZN(n6813) );
  MUX2_X1 U8535 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8670), .Z(n6808) );
  INV_X1 U8536 ( .A(n6808), .ZN(n6809) );
  MUX2_X1 U8537 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8670), .Z(n6805) );
  INV_X1 U8538 ( .A(n6805), .ZN(n6806) );
  INV_X1 U8539 ( .A(n8062), .ZN(n6804) );
  MUX2_X1 U8540 ( .A(n10439), .B(n6790), .S(n8670), .Z(n8030) );
  OAI21_X1 U8541 ( .B1(n6804), .B2(n6803), .A(n8049), .ZN(n10137) );
  XNOR2_X1 U8542 ( .A(n6805), .B(n10144), .ZN(n10138) );
  NAND2_X1 U8543 ( .A1(n10137), .A2(n10138), .ZN(n10135) );
  OAI21_X1 U8544 ( .B1(n10144), .B2(n6806), .A(n10135), .ZN(n6815) );
  XNOR2_X1 U8545 ( .A(n6808), .B(n6807), .ZN(n6816) );
  NOR2_X1 U8546 ( .A1(n6815), .A2(n6816), .ZN(n6814) );
  MUX2_X1 U8547 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8670), .Z(n6839) );
  XNOR2_X1 U8548 ( .A(n6839), .B(n6842), .ZN(n6810) );
  OAI211_X1 U8549 ( .C1(n6811), .C2(n6810), .A(n6840), .B(n10136), .ZN(n6812)
         );
  OAI211_X1 U8550 ( .C1(n8706), .C2(n4919), .A(n6813), .B(n6812), .ZN(P2_U3186) );
  AOI21_X1 U8551 ( .B1(n6816), .B2(n6815), .A(n6814), .ZN(n6827) );
  AOI21_X1 U8552 ( .B1(n5202), .B2(n6818), .A(n6817), .ZN(n6819) );
  NOR2_X1 U8553 ( .A1(n10129), .A2(n6819), .ZN(n6824) );
  AOI21_X1 U8554 ( .B1(n7235), .B2(n6821), .A(n6820), .ZN(n6822) );
  NAND2_X1 U8555 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8385) );
  OAI21_X1 U8556 ( .B1(n8666), .B2(n6822), .A(n8385), .ZN(n6823) );
  AOI211_X1 U8557 ( .C1(n8704), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6824), .B(
        n6823), .ZN(n6826) );
  NAND2_X1 U8558 ( .A1(n10143), .A2(n4671), .ZN(n6825) );
  OAI211_X1 U8559 ( .C1(n6827), .C2(n8703), .A(n6826), .B(n6825), .ZN(P2_U3185) );
  AOI21_X1 U8560 ( .B1(n7328), .B2(n6831), .A(n6979), .ZN(n6832) );
  NOR2_X1 U8561 ( .A1(n10129), .A2(n6832), .ZN(n6838) );
  AOI21_X1 U8562 ( .B1(n5248), .B2(n6835), .A(n4810), .ZN(n6836) );
  NAND2_X1 U8563 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7314) );
  OAI21_X1 U8564 ( .B1(n8666), .B2(n6836), .A(n7314), .ZN(n6837) );
  AOI211_X1 U8565 ( .C1(n8704), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6838), .B(
        n6837), .ZN(n6846) );
  INV_X1 U8566 ( .A(n6839), .ZN(n6841) );
  MUX2_X1 U8567 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8670), .Z(n6970) );
  XNOR2_X1 U8568 ( .A(n6970), .B(n6973), .ZN(n6843) );
  OAI211_X1 U8569 ( .C1(n6844), .C2(n6843), .A(n6971), .B(n10136), .ZN(n6845)
         );
  OAI211_X1 U8570 ( .C1(n8706), .C2(n6847), .A(n6846), .B(n6845), .ZN(P2_U3187) );
  NAND2_X1 U8571 ( .A1(n6855), .A2(n6853), .ZN(n6848) );
  NAND2_X1 U8572 ( .A1(n6849), .A2(n6848), .ZN(n6850) );
  AND2_X1 U8573 ( .A1(n6994), .A2(n10049), .ZN(n7000) );
  INV_X1 U8574 ( .A(n7000), .ZN(n9342) );
  NAND2_X1 U8575 ( .A1(n6993), .A2(n9482), .ZN(n9328) );
  NAND2_X1 U8576 ( .A1(n6850), .A2(n6857), .ZN(n6996) );
  OAI21_X1 U8577 ( .B1(n6850), .B2(n6857), .A(n6996), .ZN(n10060) );
  AOI21_X1 U8578 ( .B1(n6851), .B2(n10049), .A(n9750), .ZN(n6852) );
  OR2_X1 U8579 ( .A1(n6851), .A2(n10049), .ZN(n7161) );
  AND2_X1 U8580 ( .A1(n6852), .A2(n7161), .ZN(n10052) );
  NAND2_X1 U8581 ( .A1(n9483), .A2(n6853), .ZN(n9244) );
  NAND2_X1 U8582 ( .A1(n6855), .A2(n7204), .ZN(n6856) );
  INV_X1 U8583 ( .A(n6857), .ZN(n9291) );
  XNOR2_X1 U8584 ( .A(n9331), .B(n9291), .ZN(n6858) );
  AOI222_X1 U8585 ( .A1(n10116), .A2(n6858), .B1(n6529), .B2(n10105), .C1(
        n9483), .C2(n10104), .ZN(n10062) );
  INV_X1 U8586 ( .A(n10062), .ZN(n6859) );
  AOI211_X1 U8587 ( .C1(n10100), .C2(n10060), .A(n10052), .B(n6859), .ZN(n6864) );
  INV_X1 U8588 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6860) );
  OAI22_X1 U8589 ( .A1(n9948), .A2(n6993), .B1(n10119), .B2(n6860), .ZN(n6861)
         );
  INV_X1 U8590 ( .A(n6861), .ZN(n6862) );
  OAI21_X1 U8591 ( .B1(n6864), .B2(n10117), .A(n6862), .ZN(P1_U3462) );
  AOI22_X1 U8592 ( .A1(n9819), .A2(n10049), .B1(n10126), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n6863) );
  OAI21_X1 U8593 ( .B1(n6864), .B2(n10126), .A(n6863), .ZN(P1_U3525) );
  AOI22_X1 U8594 ( .A1(n7037), .A2(P1_REG1_REG_13__SCAN_IN), .B1(n6153), .B2(
        n7033), .ZN(n6868) );
  MUX2_X1 U8595 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6865), .S(n6872), .Z(n10022) );
  OAI21_X1 U8596 ( .B1(n6874), .B2(n6702), .A(n6866), .ZN(n10023) );
  NAND2_X1 U8597 ( .A1(n10022), .A2(n10023), .ZN(n10021) );
  OAI21_X1 U8598 ( .B1(n6865), .B2(n10026), .A(n10021), .ZN(n6895) );
  AOI22_X1 U8599 ( .A1(n6871), .A2(n6131), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n6899), .ZN(n6894) );
  NOR2_X1 U8600 ( .A1(n6895), .A2(n6894), .ZN(n6893) );
  AOI21_X1 U8601 ( .B1(n6899), .B2(n6131), .A(n6893), .ZN(n6867) );
  NAND2_X1 U8602 ( .A1(n6868), .A2(n6867), .ZN(n7032) );
  OAI21_X1 U8603 ( .B1(n6868), .B2(n6867), .A(n7032), .ZN(n6886) );
  INV_X1 U8604 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6869) );
  AOI22_X1 U8605 ( .A1(n7037), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n6869), .B2(
        n7033), .ZN(n6879) );
  NOR2_X1 U8606 ( .A1(n6871), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6877) );
  INV_X1 U8607 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6870) );
  AOI22_X1 U8608 ( .A1(n6871), .A2(n6870), .B1(P1_REG2_REG_12__SCAN_IN), .B2(
        n6899), .ZN(n6892) );
  INV_X1 U8609 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6876) );
  AOI22_X1 U8610 ( .A1(n6872), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n6876), .B2(
        n10026), .ZN(n10019) );
  OAI21_X1 U8611 ( .B1(n6875), .B2(n6874), .A(n6873), .ZN(n10020) );
  NAND2_X1 U8612 ( .A1(n10019), .A2(n10020), .ZN(n10018) );
  OAI21_X1 U8613 ( .B1(n6876), .B2(n10026), .A(n10018), .ZN(n6891) );
  NOR2_X1 U8614 ( .A1(n6892), .A2(n6891), .ZN(n6890) );
  NOR2_X1 U8615 ( .A1(n6877), .A2(n6890), .ZN(n6878) );
  NAND2_X1 U8616 ( .A1(n6879), .A2(n6878), .ZN(n7038) );
  OAI21_X1 U8617 ( .B1(n6879), .B2(n6878), .A(n7038), .ZN(n6883) );
  NOR2_X1 U8618 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6880), .ZN(n9152) );
  AOI21_X1 U8619 ( .B1(n10030), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9152), .ZN(
        n6882) );
  OR2_X1 U8620 ( .A1(n10027), .A2(n7033), .ZN(n6881) );
  OAI211_X1 U8621 ( .C1(n6883), .C2(n9494), .A(n6882), .B(n6881), .ZN(n6884)
         );
  INV_X1 U8622 ( .A(n6884), .ZN(n6885) );
  OAI21_X1 U8623 ( .B1(n6886), .B2(n9493), .A(n6885), .ZN(P1_U3256) );
  INV_X1 U8624 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6889) );
  INV_X1 U8625 ( .A(n7106), .ZN(n8541) );
  NAND2_X1 U8626 ( .A1(n8541), .A2(n8047), .ZN(n8192) );
  AND2_X1 U8627 ( .A1(n8193), .A2(n8192), .ZN(n8156) );
  INV_X1 U8628 ( .A(n8156), .ZN(n8044) );
  OAI21_X1 U8629 ( .B1(n8909), .B2(n8862), .A(n8044), .ZN(n6887) );
  OR2_X1 U8630 ( .A1(n5182), .A2(n7469), .ZN(n8036) );
  OAI211_X1 U8631 ( .C1(n8476), .C2(n8047), .A(n6887), .B(n8036), .ZN(n7030)
         );
  NAND2_X1 U8632 ( .A1(n10580), .A2(n7030), .ZN(n6888) );
  OAI21_X1 U8633 ( .B1(n10580), .B2(n6889), .A(n6888), .ZN(P2_U3390) );
  AOI21_X1 U8634 ( .B1(n6892), .B2(n6891), .A(n6890), .ZN(n6902) );
  AOI21_X1 U8635 ( .B1(n6895), .B2(n6894), .A(n6893), .ZN(n6896) );
  OR2_X1 U8636 ( .A1(n6896), .A2(n9493), .ZN(n6898) );
  AND2_X1 U8637 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9085) );
  AOI21_X1 U8638 ( .B1(n10030), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9085), .ZN(
        n6897) );
  OAI211_X1 U8639 ( .C1(n10027), .C2(n6899), .A(n6898), .B(n6897), .ZN(n6900)
         );
  INV_X1 U8640 ( .A(n6900), .ZN(n6901) );
  OAI21_X1 U8641 ( .B1(n6902), .B2(n9494), .A(n6901), .ZN(P1_U3255) );
  INV_X1 U8642 ( .A(n9481), .ZN(n7278) );
  INV_X1 U8643 ( .A(n10085), .ZN(n7162) );
  AOI22_X1 U8644 ( .A1(n9142), .A2(n7162), .B1(n9215), .B2(n9482), .ZN(n6903)
         );
  NAND2_X1 U8645 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10015) );
  OAI211_X1 U8646 ( .C1(n7278), .C2(n9209), .A(n6903), .B(n10015), .ZN(n6911)
         );
  INV_X1 U8647 ( .A(n6907), .ZN(n6908) );
  AOI211_X1 U8648 ( .C1(n6909), .C2(n6905), .A(n9145), .B(n6908), .ZN(n6910)
         );
  AOI211_X1 U8649 ( .C1(n7163), .C2(n9210), .A(n6911), .B(n6910), .ZN(n6912)
         );
  INV_X1 U8650 ( .A(n6912), .ZN(P1_U3230) );
  XNOR2_X1 U8651 ( .A(n7012), .B(n5183), .ZN(n7008) );
  XNOR2_X1 U8652 ( .A(n7008), .B(n8540), .ZN(n7010) );
  XOR2_X1 U8653 ( .A(n7010), .B(n7009), .Z(n6943) );
  INV_X1 U8654 ( .A(n6919), .ZN(n6917) );
  OAI21_X1 U8655 ( .B1(n6938), .B2(n6918), .A(n6917), .ZN(n6921) );
  NAND2_X1 U8656 ( .A1(n6933), .A2(n6919), .ZN(n6925) );
  AND2_X1 U8657 ( .A1(n6925), .A2(n7102), .ZN(n6920) );
  NAND2_X1 U8658 ( .A1(n6938), .A2(n6922), .ZN(n6928) );
  AND2_X1 U8659 ( .A1(n6924), .A2(n6923), .ZN(n6927) );
  NAND4_X1 U8660 ( .A1(n6928), .A2(n6927), .A3(n6926), .A4(n6925), .ZN(n6929)
         );
  NAND2_X1 U8661 ( .A1(n6929), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6931) );
  NAND2_X1 U8662 ( .A1(n6933), .A2(n8355), .ZN(n6930) );
  NAND2_X1 U8663 ( .A1(n8520), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8043) );
  INV_X1 U8664 ( .A(n8355), .ZN(n6932) );
  NOR2_X1 U8665 ( .A1(n6933), .A2(n6932), .ZN(n6936) );
  NAND2_X1 U8666 ( .A1(n6938), .A2(n6937), .ZN(n6939) );
  NOR2_X1 U8667 ( .A1(n5183), .A2(n8476), .ZN(n7176) );
  AOI22_X1 U8668 ( .A1(n8518), .A2(n8539), .B1(n8482), .B2(n7176), .ZN(n6940)
         );
  OAI21_X1 U8669 ( .B1(n7106), .B2(n8516), .A(n6940), .ZN(n6941) );
  AOI21_X1 U8670 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8043), .A(n6941), .ZN(
        n6942) );
  OAI21_X1 U8671 ( .B1(n6943), .B2(n8522), .A(n6942), .ZN(P2_U3162) );
  INV_X1 U8672 ( .A(n6944), .ZN(n6946) );
  OAI222_X1 U8673 ( .A1(P2_U3151), .A2(n8641), .B1(n9023), .B2(n6946), .C1(
        n6945), .C2(n9013), .ZN(P2_U3279) );
  INV_X1 U8674 ( .A(n7574), .ZN(n7710) );
  OAI222_X1 U8675 ( .A1(n9971), .A2(n10453), .B1(n9964), .B2(n6946), .C1(n7710), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U8676 ( .A(n6947), .ZN(n6948) );
  NAND2_X1 U8677 ( .A1(n6748), .A2(n6948), .ZN(n6949) );
  AND2_X1 U8678 ( .A1(n6950), .A2(n6949), .ZN(n10078) );
  NOR2_X1 U8679 ( .A1(n10078), .A2(n7082), .ZN(n6961) );
  INV_X1 U8680 ( .A(n10078), .ZN(n6952) );
  INV_X1 U8681 ( .A(n7083), .ZN(n6951) );
  NAND2_X1 U8682 ( .A1(n6952), .A2(n6951), .ZN(n6960) );
  OAI21_X1 U8683 ( .B1(n6954), .B2(n6748), .A(n6953), .ZN(n6958) );
  NAND2_X1 U8684 ( .A1(n9483), .A2(n10105), .ZN(n6956) );
  NAND2_X1 U8685 ( .A1(n6689), .A2(n10104), .ZN(n6955) );
  NAND2_X1 U8686 ( .A1(n6956), .A2(n6955), .ZN(n6957) );
  AOI21_X1 U8687 ( .B1(n6958), .B2(n10116), .A(n6957), .ZN(n6959) );
  NAND2_X1 U8688 ( .A1(n6960), .A2(n6959), .ZN(n10079) );
  OAI21_X1 U8689 ( .B1(n6961), .B2(n10079), .A(n10056), .ZN(n6969) );
  OAI21_X1 U8690 ( .B1(n9242), .B2(n6963), .A(n9739), .ZN(n6964) );
  OR2_X1 U8691 ( .A1(n6965), .A2(n6964), .ZN(n10076) );
  OAI22_X1 U8692 ( .A1(n9740), .A2(n10076), .B1(n6966), .B2(n9557), .ZN(n6967)
         );
  AOI21_X1 U8693 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n10063), .A(n6967), .ZN(
        n6968) );
  OAI211_X1 U8694 ( .C1(n9242), .C2(n9752), .A(n6969), .B(n6968), .ZN(P1_U3292) );
  MUX2_X1 U8695 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8670), .Z(n7179) );
  XNOR2_X1 U8696 ( .A(n7179), .B(n4904), .ZN(n6975) );
  INV_X1 U8697 ( .A(n6970), .ZN(n6972) );
  OAI21_X1 U8698 ( .B1(n6973), .B2(n6972), .A(n6971), .ZN(n6974) );
  NOR2_X1 U8699 ( .A1(n6974), .A2(n6975), .ZN(n7180) );
  AOI21_X1 U8700 ( .B1(n6975), .B2(n6974), .A(n7180), .ZN(n6992) );
  INV_X1 U8701 ( .A(n6976), .ZN(n6978) );
  XNOR2_X1 U8702 ( .A(n7184), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6977) );
  OR3_X1 U8703 ( .A1(n6979), .A2(n6978), .A3(n6977), .ZN(n6980) );
  AOI21_X1 U8704 ( .B1(n7182), .B2(n6980), .A(n10129), .ZN(n6981) );
  AOI21_X1 U8705 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(n8704), .A(n6981), .ZN(
        n6989) );
  INV_X1 U8706 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10473) );
  NOR2_X1 U8707 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10473), .ZN(n7414) );
  INV_X1 U8708 ( .A(n7414), .ZN(n6988) );
  INV_X1 U8709 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6982) );
  XNOR2_X1 U8710 ( .A(n7184), .B(n6982), .ZN(n6984) );
  AND3_X1 U8711 ( .A1(n6985), .A2(n6984), .A3(n6983), .ZN(n6986) );
  OAI21_X1 U8712 ( .B1(n7189), .B2(n6986), .A(n10149), .ZN(n6987) );
  NAND3_X1 U8713 ( .A1(n6989), .A2(n6988), .A3(n6987), .ZN(n6990) );
  AOI21_X1 U8714 ( .B1(n7184), .B2(n10143), .A(n6990), .ZN(n6991) );
  OAI21_X1 U8715 ( .B1(n6992), .B2(n8703), .A(n6991), .ZN(P2_U3188) );
  NAND2_X1 U8716 ( .A1(n6994), .A2(n6993), .ZN(n6995) );
  NAND2_X1 U8717 ( .A1(n10085), .A2(n6529), .ZN(n9347) );
  AND2_X1 U8718 ( .A1(n7162), .A2(n7022), .ZN(n7001) );
  INV_X1 U8719 ( .A(n7001), .ZN(n9343) );
  NAND2_X1 U8720 ( .A1(n10085), .A2(n7022), .ZN(n6997) );
  OR2_X1 U8721 ( .A1(n7048), .A2(n7278), .ZN(n9248) );
  NAND2_X1 U8722 ( .A1(n7048), .A2(n7278), .ZN(n9345) );
  NAND2_X1 U8723 ( .A1(n9248), .A2(n9345), .ZN(n9294) );
  OAI21_X1 U8724 ( .B1(n6998), .B2(n9294), .A(n7050), .ZN(n7081) );
  NOR2_X1 U8725 ( .A1(n7161), .A2(n7162), .ZN(n7160) );
  INV_X1 U8726 ( .A(n7048), .ZN(n7089) );
  OAI21_X1 U8727 ( .B1(n7160), .B2(n7089), .A(n9739), .ZN(n6999) );
  AND2_X1 U8728 ( .A1(n7160), .A2(n7089), .ZN(n7272) );
  NOR2_X1 U8729 ( .A1(n6999), .A2(n7272), .ZN(n7091) );
  INV_X1 U8730 ( .A(n9480), .ZN(n7051) );
  AND2_X1 U8731 ( .A1(n9347), .A2(n9328), .ZN(n9335) );
  AOI21_X2 U8732 ( .B1(n9330), .B2(n9335), .A(n7001), .ZN(n7057) );
  XOR2_X1 U8733 ( .A(n9294), .B(n7057), .Z(n7002) );
  OAI222_X1 U8734 ( .A1(n9879), .A2(n7051), .B1(n9877), .B2(n7022), .C1(n7002), 
        .C2(n10068), .ZN(n7085) );
  AOI211_X1 U8735 ( .C1(n10100), .C2(n7081), .A(n7091), .B(n7085), .ZN(n7007)
         );
  AOI22_X1 U8736 ( .A1(n9819), .A2(n7048), .B1(n10126), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n7003) );
  OAI21_X1 U8737 ( .B1(n7007), .B2(n10126), .A(n7003), .ZN(P1_U3527) );
  INV_X1 U8738 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7004) );
  OAI22_X1 U8739 ( .A1(n9948), .A2(n7089), .B1(n10119), .B2(n7004), .ZN(n7005)
         );
  INV_X1 U8740 ( .A(n7005), .ZN(n7006) );
  OAI21_X1 U8741 ( .B1(n7007), .B2(n10117), .A(n7006), .ZN(P1_U3468) );
  OAI22_X1 U8742 ( .A1(n7010), .A2(n7009), .B1(n7008), .B2(n8540), .ZN(n7146)
         );
  XNOR2_X1 U8743 ( .A(n7012), .B(n7011), .ZN(n7143) );
  XNOR2_X1 U8744 ( .A(n7143), .B(n5200), .ZN(n7145) );
  XOR2_X1 U8745 ( .A(n7146), .B(n7145), .Z(n7017) );
  NOR2_X1 U8746 ( .A1(n8516), .A2(n5182), .ZN(n7015) );
  INV_X1 U8747 ( .A(n8518), .ZN(n8508) );
  INV_X1 U8748 ( .A(n8482), .ZN(n7316) );
  NAND2_X1 U8749 ( .A1(n7013), .A2(n8037), .ZN(n10154) );
  OAI22_X1 U8750 ( .A1(n8508), .A2(n7244), .B1(n7316), .B2(n10154), .ZN(n7014)
         );
  AOI211_X1 U8751 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n8043), .A(n7015), .B(
        n7014), .ZN(n7016) );
  OAI21_X1 U8752 ( .B1(n7017), .B2(n8522), .A(n7016), .ZN(P2_U3177) );
  NAND2_X1 U8753 ( .A1(n7019), .A2(n7018), .ZN(n7021) );
  XNOR2_X1 U8754 ( .A(n7021), .B(n7020), .ZN(n7029) );
  NOR2_X1 U8755 ( .A1(n9189), .A2(n7022), .ZN(n7025) );
  OAI21_X1 U8756 ( .B1(n9209), .B2(n7051), .A(n7023), .ZN(n7024) );
  AOI211_X1 U8757 ( .C1(n7048), .C2(n9142), .A(n7025), .B(n7024), .ZN(n7028)
         );
  NAND2_X1 U8758 ( .A1(n9210), .A2(n7026), .ZN(n7027) );
  OAI211_X1 U8759 ( .C1(n7029), .C2(n9145), .A(n7028), .B(n7027), .ZN(P1_U3227) );
  NAND2_X1 U8760 ( .A1(n8928), .A2(n7030), .ZN(n7031) );
  OAI21_X1 U8761 ( .B1(n8928), .B2(n6790), .A(n7031), .ZN(P2_U3459) );
  AOI22_X1 U8762 ( .A1(n7036), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n7370), .B2(
        n7374), .ZN(n7035) );
  OAI21_X1 U8763 ( .B1(n6153), .B2(n7033), .A(n7032), .ZN(n7034) );
  NAND2_X1 U8764 ( .A1(n7035), .A2(n7034), .ZN(n7369) );
  OAI21_X1 U8765 ( .B1(n7035), .B2(n7034), .A(n7369), .ZN(n7047) );
  AOI22_X1 U8766 ( .A1(n7036), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n6173), .B2(
        n7374), .ZN(n7041) );
  NAND2_X1 U8767 ( .A1(n7037), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7039) );
  NAND2_X1 U8768 ( .A1(n7039), .A2(n7038), .ZN(n7040) );
  NAND2_X1 U8769 ( .A1(n7041), .A2(n7040), .ZN(n7373) );
  OAI21_X1 U8770 ( .B1(n7041), .B2(n7040), .A(n7373), .ZN(n7042) );
  NOR2_X1 U8771 ( .A1(n7042), .A2(n9494), .ZN(n7045) );
  NAND2_X1 U8772 ( .A1(n10030), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n7043) );
  NAND2_X1 U8773 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9029) );
  OAI211_X1 U8774 ( .C1(n10027), .C2(n7374), .A(n7043), .B(n9029), .ZN(n7044)
         );
  NOR2_X1 U8775 ( .A1(n7045), .A2(n7044), .ZN(n7046) );
  OAI21_X1 U8776 ( .B1(n7047), .B2(n9493), .A(n7046), .ZN(P1_U3257) );
  OR2_X1 U8777 ( .A1(n7048), .A2(n9481), .ZN(n7049) );
  NAND2_X1 U8778 ( .A1(n7050), .A2(n7049), .ZN(n7270) );
  NOR2_X1 U8779 ( .A1(n7274), .A2(n7051), .ZN(n7356) );
  INV_X1 U8780 ( .A(n7356), .ZN(n7058) );
  AND2_X1 U8781 ( .A1(n7274), .A2(n7051), .ZN(n7359) );
  INV_X1 U8782 ( .A(n7359), .ZN(n9350) );
  NAND2_X1 U8783 ( .A1(n7058), .A2(n9350), .ZN(n9296) );
  NAND2_X1 U8784 ( .A1(n7270), .A2(n9296), .ZN(n7269) );
  OR2_X1 U8785 ( .A1(n7274), .A2(n9480), .ZN(n7052) );
  NAND2_X1 U8786 ( .A1(n7269), .A2(n7052), .ZN(n7054) );
  XNOR2_X1 U8787 ( .A(n7355), .B(n9479), .ZN(n9349) );
  INV_X1 U8788 ( .A(n9349), .ZN(n7053) );
  NAND2_X1 U8789 ( .A1(n7054), .A2(n7053), .ZN(n7117) );
  OAI21_X1 U8790 ( .B1(n7054), .B2(n7053), .A(n7117), .ZN(n7298) );
  INV_X1 U8791 ( .A(n7274), .ZN(n10091) );
  NAND2_X1 U8792 ( .A1(n7272), .A2(n10091), .ZN(n7271) );
  AOI21_X1 U8793 ( .B1(n7271), .B2(n7355), .A(n9750), .ZN(n7055) );
  OR2_X1 U8794 ( .A1(n7271), .A2(n7355), .ZN(n7123) );
  NAND2_X1 U8795 ( .A1(n7055), .A2(n7123), .ZN(n7304) );
  AOI22_X1 U8796 ( .A1(n10104), .A2(n9480), .B1(n9478), .B2(n10105), .ZN(n7056) );
  NAND2_X1 U8797 ( .A1(n7304), .A2(n7056), .ZN(n7063) );
  NAND2_X1 U8798 ( .A1(n7057), .A2(n9345), .ZN(n7276) );
  NAND2_X1 U8799 ( .A1(n7058), .A2(n9248), .ZN(n9351) );
  INV_X1 U8800 ( .A(n9351), .ZN(n7059) );
  NAND2_X1 U8801 ( .A1(n7276), .A2(n7059), .ZN(n7060) );
  NAND2_X1 U8802 ( .A1(n7060), .A2(n9350), .ZN(n7061) );
  NAND2_X1 U8803 ( .A1(n7061), .A2(n9349), .ZN(n7120) );
  OAI21_X1 U8804 ( .B1(n7061), .B2(n9349), .A(n7120), .ZN(n7062) );
  AND2_X1 U8805 ( .A1(n7062), .A2(n10116), .ZN(n7306) );
  AOI211_X1 U8806 ( .C1(n7298), .C2(n10100), .A(n7063), .B(n7306), .ZN(n7068)
         );
  INV_X1 U8807 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7064) );
  NOR2_X1 U8808 ( .A1(n10119), .A2(n7064), .ZN(n7065) );
  AOI21_X1 U8809 ( .B1(n7355), .B2(n9936), .A(n7065), .ZN(n7066) );
  OAI21_X1 U8810 ( .B1(n7068), .B2(n10117), .A(n7066), .ZN(P1_U3474) );
  AOI22_X1 U8811 ( .A1(n7355), .A2(n9819), .B1(n10126), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7067) );
  OAI21_X1 U8812 ( .B1(n7068), .B2(n10126), .A(n7067), .ZN(P1_U3529) );
  XOR2_X1 U8813 ( .A(n7070), .B(n7071), .Z(n7077) );
  NOR2_X1 U8814 ( .A1(n9189), .A2(n7278), .ZN(n7074) );
  INV_X1 U8815 ( .A(n9479), .ZN(n7354) );
  OAI21_X1 U8816 ( .B1(n9209), .B2(n7354), .A(n7072), .ZN(n7073) );
  AOI211_X1 U8817 ( .C1(n7274), .C2(n9142), .A(n7074), .B(n7073), .ZN(n7076)
         );
  NAND2_X1 U8818 ( .A1(n9210), .A2(n7273), .ZN(n7075) );
  OAI211_X1 U8819 ( .C1(n7077), .C2(n9145), .A(n7076), .B(n7075), .ZN(P1_U3239) );
  INV_X1 U8820 ( .A(n7078), .ZN(n7080) );
  INV_X1 U8821 ( .A(n10042), .ZN(n7715) );
  OAI222_X1 U8822 ( .A1(n9971), .A2(n10319), .B1(n9964), .B2(n7080), .C1(
        P1_U3086), .C2(n7715), .ZN(P1_U3338) );
  INV_X1 U8823 ( .A(n8668), .ZN(n8640) );
  OAI222_X1 U8824 ( .A1(n8640), .A2(P2_U3151), .B1(n9023), .B2(n7080), .C1(
        n7079), .C2(n9013), .ZN(P2_U3278) );
  INV_X1 U8825 ( .A(n7081), .ZN(n7094) );
  AND2_X1 U8826 ( .A1(n7082), .A2(n7083), .ZN(n7084) );
  INV_X1 U8827 ( .A(n7085), .ZN(n7086) );
  MUX2_X1 U8828 ( .A(n7087), .B(n7086), .S(n10056), .Z(n7093) );
  OAI22_X1 U8829 ( .A1(n9752), .A2(n7089), .B1(n9557), .B2(n7088), .ZN(n7090)
         );
  AOI21_X1 U8830 ( .B1(n7091), .B2(n10053), .A(n7090), .ZN(n7092) );
  OAI211_X1 U8831 ( .C1(n7094), .C2(n9767), .A(n7093), .B(n7092), .ZN(P1_U3288) );
  XNOR2_X1 U8832 ( .A(n4847), .B(n7095), .ZN(n7173) );
  INV_X1 U8833 ( .A(n7096), .ZN(n7099) );
  NAND3_X1 U8834 ( .A1(n7099), .A2(n7098), .A3(n7097), .ZN(n7111) );
  INV_X1 U8835 ( .A(n7100), .ZN(n7101) );
  NAND2_X1 U8836 ( .A1(n10155), .A2(n8191), .ZN(n10156) );
  INV_X1 U8837 ( .A(n10156), .ZN(n7103) );
  NAND2_X1 U8838 ( .A1(n10161), .A2(n7103), .ZN(n7758) );
  OAI21_X1 U8839 ( .B1(n7105), .B2(n7095), .A(n7104), .ZN(n7109) );
  OAI22_X1 U8840 ( .A1(n7106), .A2(n8727), .B1(n5200), .B2(n7469), .ZN(n7108)
         );
  NOR2_X1 U8841 ( .A1(n7173), .A2(n7753), .ZN(n7107) );
  AOI211_X1 U8842 ( .C1(n8862), .C2(n7109), .A(n7108), .B(n7107), .ZN(n7174)
         );
  MUX2_X1 U8843 ( .A(n7110), .B(n7174), .S(n10161), .Z(n7115) );
  INV_X1 U8844 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8053) );
  OAI22_X1 U8845 ( .A1(n8856), .A2(n5183), .B1(n8053), .B2(n8854), .ZN(n7113)
         );
  INV_X1 U8846 ( .A(n7113), .ZN(n7114) );
  OAI211_X1 U8847 ( .C1(n7173), .C2(n7758), .A(n7115), .B(n7114), .ZN(P2_U3232) );
  OR2_X1 U8848 ( .A1(n7355), .A2(n9479), .ZN(n7116) );
  NAND2_X1 U8849 ( .A1(n7117), .A2(n7116), .ZN(n7118) );
  OR2_X1 U8850 ( .A1(n7285), .A2(n7609), .ZN(n9355) );
  NAND2_X1 U8851 ( .A1(n7285), .A2(n7609), .ZN(n9357) );
  NAND2_X1 U8852 ( .A1(n9355), .A2(n9357), .ZN(n7119) );
  NAND2_X1 U8853 ( .A1(n7118), .A2(n7119), .ZN(n7287) );
  OAI21_X1 U8854 ( .B1(n7118), .B2(n7119), .A(n7287), .ZN(n7209) );
  NAND2_X1 U8855 ( .A1(n7355), .A2(n7354), .ZN(n7353) );
  AOI21_X1 U8856 ( .B1(n7120), .B2(n7353), .A(n7119), .ZN(n7283) );
  AND3_X1 U8857 ( .A1(n7120), .A2(n7353), .A3(n7119), .ZN(n7121) );
  OR2_X1 U8858 ( .A1(n7283), .A2(n7121), .ZN(n7122) );
  NAND2_X1 U8859 ( .A1(n7122), .A2(n10116), .ZN(n7217) );
  AOI22_X1 U8860 ( .A1(n10104), .A2(n9479), .B1(n9477), .B2(n10105), .ZN(n7125) );
  AOI21_X1 U8861 ( .B1(n7285), .B2(n7123), .A(n9750), .ZN(n7124) );
  OR2_X1 U8862 ( .A1(n7123), .A2(n7285), .ZN(n7290) );
  NAND2_X1 U8863 ( .A1(n7124), .A2(n7290), .ZN(n7212) );
  NAND3_X1 U8864 ( .A1(n7217), .A2(n7125), .A3(n7212), .ZN(n7126) );
  AOI21_X1 U8865 ( .B1(n7209), .B2(n10100), .A(n7126), .ZN(n7131) );
  AOI22_X1 U8866 ( .A1(n7285), .A2(n9819), .B1(n10126), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7127) );
  OAI21_X1 U8867 ( .B1(n7131), .B2(n10126), .A(n7127), .ZN(P1_U3530) );
  INV_X1 U8868 ( .A(n7285), .ZN(n7519) );
  INV_X1 U8869 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7128) );
  OAI22_X1 U8870 ( .A1(n7519), .A2(n9948), .B1(n10119), .B2(n7128), .ZN(n7129)
         );
  INV_X1 U8871 ( .A(n7129), .ZN(n7130) );
  OAI21_X1 U8872 ( .B1(n7131), .B2(n10117), .A(n7130), .ZN(P1_U3477) );
  XOR2_X1 U8873 ( .A(n7134), .B(n7133), .Z(n7135) );
  XNOR2_X1 U8874 ( .A(n7132), .B(n7135), .ZN(n7141) );
  NAND2_X1 U8875 ( .A1(n9215), .A2(n9480), .ZN(n7137) );
  OAI211_X1 U8876 ( .C1(n7609), .C2(n9209), .A(n7137), .B(n7136), .ZN(n7138)
         );
  AOI21_X1 U8877 ( .B1(n7299), .B2(n9210), .A(n7138), .ZN(n7140) );
  NAND2_X1 U8878 ( .A1(n9142), .A2(n7355), .ZN(n7139) );
  OAI211_X1 U8879 ( .C1(n7141), .C2(n9145), .A(n7140), .B(n7139), .ZN(P1_U3213) );
  XNOR2_X1 U8880 ( .A(n8124), .B(n8220), .ZN(n7310) );
  XNOR2_X1 U8881 ( .A(n7310), .B(n8537), .ZN(n7150) );
  XNOR2_X1 U8882 ( .A(n7012), .B(n7477), .ZN(n7147) );
  INV_X1 U8883 ( .A(n7147), .ZN(n7148) );
  INV_X1 U8884 ( .A(n7143), .ZN(n7144) );
  XNOR2_X1 U8885 ( .A(n7147), .B(n7244), .ZN(n8383) );
  AOI21_X1 U8886 ( .B1(n7150), .B2(n7149), .A(n7311), .ZN(n7157) );
  INV_X1 U8887 ( .A(n8516), .ZN(n8506) );
  AOI22_X1 U8888 ( .A1(n8506), .A2(n8538), .B1(n8518), .B2(n7443), .ZN(n7154)
         );
  NOR2_X1 U8889 ( .A1(n8220), .A2(n8476), .ZN(n7245) );
  INV_X1 U8890 ( .A(n7151), .ZN(n7152) );
  AOI21_X1 U8891 ( .B1(n8482), .B2(n7245), .A(n7152), .ZN(n7153) );
  OAI211_X1 U8892 ( .C1(n7453), .C2(n8520), .A(n7154), .B(n7153), .ZN(n7155)
         );
  INV_X1 U8893 ( .A(n7155), .ZN(n7156) );
  OAI21_X1 U8894 ( .B1(n7157), .B2(n8522), .A(n7156), .ZN(P2_U3170) );
  OAI21_X1 U8895 ( .B1(n7159), .B2(n7165), .A(n7158), .ZN(n10088) );
  AOI211_X1 U8896 ( .C1(n7162), .C2(n7161), .A(n9750), .B(n7160), .ZN(n10083)
         );
  INV_X2 U8897 ( .A(n9557), .ZN(n10051) );
  AOI22_X1 U8898 ( .A1(n10083), .A2(n10053), .B1(n7163), .B2(n10051), .ZN(
        n7164) );
  OAI21_X1 U8899 ( .B1(n10085), .B2(n9752), .A(n7164), .ZN(n7171) );
  NAND2_X1 U8900 ( .A1(n9330), .A2(n9328), .ZN(n7166) );
  XNOR2_X1 U8901 ( .A(n7166), .B(n7165), .ZN(n7167) );
  NAND2_X1 U8902 ( .A1(n7167), .A2(n10116), .ZN(n7169) );
  AOI22_X1 U8903 ( .A1(n10105), .A2(n9481), .B1(n9482), .B2(n10104), .ZN(n7168) );
  NAND2_X1 U8904 ( .A1(n7169), .A2(n7168), .ZN(n10087) );
  MUX2_X1 U8905 ( .A(n10087), .B(P1_REG2_REG_4__SCAN_IN), .S(n10063), .Z(n7170) );
  AOI211_X1 U8906 ( .C1(n10059), .C2(n10088), .A(n7171), .B(n7170), .ZN(n7172)
         );
  INV_X1 U8907 ( .A(n7172), .ZN(P1_U3289) );
  INV_X1 U8908 ( .A(n7173), .ZN(n7177) );
  INV_X1 U8909 ( .A(n7174), .ZN(n7175) );
  AOI211_X1 U8910 ( .C1(n7840), .C2(n7177), .A(n7176), .B(n7175), .ZN(n10165)
         );
  NAND2_X1 U8911 ( .A1(n8884), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7178) );
  OAI21_X1 U8912 ( .B1(n10165), .B2(n8884), .A(n7178), .ZN(P2_U3460) );
  MUX2_X1 U8913 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8670), .Z(n7248) );
  XOR2_X1 U8914 ( .A(n7197), .B(n7248), .Z(n7249) );
  INV_X1 U8915 ( .A(n7179), .ZN(n7181) );
  AOI21_X1 U8916 ( .B1(n7184), .B2(n7181), .A(n7180), .ZN(n7250) );
  XOR2_X1 U8917 ( .A(n7249), .B(n7250), .Z(n7199) );
  NOR2_X1 U8918 ( .A1(n7186), .A2(n5299), .ZN(n7254) );
  AOI21_X1 U8919 ( .B1(n5299), .B2(n7186), .A(n7254), .ZN(n7188) );
  INV_X1 U8920 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7187) );
  OAI22_X1 U8921 ( .A1(n7188), .A2(n10129), .B1(n10141), .B2(n7187), .ZN(n7196) );
  INV_X1 U8922 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7487) );
  INV_X1 U8923 ( .A(n7192), .ZN(n7193) );
  AOI21_X1 U8924 ( .B1(n7487), .B2(n7193), .A(n4798), .ZN(n7194) );
  NAND2_X1 U8925 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7562) );
  OAI21_X1 U8926 ( .B1(n7194), .B2(n8666), .A(n7562), .ZN(n7195) );
  AOI211_X1 U8927 ( .C1(n7197), .C2(n10143), .A(n7196), .B(n7195), .ZN(n7198)
         );
  OAI21_X1 U8928 ( .B1(n7199), .B2(n8703), .A(n7198), .ZN(P2_U3189) );
  INV_X1 U8929 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7200) );
  NOR2_X1 U8930 ( .A1(n9557), .A2(n7200), .ZN(n7202) );
  AOI211_X1 U8931 ( .C1(n7203), .C2(n6736), .A(n7202), .B(n7201), .ZN(n7208)
         );
  AOI22_X1 U8932 ( .A1(n10050), .A2(n7204), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n10063), .ZN(n7207) );
  NAND2_X1 U8933 ( .A1(n7205), .A2(n10059), .ZN(n7206) );
  OAI211_X1 U8934 ( .C1(n7208), .C2(n10063), .A(n7207), .B(n7206), .ZN(
        P1_U3291) );
  NAND2_X1 U8935 ( .A1(n7209), .A2(n10059), .ZN(n7216) );
  INV_X1 U8936 ( .A(n9477), .ZN(n7514) );
  OR2_X1 U8937 ( .A1(n10063), .A2(n9879), .ZN(n9759) );
  OR2_X1 U8938 ( .A1(n10063), .A2(n9877), .ZN(n9562) );
  INV_X1 U8939 ( .A(n9562), .ZN(n9755) );
  NAND2_X1 U8940 ( .A1(n9755), .A2(n9479), .ZN(n7211) );
  AOI22_X1 U8941 ( .A1(n10063), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7516), .B2(
        n10051), .ZN(n7210) );
  OAI211_X1 U8942 ( .C1(n7514), .C2(n9759), .A(n7211), .B(n7210), .ZN(n7214)
         );
  NOR2_X1 U8943 ( .A1(n7212), .A2(n9740), .ZN(n7213) );
  AOI211_X1 U8944 ( .C1(n10050), .C2(n7285), .A(n7214), .B(n7213), .ZN(n7215)
         );
  OAI211_X1 U8945 ( .C1(n10063), .C2(n7217), .A(n7216), .B(n7215), .ZN(
        P1_U3285) );
  INV_X1 U8946 ( .A(n10154), .ZN(n7228) );
  INV_X1 U8947 ( .A(n7753), .ZN(n7226) );
  OAI22_X1 U8948 ( .A1(n5182), .A2(n8727), .B1(n7244), .B2(n7469), .ZN(n7225)
         );
  AOI21_X1 U8949 ( .B1(n7223), .B2(n7222), .A(n7467), .ZN(n7224) );
  AOI211_X1 U8950 ( .C1(n7226), .C2(n10153), .A(n7225), .B(n7224), .ZN(n7227)
         );
  INV_X1 U8951 ( .A(n7227), .ZN(n10159) );
  AOI211_X1 U8952 ( .C1(n7840), .C2(n10153), .A(n7228), .B(n10159), .ZN(n10167) );
  OR2_X1 U8953 ( .A1(n10167), .A2(n8884), .ZN(n7229) );
  OAI21_X1 U8954 ( .B1(n8928), .B2(n7230), .A(n7229), .ZN(P2_U3461) );
  XNOR2_X1 U8955 ( .A(n7231), .B(n8153), .ZN(n7480) );
  NOR2_X1 U8956 ( .A1(n7477), .A2(n8476), .ZN(n8387) );
  XNOR2_X1 U8957 ( .A(n7232), .B(n8153), .ZN(n7233) );
  OAI222_X1 U8958 ( .A1(n7469), .A2(n7323), .B1(n8727), .B2(n5200), .C1(n7467), 
        .C2(n7233), .ZN(n7476) );
  AOI211_X1 U8959 ( .C1(n7480), .C2(n8909), .A(n8387), .B(n7476), .ZN(n10169)
         );
  OR2_X1 U8960 ( .A1(n10169), .A2(n8884), .ZN(n7234) );
  OAI21_X1 U8961 ( .B1(n8928), .B2(n7235), .A(n7234), .ZN(P2_U3462) );
  INV_X1 U8962 ( .A(n7236), .ZN(n7238) );
  INV_X1 U8963 ( .A(n8696), .ZN(n8674) );
  OAI222_X1 U8964 ( .A1(n9013), .A2(n7237), .B1(n9023), .B2(n7238), .C1(
        P2_U3151), .C2(n8674), .ZN(P2_U3277) );
  INV_X1 U8965 ( .A(n9489), .ZN(n7720) );
  OAI222_X1 U8966 ( .A1(P1_U3086), .A2(n7720), .B1(n9964), .B2(n7238), .C1(
        n10338), .C2(n9971), .ZN(P1_U3337) );
  OAI21_X1 U8967 ( .B1(n7240), .B2(n8209), .A(n7239), .ZN(n7456) );
  XNOR2_X1 U8968 ( .A(n7241), .B(n8209), .ZN(n7242) );
  OAI222_X1 U8969 ( .A1(n8727), .A2(n7244), .B1(n7469), .B2(n7243), .C1(n7242), 
        .C2(n7467), .ZN(n7451) );
  AOI211_X1 U8970 ( .C1(n8909), .C2(n7456), .A(n7245), .B(n7451), .ZN(n10171)
         );
  OR2_X1 U8971 ( .A1(n10171), .A2(n8884), .ZN(n7246) );
  OAI21_X1 U8972 ( .B1(n8928), .B2(n6833), .A(n7246), .ZN(P2_U3463) );
  MUX2_X1 U8973 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8670), .Z(n7382) );
  XNOR2_X1 U8974 ( .A(n7382), .B(n7390), .ZN(n7384) );
  OAI22_X1 U8975 ( .A1(n7250), .A2(n7249), .B1(n7248), .B2(n7247), .ZN(n7385)
         );
  XOR2_X1 U8976 ( .A(n7384), .B(n7385), .Z(n7268) );
  INV_X1 U8977 ( .A(n7251), .ZN(n7253) );
  XNOR2_X1 U8978 ( .A(n7390), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7252) );
  OAI21_X1 U8979 ( .B1(n7254), .B2(n7253), .A(n7252), .ZN(n7388) );
  OR3_X1 U8980 ( .A1(n7254), .A2(n7253), .A3(n7252), .ZN(n7255) );
  AOI21_X1 U8981 ( .B1(n7388), .B2(n7255), .A(n10129), .ZN(n7266) );
  INV_X1 U8982 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7264) );
  INV_X1 U8983 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7257) );
  XNOR2_X1 U8984 ( .A(n7390), .B(n7257), .ZN(n7259) );
  AND3_X1 U8985 ( .A1(n7260), .A2(n7259), .A3(n7258), .ZN(n7261) );
  OAI21_X1 U8986 ( .B1(n4603), .B2(n7261), .A(n10149), .ZN(n7263) );
  INV_X1 U8987 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7262) );
  OR2_X1 U8988 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7262), .ZN(n7652) );
  OAI211_X1 U8989 ( .C1(n10141), .C2(n7264), .A(n7263), .B(n7652), .ZN(n7265)
         );
  AOI211_X1 U8990 ( .C1(n10143), .C2(n7390), .A(n7266), .B(n7265), .ZN(n7267)
         );
  OAI21_X1 U8991 ( .B1(n7268), .B2(n8703), .A(n7267), .ZN(P2_U3190) );
  OAI21_X1 U8992 ( .B1(n7270), .B2(n9296), .A(n7269), .ZN(n10094) );
  OAI211_X1 U8993 ( .C1(n7272), .C2(n10091), .A(n9739), .B(n7271), .ZN(n10090)
         );
  AOI22_X1 U8994 ( .A1(n10050), .A2(n7274), .B1(n7273), .B2(n10051), .ZN(n7275) );
  OAI21_X1 U8995 ( .B1(n10090), .B2(n9740), .A(n7275), .ZN(n7280) );
  AND2_X1 U8996 ( .A1(n7276), .A2(n9248), .ZN(n7358) );
  XNOR2_X1 U8997 ( .A(n7358), .B(n9296), .ZN(n7277) );
  OAI222_X1 U8998 ( .A1(n9879), .A2(n7354), .B1(n9877), .B2(n7278), .C1(n10068), .C2(n7277), .ZN(n10092) );
  MUX2_X1 U8999 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10092), .S(n10056), .Z(n7279) );
  AOI211_X1 U9000 ( .C1(n10059), .C2(n10094), .A(n7280), .B(n7279), .ZN(n7281)
         );
  INV_X1 U9001 ( .A(n7281), .ZN(P1_U3287) );
  INV_X1 U9002 ( .A(n9357), .ZN(n7282) );
  NOR2_X1 U9003 ( .A1(n7283), .A2(n7282), .ZN(n7284) );
  OR2_X2 U9004 ( .A1(n7347), .A2(n7514), .ZN(n9366) );
  NAND2_X1 U9005 ( .A1(n7347), .A2(n7514), .ZN(n9361) );
  NAND2_X1 U9006 ( .A1(n9366), .A2(n9361), .ZN(n7288) );
  XNOR2_X1 U9007 ( .A(n7284), .B(n7288), .ZN(n7341) );
  INV_X1 U9008 ( .A(n7341), .ZN(n7297) );
  OR2_X1 U9009 ( .A1(n7285), .A2(n9478), .ZN(n7286) );
  NAND2_X1 U9010 ( .A1(n7287), .A2(n7286), .ZN(n7289) );
  NAND2_X1 U9011 ( .A1(n7289), .A2(n7288), .ZN(n7349) );
  OAI21_X1 U9012 ( .B1(n7289), .B2(n7288), .A(n7349), .ZN(n7337) );
  XNOR2_X1 U9013 ( .A(n4888), .B(n7347), .ZN(n7291) );
  AOI22_X1 U9014 ( .A1(n7291), .A2(n9739), .B1(n10105), .B2(n9476), .ZN(n7338)
         );
  AOI22_X1 U9015 ( .A1(n10063), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7611), .B2(
        n10051), .ZN(n7292) );
  OAI21_X1 U9016 ( .B1(n9562), .B2(n7609), .A(n7292), .ZN(n7293) );
  AOI21_X1 U9017 ( .B1(n7347), .B2(n10050), .A(n7293), .ZN(n7294) );
  OAI21_X1 U9018 ( .B1(n7338), .B2(n9740), .A(n7294), .ZN(n7295) );
  AOI21_X1 U9019 ( .B1(n7337), .B2(n10059), .A(n7295), .ZN(n7296) );
  OAI21_X1 U9020 ( .B1(n9746), .B2(n7297), .A(n7296), .ZN(P1_U3284) );
  INV_X1 U9021 ( .A(n7298), .ZN(n7308) );
  NAND2_X1 U9022 ( .A1(n9755), .A2(n9480), .ZN(n7301) );
  AOI22_X1 U9023 ( .A1(n10063), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7299), .B2(
        n10051), .ZN(n7300) );
  OAI211_X1 U9024 ( .C1(n7609), .C2(n9759), .A(n7301), .B(n7300), .ZN(n7302)
         );
  AOI21_X1 U9025 ( .B1(n10050), .B2(n7355), .A(n7302), .ZN(n7303) );
  OAI21_X1 U9026 ( .B1(n9740), .B2(n7304), .A(n7303), .ZN(n7305) );
  AOI21_X1 U9027 ( .B1(n7306), .B2(n10056), .A(n7305), .ZN(n7307) );
  OAI21_X1 U9028 ( .B1(n7308), .B2(n9767), .A(n7307), .ZN(P1_U3286) );
  XNOR2_X1 U9029 ( .A(n8124), .B(n7309), .ZN(n7408) );
  XNOR2_X1 U9030 ( .A(n7408), .B(n7443), .ZN(n7409) );
  INV_X1 U9031 ( .A(n7310), .ZN(n7312) );
  XOR2_X1 U9032 ( .A(n7409), .B(n7410), .Z(n7319) );
  INV_X1 U9033 ( .A(n7313), .ZN(n7329) );
  NAND2_X1 U9034 ( .A1(n7330), .A2(n8037), .ZN(n7460) );
  AOI22_X1 U9035 ( .A1(n8506), .A2(n8537), .B1(n8518), .B2(n8536), .ZN(n7315)
         );
  OAI211_X1 U9036 ( .C1(n7316), .C2(n7460), .A(n7315), .B(n7314), .ZN(n7317)
         );
  AOI21_X1 U9037 ( .B1(n7329), .B2(n8510), .A(n7317), .ZN(n7318) );
  OAI21_X1 U9038 ( .B1(n7319), .B2(n8522), .A(n7318), .ZN(P2_U3167) );
  XNOR2_X1 U9039 ( .A(n7320), .B(n8158), .ZN(n7459) );
  OAI21_X1 U9040 ( .B1(n7322), .B2(n8158), .A(n7321), .ZN(n7325) );
  OAI22_X1 U9041 ( .A1(n7323), .A2(n8727), .B1(n7564), .B2(n7469), .ZN(n7324)
         );
  AOI21_X1 U9042 ( .B1(n7325), .B2(n8862), .A(n7324), .ZN(n7326) );
  OAI21_X1 U9043 ( .B1(n7459), .B2(n7753), .A(n7326), .ZN(n7461) );
  INV_X1 U9044 ( .A(n7461), .ZN(n7327) );
  MUX2_X1 U9045 ( .A(n7328), .B(n7327), .S(n10161), .Z(n7332) );
  AOI22_X1 U9046 ( .A1(n8849), .A2(n7330), .B1(n10160), .B2(n7329), .ZN(n7331)
         );
  OAI211_X1 U9047 ( .C1(n7459), .C2(n7758), .A(n7332), .B(n7331), .ZN(P2_U3228) );
  INV_X1 U9048 ( .A(n7333), .ZN(n7336) );
  OAI222_X1 U9049 ( .A1(n9971), .A2(n7334), .B1(n9964), .B2(n7336), .C1(
        P1_U3086), .C2(n6736), .ZN(P1_U3336) );
  OAI222_X1 U9050 ( .A1(n8352), .A2(P2_U3151), .B1(n9023), .B2(n7336), .C1(
        n7335), .C2(n9013), .ZN(P2_U3276) );
  NAND2_X1 U9051 ( .A1(n7337), .A2(n10100), .ZN(n7339) );
  OAI211_X1 U9052 ( .C1(n7609), .C2(n9877), .A(n7339), .B(n7338), .ZN(n7340)
         );
  AOI21_X1 U9053 ( .B1(n7341), .B2(n10116), .A(n7340), .ZN(n7346) );
  INV_X1 U9054 ( .A(n7347), .ZN(n7614) );
  INV_X1 U9055 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7342) );
  OAI22_X1 U9056 ( .A1(n7614), .A2(n9948), .B1(n10119), .B2(n7342), .ZN(n7343)
         );
  INV_X1 U9057 ( .A(n7343), .ZN(n7344) );
  OAI21_X1 U9058 ( .B1(n7346), .B2(n10117), .A(n7344), .ZN(P1_U3480) );
  AOI22_X1 U9059 ( .A1(n7347), .A2(n9819), .B1(n10126), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7345) );
  OAI21_X1 U9060 ( .B1(n7346), .B2(n10126), .A(n7345), .ZN(P1_U3531) );
  OR2_X1 U9061 ( .A1(n7347), .A2(n9477), .ZN(n7348) );
  NAND2_X1 U9062 ( .A1(n7349), .A2(n7348), .ZN(n7352) );
  INV_X1 U9063 ( .A(n9476), .ZN(n7350) );
  OR2_X1 U9064 ( .A1(n7489), .A2(n7350), .ZN(n9370) );
  NAND2_X1 U9065 ( .A1(n7489), .A2(n7350), .ZN(n9368) );
  INV_X1 U9066 ( .A(n9300), .ZN(n7351) );
  OAI21_X1 U9067 ( .B1(n7352), .B2(n7351), .A(n7491), .ZN(n7399) );
  AND2_X1 U9068 ( .A1(n9357), .A2(n7353), .ZN(n9337) );
  NOR2_X1 U9069 ( .A1(n7355), .A2(n7354), .ZN(n9353) );
  OR2_X1 U9070 ( .A1(n9340), .A2(n9353), .ZN(n9289) );
  OR2_X1 U9071 ( .A1(n9289), .A2(n7356), .ZN(n7357) );
  NAND2_X1 U9072 ( .A1(n9299), .A2(n7357), .ZN(n9250) );
  NAND3_X1 U9073 ( .A1(n9250), .A2(n9252), .A3(n9300), .ZN(n7492) );
  INV_X1 U9074 ( .A(n7492), .ZN(n7362) );
  AOI21_X1 U9075 ( .B1(n9250), .B2(n9252), .A(n9300), .ZN(n7361) );
  NOR2_X1 U9076 ( .A1(n7362), .A2(n7361), .ZN(n7407) );
  AOI22_X1 U9077 ( .A1(n10104), .A2(n9477), .B1(n9475), .B2(n10105), .ZN(n7363) );
  INV_X1 U9078 ( .A(n7489), .ZN(n7810) );
  OAI211_X1 U9079 ( .C1(n4601), .C2(n7810), .A(n9739), .B(n4531), .ZN(n7402)
         );
  OAI211_X1 U9080 ( .C1(n7407), .C2(n10068), .A(n7363), .B(n7402), .ZN(n7364)
         );
  AOI21_X1 U9081 ( .B1(n7399), .B2(n10100), .A(n7364), .ZN(n7368) );
  OAI22_X1 U9082 ( .A1(n7810), .A2(n9948), .B1(n10119), .B2(n6087), .ZN(n7365)
         );
  INV_X1 U9083 ( .A(n7365), .ZN(n7366) );
  OAI21_X1 U9084 ( .B1(n7368), .B2(n10117), .A(n7366), .ZN(P1_U3483) );
  AOI22_X1 U9085 ( .A1(n7489), .A2(n9819), .B1(n10126), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7367) );
  OAI21_X1 U9086 ( .B1(n7368), .B2(n10126), .A(n7367), .ZN(P1_U3532) );
  OAI21_X1 U9087 ( .B1(n7370), .B2(n7374), .A(n7369), .ZN(n7575) );
  XOR2_X1 U9088 ( .A(n7575), .B(n7576), .Z(n7371) );
  NAND2_X1 U9089 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7371), .ZN(n7577) );
  OAI21_X1 U9090 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n7371), .A(n7577), .ZN(
        n7380) );
  NAND2_X1 U9091 ( .A1(n10030), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7372) );
  NAND2_X1 U9092 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9208) );
  NAND2_X1 U9093 ( .A1(n7372), .A2(n9208), .ZN(n7378) );
  OAI21_X1 U9094 ( .B1(n6173), .B2(n7374), .A(n7373), .ZN(n7569) );
  XOR2_X1 U9095 ( .A(n7569), .B(n7576), .Z(n7375) );
  NAND2_X1 U9096 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n7375), .ZN(n7570) );
  OAI21_X1 U9097 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n7375), .A(n7570), .ZN(
        n7376) );
  NOR2_X1 U9098 ( .A1(n7376), .A2(n9494), .ZN(n7377) );
  AOI211_X1 U9099 ( .C1(n10041), .C2(n7576), .A(n7378), .B(n7377), .ZN(n7379)
         );
  OAI21_X1 U9100 ( .B1(n7380), .B2(n9493), .A(n7379), .ZN(P1_U3258) );
  MUX2_X1 U9101 ( .A(n7381), .B(n4655), .S(n8670), .Z(n7534) );
  XNOR2_X1 U9102 ( .A(n7534), .B(n7387), .ZN(n7537) );
  INV_X1 U9103 ( .A(n7382), .ZN(n7383) );
  XOR2_X1 U9104 ( .A(n7537), .B(n7538), .Z(n7398) );
  OAI21_X1 U9105 ( .B1(n4597), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7530), .ZN(
        n7396) );
  OAI21_X1 U9106 ( .B1(n7390), .B2(n7389), .A(n7388), .ZN(n7521) );
  XNOR2_X1 U9107 ( .A(n7521), .B(n7535), .ZN(n7391) );
  AOI21_X1 U9108 ( .B1(n7381), .B2(n7391), .A(n7520), .ZN(n7392) );
  NOR2_X1 U9109 ( .A1(n7392), .A2(n10129), .ZN(n7395) );
  AND2_X1 U9110 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7734) );
  AOI21_X1 U9111 ( .B1(n8704), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7734), .ZN(
        n7393) );
  OAI21_X1 U9112 ( .B1(n7535), .B2(n8706), .A(n7393), .ZN(n7394) );
  AOI211_X1 U9113 ( .C1(n7396), .C2(n10149), .A(n7395), .B(n7394), .ZN(n7397)
         );
  OAI21_X1 U9114 ( .B1(n7398), .B2(n8703), .A(n7397), .ZN(P2_U3191) );
  NAND2_X1 U9115 ( .A1(n7399), .A2(n10059), .ZN(n7406) );
  NAND2_X1 U9116 ( .A1(n9755), .A2(n9477), .ZN(n7401) );
  AOI22_X1 U9117 ( .A1(n10063), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n5122), .B2(
        n10051), .ZN(n7400) );
  OAI211_X1 U9118 ( .C1(n9087), .C2(n9759), .A(n7401), .B(n7400), .ZN(n7404)
         );
  NOR2_X1 U9119 ( .A1(n7402), .A2(n9740), .ZN(n7403) );
  AOI211_X1 U9120 ( .C1(n10050), .C2(n7489), .A(n7404), .B(n7403), .ZN(n7405)
         );
  OAI211_X1 U9121 ( .C1(n7407), .C2(n9746), .A(n7406), .B(n7405), .ZN(P1_U3283) );
  XNOR2_X1 U9122 ( .A(n8124), .B(n7547), .ZN(n7557) );
  XNOR2_X1 U9123 ( .A(n7557), .B(n8536), .ZN(n7412) );
  AOI211_X1 U9124 ( .C1(n7412), .C2(n7411), .A(n8522), .B(n7556), .ZN(n7418)
         );
  AOI22_X1 U9125 ( .A1(n8506), .A2(n7443), .B1(n8518), .B2(n7649), .ZN(n7416)
         );
  AND2_X1 U9126 ( .A1(n7413), .A2(n8037), .ZN(n7449) );
  AOI21_X1 U9127 ( .B1(n8482), .B2(n7449), .A(n7414), .ZN(n7415) );
  OAI211_X1 U9128 ( .C1(n7546), .C2(n8520), .A(n7416), .B(n7415), .ZN(n7417)
         );
  OR2_X1 U9129 ( .A1(n7418), .A2(n7417), .ZN(P2_U3179) );
  INV_X1 U9130 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10458) );
  INV_X1 U9131 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10415) );
  NAND2_X1 U9132 ( .A1(n7419), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7422) );
  NAND2_X1 U9133 ( .A1(n7420), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7421) );
  OAI211_X1 U9134 ( .C1(n10415), .C2(n5225), .A(n7422), .B(n7421), .ZN(n7423)
         );
  INV_X1 U9135 ( .A(n7423), .ZN(n7424) );
  NAND2_X1 U9136 ( .A1(n8710), .A2(P2_U3893), .ZN(n7426) );
  OAI21_X1 U9137 ( .B1(P2_U3893), .B2(n10458), .A(n7426), .ZN(P2_U3522) );
  XNOR2_X1 U9138 ( .A(n7427), .B(n8228), .ZN(n7484) );
  AOI22_X1 U9139 ( .A1(n8536), .A2(n8866), .B1(n8865), .B2(n8535), .ZN(n7433)
         );
  INV_X1 U9140 ( .A(n7428), .ZN(n7429) );
  OAI21_X1 U9141 ( .B1(n7429), .B2(n7441), .A(n8228), .ZN(n7431) );
  NAND3_X1 U9142 ( .A1(n7431), .A2(n8862), .A3(n7430), .ZN(n7432) );
  OAI211_X1 U9143 ( .C1(n7484), .C2(n7753), .A(n7433), .B(n7432), .ZN(n7486)
         );
  NAND2_X1 U9144 ( .A1(n7486), .A2(n10161), .ZN(n7436) );
  OAI22_X1 U9145 ( .A1(n8856), .A2(n7558), .B1(n7568), .B2(n8854), .ZN(n7434)
         );
  AOI21_X1 U9146 ( .B1(n10163), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7434), .ZN(
        n7435) );
  OAI211_X1 U9147 ( .C1(n7484), .C2(n7758), .A(n7436), .B(n7435), .ZN(P2_U3226) );
  NAND2_X1 U9148 ( .A1(n7438), .A2(n7437), .ZN(n8155) );
  INV_X1 U9149 ( .A(n8155), .ZN(n7440) );
  OAI22_X1 U9150 ( .A1(n7428), .A2(n7441), .B1(n7440), .B2(n7439), .ZN(n7442)
         );
  NAND2_X1 U9151 ( .A1(n7442), .A2(n8862), .ZN(n7445) );
  AOI22_X1 U9152 ( .A1(n8866), .A2(n7443), .B1(n7649), .B2(n8865), .ZN(n7444)
         );
  NAND2_X1 U9153 ( .A1(n7445), .A2(n7444), .ZN(n7548) );
  NAND2_X1 U9154 ( .A1(n7446), .A2(n8213), .ZN(n7447) );
  XNOR2_X1 U9155 ( .A(n7447), .B(n8155), .ZN(n7551) );
  AND2_X1 U9156 ( .A1(n7551), .A2(n8909), .ZN(n7448) );
  NAND2_X1 U9157 ( .A1(n10174), .A2(n8928), .ZN(n7450) );
  OAI21_X1 U9158 ( .B1(n8928), .B2(n6982), .A(n7450), .ZN(P2_U3465) );
  INV_X1 U9159 ( .A(n7451), .ZN(n7458) );
  NAND2_X1 U9160 ( .A1(n7753), .A2(n10156), .ZN(n7452) );
  NOR2_X1 U9161 ( .A1(n10161), .A2(n6829), .ZN(n7455) );
  OAI22_X1 U9162 ( .A1(n8856), .A2(n8220), .B1(n7453), .B2(n8854), .ZN(n7454)
         );
  AOI211_X1 U9163 ( .C1(n8872), .C2(n7456), .A(n7455), .B(n7454), .ZN(n7457)
         );
  OAI21_X1 U9164 ( .B1(n7458), .B2(n10163), .A(n7457), .ZN(P2_U3229) );
  INV_X1 U9165 ( .A(n7459), .ZN(n7463) );
  INV_X1 U9166 ( .A(n7460), .ZN(n7462) );
  AOI211_X1 U9167 ( .C1(n7840), .C2(n7463), .A(n7462), .B(n7461), .ZN(n10173)
         );
  OR2_X1 U9168 ( .A1(n10173), .A2(n8884), .ZN(n7464) );
  OAI21_X1 U9169 ( .B1(n8928), .B2(n5248), .A(n7464), .ZN(P2_U3464) );
  INV_X1 U9170 ( .A(n7649), .ZN(n8231) );
  INV_X1 U9171 ( .A(n7465), .ZN(n8233) );
  NAND2_X1 U9172 ( .A1(n8233), .A2(n8237), .ZN(n8160) );
  XNOR2_X1 U9173 ( .A(n7466), .B(n8160), .ZN(n7468) );
  OAI222_X1 U9174 ( .A1(n8727), .A2(n8231), .B1(n7469), .B2(n7886), .C1(n7468), 
        .C2(n7467), .ZN(n7632) );
  INV_X1 U9175 ( .A(n7632), .ZN(n7475) );
  XNOR2_X1 U9176 ( .A(n7470), .B(n8160), .ZN(n7633) );
  INV_X1 U9177 ( .A(n7471), .ZN(n7657) );
  AOI22_X1 U9178 ( .A1(n10163), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10160), .B2(
        n7657), .ZN(n7472) );
  OAI21_X1 U9179 ( .B1(n7647), .B2(n8856), .A(n7472), .ZN(n7473) );
  AOI21_X1 U9180 ( .B1(n7633), .B2(n8872), .A(n7473), .ZN(n7474) );
  OAI21_X1 U9181 ( .B1(n7475), .B2(n10163), .A(n7474), .ZN(P2_U3225) );
  INV_X1 U9182 ( .A(n7476), .ZN(n7482) );
  NOR2_X1 U9183 ( .A1(n10161), .A2(n5202), .ZN(n7479) );
  OAI22_X1 U9184 ( .A1(n8856), .A2(n7477), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8854), .ZN(n7478) );
  AOI211_X1 U9185 ( .C1(n7480), .C2(n8872), .A(n7479), .B(n7478), .ZN(n7481)
         );
  OAI21_X1 U9186 ( .B1(n10163), .B2(n7482), .A(n7481), .ZN(P2_U3230) );
  OAI22_X1 U9187 ( .A1(n7484), .A2(n7483), .B1(n7558), .B2(n8476), .ZN(n7485)
         );
  NOR2_X1 U9188 ( .A1(n7486), .A2(n7485), .ZN(n10176) );
  OR2_X1 U9189 ( .A1(n8928), .A2(n7487), .ZN(n7488) );
  OAI21_X1 U9190 ( .B1(n10176), .B2(n8884), .A(n7488), .ZN(P2_U3466) );
  OR2_X1 U9191 ( .A1(n7489), .A2(n9476), .ZN(n7490) );
  OR2_X1 U9192 ( .A1(n7497), .A2(n9087), .ZN(n9371) );
  NAND2_X1 U9193 ( .A1(n7497), .A2(n9087), .ZN(n9372) );
  INV_X1 U9194 ( .A(n7493), .ZN(n9301) );
  XNOR2_X1 U9195 ( .A(n7587), .B(n9301), .ZN(n7502) );
  INV_X1 U9196 ( .A(n7593), .ZN(n7595) );
  AOI211_X1 U9197 ( .C1(n7497), .C2(n4531), .A(n9750), .B(n7595), .ZN(n7503)
         );
  AND2_X2 U9198 ( .A1(n7492), .A2(n9368), .ZN(n7494) );
  NAND2_X1 U9199 ( .A1(n7494), .A2(n7493), .ZN(n7588) );
  OAI211_X1 U9200 ( .C1(n7494), .C2(n7493), .A(n7588), .B(n10116), .ZN(n7496)
         );
  AOI22_X1 U9201 ( .A1(n10104), .A2(n9476), .B1(n10103), .B2(n10105), .ZN(
        n7495) );
  NAND2_X1 U9202 ( .A1(n7496), .A2(n7495), .ZN(n7507) );
  AOI211_X1 U9203 ( .C1(n7502), .C2(n10100), .A(n7503), .B(n7507), .ZN(n7501)
         );
  AOI22_X1 U9204 ( .A1(n7497), .A2(n9819), .B1(n10126), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7498) );
  OAI21_X1 U9205 ( .B1(n7501), .B2(n10126), .A(n7498), .ZN(P1_U3533) );
  OAI22_X1 U9206 ( .A1(n9181), .A2(n9948), .B1(n10119), .B2(n6108), .ZN(n7499)
         );
  INV_X1 U9207 ( .A(n7499), .ZN(n7500) );
  OAI21_X1 U9208 ( .B1(n7501), .B2(n10117), .A(n7500), .ZN(P1_U3486) );
  INV_X1 U9209 ( .A(n7502), .ZN(n7509) );
  NAND2_X1 U9210 ( .A1(n7503), .A2(n10053), .ZN(n7505) );
  AOI22_X1 U9211 ( .A1(n10063), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9178), .B2(
        n10051), .ZN(n7504) );
  OAI211_X1 U9212 ( .C1(n9181), .C2(n9752), .A(n7505), .B(n7504), .ZN(n7506)
         );
  AOI21_X1 U9213 ( .B1(n10056), .B2(n7507), .A(n7506), .ZN(n7508) );
  OAI21_X1 U9214 ( .B1(n7509), .B2(n9767), .A(n7508), .ZN(P1_U3282) );
  OAI21_X1 U9215 ( .B1(n7511), .B2(n4598), .A(n7510), .ZN(n7512) );
  NAND2_X1 U9216 ( .A1(n7512), .A2(n9206), .ZN(n7518) );
  NOR2_X1 U9217 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6046), .ZN(n9986) );
  AOI21_X1 U9218 ( .B1(n9215), .B2(n9479), .A(n9986), .ZN(n7513) );
  OAI21_X1 U9219 ( .B1(n7514), .B2(n9209), .A(n7513), .ZN(n7515) );
  AOI21_X1 U9220 ( .B1(n7516), .B2(n9210), .A(n7515), .ZN(n7517) );
  OAI211_X1 U9221 ( .C1(n7519), .C2(n9218), .A(n7518), .B(n7517), .ZN(P1_U3221) );
  NAND2_X1 U9222 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7821), .ZN(n7522) );
  OAI21_X1 U9223 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7821), .A(n7522), .ZN(
        n7523) );
  AOI21_X1 U9224 ( .B1(n7524), .B2(n7523), .A(n7817), .ZN(n7545) );
  NOR2_X1 U9225 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7525), .ZN(n7885) );
  INV_X1 U9226 ( .A(n7885), .ZN(n7526) );
  OAI21_X1 U9227 ( .B1(n10141), .B2(n10293), .A(n7526), .ZN(n7533) );
  NAND2_X1 U9228 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7821), .ZN(n7528) );
  OAI21_X1 U9229 ( .B1(n7821), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7528), .ZN(
        n7529) );
  NAND3_X1 U9230 ( .A1(n7530), .A2(n4653), .A3(n7529), .ZN(n7531) );
  AOI21_X1 U9231 ( .B1(n4599), .B2(n7531), .A(n8666), .ZN(n7532) );
  AOI211_X1 U9232 ( .C1(n10143), .C2(n7539), .A(n7533), .B(n7532), .ZN(n7544)
         );
  INV_X1 U9233 ( .A(n7534), .ZN(n7536) );
  MUX2_X1 U9234 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8670), .Z(n7822) );
  XNOR2_X1 U9235 ( .A(n7822), .B(n7539), .ZN(n7540) );
  OAI21_X1 U9236 ( .B1(n7541), .B2(n7540), .A(n7820), .ZN(n7542) );
  NAND2_X1 U9237 ( .A1(n7542), .A2(n10136), .ZN(n7543) );
  OAI211_X1 U9238 ( .C1(n7545), .C2(n10129), .A(n7544), .B(n7543), .ZN(
        P2_U3192) );
  OAI22_X1 U9239 ( .A1(n8856), .A2(n7547), .B1(n7546), .B2(n8854), .ZN(n7550)
         );
  MUX2_X1 U9240 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7548), .S(n10161), .Z(n7549)
         );
  AOI211_X1 U9241 ( .C1(n8872), .C2(n7551), .A(n7550), .B(n7549), .ZN(n7552)
         );
  INV_X1 U9242 ( .A(n7552), .ZN(P2_U3227) );
  INV_X1 U9243 ( .A(n7553), .ZN(n7554) );
  OAI222_X1 U9244 ( .A1(n8185), .A2(P2_U3151), .B1(n9013), .B2(n5563), .C1(
        n7554), .C2(n9023), .ZN(P2_U3275) );
  OAI222_X1 U9245 ( .A1(n9971), .A2(n7555), .B1(P1_U3086), .B2(n6437), .C1(
        n9964), .C2(n7554), .ZN(P1_U3335) );
  XNOR2_X1 U9246 ( .A(n8124), .B(n7558), .ZN(n7650) );
  XNOR2_X1 U9247 ( .A(n7650), .B(n8231), .ZN(n7559) );
  OAI21_X1 U9248 ( .B1(n7560), .B2(n7559), .A(n7648), .ZN(n7561) );
  NAND2_X1 U9249 ( .A1(n7561), .A2(n8503), .ZN(n7567) );
  NAND2_X1 U9250 ( .A1(n8518), .A2(n8535), .ZN(n7563) );
  OAI211_X1 U9251 ( .C1(n7564), .C2(n8516), .A(n7563), .B(n7562), .ZN(n7565)
         );
  AOI21_X1 U9252 ( .B1(n8527), .B2(n8230), .A(n7565), .ZN(n7566) );
  OAI211_X1 U9253 ( .C1(n8520), .C2(n7568), .A(n7567), .B(n7566), .ZN(P2_U3153) );
  INV_X1 U9254 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7711) );
  AOI22_X1 U9255 ( .A1(n7574), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7711), .B2(
        n7710), .ZN(n7573) );
  NAND2_X1 U9256 ( .A1(n7576), .A2(n7569), .ZN(n7571) );
  NAND2_X1 U9257 ( .A1(n7571), .A2(n7570), .ZN(n7572) );
  NAND2_X1 U9258 ( .A1(n7573), .A2(n7572), .ZN(n7709) );
  OAI21_X1 U9259 ( .B1(n7573), .B2(n7572), .A(n7709), .ZN(n7586) );
  AOI22_X1 U9260 ( .A1(n7574), .A2(n7703), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n7710), .ZN(n7580) );
  NAND2_X1 U9261 ( .A1(n7576), .A2(n7575), .ZN(n7578) );
  NAND2_X1 U9262 ( .A1(n7578), .A2(n7577), .ZN(n7579) );
  NOR2_X1 U9263 ( .A1(n7580), .A2(n7579), .ZN(n7702) );
  AOI21_X1 U9264 ( .B1(n7580), .B2(n7579), .A(n7702), .ZN(n7581) );
  OR2_X1 U9265 ( .A1(n7581), .A2(n9493), .ZN(n7585) );
  NOR2_X1 U9266 ( .A1(n7582), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9109) );
  NOR2_X1 U9267 ( .A1(n10027), .A2(n7710), .ZN(n7583) );
  AOI211_X1 U9268 ( .C1(n10030), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9109), .B(
        n7583), .ZN(n7584) );
  OAI211_X1 U9269 ( .C1(n7586), .C2(n9494), .A(n7585), .B(n7584), .ZN(P1_U3259) );
  INV_X1 U9270 ( .A(n10103), .ZN(n9176) );
  NAND2_X1 U9271 ( .A1(n7616), .A2(n9176), .ZN(n9373) );
  XNOR2_X1 U9272 ( .A(n7615), .B(n9303), .ZN(n10101) );
  INV_X1 U9273 ( .A(n10101), .ZN(n7600) );
  OAI211_X1 U9274 ( .C1(n7590), .C2(n7589), .A(n7623), .B(n10116), .ZN(n7592)
         );
  AOI22_X1 U9275 ( .A1(n10104), .A2(n9475), .B1(n9474), .B2(n10105), .ZN(n7591) );
  NAND2_X1 U9276 ( .A1(n7592), .A2(n7591), .ZN(n10099) );
  INV_X1 U9277 ( .A(n7616), .ZN(n10097) );
  INV_X1 U9278 ( .A(n7625), .ZN(n7594) );
  OAI211_X1 U9279 ( .C1(n10097), .C2(n7595), .A(n7594), .B(n9739), .ZN(n10096)
         );
  AOI22_X1 U9280 ( .A1(n10063), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9089), .B2(
        n10051), .ZN(n7597) );
  NAND2_X1 U9281 ( .A1(n7616), .A2(n10050), .ZN(n7596) );
  OAI211_X1 U9282 ( .C1(n10096), .C2(n9740), .A(n7597), .B(n7596), .ZN(n7598)
         );
  AOI21_X1 U9283 ( .B1(n10099), .B2(n10056), .A(n7598), .ZN(n7599) );
  OAI21_X1 U9284 ( .B1(n7600), .B2(n9767), .A(n7599), .ZN(P1_U3281) );
  OAI21_X1 U9285 ( .B1(n7605), .B2(n7602), .A(n7604), .ZN(n7606) );
  NAND2_X1 U9286 ( .A1(n7606), .A2(n9206), .ZN(n7613) );
  AOI21_X1 U9287 ( .B1(n9186), .B2(n9476), .A(n7607), .ZN(n7608) );
  OAI21_X1 U9288 ( .B1(n7609), .B2(n9189), .A(n7608), .ZN(n7610) );
  AOI21_X1 U9289 ( .B1(n7611), .B2(n9210), .A(n7610), .ZN(n7612) );
  OAI211_X1 U9290 ( .C1(n7614), .C2(n9218), .A(n7613), .B(n7612), .ZN(P1_U3231) );
  NAND2_X1 U9291 ( .A1(n7615), .A2(n9303), .ZN(n7618) );
  OR2_X1 U9292 ( .A1(n7616), .A2(n10103), .ZN(n7617) );
  NAND2_X1 U9293 ( .A1(n7618), .A2(n7617), .ZN(n7759) );
  INV_X1 U9294 ( .A(n9474), .ZN(n7619) );
  OR2_X1 U9295 ( .A1(n7760), .A2(n7619), .ZN(n9379) );
  NAND2_X1 U9296 ( .A1(n7760), .A2(n7619), .ZN(n9384) );
  XOR2_X1 U9297 ( .A(n7759), .B(n9304), .Z(n10112) );
  INV_X1 U9298 ( .A(n7623), .ZN(n7620) );
  INV_X1 U9299 ( .A(n9374), .ZN(n7621) );
  OAI21_X1 U9300 ( .B1(n7620), .B2(n7621), .A(n9304), .ZN(n7624) );
  NOR2_X1 U9301 ( .A1(n9304), .A2(n7621), .ZN(n7622) );
  NAND2_X1 U9302 ( .A1(n7624), .A2(n7762), .ZN(n10115) );
  INV_X1 U9303 ( .A(n9746), .ZN(n9764) );
  INV_X1 U9304 ( .A(n7760), .ZN(n10110) );
  NAND2_X1 U9305 ( .A1(n10110), .A2(n7625), .ZN(n7766) );
  OAI211_X1 U9306 ( .C1(n10110), .C2(n7625), .A(n9739), .B(n7766), .ZN(n10108)
         );
  NAND2_X1 U9307 ( .A1(n9755), .A2(n10103), .ZN(n7627) );
  AOI22_X1 U9308 ( .A1(n10063), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9155), .B2(
        n10051), .ZN(n7626) );
  OAI211_X1 U9309 ( .C1(n9878), .C2(n9759), .A(n7627), .B(n7626), .ZN(n7628)
         );
  AOI21_X1 U9310 ( .B1(n7760), .B2(n10050), .A(n7628), .ZN(n7629) );
  OAI21_X1 U9311 ( .B1(n10108), .B2(n9740), .A(n7629), .ZN(n7630) );
  AOI21_X1 U9312 ( .B1(n10115), .B2(n9764), .A(n7630), .ZN(n7631) );
  OAI21_X1 U9313 ( .B1(n10112), .B2(n9767), .A(n7631), .ZN(P1_U3280) );
  NOR2_X1 U9314 ( .A1(n7647), .A2(n8476), .ZN(n7651) );
  AOI211_X1 U9315 ( .C1(n8909), .C2(n7633), .A(n7651), .B(n7632), .ZN(n10177)
         );
  OR2_X1 U9316 ( .A1(n10177), .A2(n8884), .ZN(n7634) );
  OAI21_X1 U9317 ( .B1(n8928), .B2(n7257), .A(n7634), .ZN(P2_U3467) );
  INV_X1 U9318 ( .A(n7635), .ZN(n7645) );
  OAI222_X1 U9319 ( .A1(P2_U3151), .A2(n7636), .B1(n9023), .B2(n7645), .C1(
        n10369), .C2(n9013), .ZN(P2_U3274) );
  XNOR2_X1 U9320 ( .A(n7637), .B(n8152), .ZN(n7781) );
  AOI22_X1 U9321 ( .A1(n8866), .A2(n8535), .B1(n8533), .B2(n8865), .ZN(n7641)
         );
  XNOR2_X1 U9322 ( .A(n7638), .B(n8152), .ZN(n7639) );
  NAND2_X1 U9323 ( .A1(n7639), .A2(n8862), .ZN(n7640) );
  OAI211_X1 U9324 ( .C1(n7781), .C2(n7753), .A(n7641), .B(n7640), .ZN(n7782)
         );
  NAND2_X1 U9325 ( .A1(n7782), .A2(n10161), .ZN(n7644) );
  OAI22_X1 U9326 ( .A1(n10161), .A2(n7381), .B1(n7738), .B2(n8854), .ZN(n7642)
         );
  AOI21_X1 U9327 ( .B1(n8849), .B2(n7732), .A(n7642), .ZN(n7643) );
  OAI211_X1 U9328 ( .C1(n7781), .C2(n7758), .A(n7644), .B(n7643), .ZN(P2_U3224) );
  INV_X1 U9329 ( .A(n9453), .ZN(n9464) );
  OAI222_X1 U9330 ( .A1(n9971), .A2(n7646), .B1(P1_U3086), .B2(n9464), .C1(
        n9964), .C2(n7645), .ZN(P1_U3334) );
  XNOR2_X1 U9331 ( .A(n8124), .B(n7647), .ZN(n7726) );
  XNOR2_X1 U9332 ( .A(n7726), .B(n7735), .ZN(n7728) );
  XOR2_X1 U9333 ( .A(n7728), .B(n7729), .Z(n7659) );
  NAND2_X1 U9334 ( .A1(n8518), .A2(n8534), .ZN(n7655) );
  NAND2_X1 U9335 ( .A1(n8482), .A2(n7651), .ZN(n7654) );
  OR2_X1 U9336 ( .A1(n8516), .A2(n8231), .ZN(n7653) );
  NAND4_X1 U9337 ( .A1(n7655), .A2(n7654), .A3(n7653), .A4(n7652), .ZN(n7656)
         );
  AOI21_X1 U9338 ( .B1(n8510), .B2(n7657), .A(n7656), .ZN(n7658) );
  OAI21_X1 U9339 ( .B1(n7659), .B2(n8522), .A(n7658), .ZN(P2_U3161) );
  INV_X1 U9340 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U9341 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7696) );
  NOR2_X1 U9342 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7693) );
  NOR2_X1 U9343 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7690) );
  NOR2_X1 U9344 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7687) );
  NOR2_X1 U9345 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7684) );
  NOR2_X1 U9346 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7681) );
  NOR2_X1 U9347 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7679) );
  INV_X1 U9348 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10482) );
  INV_X1 U9349 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7676) );
  NOR2_X1 U9350 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7674) );
  NOR2_X1 U9351 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7672) );
  NOR2_X1 U9352 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n7670) );
  NOR2_X1 U9353 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7668) );
  NOR2_X1 U9354 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7666) );
  NAND2_X1 U9355 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7664) );
  XOR2_X1 U9356 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10596) );
  NAND2_X1 U9357 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7662) );
  AOI21_X1 U9358 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10185) );
  INV_X1 U9359 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10366) );
  INV_X1 U9360 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10187) );
  NOR2_X1 U9361 ( .A1(n10366), .A2(n10187), .ZN(n10186) );
  AOI21_X1 U9362 ( .B1(n10186), .B2(P1_ADDR_REG_1__SCAN_IN), .A(
        P2_ADDR_REG_1__SCAN_IN), .ZN(n10181) );
  NOR2_X1 U9363 ( .A1(n10185), .A2(n10181), .ZN(n10594) );
  INV_X1 U9364 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7660) );
  INV_X1 U9365 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U9366 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .B1(n7660), .B2(n10414), .ZN(n10593) );
  NAND2_X1 U9367 ( .A1(n10594), .A2(n10593), .ZN(n7661) );
  NAND2_X1 U9368 ( .A1(n7662), .A2(n7661), .ZN(n10595) );
  NAND2_X1 U9369 ( .A1(n10596), .A2(n10595), .ZN(n7663) );
  NAND2_X1 U9370 ( .A1(n7664), .A2(n7663), .ZN(n10598) );
  XNOR2_X1 U9371 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10597) );
  NOR2_X1 U9372 ( .A1(n10598), .A2(n10597), .ZN(n7665) );
  NOR2_X1 U9373 ( .A1(n7666), .A2(n7665), .ZN(n10586) );
  XNOR2_X1 U9374 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10585) );
  NOR2_X1 U9375 ( .A1(n10586), .A2(n10585), .ZN(n7667) );
  NOR2_X1 U9376 ( .A1(n7668), .A2(n7667), .ZN(n10584) );
  XNOR2_X1 U9377 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10583) );
  NOR2_X1 U9378 ( .A1(n10584), .A2(n10583), .ZN(n7669) );
  NOR2_X1 U9379 ( .A1(n7670), .A2(n7669), .ZN(n10590) );
  XNOR2_X1 U9380 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10589) );
  NOR2_X1 U9381 ( .A1(n10590), .A2(n10589), .ZN(n7671) );
  NOR2_X1 U9382 ( .A1(n7672), .A2(n7671), .ZN(n10592) );
  XNOR2_X1 U9383 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10591) );
  NOR2_X1 U9384 ( .A1(n10592), .A2(n10591), .ZN(n7673) );
  NOR2_X1 U9385 ( .A1(n7674), .A2(n7673), .ZN(n10588) );
  AOI22_X1 U9386 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7676), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10482), .ZN(n10587) );
  NOR2_X1 U9387 ( .A1(n10588), .A2(n10587), .ZN(n7675) );
  AOI21_X1 U9388 ( .B1(n10482), .B2(n7676), .A(n7675), .ZN(n10207) );
  AOI22_X1 U9389 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7677), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10293), .ZN(n10206) );
  NOR2_X1 U9390 ( .A1(n10207), .A2(n10206), .ZN(n7678) );
  NOR2_X1 U9391 ( .A1(n7679), .A2(n7678), .ZN(n10205) );
  XNOR2_X1 U9392 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10204) );
  NOR2_X1 U9393 ( .A1(n10205), .A2(n10204), .ZN(n7680) );
  NOR2_X1 U9394 ( .A1(n7681), .A2(n7680), .ZN(n10203) );
  INV_X1 U9395 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7682) );
  INV_X1 U9396 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7906) );
  AOI22_X1 U9397 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7682), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7906), .ZN(n10202) );
  NOR2_X1 U9398 ( .A1(n10203), .A2(n10202), .ZN(n7683) );
  NOR2_X1 U9399 ( .A1(n7684), .A2(n7683), .ZN(n10201) );
  INV_X1 U9400 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7685) );
  INV_X1 U9401 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U9402 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n7685), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n10450), .ZN(n10200) );
  NOR2_X1 U9403 ( .A1(n10201), .A2(n10200), .ZN(n7686) );
  NOR2_X1 U9404 ( .A1(n7687), .A2(n7686), .ZN(n10199) );
  INV_X1 U9405 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7688) );
  INV_X1 U9406 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8576) );
  AOI22_X1 U9407 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n7688), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n8576), .ZN(n10198) );
  NOR2_X1 U9408 ( .A1(n10199), .A2(n10198), .ZN(n7689) );
  NOR2_X1 U9409 ( .A1(n7690), .A2(n7689), .ZN(n10197) );
  INV_X1 U9410 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7691) );
  INV_X1 U9411 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U9412 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n7691), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10485), .ZN(n10196) );
  NOR2_X1 U9413 ( .A1(n10197), .A2(n10196), .ZN(n7692) );
  NOR2_X1 U9414 ( .A1(n7693), .A2(n7692), .ZN(n10195) );
  INV_X1 U9415 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7694) );
  INV_X1 U9416 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8623) );
  AOI22_X1 U9417 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7694), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8623), .ZN(n10194) );
  NOR2_X1 U9418 ( .A1(n10195), .A2(n10194), .ZN(n7695) );
  NOR2_X1 U9419 ( .A1(n7696), .A2(n7695), .ZN(n10193) );
  AOI22_X1 U9420 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n10047), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10305), .ZN(n10192) );
  NOR2_X1 U9421 ( .A1(n10193), .A2(n10192), .ZN(n7697) );
  AOI21_X1 U9422 ( .B1(n10305), .B2(n10047), .A(n7697), .ZN(n7698) );
  AND2_X1 U9423 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7698), .ZN(n10189) );
  NOR2_X1 U9424 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10189), .ZN(n7699) );
  NOR2_X1 U9425 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7698), .ZN(n10188) );
  NOR2_X1 U9426 ( .A1(n7699), .A2(n10188), .ZN(n7701) );
  XNOR2_X1 U9427 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7700) );
  XNOR2_X1 U9428 ( .A(n7701), .B(n7700), .ZN(ADD_1068_U4) );
  AOI21_X1 U9429 ( .B1(n7710), .B2(n7703), .A(n7702), .ZN(n10033) );
  XNOR2_X1 U9430 ( .A(n10042), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10032) );
  INV_X1 U9431 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9858) );
  XNOR2_X1 U9432 ( .A(n9489), .B(n9858), .ZN(n7705) );
  NAND2_X1 U9433 ( .A1(n7715), .A2(n10307), .ZN(n7706) );
  AND2_X1 U9434 ( .A1(n7705), .A2(n7706), .ZN(n7704) );
  NAND2_X1 U9435 ( .A1(n10035), .A2(n7704), .ZN(n9491) );
  NAND2_X1 U9436 ( .A1(n9491), .A2(n10043), .ZN(n7725) );
  AOI21_X1 U9437 ( .B1(n10035), .B2(n7706), .A(n7705), .ZN(n7724) );
  INV_X1 U9438 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U9439 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9187) );
  OAI21_X1 U9440 ( .B1(n10048), .B2(n7707), .A(n9187), .ZN(n7708) );
  AOI21_X1 U9441 ( .B1(n9489), .B2(n10041), .A(n7708), .ZN(n7723) );
  OAI21_X1 U9442 ( .B1(n7711), .B2(n7710), .A(n7709), .ZN(n7712) );
  INV_X1 U9443 ( .A(n7712), .ZN(n10037) );
  INV_X1 U9444 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U9445 ( .A1(n10042), .A2(n7714), .ZN(n7713) );
  OAI21_X1 U9446 ( .B1(n10042), .B2(n7714), .A(n7713), .ZN(n10038) );
  NAND2_X1 U9447 ( .A1(n10037), .A2(n10038), .ZN(n10036) );
  NAND2_X1 U9448 ( .A1(n7715), .A2(n7714), .ZN(n7716) );
  NAND2_X1 U9449 ( .A1(n10036), .A2(n7716), .ZN(n7719) );
  NAND2_X1 U9450 ( .A1(n9489), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9486) );
  OAI21_X1 U9451 ( .B1(n9489), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9486), .ZN(
        n7717) );
  OR2_X1 U9452 ( .A1(n7719), .A2(n7717), .ZN(n9487) );
  NAND2_X1 U9453 ( .A1(n7720), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7718) );
  OAI211_X1 U9454 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n7720), .A(n7719), .B(
        n7718), .ZN(n7721) );
  NAND3_X1 U9455 ( .A1(n9487), .A2(n7721), .A3(n10039), .ZN(n7722) );
  OAI211_X1 U9456 ( .C1(n7725), .C2(n7724), .A(n7723), .B(n7722), .ZN(P1_U3261) );
  INV_X1 U9457 ( .A(n7726), .ZN(n7727) );
  XNOR2_X1 U9458 ( .A(n8124), .B(n7732), .ZN(n7860) );
  XOR2_X1 U9459 ( .A(n7886), .B(n7860), .Z(n7730) );
  OAI211_X1 U9460 ( .C1(n7731), .C2(n7730), .A(n7862), .B(n8503), .ZN(n7741)
         );
  INV_X1 U9461 ( .A(n7732), .ZN(n7733) );
  NOR2_X1 U9462 ( .A1(n7733), .A2(n8476), .ZN(n7783) );
  AOI21_X1 U9463 ( .B1(n8518), .B2(n8533), .A(n7734), .ZN(n7737) );
  OR2_X1 U9464 ( .A1(n8516), .A2(n7735), .ZN(n7736) );
  OAI211_X1 U9465 ( .C1(n8520), .C2(n7738), .A(n7737), .B(n7736), .ZN(n7739)
         );
  AOI21_X1 U9466 ( .B1(n8482), .B2(n7783), .A(n7739), .ZN(n7740) );
  NAND2_X1 U9467 ( .A1(n7741), .A2(n7740), .ZN(P2_U3171) );
  INV_X1 U9468 ( .A(n7742), .ZN(n7745) );
  OAI222_X1 U9469 ( .A1(n9971), .A2(n7743), .B1(n9964), .B2(n7745), .C1(
        P1_U3086), .C2(n9454), .ZN(P1_U3333) );
  OAI222_X1 U9470 ( .A1(n7746), .A2(P2_U3151), .B1(n9023), .B2(n7745), .C1(
        n7744), .C2(n9013), .ZN(P2_U3273) );
  INV_X1 U9471 ( .A(n7747), .ZN(n8244) );
  XNOR2_X1 U9472 ( .A(n7748), .B(n8164), .ZN(n7837) );
  AOI22_X1 U9473 ( .A1(n8866), .A2(n8534), .B1(n8532), .B2(n8865), .ZN(n7752)
         );
  XNOR2_X1 U9474 ( .A(n7749), .B(n8164), .ZN(n7750) );
  NAND2_X1 U9475 ( .A1(n7750), .A2(n8862), .ZN(n7751) );
  OAI211_X1 U9476 ( .C1(n7837), .C2(n7753), .A(n7752), .B(n7751), .ZN(n7838)
         );
  NAND2_X1 U9477 ( .A1(n7838), .A2(n10161), .ZN(n7757) );
  OAI22_X1 U9478 ( .A1(n10161), .A2(n7754), .B1(n7889), .B2(n8854), .ZN(n7755)
         );
  AOI21_X1 U9479 ( .B1(n8849), .B2(n7869), .A(n7755), .ZN(n7756) );
  OAI211_X1 U9480 ( .C1(n7837), .C2(n7758), .A(n7757), .B(n7756), .ZN(P2_U3223) );
  OR2_X1 U9481 ( .A1(n9892), .A2(n9878), .ZN(n9380) );
  NAND2_X1 U9482 ( .A1(n9892), .A2(n9878), .ZN(n9377) );
  NAND2_X1 U9483 ( .A1(n9380), .A2(n9377), .ZN(n9305) );
  OR2_X1 U9484 ( .A1(n7760), .A2(n9474), .ZN(n7761) );
  XOR2_X1 U9485 ( .A(n9305), .B(n7787), .Z(n9894) );
  INV_X1 U9486 ( .A(n9305), .ZN(n7763) );
  NAND2_X2 U9487 ( .A1(n5129), .A2(n7763), .ZN(n7797) );
  OAI211_X1 U9488 ( .C1(n5129), .C2(n7763), .A(n10116), .B(n7797), .ZN(n7765)
         );
  AOI22_X1 U9489 ( .A1(n9754), .A2(n10105), .B1(n10104), .B2(n9474), .ZN(n7764) );
  NAND2_X1 U9490 ( .A1(n7765), .A2(n7764), .ZN(n9890) );
  INV_X1 U9491 ( .A(n9892), .ZN(n7769) );
  NOR2_X2 U9492 ( .A1(n7766), .A2(n9892), .ZN(n7789) );
  AOI211_X1 U9493 ( .C1(n9892), .C2(n7766), .A(n9750), .B(n7789), .ZN(n9891)
         );
  NAND2_X1 U9494 ( .A1(n9891), .A2(n10053), .ZN(n7768) );
  AOI22_X1 U9495 ( .A1(n10063), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9032), .B2(
        n10051), .ZN(n7767) );
  OAI211_X1 U9496 ( .C1(n7769), .C2(n9752), .A(n7768), .B(n7767), .ZN(n7770)
         );
  AOI21_X1 U9497 ( .B1(n10056), .B2(n9890), .A(n7770), .ZN(n7771) );
  OAI21_X1 U9498 ( .B1(n9894), .B2(n9767), .A(n7771), .ZN(P1_U3279) );
  NAND2_X1 U9499 ( .A1(n8239), .A2(n8234), .ZN(n8166) );
  XNOR2_X1 U9500 ( .A(n7772), .B(n8166), .ZN(n7773) );
  AOI222_X1 U9501 ( .A1(n8862), .A2(n7773), .B1(n8533), .B2(n8866), .C1(n8531), 
        .C2(n8865), .ZN(n7835) );
  NAND2_X1 U9502 ( .A1(n7774), .A2(n8250), .ZN(n7775) );
  INV_X1 U9503 ( .A(n8166), .ZN(n7866) );
  XNOR2_X1 U9504 ( .A(n7775), .B(n7866), .ZN(n7833) );
  NOR2_X1 U9505 ( .A1(n7776), .A2(n8856), .ZN(n7779) );
  OAI22_X1 U9506 ( .A1(n10161), .A2(n7777), .B1(n7934), .B2(n8854), .ZN(n7778)
         );
  AOI211_X1 U9507 ( .C1(n7833), .C2(n8872), .A(n7779), .B(n7778), .ZN(n7780)
         );
  OAI21_X1 U9508 ( .B1(n7835), .B2(n10163), .A(n7780), .ZN(P2_U3222) );
  INV_X1 U9509 ( .A(n7781), .ZN(n7784) );
  AOI211_X1 U9510 ( .C1(n7840), .C2(n7784), .A(n7783), .B(n7782), .ZN(n10179)
         );
  OR2_X1 U9511 ( .A1(n10179), .A2(n8884), .ZN(n7785) );
  OAI21_X1 U9512 ( .B1(n8928), .B2(n4655), .A(n7785), .ZN(P2_U3468) );
  NAND2_X1 U9513 ( .A1(n9892), .A2(n10106), .ZN(n7786) );
  XNOR2_X1 U9514 ( .A(n9527), .B(n9754), .ZN(n7798) );
  INV_X1 U9515 ( .A(n7798), .ZN(n9306) );
  XNOR2_X1 U9516 ( .A(n9528), .B(n9306), .ZN(n9885) );
  INV_X1 U9517 ( .A(n9751), .ZN(n7790) );
  AOI211_X1 U9518 ( .C1(n9527), .C2(n7791), .A(n9750), .B(n7790), .ZN(n9881)
         );
  NOR2_X1 U9519 ( .A1(n7788), .A2(n9752), .ZN(n7796) );
  NAND2_X1 U9520 ( .A1(n9755), .A2(n10106), .ZN(n7794) );
  INV_X1 U9521 ( .A(n9211), .ZN(n7792) );
  AOI22_X1 U9522 ( .A1(n10063), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7792), .B2(
        n10051), .ZN(n7793) );
  OAI211_X1 U9523 ( .C1(n9880), .C2(n9759), .A(n7794), .B(n7793), .ZN(n7795)
         );
  AOI211_X1 U9524 ( .C1(n9881), .C2(n10053), .A(n7796), .B(n7795), .ZN(n7800)
         );
  OAI21_X1 U9525 ( .B1(n4595), .B2(n7798), .A(n9270), .ZN(n9883) );
  NAND2_X1 U9526 ( .A1(n9883), .A2(n9764), .ZN(n7799) );
  OAI211_X1 U9527 ( .C1(n9885), .C2(n9767), .A(n7800), .B(n7799), .ZN(P1_U3278) );
  OAI21_X1 U9528 ( .B1(n7803), .B2(n7801), .A(n7802), .ZN(n7804) );
  NAND2_X1 U9529 ( .A1(n7804), .A2(n9206), .ZN(n7809) );
  AOI21_X1 U9530 ( .B1(n9215), .B2(n9477), .A(n7805), .ZN(n7806) );
  OAI21_X1 U9531 ( .B1(n9087), .B2(n9209), .A(n7806), .ZN(n7807) );
  AOI21_X1 U9532 ( .B1(n5122), .B2(n9210), .A(n7807), .ZN(n7808) );
  OAI211_X1 U9533 ( .C1(n7810), .C2(n9218), .A(n7809), .B(n7808), .ZN(P1_U3217) );
  NAND2_X1 U9534 ( .A1(n7814), .A2(n7811), .ZN(n7813) );
  NAND2_X1 U9535 ( .A1(n7812), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8359) );
  OAI211_X1 U9536 ( .C1(n10354), .C2(n9013), .A(n7813), .B(n8359), .ZN(
        P2_U3272) );
  NAND2_X1 U9537 ( .A1(n7814), .A2(n9959), .ZN(n7815) );
  OAI211_X1 U9538 ( .C1(n10438), .C2(n9971), .A(n7815), .B(n9466), .ZN(
        P1_U3332) );
  AOI21_X1 U9539 ( .B1(n5383), .B2(n7816), .A(n7908), .ZN(n7832) );
  NOR2_X1 U9540 ( .A1(n7818), .A2(n7823), .ZN(n7895) );
  AOI21_X1 U9541 ( .B1(n7819), .B2(n7777), .A(n7894), .ZN(n7828) );
  NAND2_X1 U9542 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3151), .ZN(n7931) );
  MUX2_X1 U9543 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8670), .Z(n7898) );
  XNOR2_X1 U9544 ( .A(n7898), .B(n7823), .ZN(n7824) );
  NAND2_X1 U9545 ( .A1(n7824), .A2(n7825), .ZN(n7899) );
  OAI21_X1 U9546 ( .B1(n7825), .B2(n7824), .A(n7899), .ZN(n7826) );
  NAND2_X1 U9547 ( .A1(n10136), .A2(n7826), .ZN(n7827) );
  OAI211_X1 U9548 ( .C1(n10129), .C2(n7828), .A(n7931), .B(n7827), .ZN(n7830)
         );
  NOR2_X1 U9549 ( .A1(n8706), .A2(n7910), .ZN(n7829) );
  AOI211_X1 U9550 ( .C1(n8704), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7830), .B(
        n7829), .ZN(n7831) );
  OAI21_X1 U9551 ( .B1(n7832), .B2(n8666), .A(n7831), .ZN(P2_U3193) );
  AOI22_X1 U9552 ( .A1(n7833), .A2(n8909), .B1(n8037), .B2(n8246), .ZN(n7834)
         );
  NAND2_X1 U9553 ( .A1(n7835), .A2(n7834), .ZN(n10579) );
  NAND2_X1 U9554 ( .A1(n10579), .A2(n8928), .ZN(n7836) );
  OAI21_X1 U9555 ( .B1(n8928), .B2(n5383), .A(n7836), .ZN(P2_U3470) );
  INV_X1 U9556 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7842) );
  INV_X1 U9557 ( .A(n7837), .ZN(n7839) );
  NOR2_X1 U9558 ( .A1(n7865), .A2(n8476), .ZN(n7891) );
  AOI211_X1 U9559 ( .C1(n7840), .C2(n7839), .A(n7891), .B(n7838), .ZN(n10180)
         );
  OR2_X1 U9560 ( .A1(n10180), .A2(n8884), .ZN(n7841) );
  OAI21_X1 U9561 ( .B1(n8928), .B2(n7842), .A(n7841), .ZN(P2_U3469) );
  XNOR2_X1 U9562 ( .A(n7843), .B(n8256), .ZN(n7856) );
  INV_X1 U9563 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7846) );
  XNOR2_X1 U9564 ( .A(n7844), .B(n8256), .ZN(n7845) );
  AOI222_X1 U9565 ( .A1(n8862), .A2(n7845), .B1(n8530), .B2(n8865), .C1(n8532), 
        .C2(n8866), .ZN(n7851) );
  MUX2_X1 U9566 ( .A(n7846), .B(n7851), .S(n10580), .Z(n7848) );
  NAND2_X1 U9567 ( .A1(n8995), .A2(n7882), .ZN(n7847) );
  OAI211_X1 U9568 ( .C1(n7856), .C2(n9003), .A(n7848), .B(n7847), .ZN(P2_U3426) );
  MUX2_X1 U9569 ( .A(n7911), .B(n7851), .S(n8928), .Z(n7850) );
  NAND2_X1 U9570 ( .A1(n8925), .A2(n7882), .ZN(n7849) );
  OAI211_X1 U9571 ( .C1(n7856), .C2(n8930), .A(n7850), .B(n7849), .ZN(P2_U3471) );
  MUX2_X1 U9572 ( .A(n7852), .B(n7851), .S(n10161), .Z(n7855) );
  INV_X1 U9573 ( .A(n7880), .ZN(n7853) );
  AOI22_X1 U9574 ( .A1(n7882), .A2(n8849), .B1(n10160), .B2(n7853), .ZN(n7854)
         );
  OAI211_X1 U9575 ( .C1(n7856), .C2(n8882), .A(n7855), .B(n7854), .ZN(P2_U3221) );
  INV_X1 U9576 ( .A(n6416), .ZN(n7859) );
  INV_X1 U9577 ( .A(n7857), .ZN(n8077) );
  OAI222_X1 U9578 ( .A1(n7859), .A2(P1_U3086), .B1(n9964), .B2(n8077), .C1(
        n7858), .C2(n9971), .ZN(P1_U3331) );
  XOR2_X1 U9579 ( .A(n8124), .B(n8166), .Z(n7930) );
  XNOR2_X1 U9580 ( .A(n7865), .B(n8124), .ZN(n7927) );
  AND2_X1 U9581 ( .A1(n7930), .A2(n7863), .ZN(n7864) );
  NOR3_X1 U9582 ( .A1(n7865), .A2(n8124), .A3(n7868), .ZN(n7867) );
  AOI211_X1 U9583 ( .C1(n8532), .C2(n8124), .A(n7867), .B(n7866), .ZN(n7872)
         );
  NOR3_X1 U9584 ( .A1(n7869), .A2(n7868), .A3(n7142), .ZN(n7870) );
  AOI211_X1 U9585 ( .C1(n7142), .C2(n8532), .A(n7870), .B(n8166), .ZN(n7871)
         );
  XNOR2_X1 U9586 ( .A(n7882), .B(n8124), .ZN(n7944) );
  XOR2_X1 U9587 ( .A(n7948), .B(n7944), .Z(n7874) );
  NAND2_X1 U9588 ( .A1(n7875), .A2(n7874), .ZN(n7946) );
  OAI211_X1 U9589 ( .C1(n7875), .C2(n7874), .A(n7946), .B(n8503), .ZN(n7884)
         );
  INV_X1 U9590 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7876) );
  NOR2_X1 U9591 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7876), .ZN(n7903) );
  AOI21_X1 U9592 ( .B1(n8518), .B2(n8530), .A(n7903), .ZN(n7879) );
  OR2_X1 U9593 ( .A1(n8516), .A2(n7877), .ZN(n7878) );
  OAI211_X1 U9594 ( .C1(n8520), .C2(n7880), .A(n7879), .B(n7878), .ZN(n7881)
         );
  AOI21_X1 U9595 ( .B1(n8527), .B2(n7882), .A(n7881), .ZN(n7883) );
  NAND2_X1 U9596 ( .A1(n7884), .A2(n7883), .ZN(P2_U3164) );
  XNOR2_X1 U9597 ( .A(n7926), .B(n8533), .ZN(n7928) );
  XOR2_X1 U9598 ( .A(n7927), .B(n7928), .Z(n7893) );
  AOI21_X1 U9599 ( .B1(n8518), .B2(n8532), .A(n7885), .ZN(n7888) );
  OR2_X1 U9600 ( .A1(n8516), .A2(n7886), .ZN(n7887) );
  OAI211_X1 U9601 ( .C1(n8520), .C2(n7889), .A(n7888), .B(n7887), .ZN(n7890)
         );
  AOI21_X1 U9602 ( .B1(n8482), .B2(n7891), .A(n7890), .ZN(n7892) );
  OAI21_X1 U9603 ( .B1(n7893), .B2(n8522), .A(n7892), .ZN(P2_U3157) );
  NOR2_X1 U9604 ( .A1(n7895), .A2(n7894), .ZN(n7897) );
  AOI22_X1 U9605 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7917), .B1(n8551), .B2(
        n7852), .ZN(n7896) );
  NOR2_X1 U9606 ( .A1(n7897), .A2(n7896), .ZN(n8542) );
  AOI21_X1 U9607 ( .B1(n7897), .B2(n7896), .A(n8542), .ZN(n7919) );
  MUX2_X1 U9608 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8670), .Z(n8545) );
  XNOR2_X1 U9609 ( .A(n8545), .B(n7917), .ZN(n7902) );
  OR2_X1 U9610 ( .A1(n7898), .A2(n7910), .ZN(n7900) );
  NAND2_X1 U9611 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  NAND2_X1 U9612 ( .A1(n7902), .A2(n7901), .ZN(n8546) );
  OAI21_X1 U9613 ( .B1(n7902), .B2(n7901), .A(n8546), .ZN(n7904) );
  AOI21_X1 U9614 ( .B1(n10136), .B2(n7904), .A(n7903), .ZN(n7905) );
  OAI21_X1 U9615 ( .B1(n10141), .B2(n7906), .A(n7905), .ZN(n7916) );
  INV_X1 U9616 ( .A(n7907), .ZN(n7909) );
  XNOR2_X1 U9617 ( .A(n7917), .B(n7911), .ZN(n7912) );
  AOI21_X1 U9618 ( .B1(n7913), .B2(n7912), .A(n8550), .ZN(n7914) );
  NOR2_X1 U9619 ( .A1(n7914), .A2(n8666), .ZN(n7915) );
  AOI211_X1 U9620 ( .C1(n10143), .C2(n7917), .A(n7916), .B(n7915), .ZN(n7918)
         );
  OAI21_X1 U9621 ( .B1(n7919), .B2(n10129), .A(n7918), .ZN(P2_U3194) );
  INV_X1 U9622 ( .A(n5808), .ZN(n7922) );
  INV_X1 U9623 ( .A(n7920), .ZN(n7924) );
  OAI222_X1 U9624 ( .A1(n7922), .A2(P2_U3151), .B1(n9023), .B2(n7924), .C1(
        n7921), .C2(n9013), .ZN(P2_U3270) );
  OAI222_X1 U9625 ( .A1(n7925), .A2(P1_U3086), .B1(n9964), .B2(n7924), .C1(
        n7923), .C2(n9971), .ZN(P1_U3330) );
  OAI22_X1 U9626 ( .A1(n7928), .A2(n7927), .B1(n8533), .B2(n7926), .ZN(n7929)
         );
  XOR2_X1 U9627 ( .A(n7930), .B(n7929), .Z(n7937) );
  OAI21_X1 U9628 ( .B1(n8508), .B2(n7948), .A(n7931), .ZN(n7932) );
  AOI21_X1 U9629 ( .B1(n8506), .B2(n8533), .A(n7932), .ZN(n7933) );
  OAI21_X1 U9630 ( .B1(n7934), .B2(n8520), .A(n7933), .ZN(n7935) );
  AOI21_X1 U9631 ( .B1(n8527), .B2(n8246), .A(n7935), .ZN(n7936) );
  OAI21_X1 U9632 ( .B1(n7937), .B2(n8522), .A(n7936), .ZN(P2_U3176) );
  INV_X1 U9633 ( .A(n7938), .ZN(n7940) );
  INV_X1 U9634 ( .A(n7939), .ZN(n7942) );
  OAI222_X1 U9635 ( .A1(n7940), .A2(P1_U3086), .B1(n9964), .B2(n7942), .C1(
        n10451), .C2(n9971), .ZN(P1_U3329) );
  OAI222_X1 U9636 ( .A1(n7943), .A2(P2_U3151), .B1(n9023), .B2(n7942), .C1(
        n7941), .C2(n9013), .ZN(P2_U3269) );
  NAND2_X1 U9637 ( .A1(n7946), .A2(n7945), .ZN(n7981) );
  XNOR2_X1 U9638 ( .A(n7966), .B(n8124), .ZN(n7978) );
  XNOR2_X1 U9639 ( .A(n7978), .B(n8530), .ZN(n7947) );
  XNOR2_X1 U9640 ( .A(n7981), .B(n7947), .ZN(n7953) );
  AND2_X1 U9641 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8556) );
  NOR2_X1 U9642 ( .A1(n8516), .A2(n7948), .ZN(n7949) );
  AOI211_X1 U9643 ( .C1(n8518), .C2(n8867), .A(n8556), .B(n7949), .ZN(n7950)
         );
  OAI21_X1 U9644 ( .B1(n7960), .B2(n8520), .A(n7950), .ZN(n7951) );
  AOI21_X1 U9645 ( .B1(n8527), .B2(n7966), .A(n7951), .ZN(n7952) );
  OAI21_X1 U9646 ( .B1(n7953), .B2(n8522), .A(n7952), .ZN(P2_U3174) );
  NAND2_X1 U9647 ( .A1(n8263), .A2(n8266), .ZN(n8168) );
  XNOR2_X1 U9648 ( .A(n7954), .B(n8168), .ZN(n7969) );
  INV_X1 U9649 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7957) );
  XOR2_X1 U9650 ( .A(n7955), .B(n8168), .Z(n7956) );
  AOI222_X1 U9651 ( .A1(n8862), .A2(n7956), .B1(n8531), .B2(n8866), .C1(n8867), 
        .C2(n8865), .ZN(n7965) );
  MUX2_X1 U9652 ( .A(n7957), .B(n7965), .S(n10580), .Z(n7959) );
  NAND2_X1 U9653 ( .A1(n8995), .A2(n7966), .ZN(n7958) );
  OAI211_X1 U9654 ( .C1(n7969), .C2(n9003), .A(n7959), .B(n7958), .ZN(P2_U3429) );
  INV_X1 U9655 ( .A(n7965), .ZN(n7962) );
  OAI22_X1 U9656 ( .A1(n8260), .A2(n8876), .B1(n7960), .B2(n8854), .ZN(n7961)
         );
  OAI21_X1 U9657 ( .B1(n7962), .B2(n7961), .A(n10161), .ZN(n7964) );
  NAND2_X1 U9658 ( .A1(n10163), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7963) );
  OAI211_X1 U9659 ( .C1(n7969), .C2(n8882), .A(n7964), .B(n7963), .ZN(P2_U3220) );
  MUX2_X1 U9660 ( .A(n8552), .B(n7965), .S(n8928), .Z(n7968) );
  NAND2_X1 U9661 ( .A1(n7966), .A2(n8925), .ZN(n7967) );
  OAI211_X1 U9662 ( .C1(n8930), .C2(n7969), .A(n7968), .B(n7967), .ZN(P2_U3472) );
  XNOR2_X1 U9663 ( .A(n7970), .B(n8268), .ZN(n8883) );
  INV_X1 U9664 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7973) );
  XNOR2_X1 U9665 ( .A(n7971), .B(n8268), .ZN(n7972) );
  AOI222_X1 U9666 ( .A1(n8862), .A2(n7972), .B1(n8530), .B2(n8866), .C1(n8844), 
        .C2(n8865), .ZN(n8875) );
  MUX2_X1 U9667 ( .A(n7973), .B(n8875), .S(n10580), .Z(n7975) );
  NAND2_X1 U9668 ( .A1(n7982), .A2(n8995), .ZN(n7974) );
  OAI211_X1 U9669 ( .C1(n8883), .C2(n9003), .A(n7975), .B(n7974), .ZN(P2_U3432) );
  MUX2_X1 U9670 ( .A(n8581), .B(n8875), .S(n8928), .Z(n7977) );
  NAND2_X1 U9671 ( .A1(n7982), .A2(n8925), .ZN(n7976) );
  OAI211_X1 U9672 ( .C1(n8930), .C2(n8883), .A(n7977), .B(n7976), .ZN(P2_U3473) );
  INV_X1 U9673 ( .A(n7982), .ZN(n8877) );
  INV_X1 U9674 ( .A(n8527), .ZN(n8513) );
  NAND2_X1 U9675 ( .A1(n7978), .A2(n8261), .ZN(n7980) );
  INV_X1 U9676 ( .A(n7978), .ZN(n7979) );
  XNOR2_X1 U9677 ( .A(n7982), .B(n8124), .ZN(n8092) );
  XOR2_X1 U9678 ( .A(n8515), .B(n8092), .Z(n7983) );
  OAI21_X1 U9679 ( .B1(n7984), .B2(n7983), .A(n8094), .ZN(n7985) );
  NAND2_X1 U9680 ( .A1(n7985), .A2(n8503), .ZN(n7991) );
  INV_X1 U9681 ( .A(n7986), .ZN(n8879) );
  NOR2_X1 U9682 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7987), .ZN(n8573) );
  AOI21_X1 U9683 ( .B1(n8518), .B2(n8844), .A(n8573), .ZN(n7988) );
  OAI21_X1 U9684 ( .B1(n8261), .B2(n8516), .A(n7988), .ZN(n7989) );
  AOI21_X1 U9685 ( .B1(n8879), .B2(n8510), .A(n7989), .ZN(n7990) );
  OAI211_X1 U9686 ( .C1(n8877), .C2(n8513), .A(n7991), .B(n7990), .ZN(P2_U3155) );
  INV_X1 U9687 ( .A(n7993), .ZN(n7996) );
  INV_X1 U9688 ( .A(n7994), .ZN(n7995) );
  NAND2_X1 U9689 ( .A1(n7996), .A2(n7995), .ZN(n7997) );
  INV_X1 U9690 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8362) );
  INV_X1 U9691 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9965) );
  MUX2_X1 U9692 ( .A(n8362), .B(n9965), .S(n7998), .Z(n8000) );
  INV_X1 U9693 ( .A(SI_30_), .ZN(n7999) );
  NAND2_X1 U9694 ( .A1(n8000), .A2(n7999), .ZN(n8003) );
  INV_X1 U9695 ( .A(n8000), .ZN(n8001) );
  NAND2_X1 U9696 ( .A1(n8001), .A2(SI_30_), .ZN(n8002) );
  NAND2_X1 U9697 ( .A1(n8003), .A2(n8002), .ZN(n8011) );
  MUX2_X1 U9698 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n8004), .Z(n8006) );
  INV_X1 U9699 ( .A(SI_31_), .ZN(n8005) );
  XNOR2_X1 U9700 ( .A(n8006), .B(n8005), .ZN(n8007) );
  NAND2_X1 U9701 ( .A1(n9960), .A2(n6024), .ZN(n8010) );
  OR2_X1 U9702 ( .A1(n8017), .A2(n10458), .ZN(n8009) );
  INV_X1 U9703 ( .A(n9898), .ZN(n9220) );
  NAND2_X1 U9704 ( .A1(n8012), .A2(n8011), .ZN(n8013) );
  NAND2_X1 U9705 ( .A1(n8014), .A2(n8013), .ZN(n8361) );
  NAND2_X1 U9706 ( .A1(n8361), .A2(n6024), .ZN(n8016) );
  OR2_X1 U9707 ( .A1(n8017), .A2(n9965), .ZN(n8015) );
  NOR2_X2 U9708 ( .A1(n9682), .A2(n9693), .ZN(n9681) );
  NAND2_X1 U9709 ( .A1(n9663), .A2(n9681), .ZN(n9651) );
  OR2_X1 U9710 ( .A1(n9651), .A2(n9655), .ZN(n9652) );
  OR2_X2 U9711 ( .A1(n9652), .A2(n9922), .ZN(n9635) );
  NAND2_X1 U9712 ( .A1(n9012), .A2(n6024), .ZN(n8019) );
  OR2_X1 U9713 ( .A1(n8017), .A2(n9968), .ZN(n8018) );
  NOR2_X2 U9714 ( .A1(n4534), .A2(n9777), .ZN(n9554) );
  NAND2_X1 U9715 ( .A1(n9902), .A2(n9554), .ZN(n9504) );
  XNOR2_X1 U9716 ( .A(n9220), .B(n9504), .ZN(n8020) );
  NOR2_X1 U9717 ( .A1(n8020), .A2(n9750), .ZN(n8026) );
  NAND2_X1 U9718 ( .A1(n8026), .A2(n10053), .ZN(n8025) );
  INV_X1 U9719 ( .A(P1_B_REG_SCAN_IN), .ZN(n8021) );
  NOR2_X1 U9720 ( .A1(n6541), .A2(n8021), .ZN(n8022) );
  NOR2_X1 U9721 ( .A1(n9879), .A2(n8022), .ZN(n9556) );
  INV_X1 U9722 ( .A(n9768), .ZN(n8023) );
  NOR2_X1 U9723 ( .A1(n10063), .A2(n8023), .ZN(n9509) );
  AOI21_X1 U9724 ( .B1(n10063), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9509), .ZN(
        n8024) );
  OAI211_X1 U9725 ( .C1(n9898), .C2(n9752), .A(n8025), .B(n8024), .ZN(P1_U3263) );
  NOR2_X1 U9726 ( .A1(n8026), .A2(n9768), .ZN(n9895) );
  MUX2_X1 U9727 ( .A(n8027), .B(n9895), .S(n10128), .Z(n8028) );
  OAI21_X1 U9728 ( .B1(n9898), .B2(n9889), .A(n8028), .ZN(P1_U3553) );
  NAND2_X1 U9729 ( .A1(n8029), .A2(n8703), .ZN(n8032) );
  AOI22_X1 U9730 ( .A1(n8032), .A2(n8031), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n8034) );
  OAI211_X1 U9731 ( .C1(n10141), .C2(n10366), .A(n8034), .B(n8033), .ZN(
        P2_U3182) );
  AOI22_X1 U9732 ( .A1(n8849), .A2(n8035), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10160), .ZN(n8042) );
  INV_X1 U9733 ( .A(n8036), .ZN(n8040) );
  NOR3_X1 U9734 ( .A1(n8156), .A2(n8038), .A3(n8037), .ZN(n8039) );
  OAI21_X1 U9735 ( .B1(n8040), .B2(n8039), .A(n10161), .ZN(n8041) );
  OAI211_X1 U9736 ( .C1(n10161), .C2(n10439), .A(n8042), .B(n8041), .ZN(
        P2_U3233) );
  NAND2_X1 U9737 ( .A1(n8043), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8046) );
  AOI22_X1 U9738 ( .A1(n8503), .A2(n8044), .B1(n8518), .B2(n8540), .ZN(n8045)
         );
  OAI211_X1 U9739 ( .C1(n8513), .C2(n8047), .A(n8046), .B(n8045), .ZN(P2_U3172) );
  XNOR2_X1 U9740 ( .A(n8048), .B(n6802), .ZN(n8060) );
  OAI211_X1 U9741 ( .C1(n8051), .C2(n8050), .A(n10136), .B(n8049), .ZN(n8052)
         );
  OAI21_X1 U9742 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n8053), .A(n8052), .ZN(n8059) );
  INV_X1 U9743 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10182) );
  NAND2_X1 U9744 ( .A1(n8054), .A2(n7110), .ZN(n8055) );
  AND2_X1 U9745 ( .A1(n8056), .A2(n8055), .ZN(n8057) );
  OAI22_X1 U9746 ( .A1(n10141), .A2(n10182), .B1(n10129), .B2(n8057), .ZN(
        n8058) );
  AOI211_X1 U9747 ( .C1(n10149), .C2(n8060), .A(n8059), .B(n8058), .ZN(n8061)
         );
  OAI21_X1 U9748 ( .B1(n8062), .B2(n8706), .A(n8061), .ZN(P2_U3183) );
  XNOR2_X1 U9749 ( .A(n8063), .B(n8190), .ZN(n8075) );
  INV_X1 U9750 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8066) );
  INV_X1 U9751 ( .A(n8190), .ZN(n8280) );
  XNOR2_X1 U9752 ( .A(n8064), .B(n8280), .ZN(n8065) );
  AOI222_X1 U9753 ( .A1(n8862), .A2(n8065), .B1(n8529), .B2(n8865), .C1(n8864), 
        .C2(n8866), .ZN(n8071) );
  MUX2_X1 U9754 ( .A(n8066), .B(n8071), .S(n10580), .Z(n8068) );
  NAND2_X1 U9755 ( .A1(n8441), .A2(n8995), .ZN(n8067) );
  OAI211_X1 U9756 ( .C1(n8075), .C2(n9003), .A(n8068), .B(n8067), .ZN(P2_U3441) );
  MUX2_X1 U9757 ( .A(n10346), .B(n8071), .S(n8928), .Z(n8070) );
  NAND2_X1 U9758 ( .A1(n8441), .A2(n8925), .ZN(n8069) );
  OAI211_X1 U9759 ( .C1(n8930), .C2(n8075), .A(n8070), .B(n8069), .ZN(P2_U3476) );
  MUX2_X1 U9760 ( .A(n8639), .B(n8071), .S(n10161), .Z(n8074) );
  INV_X1 U9761 ( .A(n8448), .ZN(n8072) );
  AOI22_X1 U9762 ( .A1(n8441), .A2(n8849), .B1(n10160), .B2(n8072), .ZN(n8073)
         );
  OAI211_X1 U9763 ( .C1(n8075), .C2(n8882), .A(n8074), .B(n8073), .ZN(P2_U3216) );
  OAI222_X1 U9764 ( .A1(n5812), .A2(P2_U3151), .B1(n9023), .B2(n8077), .C1(
        n8076), .C2(n9013), .ZN(P2_U3271) );
  INV_X1 U9765 ( .A(n8078), .ZN(n8296) );
  NAND2_X1 U9766 ( .A1(n8293), .A2(n8296), .ZN(n8171) );
  XNOR2_X1 U9767 ( .A(n8079), .B(n8171), .ZN(n8091) );
  XNOR2_X1 U9768 ( .A(n8080), .B(n8171), .ZN(n8081) );
  AOI222_X1 U9769 ( .A1(n8862), .A2(n8081), .B1(n8529), .B2(n8866), .C1(n8810), 
        .C2(n8865), .ZN(n8087) );
  MUX2_X1 U9770 ( .A(n8082), .B(n8087), .S(n10580), .Z(n8084) );
  NAND2_X1 U9771 ( .A1(n8393), .A2(n8995), .ZN(n8083) );
  OAI211_X1 U9772 ( .C1(n8091), .C2(n9003), .A(n8084), .B(n8083), .ZN(P2_U3446) );
  MUX2_X1 U9773 ( .A(n8692), .B(n8087), .S(n8928), .Z(n8086) );
  NAND2_X1 U9774 ( .A1(n8393), .A2(n8925), .ZN(n8085) );
  OAI211_X1 U9775 ( .C1(n8930), .C2(n8091), .A(n8086), .B(n8085), .ZN(P2_U3478) );
  MUX2_X1 U9776 ( .A(n8088), .B(n8087), .S(n10161), .Z(n8090) );
  AOI22_X1 U9777 ( .A1(n8393), .A2(n8849), .B1(n10160), .B2(n8402), .ZN(n8089)
         );
  OAI211_X1 U9778 ( .C1(n8091), .C2(n8882), .A(n8090), .B(n8089), .ZN(P2_U3214) );
  XNOR2_X1 U9779 ( .A(n8978), .B(n7142), .ZN(n8117) );
  NAND2_X1 U9780 ( .A1(n8092), .A2(n8515), .ZN(n8093) );
  XNOR2_X1 U9781 ( .A(n8853), .B(n8124), .ZN(n8097) );
  XNOR2_X1 U9782 ( .A(n8097), .B(n8436), .ZN(n8524) );
  INV_X1 U9783 ( .A(n8524), .ZN(n8095) );
  XNOR2_X1 U9784 ( .A(n8440), .B(n8124), .ZN(n8096) );
  NOR2_X1 U9785 ( .A1(n8096), .A2(n8864), .ZN(n8443) );
  AOI21_X1 U9786 ( .B1(n8096), .B2(n8864), .A(n8443), .ZN(n8431) );
  INV_X1 U9787 ( .A(n8097), .ZN(n8098) );
  NAND2_X1 U9788 ( .A1(n8098), .A2(n8844), .ZN(n8432) );
  INV_X1 U9789 ( .A(n8443), .ZN(n8100) );
  NAND2_X1 U9790 ( .A1(n8429), .A2(n8100), .ZN(n8105) );
  XNOR2_X1 U9791 ( .A(n8441), .B(n8124), .ZN(n8102) );
  NAND2_X1 U9792 ( .A1(n8102), .A2(n8101), .ZN(n8485) );
  INV_X1 U9793 ( .A(n8102), .ZN(n8103) );
  NAND2_X1 U9794 ( .A1(n8103), .A2(n8845), .ZN(n8104) );
  AND2_X1 U9795 ( .A1(n8485), .A2(n8104), .ZN(n8442) );
  NAND2_X1 U9796 ( .A1(n8105), .A2(n8442), .ZN(n8445) );
  NAND2_X1 U9797 ( .A1(n8445), .A2(n8485), .ZN(n8109) );
  XNOR2_X1 U9798 ( .A(n8497), .B(n7142), .ZN(n8106) );
  NAND2_X1 U9799 ( .A1(n8106), .A2(n8447), .ZN(n8395) );
  INV_X1 U9800 ( .A(n8106), .ZN(n8107) );
  NAND2_X1 U9801 ( .A1(n8107), .A2(n8529), .ZN(n8108) );
  AND2_X1 U9802 ( .A1(n8395), .A2(n8108), .ZN(n8486) );
  XNOR2_X1 U9803 ( .A(n8393), .B(n8124), .ZN(n8110) );
  NAND2_X1 U9804 ( .A1(n8110), .A2(n8492), .ZN(n8464) );
  INV_X1 U9805 ( .A(n8110), .ZN(n8111) );
  NAND2_X1 U9806 ( .A1(n8111), .A2(n8830), .ZN(n8112) );
  AND2_X1 U9807 ( .A1(n8464), .A2(n8112), .ZN(n8396) );
  XNOR2_X1 U9808 ( .A(n8984), .B(n8124), .ZN(n8113) );
  NAND2_X1 U9809 ( .A1(n8113), .A2(n8412), .ZN(n8406) );
  INV_X1 U9810 ( .A(n8113), .ZN(n8114) );
  NAND2_X1 U9811 ( .A1(n8114), .A2(n8810), .ZN(n8115) );
  AND2_X1 U9812 ( .A1(n8406), .A2(n8115), .ZN(n8465) );
  XNOR2_X1 U9813 ( .A(n8117), .B(n8116), .ZN(n8407) );
  XNOR2_X1 U9814 ( .A(n8801), .B(n8124), .ZN(n8118) );
  INV_X1 U9815 ( .A(n8475), .ZN(n8120) );
  XNOR2_X1 U9816 ( .A(n8788), .B(n8124), .ZN(n8374) );
  XNOR2_X1 U9817 ( .A(n8965), .B(n8124), .ZN(n8122) );
  NAND2_X1 U9818 ( .A1(n8122), .A2(n8425), .ZN(n8419) );
  OAI21_X1 U9819 ( .B1(n8122), .B2(n8425), .A(n8419), .ZN(n8456) );
  AOI21_X1 U9820 ( .B1(n8374), .B2(n8795), .A(n8456), .ZN(n8123) );
  XNOR2_X1 U9821 ( .A(n8959), .B(n8124), .ZN(n8125) );
  NAND2_X1 U9822 ( .A1(n8125), .A2(n8318), .ZN(n8498) );
  INV_X1 U9823 ( .A(n8125), .ZN(n8126) );
  NAND2_X1 U9824 ( .A1(n8126), .A2(n8770), .ZN(n8127) );
  NAND2_X1 U9825 ( .A1(n8422), .A2(n8498), .ZN(n8128) );
  XNOR2_X1 U9826 ( .A(n8953), .B(n7142), .ZN(n8129) );
  XNOR2_X1 U9827 ( .A(n8129), .B(n8367), .ZN(n8499) );
  INV_X1 U9828 ( .A(n8129), .ZN(n8130) );
  NAND2_X1 U9829 ( .A1(n8130), .A2(n8367), .ZN(n8131) );
  XNOR2_X1 U9830 ( .A(n8947), .B(n8124), .ZN(n8133) );
  XNOR2_X1 U9831 ( .A(n8133), .B(n8728), .ZN(n8364) );
  INV_X1 U9832 ( .A(n8133), .ZN(n8134) );
  NAND2_X1 U9833 ( .A1(n8134), .A2(n8749), .ZN(n8135) );
  NAND2_X1 U9834 ( .A1(n8365), .A2(n8135), .ZN(n8137) );
  XNOR2_X1 U9835 ( .A(n4540), .B(n8124), .ZN(n8136) );
  XNOR2_X1 U9836 ( .A(n8137), .B(n8136), .ZN(n8144) );
  INV_X1 U9837 ( .A(n8732), .ZN(n8141) );
  OAI22_X1 U9838 ( .A1(n8728), .A2(n8516), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8138), .ZN(n8139) );
  AOI21_X1 U9839 ( .B1(n8518), .B2(n8725), .A(n8139), .ZN(n8140) );
  OAI21_X1 U9840 ( .B1(n8141), .B2(n8520), .A(n8140), .ZN(n8142) );
  AOI21_X1 U9841 ( .B1(n8329), .B2(n8527), .A(n8142), .ZN(n8143) );
  OAI21_X1 U9842 ( .B1(n8144), .B2(n8522), .A(n8143), .ZN(P2_U3160) );
  NAND2_X1 U9843 ( .A1(n9960), .A2(n5331), .ZN(n8146) );
  INV_X1 U9844 ( .A(n8886), .ZN(n8933) );
  OR2_X1 U9845 ( .A1(n8933), .A2(n8147), .ZN(n8348) );
  INV_X1 U9846 ( .A(n8348), .ZN(n8177) );
  NAND2_X1 U9847 ( .A1(n8887), .A2(n8339), .ZN(n8180) );
  INV_X1 U9848 ( .A(n8187), .ZN(n8149) );
  INV_X1 U9849 ( .A(n8150), .ZN(n8311) );
  NAND2_X1 U9850 ( .A1(n4578), .A2(n8308), .ZN(n8781) );
  INV_X1 U9851 ( .A(n8151), .ZN(n8287) );
  NAND2_X1 U9852 ( .A1(n8287), .A2(n8283), .ZN(n8829) );
  INV_X1 U9853 ( .A(n8838), .ZN(n8285) );
  NAND2_X1 U9854 ( .A1(n8839), .A2(n8285), .ZN(n8852) );
  INV_X1 U9855 ( .A(n8152), .ZN(n8163) );
  INV_X1 U9856 ( .A(n8153), .ZN(n8154) );
  NOR2_X1 U9857 ( .A1(n7095), .A2(n8154), .ZN(n8157) );
  NAND4_X1 U9858 ( .A1(n4575), .A2(n8157), .A3(n8156), .A4(n8155), .ZN(n8161)
         );
  INV_X1 U9859 ( .A(n8228), .ZN(n8159) );
  NOR4_X1 U9860 ( .A1(n8161), .A2(n8160), .A3(n8159), .A4(n8158), .ZN(n8162)
         );
  NAND3_X1 U9861 ( .A1(n8164), .A2(n8163), .A3(n8162), .ZN(n8165) );
  NOR2_X1 U9862 ( .A1(n8166), .A2(n8165), .ZN(n8167) );
  NAND3_X1 U9863 ( .A1(n8168), .A2(n8256), .A3(n8167), .ZN(n8169) );
  OR4_X1 U9864 ( .A1(n8171), .A2(n8190), .A3(n8829), .A4(n8170), .ZN(n8172) );
  NOR3_X1 U9865 ( .A1(n8781), .A2(n8794), .A3(n8173), .ZN(n8174) );
  NAND3_X1 U9866 ( .A1(n8180), .A2(n8175), .A3(n4540), .ZN(n8176) );
  NOR4_X1 U9867 ( .A1(n8177), .A2(n8335), .A3(n8326), .A4(n8176), .ZN(n8184)
         );
  NOR2_X1 U9868 ( .A1(n8178), .A2(n8334), .ZN(n8182) );
  AND2_X1 U9869 ( .A1(n8933), .A2(n8335), .ZN(n8183) );
  MUX2_X1 U9870 ( .A(n8740), .B(n8329), .S(n8344), .Z(n8331) );
  MUX2_X1 U9871 ( .A(n5790), .B(n8187), .S(n8338), .Z(n8188) );
  OR2_X1 U9872 ( .A1(n8190), .A2(n8189), .ZN(n8282) );
  NAND2_X1 U9873 ( .A1(n8192), .A2(n8191), .ZN(n8197) );
  INV_X1 U9874 ( .A(n8199), .ZN(n8195) );
  NAND3_X1 U9875 ( .A1(n8198), .A2(n8193), .A3(n8344), .ZN(n8194) );
  OAI21_X1 U9876 ( .B1(n8195), .B2(n8197), .A(n8194), .ZN(n8196) );
  OAI21_X1 U9877 ( .B1(n8357), .B2(n8197), .A(n8196), .ZN(n8201) );
  MUX2_X1 U9878 ( .A(n8199), .B(n8198), .S(n8338), .Z(n8200) );
  NAND2_X1 U9879 ( .A1(n8211), .A2(n8202), .ZN(n8205) );
  NAND2_X1 U9880 ( .A1(n8219), .A2(n8203), .ZN(n8204) );
  MUX2_X1 U9881 ( .A(n8205), .B(n8204), .S(n8344), .Z(n8206) );
  INV_X1 U9882 ( .A(n8206), .ZN(n8207) );
  NAND2_X1 U9883 ( .A1(n8208), .A2(n8207), .ZN(n8210) );
  NAND2_X1 U9884 ( .A1(n8210), .A2(n8209), .ZN(n8224) );
  INV_X1 U9885 ( .A(n8211), .ZN(n8214) );
  OAI211_X1 U9886 ( .C1(n8224), .C2(n8214), .A(n8213), .B(n8212), .ZN(n8215)
         );
  NAND3_X1 U9887 ( .A1(n8215), .A2(n8221), .A3(n8227), .ZN(n8217) );
  INV_X1 U9888 ( .A(n8219), .ZN(n8223) );
  NAND2_X1 U9889 ( .A1(n8537), .A2(n8220), .ZN(n8222) );
  OAI211_X1 U9890 ( .C1(n8224), .C2(n8223), .A(n8222), .B(n8221), .ZN(n8226)
         );
  NAND2_X1 U9891 ( .A1(n8226), .A2(n8225), .ZN(n8229) );
  NAND2_X1 U9892 ( .A1(n8231), .A2(n8230), .ZN(n8232) );
  NAND3_X1 U9893 ( .A1(n8238), .A2(n8233), .A3(n8240), .ZN(n8235) );
  AND2_X1 U9894 ( .A1(n8234), .A2(n8338), .ZN(n8243) );
  NAND4_X1 U9895 ( .A1(n8235), .A2(n8243), .A3(n8250), .A4(n8236), .ZN(n8255)
         );
  AND2_X1 U9896 ( .A1(n8239), .A2(n8344), .ZN(n8242) );
  NAND4_X1 U9897 ( .A1(n8241), .A2(n8242), .A3(n8240), .A4(n8244), .ZN(n8254)
         );
  INV_X1 U9898 ( .A(n8242), .ZN(n8251) );
  AND2_X1 U9899 ( .A1(n8532), .A2(n8338), .ZN(n8247) );
  OAI21_X1 U9900 ( .B1(n8338), .B2(n8532), .A(n8246), .ZN(n8245) );
  OAI21_X1 U9901 ( .B1(n8247), .B2(n8246), .A(n8245), .ZN(n8248) );
  OAI211_X1 U9902 ( .C1(n8251), .C2(n8250), .A(n8249), .B(n8248), .ZN(n8252)
         );
  INV_X1 U9903 ( .A(n8252), .ZN(n8253) );
  MUX2_X1 U9904 ( .A(n8258), .B(n8257), .S(n8338), .Z(n8259) );
  MUX2_X1 U9905 ( .A(n8261), .B(n8260), .S(n8338), .Z(n8262) );
  OAI21_X1 U9906 ( .B1(n8264), .B2(n8263), .A(n8262), .ZN(n8265) );
  OAI21_X1 U9907 ( .B1(n8267), .B2(n8266), .A(n8265), .ZN(n8270) );
  INV_X1 U9908 ( .A(n8268), .ZN(n8269) );
  NAND2_X1 U9909 ( .A1(n8270), .A2(n8269), .ZN(n8274) );
  MUX2_X1 U9910 ( .A(n8272), .B(n8271), .S(n8338), .Z(n8273) );
  NAND2_X1 U9911 ( .A1(n8274), .A2(n8273), .ZN(n8275) );
  INV_X1 U9912 ( .A(n8852), .ZN(n8859) );
  NAND2_X1 U9913 ( .A1(n8275), .A2(n8859), .ZN(n8286) );
  NAND3_X1 U9914 ( .A1(n8286), .A2(n8839), .A3(n5126), .ZN(n8277) );
  NAND2_X1 U9915 ( .A1(n8277), .A2(n8276), .ZN(n8281) );
  NAND2_X1 U9916 ( .A1(n8283), .A2(n8278), .ZN(n8279) );
  NAND2_X1 U9917 ( .A1(n5126), .A2(n8344), .ZN(n8284) );
  AOI21_X1 U9918 ( .B1(n8286), .B2(n8285), .A(n8284), .ZN(n8289) );
  OAI211_X1 U9919 ( .C1(n8290), .C2(n8289), .A(n8288), .B(n8287), .ZN(n8291)
         );
  NAND3_X1 U9920 ( .A1(n8292), .A2(n8296), .A3(n8291), .ZN(n8297) );
  INV_X1 U9921 ( .A(n8819), .ZN(n8816) );
  NAND3_X1 U9922 ( .A1(n8297), .A2(n8816), .A3(n8293), .ZN(n8294) );
  NAND3_X1 U9923 ( .A1(n8297), .A2(n8296), .A3(n8295), .ZN(n8300) );
  NAND2_X1 U9924 ( .A1(n4578), .A2(n8303), .ZN(n8305) );
  INV_X1 U9925 ( .A(n8801), .ZN(n8477) );
  OAI21_X1 U9926 ( .B1(n8477), .B2(n8809), .A(n8308), .ZN(n8304) );
  MUX2_X1 U9927 ( .A(n8305), .B(n8304), .S(n8344), .Z(n8306) );
  NOR2_X1 U9928 ( .A1(n8775), .A2(n8306), .ZN(n8307) );
  NAND2_X1 U9929 ( .A1(n8311), .A2(n8308), .ZN(n8309) );
  NAND2_X1 U9930 ( .A1(n8309), .A2(n8310), .ZN(n8314) );
  NAND2_X1 U9931 ( .A1(n8310), .A2(n4578), .ZN(n8312) );
  NAND2_X1 U9932 ( .A1(n8312), .A2(n8311), .ZN(n8313) );
  MUX2_X1 U9933 ( .A(n8314), .B(n8313), .S(n8344), .Z(n8315) );
  NAND2_X1 U9934 ( .A1(n8316), .A2(n8315), .ZN(n8317) );
  NAND2_X1 U9935 ( .A1(n8959), .A2(n8318), .ZN(n8320) );
  MUX2_X1 U9936 ( .A(n8320), .B(n8319), .S(n8344), .Z(n8321) );
  INV_X1 U9937 ( .A(n8322), .ZN(n8325) );
  INV_X1 U9938 ( .A(n8323), .ZN(n8324) );
  MUX2_X1 U9939 ( .A(n8325), .B(n8324), .S(n8344), .Z(n8327) );
  NOR2_X1 U9940 ( .A1(n8343), .A2(n8329), .ZN(n8337) );
  INV_X1 U9941 ( .A(n8331), .ZN(n8332) );
  NOR2_X1 U9942 ( .A1(n8333), .A2(n8332), .ZN(n8345) );
  AOI21_X1 U9943 ( .B1(n8338), .B2(n8340), .A(n8940), .ZN(n8342) );
  INV_X1 U9944 ( .A(n8343), .ZN(n8347) );
  NAND2_X1 U9945 ( .A1(n5130), .A2(n8344), .ZN(n8346) );
  AOI211_X1 U9946 ( .C1(n8368), .C2(n8347), .A(n8346), .B(n8345), .ZN(n8349)
         );
  XNOR2_X1 U9947 ( .A(n8353), .B(n8352), .ZN(n8360) );
  NAND3_X1 U9948 ( .A1(n8355), .A2(n8354), .A3(n8670), .ZN(n8356) );
  OAI211_X1 U9949 ( .C1(n8357), .C2(n8359), .A(n8356), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8358) );
  OAI21_X1 U9950 ( .B1(n8360), .B2(n8359), .A(n8358), .ZN(P2_U3296) );
  INV_X1 U9951 ( .A(n8361), .ZN(n9963) );
  OAI222_X1 U9952 ( .A1(n8363), .A2(P2_U3151), .B1(n9023), .B2(n9963), .C1(
        n8362), .C2(n9013), .ZN(P2_U3265) );
  INV_X1 U9953 ( .A(n8947), .ZN(n8373) );
  NAND2_X1 U9954 ( .A1(n8366), .A2(n8365), .ZN(n8372) );
  NOR2_X1 U9955 ( .A1(n8367), .A2(n8516), .ZN(n8370) );
  INV_X1 U9956 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10389) );
  OAI22_X1 U9957 ( .A1(n8368), .A2(n8508), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10389), .ZN(n8369) );
  AOI211_X1 U9958 ( .C1(n8743), .C2(n8510), .A(n8370), .B(n8369), .ZN(n8371)
         );
  OAI211_X1 U9959 ( .C1(n8373), .C2(n8513), .A(n8372), .B(n8371), .ZN(P2_U3154) );
  NOR2_X1 U9960 ( .A1(n4536), .A2(n8374), .ZN(n8454) );
  AOI21_X1 U9961 ( .B1(n4536), .B2(n8374), .A(n8454), .ZN(n8375) );
  NAND2_X1 U9962 ( .A1(n8375), .A2(n8480), .ZN(n8457) );
  OAI21_X1 U9963 ( .B1(n8480), .B2(n8375), .A(n8457), .ZN(n8376) );
  NAND2_X1 U9964 ( .A1(n8376), .A2(n8503), .ZN(n8381) );
  INV_X1 U9965 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8377) );
  OAI22_X1 U9966 ( .A1(n8516), .A2(n8413), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8377), .ZN(n8379) );
  NOR2_X1 U9967 ( .A1(n8508), .A2(n8425), .ZN(n8378) );
  AOI211_X1 U9968 ( .C1(n8786), .C2(n8510), .A(n8379), .B(n8378), .ZN(n8380)
         );
  OAI211_X1 U9969 ( .C1(n8788), .C2(n8513), .A(n8381), .B(n8380), .ZN(P2_U3156) );
  OAI211_X1 U9970 ( .C1(n8384), .C2(n8383), .A(n8382), .B(n8503), .ZN(n8392)
         );
  INV_X1 U9971 ( .A(n8385), .ZN(n8386) );
  AOI21_X1 U9972 ( .B1(n8482), .B2(n8387), .A(n8386), .ZN(n8391) );
  AOI22_X1 U9973 ( .A1(n8506), .A2(n8539), .B1(n8518), .B2(n8537), .ZN(n8390)
         );
  NAND2_X1 U9974 ( .A1(n8510), .A2(n8388), .ZN(n8389) );
  NAND4_X1 U9975 ( .A1(n8392), .A2(n8391), .A3(n8390), .A4(n8389), .ZN(
        P2_U3158) );
  INV_X1 U9976 ( .A(n8393), .ZN(n8405) );
  INV_X1 U9977 ( .A(n8394), .ZN(n8489) );
  INV_X1 U9978 ( .A(n8395), .ZN(n8397) );
  NOR3_X1 U9979 ( .A1(n8489), .A2(n8397), .A3(n8396), .ZN(n8399) );
  INV_X1 U9980 ( .A(n8398), .ZN(n8466) );
  OAI21_X1 U9981 ( .B1(n8399), .B2(n8466), .A(n8503), .ZN(n8404) );
  NAND2_X1 U9982 ( .A1(n8518), .A2(n8810), .ZN(n8400) );
  NAND2_X1 U9983 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8702) );
  OAI211_X1 U9984 ( .C1(n8447), .C2(n8516), .A(n8400), .B(n8702), .ZN(n8401)
         );
  AOI21_X1 U9985 ( .B1(n8510), .B2(n8402), .A(n8401), .ZN(n8403) );
  OAI211_X1 U9986 ( .C1(n8405), .C2(n8513), .A(n8404), .B(n8403), .ZN(P2_U3159) );
  INV_X1 U9987 ( .A(n8978), .ZN(n8418) );
  NOR3_X1 U9988 ( .A1(n4537), .A2(n5097), .A3(n8407), .ZN(n8410) );
  INV_X1 U9989 ( .A(n8408), .ZN(n8409) );
  OAI21_X1 U9990 ( .B1(n8410), .B2(n8409), .A(n8503), .ZN(n8417) );
  INV_X1 U9991 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8411) );
  OAI22_X1 U9992 ( .A1(n8516), .A2(n8412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8411), .ZN(n8415) );
  NOR2_X1 U9993 ( .A1(n8508), .A2(n8413), .ZN(n8414) );
  AOI211_X1 U9994 ( .C1(n8813), .C2(n8510), .A(n8415), .B(n8414), .ZN(n8416)
         );
  OAI211_X1 U9995 ( .C1(n8418), .C2(n8513), .A(n8417), .B(n8416), .ZN(P2_U3163) );
  INV_X1 U9996 ( .A(n8959), .ZN(n8754) );
  INV_X1 U9997 ( .A(n8419), .ZN(n8421) );
  NOR3_X1 U9998 ( .A1(n4535), .A2(n8421), .A3(n8420), .ZN(n8423) );
  INV_X1 U9999 ( .A(n8422), .ZN(n8501) );
  OAI21_X1 U10000 ( .B1(n8423), .B2(n8501), .A(n8503), .ZN(n8428) );
  AOI22_X1 U10001 ( .A1(n8758), .A2(n8518), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8424) );
  OAI21_X1 U10002 ( .B1(n8425), .B2(n8516), .A(n8424), .ZN(n8426) );
  AOI21_X1 U10003 ( .B1(n8762), .B2(n8510), .A(n8426), .ZN(n8427) );
  OAI211_X1 U10004 ( .C1(n8754), .C2(n8513), .A(n8428), .B(n8427), .ZN(
        P2_U3165) );
  INV_X1 U10005 ( .A(n8429), .ZN(n8444) );
  AOI21_X1 U10006 ( .B1(n8430), .B2(n8432), .A(n8431), .ZN(n8433) );
  OAI21_X1 U10007 ( .B1(n8444), .B2(n8433), .A(n8503), .ZN(n8439) );
  INV_X1 U10008 ( .A(n8434), .ZN(n8848) );
  AND2_X1 U10009 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8620) );
  AOI21_X1 U10010 ( .B1(n8518), .B2(n8845), .A(n8620), .ZN(n8435) );
  OAI21_X1 U10011 ( .B1(n8436), .B2(n8516), .A(n8435), .ZN(n8437) );
  AOI21_X1 U10012 ( .B1(n8848), .B2(n8510), .A(n8437), .ZN(n8438) );
  OAI211_X1 U10013 ( .C1(n8440), .C2(n8513), .A(n8439), .B(n8438), .ZN(
        P2_U3166) );
  INV_X1 U10014 ( .A(n8441), .ZN(n8453) );
  NOR3_X1 U10015 ( .A1(n8444), .A2(n8443), .A3(n8442), .ZN(n8446) );
  INV_X1 U10016 ( .A(n8445), .ZN(n8488) );
  OAI21_X1 U10017 ( .B1(n8446), .B2(n8488), .A(n8503), .ZN(n8452) );
  NAND2_X1 U10018 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8649) );
  OAI21_X1 U10019 ( .B1(n8508), .B2(n8447), .A(n8649), .ZN(n8450) );
  NOR2_X1 U10020 ( .A1(n8520), .A2(n8448), .ZN(n8449) );
  AOI211_X1 U10021 ( .C1(n8506), .C2(n8864), .A(n8450), .B(n8449), .ZN(n8451)
         );
  OAI211_X1 U10022 ( .C1(n8453), .C2(n8513), .A(n8452), .B(n8451), .ZN(
        P2_U3168) );
  INV_X1 U10023 ( .A(n8965), .ZN(n8463) );
  INV_X1 U10024 ( .A(n8454), .ZN(n8455) );
  AND3_X1 U10025 ( .A1(n8457), .A2(n8456), .A3(n8455), .ZN(n8458) );
  AOI22_X1 U10026 ( .A1(n8518), .A2(n8770), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8459) );
  OAI21_X1 U10027 ( .B1(n8480), .B2(n8516), .A(n8459), .ZN(n8460) );
  AOI21_X1 U10028 ( .B1(n8772), .B2(n8510), .A(n8460), .ZN(n8461) );
  OAI211_X1 U10029 ( .C1(n8463), .C2(n8513), .A(n8462), .B(n8461), .ZN(
        P2_U3169) );
  INV_X1 U10030 ( .A(n8984), .ZN(n8472) );
  NOR3_X1 U10031 ( .A1(n8466), .A2(n5098), .A3(n8465), .ZN(n8467) );
  OAI21_X1 U10032 ( .B1(n8467), .B2(n4537), .A(n8503), .ZN(n8471) );
  AOI22_X1 U10033 ( .A1(n8518), .A2(n8821), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8468) );
  OAI21_X1 U10034 ( .B1(n8492), .B2(n8516), .A(n8468), .ZN(n8469) );
  AOI21_X1 U10035 ( .B1(n8824), .B2(n8510), .A(n8469), .ZN(n8470) );
  OAI211_X1 U10036 ( .C1(n8472), .C2(n8513), .A(n8471), .B(n8470), .ZN(
        P2_U3173) );
  INV_X1 U10037 ( .A(n8473), .ZN(n8474) );
  AOI21_X1 U10038 ( .B1(n8809), .B2(n8475), .A(n8474), .ZN(n8484) );
  NOR2_X1 U10039 ( .A1(n8477), .A2(n8476), .ZN(n8912) );
  NAND2_X1 U10040 ( .A1(n8510), .A2(n8797), .ZN(n8479) );
  AOI22_X1 U10041 ( .A1(n8506), .A2(n8821), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8478) );
  OAI211_X1 U10042 ( .C1(n8480), .C2(n8508), .A(n8479), .B(n8478), .ZN(n8481)
         );
  AOI21_X1 U10043 ( .B1(n8912), .B2(n8482), .A(n8481), .ZN(n8483) );
  OAI21_X1 U10044 ( .B1(n8484), .B2(n8522), .A(n8483), .ZN(P2_U3175) );
  INV_X1 U10045 ( .A(n8485), .ZN(n8487) );
  NOR3_X1 U10046 ( .A1(n8488), .A2(n8487), .A3(n8486), .ZN(n8490) );
  OAI21_X1 U10047 ( .B1(n8490), .B2(n8489), .A(n8503), .ZN(n8496) );
  NAND2_X1 U10048 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8676) );
  OAI21_X1 U10049 ( .B1(n8508), .B2(n8492), .A(n8676), .ZN(n8494) );
  NOR2_X1 U10050 ( .A1(n8520), .A2(n8833), .ZN(n8493) );
  AOI211_X1 U10051 ( .C1(n8506), .C2(n8845), .A(n8494), .B(n8493), .ZN(n8495)
         );
  OAI211_X1 U10052 ( .C1(n8497), .C2(n8513), .A(n8496), .B(n8495), .ZN(
        P2_U3178) );
  INV_X1 U10053 ( .A(n8953), .ZN(n8514) );
  INV_X1 U10054 ( .A(n8498), .ZN(n8500) );
  NOR3_X1 U10055 ( .A1(n8501), .A2(n8500), .A3(n8499), .ZN(n8505) );
  INV_X1 U10056 ( .A(n8502), .ZN(n8504) );
  OAI21_X1 U10057 ( .B1(n8505), .B2(n8504), .A(n8503), .ZN(n8512) );
  AOI22_X1 U10058 ( .A1(n8506), .A2(n8770), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8507) );
  OAI21_X1 U10059 ( .B1(n8728), .B2(n8508), .A(n8507), .ZN(n8509) );
  AOI21_X1 U10060 ( .B1(n8752), .B2(n8510), .A(n8509), .ZN(n8511) );
  OAI211_X1 U10061 ( .C1(n8514), .C2(n8513), .A(n8512), .B(n8511), .ZN(
        P2_U3180) );
  AND2_X1 U10062 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8602) );
  NOR2_X1 U10063 ( .A1(n8516), .A2(n8515), .ZN(n8517) );
  AOI211_X1 U10064 ( .C1(n8518), .C2(n8864), .A(n8602), .B(n8517), .ZN(n8519)
         );
  OAI21_X1 U10065 ( .B1(n8855), .B2(n8520), .A(n8519), .ZN(n8526) );
  INV_X1 U10066 ( .A(n8430), .ZN(n8521) );
  AOI211_X1 U10067 ( .C1(n8524), .C2(n8523), .A(n8522), .B(n8521), .ZN(n8525)
         );
  AOI211_X1 U10068 ( .C1(n8527), .C2(n8853), .A(n8526), .B(n8525), .ZN(n8528)
         );
  INV_X1 U10069 ( .A(n8528), .ZN(P2_U3181) );
  MUX2_X1 U10070 ( .A(n8340), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8679), .Z(
        P2_U3521) );
  MUX2_X1 U10071 ( .A(n8725), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8679), .Z(
        P2_U3520) );
  MUX2_X1 U10072 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8740), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10073 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8749), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10074 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8758), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10075 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8770), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10076 ( .A(n8783), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8679), .Z(
        P2_U3515) );
  MUX2_X1 U10077 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8795), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10078 ( .A(n8809), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8679), .Z(
        P2_U3513) );
  MUX2_X1 U10079 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8821), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10080 ( .A(n8810), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8679), .Z(
        P2_U3511) );
  MUX2_X1 U10081 ( .A(n8830), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8679), .Z(
        P2_U3510) );
  MUX2_X1 U10082 ( .A(n8529), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8679), .Z(
        P2_U3509) );
  MUX2_X1 U10083 ( .A(n8845), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8679), .Z(
        P2_U3508) );
  MUX2_X1 U10084 ( .A(n8864), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8679), .Z(
        P2_U3507) );
  MUX2_X1 U10085 ( .A(n8844), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8679), .Z(
        P2_U3506) );
  MUX2_X1 U10086 ( .A(n8867), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8679), .Z(
        P2_U3505) );
  MUX2_X1 U10087 ( .A(n8530), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8679), .Z(
        P2_U3504) );
  MUX2_X1 U10088 ( .A(n8531), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8679), .Z(
        P2_U3503) );
  MUX2_X1 U10089 ( .A(n8532), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8679), .Z(
        P2_U3502) );
  MUX2_X1 U10090 ( .A(n8533), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8679), .Z(
        P2_U3501) );
  MUX2_X1 U10091 ( .A(n8534), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8679), .Z(
        P2_U3500) );
  MUX2_X1 U10092 ( .A(n8535), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8679), .Z(
        P2_U3499) );
  MUX2_X1 U10093 ( .A(n8536), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8679), .Z(
        P2_U3497) );
  MUX2_X1 U10094 ( .A(n8537), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8679), .Z(
        P2_U3495) );
  MUX2_X1 U10095 ( .A(n8538), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8679), .Z(
        P2_U3494) );
  MUX2_X1 U10096 ( .A(n8539), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8679), .Z(
        P2_U3493) );
  MUX2_X1 U10097 ( .A(n8540), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8679), .Z(
        P2_U3492) );
  MUX2_X1 U10098 ( .A(n8541), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8679), .Z(
        P2_U3491) );
  AOI21_X1 U10099 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8551), .A(n8542), .ZN(
        n8562) );
  AOI21_X1 U10100 ( .B1(n8544), .B2(n8543), .A(n8563), .ZN(n8561) );
  MUX2_X1 U10101 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8670), .Z(n8567) );
  XNOR2_X1 U10102 ( .A(n8567), .B(n8578), .ZN(n8549) );
  OR2_X1 U10103 ( .A1(n8545), .A2(n8551), .ZN(n8547) );
  NAND2_X1 U10104 ( .A1(n8547), .A2(n8546), .ZN(n8548) );
  NAND2_X1 U10105 ( .A1(n8549), .A2(n8548), .ZN(n8569) );
  OAI21_X1 U10106 ( .B1(n8549), .B2(n8548), .A(n8569), .ZN(n8557) );
  AOI21_X1 U10107 ( .B1(n8553), .B2(n8552), .A(n8579), .ZN(n8554) );
  NOR2_X1 U10108 ( .A1(n8666), .A2(n8554), .ZN(n8555) );
  AOI211_X1 U10109 ( .C1(n10136), .C2(n8557), .A(n8556), .B(n8555), .ZN(n8558)
         );
  OAI21_X1 U10110 ( .B1(n10450), .B2(n10141), .A(n8558), .ZN(n8559) );
  AOI21_X1 U10111 ( .B1(n8578), .B2(n10143), .A(n8559), .ZN(n8560) );
  OAI21_X1 U10112 ( .B1(n8561), .B2(n10129), .A(n8560), .ZN(P2_U3195) );
  NOR2_X1 U10113 ( .A1(n8578), .A2(n8562), .ZN(n8564) );
  AOI22_X1 U10114 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8587), .B1(n8597), .B2(
        n8565), .ZN(n8566) );
  AOI21_X1 U10115 ( .B1(n4590), .B2(n8566), .A(n8590), .ZN(n8589) );
  MUX2_X1 U10116 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8670), .Z(n8592) );
  XNOR2_X1 U10117 ( .A(n8592), .B(n8587), .ZN(n8572) );
  INV_X1 U10118 ( .A(n8567), .ZN(n8568) );
  NAND2_X1 U10119 ( .A1(n8578), .A2(n8568), .ZN(n8570) );
  NAND2_X1 U10120 ( .A1(n8570), .A2(n8569), .ZN(n8571) );
  NAND2_X1 U10121 ( .A1(n8572), .A2(n8571), .ZN(n8593) );
  OAI21_X1 U10122 ( .B1(n8572), .B2(n8571), .A(n8593), .ZN(n8574) );
  AOI21_X1 U10123 ( .B1(n10136), .B2(n8574), .A(n8573), .ZN(n8575) );
  OAI21_X1 U10124 ( .B1(n10141), .B2(n8576), .A(n8575), .ZN(n8586) );
  NOR2_X1 U10125 ( .A1(n8578), .A2(n8577), .ZN(n8580) );
  XNOR2_X1 U10126 ( .A(n8587), .B(n8581), .ZN(n8582) );
  AOI21_X1 U10127 ( .B1(n8583), .B2(n8582), .A(n4591), .ZN(n8584) );
  NOR2_X1 U10128 ( .A1(n8584), .A2(n8666), .ZN(n8585) );
  AOI211_X1 U10129 ( .C1(n10143), .C2(n8587), .A(n8586), .B(n8585), .ZN(n8588)
         );
  OAI21_X1 U10130 ( .B1(n8589), .B2(n10129), .A(n8588), .ZN(P2_U3196) );
  NOR2_X1 U10131 ( .A1(n10421), .A2(n8591), .ZN(n8609) );
  AOI21_X1 U10132 ( .B1(n10421), .B2(n8591), .A(n8609), .ZN(n8607) );
  MUX2_X1 U10133 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8670), .Z(n8615) );
  XNOR2_X1 U10134 ( .A(n8625), .B(n8615), .ZN(n8596) );
  OR2_X1 U10135 ( .A1(n8592), .A2(n8597), .ZN(n8594) );
  NAND2_X1 U10136 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  NAND2_X1 U10137 ( .A1(n8596), .A2(n8595), .ZN(n8616) );
  OAI21_X1 U10138 ( .B1(n8596), .B2(n8595), .A(n8616), .ZN(n8603) );
  AOI21_X1 U10139 ( .B1(n8599), .B2(n8598), .A(n8626), .ZN(n8600) );
  NOR2_X1 U10140 ( .A1(n8666), .A2(n8600), .ZN(n8601) );
  AOI211_X1 U10141 ( .C1(n10136), .C2(n8603), .A(n8602), .B(n8601), .ZN(n8604)
         );
  OAI21_X1 U10142 ( .B1(n10485), .B2(n10141), .A(n8604), .ZN(n8605) );
  AOI21_X1 U10143 ( .B1(n8625), .B2(n10143), .A(n8605), .ZN(n8606) );
  OAI21_X1 U10144 ( .B1(n8607), .B2(n10129), .A(n8606), .ZN(P2_U3197) );
  NOR2_X1 U10145 ( .A1(n8625), .A2(n8608), .ZN(n8610) );
  NAND2_X1 U10146 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8641), .ZN(n8611) );
  OAI21_X1 U10147 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8641), .A(n8611), .ZN(
        n8612) );
  AOI21_X1 U10148 ( .B1(n8613), .B2(n8612), .A(n8635), .ZN(n8634) );
  MUX2_X1 U10149 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8670), .Z(n8642) );
  XNOR2_X1 U10150 ( .A(n8642), .B(n8632), .ZN(n8619) );
  OR2_X1 U10151 ( .A1(n8615), .A2(n8614), .ZN(n8617) );
  NAND2_X1 U10152 ( .A1(n8617), .A2(n8616), .ZN(n8618) );
  NAND2_X1 U10153 ( .A1(n8619), .A2(n8618), .ZN(n8643) );
  OAI21_X1 U10154 ( .B1(n8619), .B2(n8618), .A(n8643), .ZN(n8621) );
  AOI21_X1 U10155 ( .B1(n10136), .B2(n8621), .A(n8620), .ZN(n8622) );
  OAI21_X1 U10156 ( .B1(n10141), .B2(n8623), .A(n8622), .ZN(n8631) );
  XNOR2_X1 U10157 ( .A(n8641), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8627) );
  AOI21_X1 U10158 ( .B1(n8628), .B2(n8627), .A(n8637), .ZN(n8629) );
  NOR2_X1 U10159 ( .A1(n8629), .A2(n8666), .ZN(n8630) );
  AOI211_X1 U10160 ( .C1(n10143), .C2(n8632), .A(n8631), .B(n8630), .ZN(n8633)
         );
  OAI21_X1 U10161 ( .B1(n8634), .B2(n10129), .A(n8633), .ZN(P2_U3198) );
  AOI21_X1 U10162 ( .B1(n8639), .B2(n8636), .A(n8656), .ZN(n8654) );
  NOR2_X1 U10163 ( .A1(n10141), .A2(n10305), .ZN(n8652) );
  NOR2_X1 U10164 ( .A1(n10346), .A2(n8638), .ZN(n8662) );
  AOI21_X1 U10165 ( .B1(n8638), .B2(n10346), .A(n8662), .ZN(n8650) );
  MUX2_X1 U10166 ( .A(n8639), .B(n10346), .S(n8670), .Z(n8669) );
  XNOR2_X1 U10167 ( .A(n8669), .B(n8640), .ZN(n8646) );
  OR2_X1 U10168 ( .A1(n8642), .A2(n8641), .ZN(n8644) );
  OAI21_X1 U10169 ( .B1(n8646), .B2(n8645), .A(n8667), .ZN(n8647) );
  NAND2_X1 U10170 ( .A1(n10136), .A2(n8647), .ZN(n8648) );
  OAI211_X1 U10171 ( .C1(n8666), .C2(n8650), .A(n8649), .B(n8648), .ZN(n8651)
         );
  AOI211_X1 U10172 ( .C1(n10143), .C2(n8668), .A(n8652), .B(n8651), .ZN(n8653)
         );
  OAI21_X1 U10173 ( .B1(n8654), .B2(n10129), .A(n8653), .ZN(P2_U3199) );
  NOR2_X1 U10174 ( .A1(n8668), .A2(n8655), .ZN(n8657) );
  NAND2_X1 U10175 ( .A1(n8674), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8687) );
  OAI21_X1 U10176 ( .B1(n8674), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8687), .ZN(
        n8658) );
  NOR2_X1 U10177 ( .A1(n8668), .A2(n8660), .ZN(n8661) );
  NAND2_X1 U10178 ( .A1(n8674), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8689) );
  OAI21_X1 U10179 ( .B1(n8674), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8689), .ZN(
        n8663) );
  NOR2_X1 U10180 ( .A1(n8664), .A2(n8663), .ZN(n8691) );
  AOI21_X1 U10181 ( .B1(n8664), .B2(n8663), .A(n8691), .ZN(n8665) );
  INV_X1 U10182 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10190) );
  MUX2_X1 U10183 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8670), .Z(n8671) );
  NOR2_X1 U10184 ( .A1(n8672), .A2(n8671), .ZN(n8694) );
  INV_X1 U10185 ( .A(n8694), .ZN(n8673) );
  NAND2_X1 U10186 ( .A1(n8672), .A2(n8671), .ZN(n8695) );
  NAND2_X1 U10187 ( .A1(n8673), .A2(n8695), .ZN(n8678) );
  NAND3_X1 U10188 ( .A1(n10136), .A2(n8674), .A3(n8678), .ZN(n8675) );
  OAI211_X1 U10189 ( .C1(n10141), .C2(n10190), .A(n8676), .B(n8675), .ZN(n8677) );
  INV_X1 U10190 ( .A(n8677), .ZN(n8682) );
  OAI21_X1 U10191 ( .B1(n8679), .B2(n8678), .A(n8706), .ZN(n8680) );
  NAND2_X1 U10192 ( .A1(n8682), .A2(n8681), .ZN(n8683) );
  OAI21_X1 U10193 ( .B1(n8686), .B2(n10129), .A(n8685), .ZN(P2_U3200) );
  INV_X1 U10194 ( .A(n8687), .ZN(n8688) );
  MUX2_X1 U10195 ( .A(n8088), .B(P2_REG2_REG_19__SCAN_IN), .S(n8693), .Z(n8699) );
  INV_X1 U10196 ( .A(n8689), .ZN(n8690) );
  XNOR2_X1 U10197 ( .A(n8693), .B(n8692), .ZN(n8697) );
  INV_X1 U10198 ( .A(n8697), .ZN(n8700) );
  MUX2_X1 U10199 ( .A(n8700), .B(n8699), .S(n8698), .Z(n8701) );
  OAI21_X1 U10200 ( .B1(n8352), .B2(n8706), .A(n8705), .ZN(n8707) );
  INV_X1 U10201 ( .A(n8708), .ZN(n8709) );
  NAND2_X1 U10202 ( .A1(n8710), .A2(n8709), .ZN(n8934) );
  INV_X1 U10203 ( .A(n8711), .ZN(n8712) );
  NAND2_X1 U10204 ( .A1(n8712), .A2(n10160), .ZN(n8718) );
  OAI21_X1 U10205 ( .B1(n10163), .B2(n8934), .A(n8718), .ZN(n8714) );
  AOI21_X1 U10206 ( .B1(n10163), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8714), .ZN(
        n8713) );
  OAI21_X1 U10207 ( .B1(n8886), .B2(n8856), .A(n8713), .ZN(P2_U3202) );
  AOI21_X1 U10208 ( .B1(n10163), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8714), .ZN(
        n8715) );
  OAI21_X1 U10209 ( .B1(n8940), .B2(n8856), .A(n8715), .ZN(P2_U3203) );
  INV_X1 U10210 ( .A(n8716), .ZN(n8723) );
  NAND2_X1 U10211 ( .A1(n10163), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8717) );
  OAI211_X1 U10212 ( .C1(n8719), .C2(n8856), .A(n8718), .B(n8717), .ZN(n8720)
         );
  AOI21_X1 U10213 ( .B1(n8721), .B2(n8872), .A(n8720), .ZN(n8722) );
  OAI21_X1 U10214 ( .B1(n8723), .B2(n10163), .A(n8722), .ZN(P2_U3204) );
  XNOR2_X1 U10215 ( .A(n8724), .B(n4540), .ZN(n8730) );
  NAND2_X1 U10216 ( .A1(n8725), .A2(n8865), .ZN(n8726) );
  OAI21_X1 U10217 ( .B1(n8728), .B2(n8727), .A(n8726), .ZN(n8729) );
  XNOR2_X1 U10218 ( .A(n8731), .B(n4540), .ZN(n8892) );
  AOI22_X1 U10219 ( .A1(n10163), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8732), 
        .B2(n10160), .ZN(n8733) );
  OAI21_X1 U10220 ( .B1(n8944), .B2(n8856), .A(n8733), .ZN(n8734) );
  AOI21_X1 U10221 ( .B1(n8892), .B2(n8872), .A(n8734), .ZN(n8735) );
  OAI21_X1 U10222 ( .B1(n8894), .B2(n10163), .A(n8735), .ZN(P2_U3205) );
  OAI21_X1 U10223 ( .B1(n4549), .B2(n8737), .A(n8736), .ZN(n8950) );
  INV_X1 U10224 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8742) );
  XNOR2_X1 U10225 ( .A(n8739), .B(n8738), .ZN(n8741) );
  AOI222_X1 U10226 ( .A1(n8862), .A2(n8741), .B1(n8758), .B2(n8866), .C1(n8740), .C2(n8865), .ZN(n8945) );
  MUX2_X1 U10227 ( .A(n8742), .B(n8945), .S(n10161), .Z(n8745) );
  AOI22_X1 U10228 ( .A1(n8947), .A2(n8849), .B1(n10160), .B2(n8743), .ZN(n8744) );
  OAI211_X1 U10229 ( .C1(n8950), .C2(n8882), .A(n8745), .B(n8744), .ZN(
        P2_U3206) );
  XNOR2_X1 U10230 ( .A(n8746), .B(n8748), .ZN(n8956) );
  XOR2_X1 U10231 ( .A(n8748), .B(n8747), .Z(n8750) );
  AOI222_X1 U10232 ( .A1(n8862), .A2(n8750), .B1(n8770), .B2(n8866), .C1(n8749), .C2(n8865), .ZN(n8951) );
  AOI22_X1 U10233 ( .A1(n8953), .A2(n8849), .B1(n10160), .B2(n8752), .ZN(n8753) );
  NOR2_X1 U10234 ( .A1(n8754), .A2(n8876), .ZN(n8761) );
  OAI21_X1 U10235 ( .B1(n8757), .B2(n8756), .A(n8755), .ZN(n8759) );
  AOI222_X1 U10236 ( .A1(n8862), .A2(n8759), .B1(n8783), .B2(n8866), .C1(n8758), .C2(n8865), .ZN(n8957) );
  INV_X1 U10237 ( .A(n8957), .ZN(n8760) );
  AOI211_X1 U10238 ( .C1(n10160), .C2(n8762), .A(n8761), .B(n8760), .ZN(n8768)
         );
  OAI21_X1 U10239 ( .B1(n8765), .B2(n8764), .A(n8763), .ZN(n8962) );
  INV_X1 U10240 ( .A(n8962), .ZN(n8766) );
  AOI22_X1 U10241 ( .A1(n8766), .A2(n8872), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10163), .ZN(n8767) );
  OAI21_X1 U10242 ( .B1(n8768), .B2(n10163), .A(n8767), .ZN(P2_U3208) );
  XNOR2_X1 U10243 ( .A(n8769), .B(n8775), .ZN(n8771) );
  AOI222_X1 U10244 ( .A1(n8862), .A2(n8771), .B1(n8795), .B2(n8866), .C1(n8770), .C2(n8865), .ZN(n8963) );
  INV_X1 U10245 ( .A(n8876), .ZN(n8773) );
  AOI22_X1 U10246 ( .A1(n8965), .A2(n8773), .B1(n10160), .B2(n8772), .ZN(n8774) );
  AOI21_X1 U10247 ( .B1(n8963), .B2(n8774), .A(n10163), .ZN(n8779) );
  XNOR2_X1 U10248 ( .A(n8776), .B(n8775), .ZN(n8968) );
  INV_X1 U10249 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8777) );
  OAI22_X1 U10250 ( .A1(n8968), .A2(n8882), .B1(n8777), .B2(n10161), .ZN(n8778) );
  OR2_X1 U10251 ( .A1(n8779), .A2(n8778), .ZN(P2_U3209) );
  XOR2_X1 U10252 ( .A(n8781), .B(n8780), .Z(n8974) );
  XNOR2_X1 U10253 ( .A(n8782), .B(n8781), .ZN(n8784) );
  AOI222_X1 U10254 ( .A1(n8862), .A2(n8784), .B1(n8809), .B2(n8866), .C1(n8783), .C2(n8865), .ZN(n8969) );
  MUX2_X1 U10255 ( .A(n8785), .B(n8969), .S(n10161), .Z(n8791) );
  INV_X1 U10256 ( .A(n8786), .ZN(n8787) );
  OAI22_X1 U10257 ( .A1(n8788), .A2(n8856), .B1(n8787), .B2(n8854), .ZN(n8789)
         );
  INV_X1 U10258 ( .A(n8789), .ZN(n8790) );
  OAI211_X1 U10259 ( .C1(n8974), .C2(n8882), .A(n8791), .B(n8790), .ZN(
        P2_U3210) );
  OAI21_X1 U10260 ( .B1(n8794), .B2(n8793), .A(n8792), .ZN(n8796) );
  AOI222_X1 U10261 ( .A1(n8862), .A2(n8796), .B1(n8821), .B2(n8866), .C1(n8795), .C2(n8865), .ZN(n8915) );
  INV_X1 U10262 ( .A(n8797), .ZN(n8798) );
  OAI22_X1 U10263 ( .A1(n10161), .A2(n8799), .B1(n8798), .B2(n8854), .ZN(n8800) );
  AOI21_X1 U10264 ( .B1(n8801), .B2(n8849), .A(n8800), .ZN(n8805) );
  OR2_X1 U10265 ( .A1(n8803), .A2(n8802), .ZN(n8911) );
  NAND3_X1 U10266 ( .A1(n8911), .A2(n8872), .A3(n8910), .ZN(n8804) );
  OAI211_X1 U10267 ( .C1(n8915), .C2(n10163), .A(n8805), .B(n8804), .ZN(
        P2_U3211) );
  XNOR2_X1 U10268 ( .A(n8806), .B(n8807), .ZN(n8981) );
  INV_X1 U10269 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8812) );
  XNOR2_X1 U10270 ( .A(n8808), .B(n8807), .ZN(n8811) );
  AOI222_X1 U10271 ( .A1(n8862), .A2(n8811), .B1(n8810), .B2(n8866), .C1(n8809), .C2(n8865), .ZN(n8976) );
  MUX2_X1 U10272 ( .A(n8812), .B(n8976), .S(n10161), .Z(n8815) );
  AOI22_X1 U10273 ( .A1(n8978), .A2(n8849), .B1(n10160), .B2(n8813), .ZN(n8814) );
  OAI211_X1 U10274 ( .C1(n8981), .C2(n8882), .A(n8815), .B(n8814), .ZN(
        P2_U3212) );
  XNOR2_X1 U10275 ( .A(n8817), .B(n8816), .ZN(n8987) );
  INV_X1 U10276 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8823) );
  OAI21_X1 U10277 ( .B1(n8820), .B2(n8819), .A(n8818), .ZN(n8822) );
  AOI222_X1 U10278 ( .A1(n8862), .A2(n8822), .B1(n8821), .B2(n8865), .C1(n8830), .C2(n8866), .ZN(n8982) );
  MUX2_X1 U10279 ( .A(n8823), .B(n8982), .S(n10161), .Z(n8826) );
  AOI22_X1 U10280 ( .A1(n8984), .A2(n8849), .B1(n10160), .B2(n8824), .ZN(n8825) );
  OAI211_X1 U10281 ( .C1(n8987), .C2(n8882), .A(n8826), .B(n8825), .ZN(
        P2_U3213) );
  XOR2_X1 U10282 ( .A(n8829), .B(n8827), .Z(n8992) );
  XOR2_X1 U10283 ( .A(n8828), .B(n8829), .Z(n8831) );
  AOI222_X1 U10284 ( .A1(n8862), .A2(n8831), .B1(n8845), .B2(n8866), .C1(n8830), .C2(n8865), .ZN(n8988) );
  MUX2_X1 U10285 ( .A(n8832), .B(n8988), .S(n10161), .Z(n8836) );
  INV_X1 U10286 ( .A(n8833), .ZN(n8834) );
  AOI22_X1 U10287 ( .A1(n8989), .A2(n8849), .B1(n10160), .B2(n8834), .ZN(n8835) );
  OAI211_X1 U10288 ( .C1(n8992), .C2(n8882), .A(n8836), .B(n8835), .ZN(
        P2_U3215) );
  OR2_X1 U10289 ( .A1(n8837), .A2(n8838), .ZN(n8840) );
  NAND2_X1 U10290 ( .A1(n8840), .A2(n8839), .ZN(n8841) );
  XOR2_X1 U10291 ( .A(n8842), .B(n8841), .Z(n8999) );
  XOR2_X1 U10292 ( .A(n8843), .B(n8842), .Z(n8846) );
  AOI222_X1 U10293 ( .A1(n8862), .A2(n8846), .B1(n8845), .B2(n8865), .C1(n8844), .C2(n8866), .ZN(n8993) );
  MUX2_X1 U10294 ( .A(n8847), .B(n8993), .S(n10161), .Z(n8851) );
  AOI22_X1 U10295 ( .A1(n8996), .A2(n8849), .B1(n10160), .B2(n8848), .ZN(n8850) );
  OAI211_X1 U10296 ( .C1(n8999), .C2(n8882), .A(n8851), .B(n8850), .ZN(
        P2_U3217) );
  XNOR2_X1 U10297 ( .A(n8837), .B(n8852), .ZN(n9004) );
  INV_X1 U10298 ( .A(n9004), .ZN(n8873) );
  INV_X1 U10299 ( .A(n8853), .ZN(n9002) );
  OAI22_X1 U10300 ( .A1(n9002), .A2(n8856), .B1(n8855), .B2(n8854), .ZN(n8871)
         );
  INV_X1 U10301 ( .A(n8858), .ZN(n8860) );
  NAND2_X1 U10302 ( .A1(n8860), .A2(n8859), .ZN(n8861) );
  OAI211_X1 U10303 ( .C1(n8863), .C2(n4977), .A(n8862), .B(n8861), .ZN(n8869)
         );
  AOI22_X1 U10304 ( .A1(n8867), .A2(n8866), .B1(n8865), .B2(n8864), .ZN(n8868)
         );
  NAND2_X1 U10305 ( .A1(n8869), .A2(n8868), .ZN(n9000) );
  MUX2_X1 U10306 ( .A(P2_REG2_REG_15__SCAN_IN), .B(n9000), .S(n10161), .Z(
        n8870) );
  AOI211_X1 U10307 ( .C1(n8873), .C2(n8872), .A(n8871), .B(n8870), .ZN(n8874)
         );
  INV_X1 U10308 ( .A(n8874), .ZN(P2_U3218) );
  OAI21_X1 U10309 ( .B1(n8877), .B2(n8876), .A(n8875), .ZN(n8878) );
  NAND2_X1 U10310 ( .A1(n8878), .A2(n10161), .ZN(n8881) );
  AOI22_X1 U10311 ( .A1(n10163), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n10160), 
        .B2(n8879), .ZN(n8880) );
  OAI211_X1 U10312 ( .C1(n8883), .C2(n8882), .A(n8881), .B(n8880), .ZN(
        P2_U3219) );
  NOR2_X1 U10313 ( .A1(n8934), .A2(n8884), .ZN(n8888) );
  AOI21_X1 U10314 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n8884), .A(n8888), .ZN(
        n8885) );
  OAI21_X1 U10315 ( .B1(n8886), .B2(n8929), .A(n8885), .ZN(P2_U3490) );
  INV_X1 U10316 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U10317 ( .A1(n8887), .A2(n8925), .ZN(n8890) );
  INV_X1 U10318 ( .A(n8888), .ZN(n8889) );
  OAI211_X1 U10319 ( .C1(n8928), .C2(n8891), .A(n8890), .B(n8889), .ZN(
        P2_U3489) );
  NAND2_X1 U10320 ( .A1(n8892), .A2(n8909), .ZN(n8893) );
  NAND2_X1 U10321 ( .A1(n8894), .A2(n8893), .ZN(n8941) );
  INV_X1 U10322 ( .A(n8895), .ZN(n8896) );
  OAI21_X1 U10323 ( .B1(n8944), .B2(n8929), .A(n8896), .ZN(P2_U3487) );
  MUX2_X1 U10324 ( .A(n10399), .B(n8945), .S(n8928), .Z(n8898) );
  NAND2_X1 U10325 ( .A1(n8947), .A2(n8925), .ZN(n8897) );
  OAI211_X1 U10326 ( .C1(n8950), .C2(n8930), .A(n8898), .B(n8897), .ZN(
        P2_U3486) );
  INV_X1 U10327 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8899) );
  MUX2_X1 U10328 ( .A(n8899), .B(n8951), .S(n8928), .Z(n8901) );
  NAND2_X1 U10329 ( .A1(n8953), .A2(n8925), .ZN(n8900) );
  OAI211_X1 U10330 ( .C1(n8956), .C2(n8930), .A(n8901), .B(n8900), .ZN(
        P2_U3485) );
  MUX2_X1 U10331 ( .A(n10400), .B(n8957), .S(n8928), .Z(n8903) );
  NAND2_X1 U10332 ( .A1(n8959), .A2(n8925), .ZN(n8902) );
  OAI211_X1 U10333 ( .C1(n8930), .C2(n8962), .A(n8903), .B(n8902), .ZN(
        P2_U3484) );
  MUX2_X1 U10334 ( .A(n10295), .B(n8963), .S(n8928), .Z(n8905) );
  NAND2_X1 U10335 ( .A1(n8965), .A2(n8925), .ZN(n8904) );
  OAI211_X1 U10336 ( .C1(n8930), .C2(n8968), .A(n8905), .B(n8904), .ZN(
        P2_U3483) );
  INV_X1 U10337 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8906) );
  MUX2_X1 U10338 ( .A(n8906), .B(n8969), .S(n8928), .Z(n8908) );
  NAND2_X1 U10339 ( .A1(n8971), .A2(n8925), .ZN(n8907) );
  OAI211_X1 U10340 ( .C1(n8974), .C2(n8930), .A(n8908), .B(n8907), .ZN(
        P2_U3482) );
  NAND3_X1 U10341 ( .A1(n8911), .A2(n8910), .A3(n8909), .ZN(n8914) );
  INV_X1 U10342 ( .A(n8912), .ZN(n8913) );
  NAND3_X1 U10343 ( .A1(n8915), .A2(n8914), .A3(n8913), .ZN(n8975) );
  MUX2_X1 U10344 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8975), .S(n8928), .Z(
        P2_U3481) );
  INV_X1 U10345 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8916) );
  MUX2_X1 U10346 ( .A(n8916), .B(n8976), .S(n8928), .Z(n8918) );
  NAND2_X1 U10347 ( .A1(n8978), .A2(n8925), .ZN(n8917) );
  OAI211_X1 U10348 ( .C1(n8930), .C2(n8981), .A(n8918), .B(n8917), .ZN(
        P2_U3480) );
  INV_X1 U10349 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8919) );
  MUX2_X1 U10350 ( .A(n8919), .B(n8982), .S(n8928), .Z(n8921) );
  NAND2_X1 U10351 ( .A1(n8984), .A2(n8925), .ZN(n8920) );
  OAI211_X1 U10352 ( .C1(n8987), .C2(n8930), .A(n8921), .B(n8920), .ZN(
        P2_U3479) );
  MUX2_X1 U10353 ( .A(n8922), .B(n8988), .S(n8928), .Z(n8924) );
  NAND2_X1 U10354 ( .A1(n8989), .A2(n8925), .ZN(n8923) );
  OAI211_X1 U10355 ( .C1(n8992), .C2(n8930), .A(n8924), .B(n8923), .ZN(
        P2_U3477) );
  MUX2_X1 U10356 ( .A(n10489), .B(n8993), .S(n8928), .Z(n8927) );
  NAND2_X1 U10357 ( .A1(n8996), .A2(n8925), .ZN(n8926) );
  OAI211_X1 U10358 ( .C1(n8999), .C2(n8930), .A(n8927), .B(n8926), .ZN(
        P2_U3475) );
  MUX2_X1 U10359 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9000), .S(n8928), .Z(n8932) );
  OAI22_X1 U10360 ( .A1(n9004), .A2(n8930), .B1(n9002), .B2(n8929), .ZN(n8931)
         );
  OR2_X1 U10361 ( .A1(n8932), .A2(n8931), .ZN(P2_U3474) );
  INV_X1 U10362 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U10363 ( .A1(n8933), .A2(n8995), .ZN(n8936) );
  INV_X1 U10364 ( .A(n8934), .ZN(n8935) );
  NAND2_X1 U10365 ( .A1(n8935), .A2(n10580), .ZN(n8938) );
  OAI211_X1 U10366 ( .C1(n8937), .C2(n10580), .A(n8936), .B(n8938), .ZN(
        P2_U3458) );
  NAND2_X1 U10367 ( .A1(n10578), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8939) );
  OAI211_X1 U10368 ( .C1(n8940), .C2(n9001), .A(n8939), .B(n8938), .ZN(
        P2_U3457) );
  INV_X1 U10369 ( .A(n8942), .ZN(n8943) );
  OAI21_X1 U10370 ( .B1(n8944), .B2(n9001), .A(n8943), .ZN(P2_U3455) );
  INV_X1 U10371 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8946) );
  MUX2_X1 U10372 ( .A(n8946), .B(n8945), .S(n10580), .Z(n8949) );
  NAND2_X1 U10373 ( .A1(n8947), .A2(n8995), .ZN(n8948) );
  OAI211_X1 U10374 ( .C1(n8950), .C2(n9003), .A(n8949), .B(n8948), .ZN(
        P2_U3454) );
  INV_X1 U10375 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8952) );
  MUX2_X1 U10376 ( .A(n8952), .B(n8951), .S(n10580), .Z(n8955) );
  NAND2_X1 U10377 ( .A1(n8953), .A2(n8995), .ZN(n8954) );
  OAI211_X1 U10378 ( .C1(n8956), .C2(n9003), .A(n8955), .B(n8954), .ZN(
        P2_U3453) );
  INV_X1 U10379 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8958) );
  MUX2_X1 U10380 ( .A(n8958), .B(n8957), .S(n10580), .Z(n8961) );
  NAND2_X1 U10381 ( .A1(n8959), .A2(n8995), .ZN(n8960) );
  OAI211_X1 U10382 ( .C1(n8962), .C2(n9003), .A(n8961), .B(n8960), .ZN(
        P2_U3452) );
  INV_X1 U10383 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8964) );
  MUX2_X1 U10384 ( .A(n8964), .B(n8963), .S(n10580), .Z(n8967) );
  NAND2_X1 U10385 ( .A1(n8965), .A2(n8995), .ZN(n8966) );
  OAI211_X1 U10386 ( .C1(n8968), .C2(n9003), .A(n8967), .B(n8966), .ZN(
        P2_U3451) );
  INV_X1 U10387 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8970) );
  MUX2_X1 U10388 ( .A(n8970), .B(n8969), .S(n10580), .Z(n8973) );
  NAND2_X1 U10389 ( .A1(n8971), .A2(n8995), .ZN(n8972) );
  OAI211_X1 U10390 ( .C1(n8974), .C2(n9003), .A(n8973), .B(n8972), .ZN(
        P2_U3450) );
  MUX2_X1 U10391 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8975), .S(n10580), .Z(
        P2_U3449) );
  INV_X1 U10392 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8977) );
  MUX2_X1 U10393 ( .A(n8977), .B(n8976), .S(n10580), .Z(n8980) );
  NAND2_X1 U10394 ( .A1(n8978), .A2(n8995), .ZN(n8979) );
  OAI211_X1 U10395 ( .C1(n8981), .C2(n9003), .A(n8980), .B(n8979), .ZN(
        P2_U3448) );
  INV_X1 U10396 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8983) );
  MUX2_X1 U10397 ( .A(n8983), .B(n8982), .S(n10580), .Z(n8986) );
  NAND2_X1 U10398 ( .A1(n8984), .A2(n8995), .ZN(n8985) );
  OAI211_X1 U10399 ( .C1(n8987), .C2(n9003), .A(n8986), .B(n8985), .ZN(
        P2_U3447) );
  MUX2_X1 U10400 ( .A(n10285), .B(n8988), .S(n10580), .Z(n8991) );
  NAND2_X1 U10401 ( .A1(n8989), .A2(n8995), .ZN(n8990) );
  OAI211_X1 U10402 ( .C1(n8992), .C2(n9003), .A(n8991), .B(n8990), .ZN(
        P2_U3444) );
  INV_X1 U10403 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8994) );
  MUX2_X1 U10404 ( .A(n8994), .B(n8993), .S(n10580), .Z(n8998) );
  NAND2_X1 U10405 ( .A1(n8996), .A2(n8995), .ZN(n8997) );
  OAI211_X1 U10406 ( .C1(n8999), .C2(n9003), .A(n8998), .B(n8997), .ZN(
        P2_U3438) );
  MUX2_X1 U10407 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9000), .S(n10580), .Z(
        n9006) );
  OAI22_X1 U10408 ( .A1(n9004), .A2(n9003), .B1(n9002), .B2(n9001), .ZN(n9005)
         );
  OR2_X1 U10409 ( .A1(n9006), .A2(n9005), .ZN(P2_U3435) );
  INV_X1 U10410 ( .A(n9960), .ZN(n9011) );
  NOR4_X1 U10411 ( .A1(n9008), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9007), .ZN(n9009) );
  AOI21_X1 U10412 ( .B1(n9021), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9009), .ZN(
        n9010) );
  OAI21_X1 U10413 ( .B1(n9011), .B2(n9023), .A(n9010), .ZN(P2_U3264) );
  INV_X1 U10414 ( .A(n9012), .ZN(n9966) );
  OAI222_X1 U10415 ( .A1(P2_U3151), .A2(n9015), .B1(n9023), .B2(n9966), .C1(
        n9014), .C2(n9013), .ZN(P2_U3266) );
  INV_X1 U10416 ( .A(n9016), .ZN(n9969) );
  AOI21_X1 U10417 ( .B1(n9021), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9017), .ZN(
        n9018) );
  OAI21_X1 U10418 ( .B1(n9969), .B2(n9023), .A(n9018), .ZN(P2_U3267) );
  INV_X1 U10419 ( .A(n9019), .ZN(n9972) );
  AOI21_X1 U10420 ( .B1(n9021), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n9020), .ZN(
        n9022) );
  OAI21_X1 U10421 ( .B1(n9972), .B2(n9023), .A(n9022), .ZN(P2_U3268) );
  INV_X1 U10422 ( .A(n9025), .ZN(n9026) );
  AOI21_X1 U10423 ( .B1(n9028), .B2(n9027), .A(n9026), .ZN(n9035) );
  INV_X1 U10424 ( .A(n9754), .ZN(n9868) );
  NAND2_X1 U10425 ( .A1(n9215), .A2(n9474), .ZN(n9030) );
  OAI211_X1 U10426 ( .C1(n9868), .C2(n9209), .A(n9030), .B(n9029), .ZN(n9031)
         );
  AOI21_X1 U10427 ( .B1(n9032), .B2(n9210), .A(n9031), .ZN(n9034) );
  NAND2_X1 U10428 ( .A1(n9892), .A2(n9142), .ZN(n9033) );
  OAI211_X1 U10429 ( .C1(n9035), .C2(n9145), .A(n9034), .B(n9033), .ZN(
        P1_U3215) );
  INV_X1 U10430 ( .A(n9036), .ZN(n9038) );
  NAND2_X1 U10431 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  XNOR2_X1 U10432 ( .A(n9040), .B(n9039), .ZN(n9045) );
  NAND2_X1 U10433 ( .A1(n9210), .A2(n9647), .ZN(n9042) );
  AOI22_X1 U10434 ( .A1(n9186), .A2(n9821), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9041) );
  OAI211_X1 U10435 ( .C1(n9680), .C2(n9189), .A(n9042), .B(n9041), .ZN(n9043)
         );
  AOI21_X1 U10436 ( .B1(n9655), .B2(n9142), .A(n9043), .ZN(n9044) );
  OAI21_X1 U10437 ( .B1(n9045), .B2(n9145), .A(n9044), .ZN(P1_U3216) );
  XNOR2_X1 U10438 ( .A(n9046), .B(n9047), .ZN(n9183) );
  NAND2_X1 U10439 ( .A1(n9183), .A2(n9184), .ZN(n9182) );
  INV_X1 U10440 ( .A(n9046), .ZN(n9048) );
  NAND2_X1 U10441 ( .A1(n9048), .A2(n9047), .ZN(n9051) );
  AND2_X1 U10442 ( .A1(n9182), .A2(n9051), .ZN(n9053) );
  XNOR2_X1 U10443 ( .A(n9050), .B(n9049), .ZN(n9052) );
  NAND3_X1 U10444 ( .A1(n9182), .A2(n9052), .A3(n9051), .ZN(n9136) );
  OAI211_X1 U10445 ( .C1(n9053), .C2(n9052), .A(n9206), .B(n9136), .ZN(n9057)
         );
  NAND2_X1 U10446 ( .A1(n9186), .A2(n9287), .ZN(n9054) );
  NAND2_X1 U10447 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9485) );
  OAI211_X1 U10448 ( .C1(n9860), .C2(n9189), .A(n9054), .B(n9485), .ZN(n9055)
         );
  AOI21_X1 U10449 ( .B1(n9705), .B2(n9210), .A(n9055), .ZN(n9056) );
  OAI211_X1 U10450 ( .C1(n4896), .C2(n9218), .A(n9057), .B(n9056), .ZN(
        P1_U3219) );
  AOI22_X1 U10451 ( .A1(n9142), .A2(n10074), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9058), .ZN(n9065) );
  AOI22_X1 U10452 ( .A1(n9215), .A2(n6689), .B1(n9186), .B2(n9483), .ZN(n9064)
         );
  OAI21_X1 U10453 ( .B1(n9059), .B2(n9061), .A(n9060), .ZN(n9062) );
  NAND2_X1 U10454 ( .A1(n9062), .A2(n9206), .ZN(n9063) );
  NAND3_X1 U10455 ( .A1(n9065), .A2(n9064), .A3(n9063), .ZN(P1_U3222) );
  INV_X1 U10456 ( .A(n9068), .ZN(n9069) );
  AOI21_X1 U10457 ( .B1(n9070), .B2(n9067), .A(n9069), .ZN(n9076) );
  INV_X1 U10458 ( .A(n9287), .ZN(n9845) );
  NOR2_X1 U10459 ( .A1(n9189), .A2(n9845), .ZN(n9073) );
  OAI22_X1 U10460 ( .A1(n9209), .A2(n9680), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9071), .ZN(n9072) );
  AOI211_X1 U10461 ( .C1(n9683), .C2(n9210), .A(n9073), .B(n9072), .ZN(n9075)
         );
  NAND2_X1 U10462 ( .A1(n9682), .A2(n9142), .ZN(n9074) );
  OAI211_X1 U10463 ( .C1(n9076), .C2(n9145), .A(n9075), .B(n9074), .ZN(
        P1_U3223) );
  INV_X1 U10464 ( .A(n9077), .ZN(n9172) );
  INV_X1 U10465 ( .A(n9078), .ZN(n9080) );
  NOR3_X1 U10466 ( .A1(n9172), .A2(n9080), .A3(n9079), .ZN(n9084) );
  INV_X1 U10467 ( .A(n9082), .ZN(n9083) );
  OAI21_X1 U10468 ( .B1(n9084), .B2(n9083), .A(n9206), .ZN(n9091) );
  AOI21_X1 U10469 ( .B1(n9186), .B2(n9474), .A(n9085), .ZN(n9086) );
  OAI21_X1 U10470 ( .B1(n9087), .B2(n9189), .A(n9086), .ZN(n9088) );
  AOI21_X1 U10471 ( .B1(n9089), .B2(n9210), .A(n9088), .ZN(n9090) );
  OAI211_X1 U10472 ( .C1(n10097), .C2(n9218), .A(n9091), .B(n9090), .ZN(
        P1_U3224) );
  AOI21_X1 U10473 ( .B1(n9093), .B2(n9092), .A(n9196), .ZN(n9098) );
  INV_X1 U10474 ( .A(n9821), .ZN(n9650) );
  NAND2_X1 U10475 ( .A1(n9210), .A2(n9613), .ZN(n9095) );
  AOI22_X1 U10476 ( .A1(n9186), .A2(n9806), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9094) );
  OAI211_X1 U10477 ( .C1(n9650), .C2(n9189), .A(n9095), .B(n9094), .ZN(n9096)
         );
  AOI21_X1 U10478 ( .B1(n9622), .B2(n9142), .A(n9096), .ZN(n9097) );
  OAI21_X1 U10479 ( .B1(n9098), .B2(n9145), .A(n9097), .ZN(P1_U3225) );
  INV_X1 U10480 ( .A(n9100), .ZN(n9102) );
  NOR2_X1 U10481 ( .A1(n9102), .A2(n9101), .ZN(n9103) );
  AOI21_X1 U10482 ( .B1(n9102), .B2(n9101), .A(n9103), .ZN(n9204) );
  NAND2_X1 U10483 ( .A1(n9204), .A2(n9205), .ZN(n9203) );
  INV_X1 U10484 ( .A(n9103), .ZN(n9104) );
  NAND2_X1 U10485 ( .A1(n9203), .A2(n9104), .ZN(n9108) );
  NAND2_X1 U10486 ( .A1(n9106), .A2(n9105), .ZN(n9107) );
  XNOR2_X1 U10487 ( .A(n9108), .B(n9107), .ZN(n9114) );
  NAND2_X1 U10488 ( .A1(n9210), .A2(n9756), .ZN(n9111) );
  INV_X1 U10489 ( .A(n9869), .ZN(n9531) );
  AOI21_X1 U10490 ( .B1(n9531), .B2(n9186), .A(n9109), .ZN(n9110) );
  OAI211_X1 U10491 ( .C1(n9868), .C2(n9189), .A(n9111), .B(n9110), .ZN(n9112)
         );
  AOI21_X1 U10492 ( .B1(n9872), .B2(n9142), .A(n9112), .ZN(n9113) );
  OAI21_X1 U10493 ( .B1(n9114), .B2(n9145), .A(n9113), .ZN(P1_U3226) );
  XNOR2_X1 U10494 ( .A(n9116), .B(n9115), .ZN(n9117) );
  XNOR2_X1 U10495 ( .A(n9118), .B(n9117), .ZN(n9123) );
  NAND2_X1 U10496 ( .A1(n9215), .A2(n9735), .ZN(n9119) );
  NAND2_X1 U10497 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10045)
         );
  OAI211_X1 U10498 ( .C1(n9860), .C2(n9209), .A(n9119), .B(n10045), .ZN(n9121)
         );
  NOR2_X1 U10499 ( .A1(n9944), .A2(n9218), .ZN(n9120) );
  AOI211_X1 U10500 ( .C1(n5123), .C2(n9210), .A(n9121), .B(n9120), .ZN(n9122)
         );
  OAI21_X1 U10501 ( .B1(n9123), .B2(n9145), .A(n9122), .ZN(P1_U3228) );
  AOI21_X1 U10502 ( .B1(n9126), .B2(n9125), .A(n9124), .ZN(n9132) );
  INV_X1 U10503 ( .A(n9631), .ZN(n9666) );
  NOR2_X1 U10504 ( .A1(n9189), .A2(n9666), .ZN(n9129) );
  OAI22_X1 U10505 ( .A1(n9209), .A2(n9549), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9127), .ZN(n9128) );
  AOI211_X1 U10506 ( .C1(n9636), .C2(n9210), .A(n9129), .B(n9128), .ZN(n9131)
         );
  NAND2_X1 U10507 ( .A1(n9922), .A2(n9142), .ZN(n9130) );
  OAI211_X1 U10508 ( .C1(n9132), .C2(n9145), .A(n9131), .B(n9130), .ZN(
        P1_U3229) );
  NAND2_X1 U10509 ( .A1(n9134), .A2(n9133), .ZN(n9138) );
  NAND2_X1 U10510 ( .A1(n9136), .A2(n9135), .ZN(n9137) );
  XOR2_X1 U10511 ( .A(n9138), .B(n9137), .Z(n9146) );
  INV_X1 U10512 ( .A(n9537), .ZN(n9724) );
  NOR2_X1 U10513 ( .A1(n9189), .A2(n9724), .ZN(n9141) );
  OAI22_X1 U10514 ( .A1(n9209), .A2(n9692), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9139), .ZN(n9140) );
  AOI211_X1 U10515 ( .C1(n9695), .C2(n9210), .A(n9141), .B(n9140), .ZN(n9144)
         );
  NAND2_X1 U10516 ( .A1(n9842), .A2(n9142), .ZN(n9143) );
  OAI211_X1 U10517 ( .C1(n9146), .C2(n9145), .A(n9144), .B(n9143), .ZN(
        P1_U3233) );
  OAI21_X1 U10518 ( .B1(n9150), .B2(n9148), .A(n9149), .ZN(n9151) );
  NAND2_X1 U10519 ( .A1(n9151), .A2(n9206), .ZN(n9157) );
  AOI21_X1 U10520 ( .B1(n9186), .B2(n10106), .A(n9152), .ZN(n9153) );
  OAI21_X1 U10521 ( .B1(n9176), .B2(n9189), .A(n9153), .ZN(n9154) );
  AOI21_X1 U10522 ( .B1(n9155), .B2(n9210), .A(n9154), .ZN(n9156) );
  OAI211_X1 U10523 ( .C1(n10110), .C2(n9218), .A(n9157), .B(n9156), .ZN(
        P1_U3234) );
  INV_X1 U10524 ( .A(n9158), .ZN(n9160) );
  NAND2_X1 U10525 ( .A1(n9160), .A2(n9159), .ZN(n9162) );
  XNOR2_X1 U10526 ( .A(n9162), .B(n9161), .ZN(n9163) );
  NAND2_X1 U10527 ( .A1(n9163), .A2(n9206), .ZN(n9168) );
  NOR2_X1 U10528 ( .A1(n9189), .A2(n9692), .ZN(n9166) );
  OAI22_X1 U10529 ( .A1(n9209), .A2(n9666), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9164), .ZN(n9165) );
  AOI211_X1 U10530 ( .C1(n9661), .C2(n9210), .A(n9166), .B(n9165), .ZN(n9167)
         );
  OAI211_X1 U10531 ( .C1(n9663), .C2(n9218), .A(n9168), .B(n9167), .ZN(
        P1_U3235) );
  INV_X1 U10532 ( .A(n7802), .ZN(n9171) );
  NOR3_X1 U10533 ( .A1(n9171), .A2(n5015), .A3(n9170), .ZN(n9173) );
  OAI21_X1 U10534 ( .B1(n9173), .B2(n9172), .A(n9206), .ZN(n9180) );
  INV_X1 U10535 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9174) );
  NOR2_X1 U10536 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9174), .ZN(n10029) );
  AOI21_X1 U10537 ( .B1(n9215), .B2(n9476), .A(n10029), .ZN(n9175) );
  OAI21_X1 U10538 ( .B1(n9176), .B2(n9209), .A(n9175), .ZN(n9177) );
  AOI21_X1 U10539 ( .B1(n9178), .B2(n9210), .A(n9177), .ZN(n9179) );
  OAI211_X1 U10540 ( .C1(n9181), .C2(n9218), .A(n9180), .B(n9179), .ZN(
        P1_U3236) );
  OAI21_X1 U10541 ( .B1(n9184), .B2(n9183), .A(n9182), .ZN(n9185) );
  NAND2_X1 U10542 ( .A1(n9185), .A2(n9206), .ZN(n9192) );
  NAND2_X1 U10543 ( .A1(n9186), .A2(n9537), .ZN(n9188) );
  OAI211_X1 U10544 ( .C1(n9869), .C2(n9189), .A(n9188), .B(n9187), .ZN(n9190)
         );
  AOI21_X1 U10545 ( .B1(n9717), .B2(n9210), .A(n9190), .ZN(n9191) );
  OAI211_X1 U10546 ( .C1(n9940), .C2(n9218), .A(n9192), .B(n9191), .ZN(
        P1_U3238) );
  INV_X1 U10547 ( .A(n9193), .ZN(n9198) );
  OAI21_X1 U10548 ( .B1(n9196), .B2(n9195), .A(n9194), .ZN(n9197) );
  NAND3_X1 U10549 ( .A1(n9198), .A2(n9206), .A3(n9197), .ZN(n9202) );
  AOI22_X1 U10550 ( .A1(n9215), .A2(n9798), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9199) );
  OAI21_X1 U10551 ( .B1(n9602), .B2(n9209), .A(n9199), .ZN(n9200) );
  AOI21_X1 U10552 ( .B1(n9599), .B2(n9210), .A(n9200), .ZN(n9201) );
  OAI211_X1 U10553 ( .C1(n9915), .C2(n9218), .A(n9202), .B(n9201), .ZN(
        P1_U3240) );
  OAI21_X1 U10554 ( .B1(n9205), .B2(n9204), .A(n9203), .ZN(n9207) );
  NAND2_X1 U10555 ( .A1(n9207), .A2(n9206), .ZN(n9217) );
  OAI21_X1 U10556 ( .B1(n9209), .B2(n9880), .A(n9208), .ZN(n9214) );
  INV_X1 U10557 ( .A(n9210), .ZN(n9212) );
  NOR2_X1 U10558 ( .A1(n9212), .A2(n9211), .ZN(n9213) );
  AOI211_X1 U10559 ( .C1(n9215), .C2(n10106), .A(n9214), .B(n9213), .ZN(n9216)
         );
  OAI211_X1 U10560 ( .C1(n7788), .C2(n9218), .A(n9217), .B(n9216), .ZN(
        P1_U3241) );
  NOR4_X1 U10561 ( .A1(n9219), .A2(n9877), .A3(n6541), .A4(n9459), .ZN(n9473)
         );
  OAI21_X1 U10562 ( .B1(n9466), .B2(n9465), .A(P1_B_REG_SCAN_IN), .ZN(n9472)
         );
  INV_X1 U10563 ( .A(n9280), .ZN(n9448) );
  INV_X1 U10564 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9223) );
  INV_X1 U10565 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9770) );
  OR2_X1 U10566 ( .A1(n5975), .A2(n9770), .ZN(n9222) );
  INV_X1 U10567 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9900) );
  OR2_X1 U10568 ( .A1(n6086), .A2(n9900), .ZN(n9221) );
  OAI211_X1 U10569 ( .C1(n9224), .C2(n9223), .A(n9222), .B(n9221), .ZN(n9555)
         );
  INV_X1 U10570 ( .A(n9555), .ZN(n9447) );
  NOR2_X1 U10571 ( .A1(n9507), .A2(n9447), .ZN(n9281) );
  INV_X1 U10572 ( .A(n9281), .ZN(n9225) );
  NAND2_X1 U10573 ( .A1(n9578), .A2(n9774), .ZN(n9524) );
  NAND2_X1 U10574 ( .A1(n9591), .A2(n9602), .ZN(n9521) );
  OR2_X1 U10575 ( .A1(n9591), .A2(n9602), .ZN(n9437) );
  OR2_X1 U10576 ( .A1(n9233), .A2(n9616), .ZN(n9321) );
  NAND2_X1 U10577 ( .A1(n9437), .A2(n9321), .ZN(n9237) );
  OR2_X1 U10578 ( .A1(n9622), .A2(n9549), .ZN(n9320) );
  OR2_X1 U10579 ( .A1(n9922), .A2(n9650), .ZN(n9518) );
  NAND2_X1 U10580 ( .A1(n9417), .A2(n9515), .ZN(n9326) );
  NAND2_X1 U10581 ( .A1(n9655), .A2(n9666), .ZN(n9517) );
  NAND2_X1 U10582 ( .A1(n9326), .A2(n9517), .ZN(n9226) );
  NAND2_X1 U10583 ( .A1(n9518), .A2(n9226), .ZN(n9227) );
  NAND2_X1 U10584 ( .A1(n9922), .A2(n9650), .ZN(n9422) );
  NAND2_X1 U10585 ( .A1(n9227), .A2(n9422), .ZN(n9228) );
  AND2_X1 U10586 ( .A1(n9228), .A2(n9320), .ZN(n9234) );
  OR2_X1 U10587 ( .A1(n9682), .A2(n9692), .ZN(n9404) );
  AND2_X1 U10588 ( .A1(n9842), .A2(n9845), .ZN(n9405) );
  NAND2_X1 U10589 ( .A1(n9404), .A2(n9405), .ZN(n9229) );
  NAND2_X1 U10590 ( .A1(n9682), .A2(n9692), .ZN(n9411) );
  AND2_X1 U10591 ( .A1(n9229), .A2(n9411), .ZN(n9514) );
  NAND2_X1 U10592 ( .A1(n9831), .A2(n9680), .ZN(n9286) );
  AND2_X1 U10593 ( .A1(n9517), .A2(n9286), .ZN(n9324) );
  NAND3_X1 U10594 ( .A1(n9422), .A2(n9514), .A3(n9324), .ZN(n9230) );
  AND2_X1 U10595 ( .A1(n9622), .A2(n9549), .ZN(n9312) );
  AOI21_X1 U10596 ( .B1(n9234), .B2(n9230), .A(n9312), .ZN(n9231) );
  NOR2_X1 U10597 ( .A1(n9237), .A2(n9231), .ZN(n9232) );
  AND2_X1 U10598 ( .A1(n9233), .A2(n9616), .ZN(n9285) );
  INV_X1 U10599 ( .A(n9234), .ZN(n9235) );
  OR2_X1 U10600 ( .A1(n9842), .A2(n9845), .ZN(n9674) );
  NAND2_X1 U10601 ( .A1(n9404), .A2(n9674), .ZN(n9513) );
  NOR2_X1 U10602 ( .A1(n9235), .A2(n9513), .ZN(n9240) );
  INV_X1 U10603 ( .A(n9236), .ZN(n9238) );
  AND2_X1 U10604 ( .A1(n9907), .A2(n9789), .ZN(n9284) );
  AOI21_X1 U10605 ( .B1(n9238), .B2(n9237), .A(n9284), .ZN(n9239) );
  OR2_X1 U10606 ( .A1(n9575), .A2(n9777), .ZN(n9441) );
  OR2_X1 U10607 ( .A1(n9534), .A2(n9860), .ZN(n9288) );
  OR2_X1 U10608 ( .A1(n9743), .A2(n9869), .ZN(n9719) );
  AND2_X1 U10609 ( .A1(n9288), .A2(n9719), .ZN(n9399) );
  NAND2_X1 U10610 ( .A1(n9872), .A2(n9880), .ZN(n9392) );
  NAND2_X1 U10611 ( .A1(n9527), .A2(n9868), .ZN(n9269) );
  NAND2_X1 U10612 ( .A1(n9392), .A2(n9269), .ZN(n9391) );
  INV_X1 U10613 ( .A(n9377), .ZN(n9241) );
  OR2_X1 U10614 ( .A1(n9391), .A2(n9241), .ZN(n9394) );
  INV_X1 U10615 ( .A(n9394), .ZN(n9259) );
  AND2_X1 U10616 ( .A1(n9380), .A2(n9379), .ZN(n9393) );
  INV_X1 U10617 ( .A(n9335), .ZN(n9247) );
  NAND4_X1 U10618 ( .A1(n9453), .A2(n9245), .A3(n9244), .A4(n9243), .ZN(n9246)
         );
  NOR2_X1 U10619 ( .A1(n9247), .A2(n9246), .ZN(n9249) );
  AND2_X1 U10620 ( .A1(n9249), .A2(n9248), .ZN(n9251) );
  OAI211_X1 U10621 ( .C1(n9252), .C2(n9251), .A(n9370), .B(n9250), .ZN(n9254)
         );
  NAND2_X1 U10622 ( .A1(n9372), .A2(n9368), .ZN(n9362) );
  INV_X1 U10623 ( .A(n9362), .ZN(n9253) );
  AND2_X1 U10624 ( .A1(n9254), .A2(n9253), .ZN(n9255) );
  NAND2_X1 U10625 ( .A1(n9374), .A2(n9371), .ZN(n9364) );
  OAI211_X1 U10626 ( .C1(n9255), .C2(n9364), .A(n9384), .B(n9373), .ZN(n9256)
         );
  NAND2_X1 U10627 ( .A1(n9393), .A2(n9256), .ZN(n9258) );
  OR2_X1 U10628 ( .A1(n9527), .A2(n9868), .ZN(n9257) );
  NAND2_X1 U10629 ( .A1(n9390), .A2(n9257), .ZN(n9383) );
  AOI22_X1 U10630 ( .A1(n9259), .A2(n9258), .B1(n9392), .B2(n9383), .ZN(n9261)
         );
  NAND2_X1 U10631 ( .A1(n9534), .A2(n9860), .ZN(n9400) );
  AND2_X1 U10632 ( .A1(n9743), .A2(n9869), .ZN(n9272) );
  AND2_X1 U10633 ( .A1(n9400), .A2(n9273), .ZN(n9408) );
  INV_X1 U10634 ( .A(n9408), .ZN(n9260) );
  AOI21_X1 U10635 ( .B1(n9399), .B2(n9261), .A(n9260), .ZN(n9262) );
  OR2_X1 U10636 ( .A1(n9935), .A2(n9724), .ZN(n9327) );
  NAND2_X1 U10637 ( .A1(n9327), .A2(n9288), .ZN(n9412) );
  NAND2_X1 U10638 ( .A1(n9935), .A2(n9724), .ZN(n9406) );
  OAI21_X1 U10639 ( .B1(n9262), .B2(n9412), .A(n9406), .ZN(n9263) );
  NOR2_X1 U10640 ( .A1(n9268), .A2(n9263), .ZN(n9265) );
  NAND2_X1 U10641 ( .A1(n9507), .A2(n9447), .ZN(n9316) );
  NAND2_X1 U10642 ( .A1(n9777), .A2(n9575), .ZN(n9442) );
  NAND2_X1 U10643 ( .A1(n9316), .A2(n9442), .ZN(n9278) );
  INV_X1 U10644 ( .A(n9278), .ZN(n9264) );
  OAI21_X1 U10645 ( .B1(n9275), .B2(n9265), .A(n9264), .ZN(n9266) );
  NAND2_X1 U10646 ( .A1(n4564), .A2(n9266), .ZN(n9267) );
  AND2_X1 U10647 ( .A1(n9898), .A2(n9280), .ZN(n9318) );
  INV_X1 U10648 ( .A(n9318), .ZN(n9469) );
  NAND2_X1 U10649 ( .A1(n9267), .A2(n9469), .ZN(n9458) );
  INV_X1 U10650 ( .A(n9268), .ZN(n9276) );
  NAND2_X1 U10651 ( .A1(n9271), .A2(n9392), .ZN(n9732) );
  INV_X1 U10652 ( .A(n9406), .ZN(n9274) );
  AOI21_X1 U10653 ( .B1(n9276), .B2(n9512), .A(n9275), .ZN(n9277) );
  AOI21_X1 U10654 ( .B1(n9281), .B2(n9280), .A(n9279), .ZN(n9283) );
  OAI211_X1 U10655 ( .C1(n9283), .C2(n9318), .A(n9282), .B(n9462), .ZN(n9319)
         );
  NAND2_X1 U10656 ( .A1(n9441), .A2(n9442), .ZN(n9525) );
  NAND2_X1 U10657 ( .A1(n9436), .A2(n9524), .ZN(n9569) );
  NAND2_X1 U10658 ( .A1(n9437), .A2(n9521), .ZN(n9582) );
  INV_X1 U10659 ( .A(n9285), .ZN(n9520) );
  NAND2_X1 U10660 ( .A1(n9321), .A2(n9520), .ZN(n9551) );
  NAND2_X1 U10661 ( .A1(n9417), .A2(n9517), .ZN(n9516) );
  XNOR2_X1 U10662 ( .A(n9682), .B(n9692), .ZN(n9677) );
  OR2_X1 U10663 ( .A1(n9842), .A2(n9287), .ZN(n9539) );
  NAND2_X1 U10664 ( .A1(n9842), .A2(n9287), .ZN(n9541) );
  NAND2_X1 U10665 ( .A1(n9539), .A2(n9541), .ZN(n9690) );
  NAND2_X1 U10666 ( .A1(n9719), .A2(n9273), .ZN(n9731) );
  INV_X1 U10667 ( .A(n9289), .ZN(n9298) );
  AND4_X1 U10668 ( .A1(n9291), .A2(n10067), .A3(n9290), .A4(n9464), .ZN(n9293)
         );
  NAND3_X1 U10669 ( .A1(n9293), .A2(n9292), .A3(n6748), .ZN(n9295) );
  NOR3_X1 U10670 ( .A1(n9296), .A2(n9295), .A3(n9294), .ZN(n9297) );
  NAND4_X1 U10671 ( .A1(n9300), .A2(n9299), .A3(n9298), .A4(n9297), .ZN(n9302)
         );
  OR4_X1 U10672 ( .A1(n9304), .A2(n9303), .A3(n9302), .A4(n9301), .ZN(n9307)
         );
  INV_X1 U10673 ( .A(n9762), .ZN(n9748) );
  OR4_X1 U10674 ( .A1(n9307), .A2(n9748), .A3(n9306), .A4(n9305), .ZN(n9308)
         );
  NOR2_X1 U10675 ( .A1(n9731), .A2(n9308), .ZN(n9309) );
  NAND4_X1 U10676 ( .A1(n9690), .A2(n9710), .A3(n9721), .A4(n9309), .ZN(n9310)
         );
  NOR4_X1 U10677 ( .A1(n9516), .A2(n9664), .A3(n9677), .A4(n9310), .ZN(n9311)
         );
  NAND2_X1 U10678 ( .A1(n9629), .A2(n9311), .ZN(n9313) );
  NAND2_X1 U10679 ( .A1(n9320), .A2(n9519), .ZN(n9612) );
  OR4_X1 U10680 ( .A1(n9582), .A2(n9551), .A3(n9313), .A4(n9612), .ZN(n9314)
         );
  NOR2_X1 U10681 ( .A1(n9569), .A2(n9314), .ZN(n9315) );
  NAND2_X1 U10682 ( .A1(n9316), .A2(n9315), .ZN(n9317) );
  INV_X1 U10683 ( .A(n9463), .ZN(n9444) );
  NAND2_X1 U10684 ( .A1(n9520), .A2(n9519), .ZN(n9428) );
  OR3_X1 U10685 ( .A1(n9438), .A2(n9463), .A3(n9428), .ZN(n9427) );
  OR2_X1 U10686 ( .A1(n9428), .A2(n9320), .ZN(n9322) );
  NAND2_X1 U10687 ( .A1(n9322), .A2(n9321), .ZN(n9433) );
  INV_X1 U10688 ( .A(n9437), .ZN(n9323) );
  OR3_X1 U10689 ( .A1(n9433), .A2(n9323), .A3(n9444), .ZN(n9426) );
  INV_X1 U10690 ( .A(n9324), .ZN(n9325) );
  MUX2_X1 U10691 ( .A(n9326), .B(n9325), .S(n9463), .Z(n9420) );
  AND2_X1 U10692 ( .A1(n9327), .A2(n9444), .ZN(n9403) );
  NAND2_X1 U10693 ( .A1(n9328), .A2(n9444), .ZN(n9329) );
  OR2_X1 U10694 ( .A1(n9331), .A2(n9463), .ZN(n9332) );
  NAND2_X1 U10695 ( .A1(n9333), .A2(n9332), .ZN(n9344) );
  NAND2_X1 U10696 ( .A1(n9345), .A2(n9343), .ZN(n9334) );
  AOI21_X1 U10697 ( .B1(n9344), .B2(n9335), .A(n9334), .ZN(n9336) );
  OAI21_X1 U10698 ( .B1(n9336), .B2(n9351), .A(n9350), .ZN(n9339) );
  INV_X1 U10699 ( .A(n9337), .ZN(n9338) );
  AOI21_X1 U10700 ( .B1(n9339), .B2(n9349), .A(n9338), .ZN(n9341) );
  OR2_X1 U10701 ( .A1(n9341), .A2(n9340), .ZN(n9360) );
  NAND3_X1 U10702 ( .A1(n9344), .A2(n9343), .A3(n9342), .ZN(n9348) );
  INV_X1 U10703 ( .A(n9345), .ZN(n9346) );
  AOI21_X1 U10704 ( .B1(n9348), .B2(n9347), .A(n9346), .ZN(n9352) );
  OAI211_X1 U10705 ( .C1(n9352), .C2(n9351), .A(n9350), .B(n9349), .ZN(n9356)
         );
  INV_X1 U10706 ( .A(n9353), .ZN(n9354) );
  NAND3_X1 U10707 ( .A1(n9356), .A2(n9355), .A3(n9354), .ZN(n9358) );
  NAND3_X1 U10708 ( .A1(n9358), .A2(n9361), .A3(n9357), .ZN(n9359) );
  MUX2_X1 U10709 ( .A(n9360), .B(n9359), .S(n9444), .Z(n9367) );
  NAND2_X1 U10710 ( .A1(n9367), .A2(n9361), .ZN(n9363) );
  AOI21_X1 U10711 ( .B1(n9363), .B2(n9370), .A(n9362), .ZN(n9365) );
  OAI21_X1 U10712 ( .B1(n9365), .B2(n9364), .A(n9373), .ZN(n9376) );
  NAND2_X1 U10713 ( .A1(n9367), .A2(n9366), .ZN(n9369) );
  MUX2_X1 U10714 ( .A(n9376), .B(n9375), .S(n9444), .Z(n9385) );
  NAND2_X1 U10715 ( .A1(n9377), .A2(n9384), .ZN(n9378) );
  AOI21_X1 U10716 ( .B1(n9385), .B2(n9379), .A(n9378), .ZN(n9382) );
  INV_X1 U10717 ( .A(n9380), .ZN(n9381) );
  NOR3_X1 U10718 ( .A1(n9383), .A2(n9382), .A3(n9381), .ZN(n9388) );
  NAND2_X1 U10719 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  OAI21_X1 U10720 ( .B1(n9394), .B2(n9386), .A(n9390), .ZN(n9387) );
  NOR2_X1 U10721 ( .A1(n9527), .A2(n9463), .ZN(n9389) );
  AOI21_X1 U10722 ( .B1(n9391), .B2(n9390), .A(n9389), .ZN(n9397) );
  AOI21_X1 U10723 ( .B1(n9392), .B2(n9754), .A(n9463), .ZN(n9396) );
  OR3_X1 U10724 ( .A1(n9394), .A2(n9393), .A3(n9463), .ZN(n9395) );
  OAI21_X1 U10725 ( .B1(n9397), .B2(n9396), .A(n9395), .ZN(n9398) );
  INV_X1 U10726 ( .A(n9731), .ZN(n9733) );
  NAND3_X1 U10727 ( .A1(n9401), .A2(n9406), .A3(n9400), .ZN(n9402) );
  INV_X1 U10728 ( .A(n9405), .ZN(n9676) );
  AND2_X1 U10729 ( .A1(n9406), .A2(n9463), .ZN(n9407) );
  OAI211_X1 U10730 ( .C1(n9412), .C2(n9408), .A(n9676), .B(n9407), .ZN(n9409)
         );
  INV_X1 U10731 ( .A(n9409), .ZN(n9410) );
  OAI211_X1 U10732 ( .C1(n9413), .C2(n9412), .A(n9411), .B(n9410), .ZN(n9416)
         );
  OAI21_X1 U10733 ( .B1(n9692), .B2(n9674), .A(n9682), .ZN(n9415) );
  AOI21_X1 U10734 ( .B1(n9674), .B2(n9692), .A(n9444), .ZN(n9414) );
  MUX2_X1 U10735 ( .A(n9517), .B(n9417), .S(n9463), .Z(n9418) );
  OAI21_X1 U10736 ( .B1(n9420), .B2(n9419), .A(n9418), .ZN(n9421) );
  NAND2_X1 U10737 ( .A1(n9421), .A2(n9629), .ZN(n9424) );
  MUX2_X1 U10738 ( .A(n9422), .B(n9518), .S(n9463), .Z(n9423) );
  NAND2_X1 U10739 ( .A1(n9424), .A2(n9423), .ZN(n9425) );
  AOI21_X1 U10740 ( .B1(n9427), .B2(n9426), .A(n9425), .ZN(n9435) );
  NAND3_X1 U10741 ( .A1(n9437), .A2(n9463), .A3(n9428), .ZN(n9432) );
  INV_X1 U10742 ( .A(n9438), .ZN(n9429) );
  NAND3_X1 U10743 ( .A1(n9429), .A2(n9433), .A3(n9444), .ZN(n9431) );
  NAND2_X1 U10744 ( .A1(n9438), .A2(n9463), .ZN(n9430) );
  OAI211_X1 U10745 ( .C1(n9433), .C2(n9432), .A(n9431), .B(n9430), .ZN(n9434)
         );
  OAI21_X1 U10746 ( .B1(n9438), .B2(n9437), .A(n9436), .ZN(n9439) );
  NAND2_X1 U10747 ( .A1(n9439), .A2(n9444), .ZN(n9440) );
  INV_X1 U10748 ( .A(n9525), .ZN(n9552) );
  MUX2_X1 U10749 ( .A(n9442), .B(n9441), .S(n9444), .Z(n9443) );
  MUX2_X1 U10750 ( .A(n9444), .B(n9446), .S(n9507), .Z(n9445) );
  NOR3_X2 U10751 ( .A1(n9445), .A2(n9898), .A3(n9447), .ZN(n9452) );
  MUX2_X1 U10752 ( .A(n9446), .B(n9463), .S(n9507), .Z(n9450) );
  OAI21_X1 U10753 ( .B1(n9448), .B2(n9447), .A(n9469), .ZN(n9449) );
  AOI21_X1 U10754 ( .B1(n9450), .B2(n9462), .A(n9449), .ZN(n9451) );
  NOR2_X1 U10755 ( .A1(n9452), .A2(n9451), .ZN(n9460) );
  OAI21_X1 U10756 ( .B1(n9460), .B2(n9454), .A(n9453), .ZN(n9455) );
  AOI21_X1 U10757 ( .B1(n9458), .B2(n9456), .A(n9466), .ZN(n9457) );
  INV_X1 U10758 ( .A(n9460), .ZN(n9461) );
  OAI21_X1 U10759 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(n9468) );
  NOR4_X1 U10760 ( .A1(n9466), .A2(n9465), .A3(n9464), .A4(n6437), .ZN(n9467)
         );
  OAI211_X1 U10761 ( .C1(n6736), .C2(n9469), .A(n9468), .B(n9467), .ZN(n9470)
         );
  OAI211_X1 U10762 ( .C1(n9473), .C2(n9472), .A(n9471), .B(n9470), .ZN(
        P1_U3242) );
  MUX2_X1 U10763 ( .A(n9555), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9484), .Z(
        P1_U3584) );
  MUX2_X1 U10764 ( .A(n9781), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9484), .Z(
        P1_U3583) );
  MUX2_X1 U10765 ( .A(n9789), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9484), .Z(
        P1_U3582) );
  MUX2_X1 U10766 ( .A(n9797), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9484), .Z(
        P1_U3581) );
  MUX2_X1 U10767 ( .A(n9806), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9484), .Z(
        P1_U3580) );
  MUX2_X1 U10768 ( .A(n9798), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9484), .Z(
        P1_U3579) );
  MUX2_X1 U10769 ( .A(n9821), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9484), .Z(
        P1_U3578) );
  MUX2_X1 U10770 ( .A(n9631), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9484), .Z(
        P1_U3577) );
  MUX2_X1 U10771 ( .A(n9822), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9484), .Z(
        P1_U3576) );
  MUX2_X1 U10772 ( .A(n9542), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9484), .Z(
        P1_U3575) );
  MUX2_X1 U10773 ( .A(n9537), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9484), .Z(
        P1_U3573) );
  MUX2_X1 U10774 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9704), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10775 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9531), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10776 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9735), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10777 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9754), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10778 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10106), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10779 ( .A(n9474), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9484), .Z(
        P1_U3567) );
  MUX2_X1 U10780 ( .A(n10103), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9484), .Z(
        P1_U3566) );
  MUX2_X1 U10781 ( .A(n9475), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9484), .Z(
        P1_U3565) );
  MUX2_X1 U10782 ( .A(n9476), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9484), .Z(
        P1_U3564) );
  MUX2_X1 U10783 ( .A(n9477), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9484), .Z(
        P1_U3563) );
  MUX2_X1 U10784 ( .A(n9478), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9484), .Z(
        P1_U3562) );
  MUX2_X1 U10785 ( .A(n9479), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9484), .Z(
        P1_U3561) );
  MUX2_X1 U10786 ( .A(n9480), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9484), .Z(
        P1_U3560) );
  MUX2_X1 U10787 ( .A(n9481), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9484), .Z(
        P1_U3559) );
  MUX2_X1 U10788 ( .A(n9482), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9484), .Z(
        P1_U3557) );
  MUX2_X1 U10789 ( .A(n9483), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9484), .Z(
        P1_U3556) );
  MUX2_X1 U10790 ( .A(n6689), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9484), .Z(
        P1_U3554) );
  INV_X1 U10791 ( .A(n9485), .ZN(n9502) );
  NAND2_X1 U10792 ( .A1(n9487), .A2(n9486), .ZN(n9488) );
  XNOR2_X1 U10793 ( .A(n9488), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U10794 ( .A1(n9489), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U10795 ( .A1(n9491), .A2(n9490), .ZN(n9492) );
  XNOR2_X1 U10796 ( .A(n9492), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9496) );
  OAI22_X1 U10797 ( .A1(n9495), .A2(n9494), .B1(n9496), .B2(n9493), .ZN(n9500)
         );
  NAND2_X1 U10798 ( .A1(n9495), .A2(n10039), .ZN(n9498) );
  NAND2_X1 U10799 ( .A1(n9496), .A2(n10043), .ZN(n9497) );
  NAND3_X1 U10800 ( .A1(n9498), .A2(n9497), .A3(n10027), .ZN(n9499) );
  MUX2_X1 U10801 ( .A(n9500), .B(n9499), .S(n6264), .Z(n9501) );
  AOI211_X1 U10802 ( .C1(P1_ADDR_REG_19__SCAN_IN), .C2(n10030), .A(n9502), .B(
        n9501), .ZN(n9503) );
  INV_X1 U10803 ( .A(n9503), .ZN(P1_U3262) );
  INV_X1 U10804 ( .A(n9554), .ZN(n9506) );
  INV_X1 U10805 ( .A(n9504), .ZN(n9505) );
  AOI211_X1 U10806 ( .C1(n9507), .C2(n9506), .A(n9750), .B(n9505), .ZN(n9769)
         );
  NAND2_X1 U10807 ( .A1(n9769), .A2(n10053), .ZN(n9511) );
  AND2_X1 U10808 ( .A1(n10063), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9508) );
  NOR2_X1 U10809 ( .A1(n9509), .A2(n9508), .ZN(n9510) );
  OAI211_X1 U10810 ( .C1(n9902), .C2(n9752), .A(n9511), .B(n9510), .ZN(
        P1_U3264) );
  INV_X1 U10811 ( .A(n9516), .ZN(n9646) );
  NAND2_X1 U10812 ( .A1(n9643), .A2(n9646), .ZN(n9642) );
  AND2_X2 U10813 ( .A1(n9642), .A2(n9517), .ZN(n9630) );
  NAND2_X1 U10814 ( .A1(n9630), .A2(n9629), .ZN(n9628) );
  INV_X1 U10815 ( .A(n9612), .ZN(n9609) );
  NAND2_X1 U10816 ( .A1(n9608), .A2(n9519), .ZN(n9595) );
  INV_X1 U10817 ( .A(n9551), .ZN(n9597) );
  NAND2_X1 U10818 ( .A1(n9595), .A2(n9597), .ZN(n9594) );
  INV_X1 U10819 ( .A(n9582), .ZN(n9523) );
  INV_X1 U10820 ( .A(n9521), .ZN(n9522) );
  OAI21_X1 U10821 ( .B1(n9567), .B2(n9569), .A(n9524), .ZN(n9526) );
  XNOR2_X1 U10822 ( .A(n9526), .B(n9525), .ZN(n9778) );
  NAND2_X1 U10823 ( .A1(n4518), .A2(n9748), .ZN(n9747) );
  NAND2_X1 U10824 ( .A1(n9872), .A2(n9735), .ZN(n9529) );
  NAND2_X1 U10825 ( .A1(n9747), .A2(n9529), .ZN(n9734) );
  AND2_X1 U10826 ( .A1(n9743), .A2(n9531), .ZN(n9530) );
  OR2_X1 U10827 ( .A1(n9743), .A2(n9531), .ZN(n9532) );
  NOR2_X1 U10828 ( .A1(n9534), .A2(n9704), .ZN(n9533) );
  NAND2_X1 U10829 ( .A1(n9534), .A2(n9704), .ZN(n9535) );
  INV_X1 U10830 ( .A(n9701), .ZN(n9536) );
  OR2_X1 U10831 ( .A1(n9935), .A2(n9537), .ZN(n9538) );
  INV_X1 U10832 ( .A(n9539), .ZN(n9540) );
  AND2_X1 U10833 ( .A1(n9682), .A2(n9542), .ZN(n9543) );
  OAI22_X1 U10834 ( .A1(n9673), .A2(n9543), .B1(n9542), .B2(n9682), .ZN(n9658)
         );
  NOR2_X1 U10835 ( .A1(n9831), .A2(n9822), .ZN(n9545) );
  NAND2_X1 U10836 ( .A1(n9831), .A2(n9822), .ZN(n9544) );
  OAI21_X1 U10837 ( .B1(n9658), .B2(n9545), .A(n9544), .ZN(n9645) );
  AND2_X1 U10838 ( .A1(n9655), .A2(n9631), .ZN(n9546) );
  OR2_X1 U10839 ( .A1(n9655), .A2(n9631), .ZN(n9547) );
  NAND2_X1 U10840 ( .A1(n9550), .A2(n5117), .ZN(n9598) );
  NAND2_X1 U10841 ( .A1(n9772), .A2(n10059), .ZN(n9565) );
  AOI211_X1 U10842 ( .C1(n4534), .C2(n9777), .A(n9554), .B(n9750), .ZN(n9775)
         );
  NAND2_X1 U10843 ( .A1(n9777), .A2(n10050), .ZN(n9561) );
  NAND2_X1 U10844 ( .A1(n9556), .A2(n9555), .ZN(n9773) );
  OAI22_X1 U10845 ( .A1(n10063), .A2(n9773), .B1(n9558), .B2(n9557), .ZN(n9559) );
  AOI21_X1 U10846 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n10063), .A(n9559), .ZN(
        n9560) );
  OAI211_X1 U10847 ( .C1(n9774), .C2(n9562), .A(n9561), .B(n9560), .ZN(n9563)
         );
  AOI21_X1 U10848 ( .B1(n9775), .B2(n10053), .A(n9563), .ZN(n9564) );
  OAI211_X1 U10849 ( .C1(n9778), .C2(n9746), .A(n9565), .B(n9564), .ZN(
        P1_U3356) );
  INV_X1 U10850 ( .A(n9569), .ZN(n9566) );
  XNOR2_X1 U10851 ( .A(n9567), .B(n9566), .ZN(n9784) );
  OAI21_X1 U10852 ( .B1(n9570), .B2(n9569), .A(n9568), .ZN(n9571) );
  INV_X1 U10853 ( .A(n9571), .ZN(n9786) );
  NAND2_X1 U10854 ( .A1(n9786), .A2(n10059), .ZN(n9580) );
  NAND2_X1 U10855 ( .A1(n9755), .A2(n9797), .ZN(n9574) );
  AOI22_X1 U10856 ( .A1(n10063), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9572), 
        .B2(n10051), .ZN(n9573) );
  OAI211_X1 U10857 ( .C1(n9575), .C2(n9759), .A(n9574), .B(n9573), .ZN(n9577)
         );
  OAI211_X1 U10858 ( .C1(n9907), .C2(n9587), .A(n9739), .B(n4534), .ZN(n9782)
         );
  NOR2_X1 U10859 ( .A1(n9782), .A2(n9740), .ZN(n9576) );
  AOI211_X1 U10860 ( .C1(n10050), .C2(n9578), .A(n9577), .B(n9576), .ZN(n9579)
         );
  OAI211_X1 U10861 ( .C1(n9746), .C2(n9784), .A(n9580), .B(n9579), .ZN(
        P1_U3265) );
  XNOR2_X1 U10862 ( .A(n9581), .B(n9582), .ZN(n9792) );
  XNOR2_X1 U10863 ( .A(n9583), .B(n9582), .ZN(n9794) );
  NAND2_X1 U10864 ( .A1(n9794), .A2(n10059), .ZN(n9593) );
  NAND2_X1 U10865 ( .A1(n9755), .A2(n9806), .ZN(n9586) );
  AOI22_X1 U10866 ( .A1(n10063), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9584), 
        .B2(n10051), .ZN(n9585) );
  OAI211_X1 U10867 ( .C1(n9774), .C2(n9759), .A(n9586), .B(n9585), .ZN(n9590)
         );
  INV_X1 U10868 ( .A(n9587), .ZN(n9588) );
  OAI211_X1 U10869 ( .C1(n9911), .C2(n4893), .A(n9588), .B(n9739), .ZN(n9790)
         );
  NOR2_X1 U10870 ( .A1(n9790), .A2(n9740), .ZN(n9589) );
  AOI211_X1 U10871 ( .C1(n10050), .C2(n9591), .A(n9590), .B(n9589), .ZN(n9592)
         );
  OAI211_X1 U10872 ( .C1(n9746), .C2(n9792), .A(n9593), .B(n9592), .ZN(
        P1_U3266) );
  OAI21_X1 U10873 ( .B1(n9595), .B2(n9597), .A(n9594), .ZN(n9596) );
  INV_X1 U10874 ( .A(n9596), .ZN(n9801) );
  XNOR2_X1 U10875 ( .A(n9598), .B(n9597), .ZN(n9803) );
  NAND2_X1 U10876 ( .A1(n9803), .A2(n10059), .ZN(n9607) );
  NAND2_X1 U10877 ( .A1(n9755), .A2(n9798), .ZN(n9601) );
  AOI22_X1 U10878 ( .A1(n10063), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9599), 
        .B2(n10051), .ZN(n9600) );
  OAI211_X1 U10879 ( .C1(n9602), .C2(n9759), .A(n9601), .B(n9600), .ZN(n9605)
         );
  OAI211_X1 U10880 ( .C1(n9915), .C2(n9617), .A(n9603), .B(n9739), .ZN(n9799)
         );
  NOR2_X1 U10881 ( .A1(n9799), .A2(n9740), .ZN(n9604) );
  AOI211_X1 U10882 ( .C1(n10050), .C2(n9233), .A(n9605), .B(n9604), .ZN(n9606)
         );
  OAI211_X1 U10883 ( .C1(n9801), .C2(n9746), .A(n9607), .B(n9606), .ZN(
        P1_U3267) );
  OAI21_X1 U10884 ( .B1(n9610), .B2(n9609), .A(n9608), .ZN(n9611) );
  INV_X1 U10885 ( .A(n9611), .ZN(n9809) );
  XNOR2_X1 U10886 ( .A(n4545), .B(n9612), .ZN(n9811) );
  NAND2_X1 U10887 ( .A1(n9811), .A2(n10059), .ZN(n9624) );
  NAND2_X1 U10888 ( .A1(n9755), .A2(n9821), .ZN(n9615) );
  AOI22_X1 U10889 ( .A1(n10063), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9613), 
        .B2(n10051), .ZN(n9614) );
  OAI211_X1 U10890 ( .C1(n9616), .C2(n9759), .A(n9615), .B(n9614), .ZN(n9621)
         );
  INV_X1 U10891 ( .A(n9635), .ZN(n9619) );
  INV_X1 U10892 ( .A(n9617), .ZN(n9618) );
  OAI211_X1 U10893 ( .C1(n9919), .C2(n9619), .A(n9618), .B(n9739), .ZN(n9807)
         );
  NOR2_X1 U10894 ( .A1(n9807), .A2(n9740), .ZN(n9620) );
  AOI211_X1 U10895 ( .C1(n10050), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9623)
         );
  OAI211_X1 U10896 ( .C1(n9809), .C2(n9746), .A(n9624), .B(n9623), .ZN(
        P1_U3268) );
  AND2_X1 U10897 ( .A1(n9625), .A2(n9629), .ZN(n9626) );
  OR2_X1 U10898 ( .A1(n9627), .A2(n9626), .ZN(n9817) );
  OAI211_X1 U10899 ( .C1(n9630), .C2(n9629), .A(n9628), .B(n10116), .ZN(n9633)
         );
  AOI22_X1 U10900 ( .A1(n10104), .A2(n9631), .B1(n9798), .B2(n10105), .ZN(
        n9632) );
  NAND2_X1 U10901 ( .A1(n9633), .A2(n9632), .ZN(n9815) );
  INV_X1 U10902 ( .A(n9922), .ZN(n9639) );
  AOI21_X1 U10903 ( .B1(n9922), .B2(n9652), .A(n9750), .ZN(n9634) );
  AND2_X1 U10904 ( .A1(n9635), .A2(n9634), .ZN(n9814) );
  NAND2_X1 U10905 ( .A1(n9814), .A2(n10053), .ZN(n9638) );
  AOI22_X1 U10906 ( .A1(n10063), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9636), 
        .B2(n10051), .ZN(n9637) );
  OAI211_X1 U10907 ( .C1(n9639), .C2(n9752), .A(n9638), .B(n9637), .ZN(n9640)
         );
  AOI21_X1 U10908 ( .B1(n9815), .B2(n10056), .A(n9640), .ZN(n9641) );
  OAI21_X1 U10909 ( .B1(n9817), .B2(n9767), .A(n9641), .ZN(P1_U3269) );
  OAI21_X1 U10910 ( .B1(n9643), .B2(n9646), .A(n9642), .ZN(n9644) );
  INV_X1 U10911 ( .A(n9644), .ZN(n9825) );
  XNOR2_X1 U10912 ( .A(n9645), .B(n9646), .ZN(n9827) );
  NAND2_X1 U10913 ( .A1(n9827), .A2(n10059), .ZN(n9657) );
  NAND2_X1 U10914 ( .A1(n9755), .A2(n9822), .ZN(n9649) );
  AOI22_X1 U10915 ( .A1(n10063), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9647), 
        .B2(n10051), .ZN(n9648) );
  OAI211_X1 U10916 ( .C1(n9650), .C2(n9759), .A(n9649), .B(n9648), .ZN(n9654)
         );
  INV_X1 U10917 ( .A(n9651), .ZN(n9659) );
  INV_X1 U10918 ( .A(n9655), .ZN(n9926) );
  OAI211_X1 U10919 ( .C1(n9659), .C2(n9926), .A(n9739), .B(n9652), .ZN(n9823)
         );
  NOR2_X1 U10920 ( .A1(n9823), .A2(n9740), .ZN(n9653) );
  AOI211_X1 U10921 ( .C1(n10050), .C2(n9655), .A(n9654), .B(n9653), .ZN(n9656)
         );
  OAI211_X1 U10922 ( .C1(n9825), .C2(n9746), .A(n9657), .B(n9656), .ZN(
        P1_U3270) );
  XOR2_X1 U10923 ( .A(n9664), .B(n9658), .Z(n9834) );
  INV_X1 U10924 ( .A(n9681), .ZN(n9660) );
  AOI211_X1 U10925 ( .C1(n9831), .C2(n9660), .A(n9750), .B(n9659), .ZN(n9830)
         );
  AOI22_X1 U10926 ( .A1(n10063), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9661), 
        .B2(n10051), .ZN(n9662) );
  OAI21_X1 U10927 ( .B1(n9663), .B2(n9752), .A(n9662), .ZN(n9671) );
  AOI21_X1 U10928 ( .B1(n9665), .B2(n9664), .A(n10068), .ZN(n9669) );
  OAI22_X1 U10929 ( .A1(n9692), .A2(n9877), .B1(n9666), .B2(n9879), .ZN(n9667)
         );
  AOI21_X1 U10930 ( .B1(n9669), .B2(n9668), .A(n9667), .ZN(n9833) );
  NOR2_X1 U10931 ( .A1(n9833), .A2(n10063), .ZN(n9670) );
  AOI211_X1 U10932 ( .C1(n9830), .C2(n10053), .A(n9671), .B(n9670), .ZN(n9672)
         );
  OAI21_X1 U10933 ( .B1(n9834), .B2(n9767), .A(n9672), .ZN(P1_U3271) );
  XOR2_X1 U10934 ( .A(n9673), .B(n9677), .Z(n9837) );
  INV_X1 U10935 ( .A(n9837), .ZN(n9688) );
  INV_X1 U10936 ( .A(n9674), .ZN(n9675) );
  AOI21_X1 U10937 ( .B1(n9512), .B2(n9676), .A(n9675), .ZN(n9678) );
  XNOR2_X1 U10938 ( .A(n9678), .B(n9677), .ZN(n9679) );
  OAI222_X1 U10939 ( .A1(n9877), .A2(n9845), .B1(n9879), .B2(n9680), .C1(n9679), .C2(n10068), .ZN(n9835) );
  INV_X1 U10940 ( .A(n9682), .ZN(n9931) );
  AOI211_X1 U10941 ( .C1(n9682), .C2(n9693), .A(n9750), .B(n9681), .ZN(n9836)
         );
  NAND2_X1 U10942 ( .A1(n9836), .A2(n10053), .ZN(n9685) );
  AOI22_X1 U10943 ( .A1(n10063), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9683), 
        .B2(n10051), .ZN(n9684) );
  OAI211_X1 U10944 ( .C1(n9931), .C2(n9752), .A(n9685), .B(n9684), .ZN(n9686)
         );
  AOI21_X1 U10945 ( .B1(n10056), .B2(n9835), .A(n9686), .ZN(n9687) );
  OAI21_X1 U10946 ( .B1(n9688), .B2(n9767), .A(n9687), .ZN(P1_U3272) );
  XNOR2_X1 U10947 ( .A(n9689), .B(n9690), .ZN(n9844) );
  XNOR2_X1 U10948 ( .A(n9512), .B(n9690), .ZN(n9691) );
  OAI222_X1 U10949 ( .A1(n9877), .A2(n9724), .B1(n9879), .B2(n9692), .C1(
        n10068), .C2(n9691), .ZN(n9840) );
  INV_X1 U10950 ( .A(n9842), .ZN(n9698) );
  INV_X1 U10951 ( .A(n9693), .ZN(n9694) );
  AOI211_X1 U10952 ( .C1(n9842), .C2(n9702), .A(n9750), .B(n9694), .ZN(n9841)
         );
  NAND2_X1 U10953 ( .A1(n9841), .A2(n10053), .ZN(n9697) );
  AOI22_X1 U10954 ( .A1(n10063), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9695), 
        .B2(n10051), .ZN(n9696) );
  OAI211_X1 U10955 ( .C1(n9698), .C2(n9752), .A(n9697), .B(n9696), .ZN(n9699)
         );
  AOI21_X1 U10956 ( .B1(n9840), .B2(n10056), .A(n9699), .ZN(n9700) );
  OAI21_X1 U10957 ( .B1(n9844), .B2(n9767), .A(n9700), .ZN(P1_U3273) );
  XOR2_X1 U10958 ( .A(n9710), .B(n9701), .Z(n9850) );
  INV_X1 U10959 ( .A(n9702), .ZN(n9703) );
  AOI211_X1 U10960 ( .C1(n9935), .C2(n9715), .A(n9750), .B(n9703), .ZN(n9846)
         );
  NOR2_X1 U10961 ( .A1(n4896), .A2(n9752), .ZN(n9709) );
  NAND2_X1 U10962 ( .A1(n9755), .A2(n9704), .ZN(n9707) );
  AOI22_X1 U10963 ( .A1(n10063), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9705), 
        .B2(n10051), .ZN(n9706) );
  OAI211_X1 U10964 ( .C1(n9845), .C2(n9759), .A(n9707), .B(n9706), .ZN(n9708)
         );
  AOI211_X1 U10965 ( .C1(n9846), .C2(n10053), .A(n9709), .B(n9708), .ZN(n9713)
         );
  XNOR2_X1 U10966 ( .A(n9711), .B(n9710), .ZN(n9848) );
  NAND2_X1 U10967 ( .A1(n9848), .A2(n9764), .ZN(n9712) );
  OAI211_X1 U10968 ( .C1(n9850), .C2(n9767), .A(n9713), .B(n9712), .ZN(
        P1_U3274) );
  XNOR2_X1 U10969 ( .A(n9714), .B(n9721), .ZN(n9856) );
  INV_X1 U10970 ( .A(n9738), .ZN(n9716) );
  OAI211_X1 U10971 ( .C1(n9716), .C2(n9940), .A(n9739), .B(n9715), .ZN(n9854)
         );
  INV_X1 U10972 ( .A(n9854), .ZN(n9729) );
  AOI22_X1 U10973 ( .A1(n10063), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9717), 
        .B2(n10051), .ZN(n9718) );
  OAI21_X1 U10974 ( .B1(n9940), .B2(n9752), .A(n9718), .ZN(n9728) );
  NAND2_X1 U10975 ( .A1(n9720), .A2(n9719), .ZN(n9723) );
  INV_X1 U10976 ( .A(n9721), .ZN(n9722) );
  XNOR2_X1 U10977 ( .A(n9723), .B(n9722), .ZN(n9726) );
  OAI22_X1 U10978 ( .A1(n9869), .A2(n9877), .B1(n9724), .B2(n9879), .ZN(n9725)
         );
  AOI21_X1 U10979 ( .B1(n9726), .B2(n10116), .A(n9725), .ZN(n9855) );
  NOR2_X1 U10980 ( .A1(n9855), .A2(n10063), .ZN(n9727) );
  AOI211_X1 U10981 ( .C1(n9729), .C2(n10053), .A(n9728), .B(n9727), .ZN(n9730)
         );
  OAI21_X1 U10982 ( .B1(n9856), .B2(n9767), .A(n9730), .ZN(P1_U3275) );
  XNOR2_X1 U10983 ( .A(n9732), .B(n9731), .ZN(n9864) );
  XNOR2_X1 U10984 ( .A(n9734), .B(n9733), .ZN(n9866) );
  NAND2_X1 U10985 ( .A1(n9866), .A2(n10059), .ZN(n9745) );
  NAND2_X1 U10986 ( .A1(n9755), .A2(n9735), .ZN(n9737) );
  AOI22_X1 U10987 ( .A1(n10063), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n5123), 
        .B2(n10051), .ZN(n9736) );
  OAI211_X1 U10988 ( .C1(n9860), .C2(n9759), .A(n9737), .B(n9736), .ZN(n9742)
         );
  OAI211_X1 U10989 ( .C1(n9944), .C2(n9749), .A(n9739), .B(n9738), .ZN(n9862)
         );
  NOR2_X1 U10990 ( .A1(n9862), .A2(n9740), .ZN(n9741) );
  AOI211_X1 U10991 ( .C1(n10050), .C2(n9743), .A(n9742), .B(n9741), .ZN(n9744)
         );
  OAI211_X1 U10992 ( .C1(n9864), .C2(n9746), .A(n9745), .B(n9744), .ZN(
        P1_U3276) );
  OAI21_X1 U10993 ( .B1(n4518), .B2(n9748), .A(n9747), .ZN(n9876) );
  AOI211_X1 U10994 ( .C1(n9872), .C2(n9751), .A(n9750), .B(n9749), .ZN(n9870)
         );
  INV_X1 U10995 ( .A(n9872), .ZN(n9753) );
  NOR2_X1 U10996 ( .A1(n9753), .A2(n9752), .ZN(n9761) );
  NAND2_X1 U10997 ( .A1(n9755), .A2(n9754), .ZN(n9758) );
  AOI22_X1 U10998 ( .A1(n10063), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9756), 
        .B2(n10051), .ZN(n9757) );
  OAI211_X1 U10999 ( .C1(n9869), .C2(n9759), .A(n9758), .B(n9757), .ZN(n9760)
         );
  AOI211_X1 U11000 ( .C1(n9870), .C2(n10053), .A(n9761), .B(n9760), .ZN(n9766)
         );
  XNOR2_X1 U11001 ( .A(n9763), .B(n9762), .ZN(n9873) );
  NAND2_X1 U11002 ( .A1(n9873), .A2(n9764), .ZN(n9765) );
  OAI211_X1 U11003 ( .C1(n9876), .C2(n9767), .A(n9766), .B(n9765), .ZN(
        P1_U3277) );
  NOR2_X1 U11004 ( .A1(n9769), .A2(n9768), .ZN(n9899) );
  MUX2_X1 U11005 ( .A(n9770), .B(n9899), .S(n10128), .Z(n9771) );
  OAI21_X1 U11006 ( .B1(n9902), .B2(n9889), .A(n9771), .ZN(P1_U3552) );
  NAND2_X1 U11007 ( .A1(n9772), .A2(n10100), .ZN(n9780) );
  OAI21_X1 U11008 ( .B1(n9774), .B2(n9877), .A(n9773), .ZN(n9776) );
  AOI211_X1 U11009 ( .C1(n10082), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9779)
         );
  MUX2_X1 U11010 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9903), .S(n10128), .Z(
        P1_U3551) );
  AOI22_X1 U11011 ( .A1(n10104), .A2(n9797), .B1(n9781), .B2(n10105), .ZN(
        n9783) );
  OAI211_X1 U11012 ( .C1(n9784), .C2(n10068), .A(n9783), .B(n9782), .ZN(n9785)
         );
  MUX2_X1 U11013 ( .A(n9787), .B(n9904), .S(n10128), .Z(n9788) );
  INV_X1 U11014 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9795) );
  AOI22_X1 U11015 ( .A1(n10104), .A2(n9806), .B1(n9789), .B2(n10105), .ZN(
        n9791) );
  OAI211_X1 U11016 ( .C1(n9792), .C2(n10068), .A(n9791), .B(n9790), .ZN(n9793)
         );
  AOI21_X1 U11017 ( .B1(n9794), .B2(n10100), .A(n9793), .ZN(n9908) );
  MUX2_X1 U11018 ( .A(n9795), .B(n9908), .S(n10128), .Z(n9796) );
  OAI21_X1 U11019 ( .B1(n9911), .B2(n9889), .A(n9796), .ZN(P1_U3549) );
  INV_X1 U11020 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9804) );
  AOI22_X1 U11021 ( .A1(n10104), .A2(n9798), .B1(n9797), .B2(n10105), .ZN(
        n9800) );
  OAI211_X1 U11022 ( .C1(n9801), .C2(n10068), .A(n9800), .B(n9799), .ZN(n9802)
         );
  AOI21_X1 U11023 ( .B1(n9803), .B2(n10100), .A(n9802), .ZN(n9912) );
  MUX2_X1 U11024 ( .A(n9804), .B(n9912), .S(n10128), .Z(n9805) );
  OAI21_X1 U11025 ( .B1(n9915), .B2(n9889), .A(n9805), .ZN(P1_U3548) );
  INV_X1 U11026 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9812) );
  AOI22_X1 U11027 ( .A1(n10105), .A2(n9806), .B1(n9821), .B2(n10104), .ZN(
        n9808) );
  OAI211_X1 U11028 ( .C1(n9809), .C2(n10068), .A(n9808), .B(n9807), .ZN(n9810)
         );
  AOI21_X1 U11029 ( .B1(n9811), .B2(n10100), .A(n9810), .ZN(n9916) );
  MUX2_X1 U11030 ( .A(n9812), .B(n9916), .S(n10128), .Z(n9813) );
  OAI21_X1 U11031 ( .B1(n9919), .B2(n9889), .A(n9813), .ZN(P1_U3547) );
  NOR2_X1 U11032 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  OAI21_X1 U11033 ( .B1(n9817), .B2(n10111), .A(n9816), .ZN(n9920) );
  MUX2_X1 U11034 ( .A(n9920), .B(P1_REG1_REG_24__SCAN_IN), .S(n10126), .Z(
        n9818) );
  AOI21_X1 U11035 ( .B1(n9819), .B2(n9922), .A(n9818), .ZN(n9820) );
  INV_X1 U11036 ( .A(n9820), .ZN(P1_U3546) );
  INV_X1 U11037 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U11038 ( .A1(n10104), .A2(n9822), .B1(n9821), .B2(n10105), .ZN(
        n9824) );
  OAI211_X1 U11039 ( .C1(n9825), .C2(n10068), .A(n9824), .B(n9823), .ZN(n9826)
         );
  AOI21_X1 U11040 ( .B1(n9827), .B2(n10100), .A(n9826), .ZN(n9924) );
  MUX2_X1 U11041 ( .A(n9828), .B(n9924), .S(n10128), .Z(n9829) );
  OAI21_X1 U11042 ( .B1(n9926), .B2(n9889), .A(n9829), .ZN(P1_U3545) );
  AOI21_X1 U11043 ( .B1(n10082), .B2(n9831), .A(n9830), .ZN(n9832) );
  OAI211_X1 U11044 ( .C1(n9834), .C2(n10111), .A(n9833), .B(n9832), .ZN(n9927)
         );
  MUX2_X1 U11045 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9927), .S(n10128), .Z(
        P1_U3544) );
  INV_X1 U11046 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9838) );
  AOI211_X1 U11047 ( .C1(n9837), .C2(n10100), .A(n9836), .B(n9835), .ZN(n9928)
         );
  MUX2_X1 U11048 ( .A(n9838), .B(n9928), .S(n10128), .Z(n9839) );
  OAI21_X1 U11049 ( .B1(n9931), .B2(n9889), .A(n9839), .ZN(P1_U3543) );
  AOI211_X1 U11050 ( .C1(n10082), .C2(n9842), .A(n9841), .B(n9840), .ZN(n9843)
         );
  OAI21_X1 U11051 ( .B1(n10111), .B2(n9844), .A(n9843), .ZN(n9932) );
  MUX2_X1 U11052 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9932), .S(n10128), .Z(
        P1_U3542) );
  OAI22_X1 U11053 ( .A1(n9860), .A2(n9877), .B1(n9845), .B2(n9879), .ZN(n9847)
         );
  AOI211_X1 U11054 ( .C1(n9848), .C2(n10116), .A(n9847), .B(n9846), .ZN(n9849)
         );
  OAI21_X1 U11055 ( .B1(n9850), .B2(n10111), .A(n9849), .ZN(n9933) );
  INV_X1 U11056 ( .A(n9933), .ZN(n9851) );
  MUX2_X1 U11057 ( .A(n9852), .B(n9851), .S(n10128), .Z(n9853) );
  OAI21_X1 U11058 ( .B1(n4896), .B2(n9889), .A(n9853), .ZN(P1_U3541) );
  OAI211_X1 U11059 ( .C1(n9856), .C2(n10111), .A(n9855), .B(n9854), .ZN(n9857)
         );
  INV_X1 U11060 ( .A(n9857), .ZN(n9938) );
  MUX2_X1 U11061 ( .A(n9858), .B(n9938), .S(n10128), .Z(n9859) );
  OAI21_X1 U11062 ( .B1(n9940), .B2(n9889), .A(n9859), .ZN(P1_U3540) );
  OAI22_X1 U11063 ( .A1(n9860), .A2(n9879), .B1(n9880), .B2(n9877), .ZN(n9861)
         );
  INV_X1 U11064 ( .A(n9861), .ZN(n9863) );
  OAI211_X1 U11065 ( .C1(n9864), .C2(n10068), .A(n9863), .B(n9862), .ZN(n9865)
         );
  AOI21_X1 U11066 ( .B1(n9866), .B2(n10100), .A(n9865), .ZN(n9941) );
  MUX2_X1 U11067 ( .A(n10307), .B(n9941), .S(n10128), .Z(n9867) );
  OAI21_X1 U11068 ( .B1(n9944), .B2(n9889), .A(n9867), .ZN(P1_U3539) );
  OAI22_X1 U11069 ( .A1(n9869), .A2(n9879), .B1(n9868), .B2(n9877), .ZN(n9871)
         );
  AOI211_X1 U11070 ( .C1(n10082), .C2(n9872), .A(n9871), .B(n9870), .ZN(n9875)
         );
  NAND2_X1 U11071 ( .A1(n9873), .A2(n10116), .ZN(n9874) );
  OAI211_X1 U11072 ( .C1(n9876), .C2(n10111), .A(n9875), .B(n9874), .ZN(n9945)
         );
  MUX2_X1 U11073 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9945), .S(n10128), .Z(
        P1_U3538) );
  OAI22_X1 U11074 ( .A1(n9880), .A2(n9879), .B1(n9878), .B2(n9877), .ZN(n9882)
         );
  AOI211_X1 U11075 ( .C1(n10116), .C2(n9883), .A(n9882), .B(n9881), .ZN(n9884)
         );
  OAI21_X1 U11076 ( .B1(n9885), .B2(n10111), .A(n9884), .ZN(n9886) );
  INV_X1 U11077 ( .A(n9886), .ZN(n9946) );
  MUX2_X1 U11078 ( .A(n9887), .B(n9946), .S(n10128), .Z(n9888) );
  OAI21_X1 U11079 ( .B1(n7788), .B2(n9889), .A(n9888), .ZN(P1_U3537) );
  AOI211_X1 U11080 ( .C1(n10082), .C2(n9892), .A(n9891), .B(n9890), .ZN(n9893)
         );
  OAI21_X1 U11081 ( .B1(n9894), .B2(n10111), .A(n9893), .ZN(n9949) );
  MUX2_X1 U11082 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9949), .S(n10128), .Z(
        P1_U3536) );
  MUX2_X1 U11083 ( .A(n9896), .B(n9895), .S(n10119), .Z(n9897) );
  OAI21_X1 U11084 ( .B1(n9898), .B2(n9948), .A(n9897), .ZN(P1_U3521) );
  MUX2_X1 U11085 ( .A(n9900), .B(n9899), .S(n10119), .Z(n9901) );
  OAI21_X1 U11086 ( .B1(n9902), .B2(n9948), .A(n9901), .ZN(P1_U3520) );
  INV_X1 U11087 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9905) );
  MUX2_X1 U11088 ( .A(n9905), .B(n9904), .S(n10119), .Z(n9906) );
  INV_X1 U11089 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9909) );
  MUX2_X1 U11090 ( .A(n9909), .B(n9908), .S(n10119), .Z(n9910) );
  OAI21_X1 U11091 ( .B1(n9911), .B2(n9948), .A(n9910), .ZN(P1_U3517) );
  INV_X1 U11092 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9913) );
  MUX2_X1 U11093 ( .A(n9913), .B(n9912), .S(n10119), .Z(n9914) );
  OAI21_X1 U11094 ( .B1(n9915), .B2(n9948), .A(n9914), .ZN(P1_U3516) );
  INV_X1 U11095 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9917) );
  MUX2_X1 U11096 ( .A(n9917), .B(n9916), .S(n10119), .Z(n9918) );
  OAI21_X1 U11097 ( .B1(n9919), .B2(n9948), .A(n9918), .ZN(P1_U3515) );
  MUX2_X1 U11098 ( .A(n9920), .B(P1_REG0_REG_24__SCAN_IN), .S(n10117), .Z(
        n9921) );
  AOI21_X1 U11099 ( .B1(n9936), .B2(n9922), .A(n9921), .ZN(n9923) );
  INV_X1 U11100 ( .A(n9923), .ZN(P1_U3514) );
  MUX2_X1 U11101 ( .A(n10409), .B(n9924), .S(n10119), .Z(n9925) );
  OAI21_X1 U11102 ( .B1(n9926), .B2(n9948), .A(n9925), .ZN(P1_U3513) );
  MUX2_X1 U11103 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9927), .S(n10119), .Z(
        P1_U3512) );
  INV_X1 U11104 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9929) );
  MUX2_X1 U11105 ( .A(n9929), .B(n9928), .S(n10119), .Z(n9930) );
  OAI21_X1 U11106 ( .B1(n9931), .B2(n9948), .A(n9930), .ZN(P1_U3511) );
  MUX2_X1 U11107 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9932), .S(n10119), .Z(
        P1_U3510) );
  MUX2_X1 U11108 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9933), .S(n10119), .Z(
        n9934) );
  AOI21_X1 U11109 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9937) );
  INV_X1 U11110 ( .A(n9937), .ZN(P1_U3509) );
  MUX2_X1 U11111 ( .A(n10457), .B(n9938), .S(n10119), .Z(n9939) );
  OAI21_X1 U11112 ( .B1(n9940), .B2(n9948), .A(n9939), .ZN(P1_U3507) );
  INV_X1 U11113 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9942) );
  MUX2_X1 U11114 ( .A(n9942), .B(n9941), .S(n10119), .Z(n9943) );
  OAI21_X1 U11115 ( .B1(n9944), .B2(n9948), .A(n9943), .ZN(P1_U3504) );
  MUX2_X1 U11116 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9945), .S(n10119), .Z(
        P1_U3501) );
  INV_X1 U11117 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10424) );
  MUX2_X1 U11118 ( .A(n10424), .B(n9946), .S(n10119), .Z(n9947) );
  OAI21_X1 U11119 ( .B1(n7788), .B2(n9948), .A(n9947), .ZN(P1_U3498) );
  MUX2_X1 U11120 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9949), .S(n10119), .Z(
        P1_U3495) );
  MUX2_X1 U11121 ( .A(P1_D_REG_1__SCAN_IN), .B(n9952), .S(n10065), .Z(P1_U3440) );
  MUX2_X1 U11122 ( .A(P1_D_REG_0__SCAN_IN), .B(n9953), .S(n10065), .Z(P1_U3439) );
  NOR2_X1 U11123 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n9955) );
  NAND4_X1 U11124 ( .A1(n9955), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .A4(n9954), .ZN(n9956) );
  OAI22_X1 U11125 ( .A1(n9957), .A2(n9956), .B1(n10458), .B2(n9971), .ZN(n9958) );
  AOI21_X1 U11126 ( .B1(n9960), .B2(n9959), .A(n9958), .ZN(n9961) );
  INV_X1 U11127 ( .A(n9961), .ZN(P1_U3324) );
  OAI222_X1 U11128 ( .A1(n9965), .A2(n9971), .B1(n9964), .B2(n9963), .C1(
        P1_U3086), .C2(n9962), .ZN(P1_U3325) );
  OAI222_X1 U11129 ( .A1(n9971), .A2(n9968), .B1(P1_U3086), .B2(n9967), .C1(
        n9964), .C2(n9966), .ZN(P1_U3326) );
  OAI222_X1 U11130 ( .A1(n9971), .A2(n9970), .B1(P1_U3086), .B2(n6443), .C1(
        n9964), .C2(n9969), .ZN(P1_U3327) );
  OAI222_X1 U11131 ( .A1(n9971), .A2(n9973), .B1(P1_U3086), .B2(n6541), .C1(
        n9964), .C2(n9972), .ZN(P1_U3328) );
  INV_X1 U11132 ( .A(n9974), .ZN(n9975) );
  MUX2_X1 U11133 ( .A(n9975), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI211_X1 U11134 ( .C1(n9978), .C2(n9977), .A(n10043), .B(n9976), .ZN(n9983)
         );
  OAI211_X1 U11135 ( .C1(n9981), .C2(n9980), .A(n10039), .B(n9979), .ZN(n9982)
         );
  OAI211_X1 U11136 ( .C1(n10027), .C2(n9984), .A(n9983), .B(n9982), .ZN(n9985)
         );
  AOI211_X1 U11137 ( .C1(n10030), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9986), .B(
        n9985), .ZN(n9987) );
  INV_X1 U11138 ( .A(n9987), .ZN(P1_U3251) );
  XNOR2_X1 U11139 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11140 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11141 ( .A(n9988), .ZN(n9993) );
  NAND2_X1 U11142 ( .A1(n6541), .A2(n6545), .ZN(n9991) );
  NAND2_X1 U11143 ( .A1(n9989), .A2(n9991), .ZN(n9990) );
  MUX2_X1 U11144 ( .A(n9991), .B(n9990), .S(P1_IR_REG_0__SCAN_IN), .Z(n9992)
         );
  NAND2_X1 U11145 ( .A1(n9993), .A2(n9992), .ZN(n9995) );
  AOI22_X1 U11146 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10030), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9994) );
  OAI21_X1 U11147 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(P1_U3243) );
  INV_X1 U11148 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10017) );
  MUX2_X1 U11149 ( .A(n6567), .B(P1_REG1_REG_4__SCAN_IN), .S(n10003), .Z(n9999) );
  INV_X1 U11150 ( .A(n9997), .ZN(n9998) );
  NAND2_X1 U11151 ( .A1(n9999), .A2(n9998), .ZN(n10001) );
  OAI211_X1 U11152 ( .C1(n10002), .C2(n10001), .A(n10043), .B(n10000), .ZN(
        n10011) );
  MUX2_X1 U11153 ( .A(n6577), .B(P1_REG2_REG_4__SCAN_IN), .S(n10003), .Z(
        n10006) );
  INV_X1 U11154 ( .A(n10004), .ZN(n10005) );
  NAND2_X1 U11155 ( .A1(n10006), .A2(n10005), .ZN(n10008) );
  OAI211_X1 U11156 ( .C1(n10009), .C2(n10008), .A(n10039), .B(n10007), .ZN(
        n10010) );
  OAI211_X1 U11157 ( .C1(n10027), .C2(n10012), .A(n10011), .B(n10010), .ZN(
        n10013) );
  NOR2_X1 U11158 ( .A1(n10014), .A2(n10013), .ZN(n10016) );
  OAI211_X1 U11159 ( .C1(n10017), .C2(n10048), .A(n10016), .B(n10015), .ZN(
        P1_U3247) );
  OAI211_X1 U11160 ( .C1(n10020), .C2(n10019), .A(n10039), .B(n10018), .ZN(
        n10025) );
  OAI211_X1 U11161 ( .C1(n10023), .C2(n10022), .A(n10043), .B(n10021), .ZN(
        n10024) );
  OAI211_X1 U11162 ( .C1(n10027), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10028) );
  AOI211_X1 U11163 ( .C1(n10030), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10029), 
        .B(n10028), .ZN(n10031) );
  INV_X1 U11164 ( .A(n10031), .ZN(P1_U3254) );
  NAND2_X1 U11165 ( .A1(n10033), .A2(n10032), .ZN(n10034) );
  NAND2_X1 U11166 ( .A1(n10035), .A2(n10034), .ZN(n10044) );
  OAI21_X1 U11167 ( .B1(n10038), .B2(n10037), .A(n10036), .ZN(n10040) );
  AOI222_X1 U11168 ( .A1(n10044), .A2(n10043), .B1(n10042), .B2(n10041), .C1(
        n10040), .C2(n10039), .ZN(n10046) );
  OAI211_X1 U11169 ( .C1(n10048), .C2(n10047), .A(n10046), .B(n10045), .ZN(
        P1_U3260) );
  NAND2_X1 U11170 ( .A1(n10050), .A2(n10049), .ZN(n10055) );
  AOI22_X1 U11171 ( .A1(n10053), .A2(n10052), .B1(n10051), .B2(n5954), .ZN(
        n10054) );
  OAI211_X1 U11172 ( .C1(n10057), .C2(n10056), .A(n10055), .B(n10054), .ZN(
        n10058) );
  AOI21_X1 U11173 ( .B1(n10060), .B2(n10059), .A(n10058), .ZN(n10061) );
  OAI21_X1 U11174 ( .B1(n10063), .B2(n10062), .A(n10061), .ZN(P1_U3290) );
  AND2_X1 U11175 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10066), .ZN(P1_U3294) );
  NOR2_X1 U11176 ( .A1(n10065), .A2(n10335), .ZN(P1_U3295) );
  AND2_X1 U11177 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10066), .ZN(P1_U3296) );
  NOR2_X1 U11178 ( .A1(n10065), .A2(n10064), .ZN(P1_U3297) );
  NOR2_X1 U11179 ( .A1(n10065), .A2(n10316), .ZN(P1_U3298) );
  AND2_X1 U11180 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10066), .ZN(P1_U3299) );
  AND2_X1 U11181 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10066), .ZN(P1_U3300) );
  AND2_X1 U11182 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10066), .ZN(P1_U3301) );
  AND2_X1 U11183 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10066), .ZN(P1_U3302) );
  INV_X1 U11184 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10475) );
  NOR2_X1 U11185 ( .A1(n10065), .A2(n10475), .ZN(P1_U3303) );
  AND2_X1 U11186 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10066), .ZN(P1_U3304) );
  AND2_X1 U11187 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10066), .ZN(P1_U3305) );
  NOR2_X1 U11188 ( .A1(n10065), .A2(n10272), .ZN(P1_U3306) );
  AND2_X1 U11189 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10066), .ZN(P1_U3307) );
  AND2_X1 U11190 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10066), .ZN(P1_U3308) );
  AND2_X1 U11191 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10066), .ZN(P1_U3309) );
  AND2_X1 U11192 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10066), .ZN(P1_U3310) );
  AND2_X1 U11193 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10066), .ZN(P1_U3311) );
  AND2_X1 U11194 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10066), .ZN(P1_U3312) );
  AND2_X1 U11195 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10066), .ZN(P1_U3313) );
  INV_X1 U11196 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10466) );
  NOR2_X1 U11197 ( .A1(n10065), .A2(n10466), .ZN(P1_U3314) );
  AND2_X1 U11198 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10066), .ZN(P1_U3315) );
  AND2_X1 U11199 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10066), .ZN(P1_U3316) );
  AND2_X1 U11200 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10066), .ZN(P1_U3317) );
  AND2_X1 U11201 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10066), .ZN(P1_U3318) );
  AND2_X1 U11202 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10066), .ZN(P1_U3319) );
  AND2_X1 U11203 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10066), .ZN(P1_U3320) );
  AND2_X1 U11204 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10066), .ZN(P1_U3321) );
  AND2_X1 U11205 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10066), .ZN(P1_U3322) );
  AND2_X1 U11206 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10066), .ZN(P1_U3323) );
  AOI21_X1 U11207 ( .B1(n10111), .B2(n10068), .A(n10067), .ZN(n10072) );
  INV_X1 U11208 ( .A(n10069), .ZN(n10070) );
  NOR3_X1 U11209 ( .A1(n10072), .A2(n10071), .A3(n10070), .ZN(n10120) );
  INV_X1 U11210 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U11211 ( .A1(n10119), .A2(n10120), .B1(n10073), .B2(n10117), .ZN(
        P1_U3453) );
  NAND2_X1 U11212 ( .A1(n10082), .A2(n10074), .ZN(n10075) );
  OAI211_X1 U11213 ( .C1(n10078), .C2(n10077), .A(n10076), .B(n10075), .ZN(
        n10080) );
  NOR2_X1 U11214 ( .A1(n10080), .A2(n10079), .ZN(n10121) );
  INV_X1 U11215 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10081) );
  AOI22_X1 U11216 ( .A1(n10119), .A2(n10121), .B1(n10081), .B2(n10117), .ZN(
        P1_U3456) );
  INV_X1 U11217 ( .A(n10082), .ZN(n10109) );
  INV_X1 U11218 ( .A(n10083), .ZN(n10084) );
  OAI21_X1 U11219 ( .B1(n10085), .B2(n10109), .A(n10084), .ZN(n10086) );
  AOI211_X1 U11220 ( .C1(n10100), .C2(n10088), .A(n10087), .B(n10086), .ZN(
        n10122) );
  INV_X1 U11221 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U11222 ( .A1(n10119), .A2(n10122), .B1(n10089), .B2(n10117), .ZN(
        P1_U3465) );
  OAI21_X1 U11223 ( .B1(n10091), .B2(n10109), .A(n10090), .ZN(n10093) );
  AOI211_X1 U11224 ( .C1(n10100), .C2(n10094), .A(n10093), .B(n10092), .ZN(
        n10124) );
  INV_X1 U11225 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U11226 ( .A1(n10119), .A2(n10124), .B1(n10095), .B2(n10117), .ZN(
        P1_U3471) );
  OAI21_X1 U11227 ( .B1(n10097), .B2(n10109), .A(n10096), .ZN(n10098) );
  AOI211_X1 U11228 ( .C1(n10101), .C2(n10100), .A(n10099), .B(n10098), .ZN(
        n10125) );
  INV_X1 U11229 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10102) );
  AOI22_X1 U11230 ( .A1(n10119), .A2(n10125), .B1(n10102), .B2(n10117), .ZN(
        P1_U3489) );
  AOI22_X1 U11231 ( .A1(n10106), .A2(n10105), .B1(n10104), .B2(n10103), .ZN(
        n10107) );
  OAI211_X1 U11232 ( .C1(n10110), .C2(n10109), .A(n10108), .B(n10107), .ZN(
        n10114) );
  NOR2_X1 U11233 ( .A1(n10112), .A2(n10111), .ZN(n10113) );
  AOI211_X1 U11234 ( .C1(n10116), .C2(n10115), .A(n10114), .B(n10113), .ZN(
        n10127) );
  INV_X1 U11235 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U11236 ( .A1(n10119), .A2(n10127), .B1(n10118), .B2(n10117), .ZN(
        P1_U3492) );
  AOI22_X1 U11237 ( .A1(n10128), .A2(n10120), .B1(n6545), .B2(n10126), .ZN(
        P1_U3522) );
  AOI22_X1 U11238 ( .A1(n10128), .A2(n10121), .B1(n5911), .B2(n10126), .ZN(
        P1_U3523) );
  AOI22_X1 U11239 ( .A1(n10128), .A2(n10122), .B1(n6567), .B2(n10126), .ZN(
        P1_U3526) );
  AOI22_X1 U11240 ( .A1(n10128), .A2(n10124), .B1(n10123), .B2(n10126), .ZN(
        P1_U3528) );
  AOI22_X1 U11241 ( .A1(n10128), .A2(n10125), .B1(n6131), .B2(n10126), .ZN(
        P1_U3534) );
  AOI22_X1 U11242 ( .A1(n10128), .A2(n10127), .B1(n6153), .B2(n10126), .ZN(
        P1_U3535) );
  INV_X1 U11243 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10152) );
  INV_X1 U11244 ( .A(n10129), .ZN(n10134) );
  OAI21_X1 U11245 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(n10133) );
  NAND2_X1 U11246 ( .A1(n10134), .A2(n10133), .ZN(n10140) );
  OAI211_X1 U11247 ( .C1(n10138), .C2(n10137), .A(n10136), .B(n10135), .ZN(
        n10139) );
  OAI211_X1 U11248 ( .C1(n10141), .C2(n10414), .A(n10140), .B(n10139), .ZN(
        n10142) );
  AOI21_X1 U11249 ( .B1(n10144), .B2(n10143), .A(n10142), .ZN(n10151) );
  OAI21_X1 U11250 ( .B1(n10147), .B2(n10146), .A(n10145), .ZN(n10148) );
  NAND2_X1 U11251 ( .A1(n10149), .A2(n10148), .ZN(n10150) );
  OAI211_X1 U11252 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10152), .A(n10151), .B(
        n10150), .ZN(P2_U3184) );
  INV_X1 U11253 ( .A(n10153), .ZN(n10157) );
  OAI22_X1 U11254 ( .A1(n10157), .A2(n10156), .B1(n10155), .B2(n10154), .ZN(
        n10158) );
  AOI211_X1 U11255 ( .C1(n10160), .C2(P2_REG3_REG_2__SCAN_IN), .A(n10159), .B(
        n10158), .ZN(n10162) );
  AOI22_X1 U11256 ( .A1(n10163), .A2(n6780), .B1(n10162), .B2(n10161), .ZN(
        P2_U3231) );
  INV_X1 U11257 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U11258 ( .A1(n10580), .A2(n10165), .B1(n10164), .B2(n10578), .ZN(
        P2_U3393) );
  INV_X1 U11259 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U11260 ( .A1(n10580), .A2(n10167), .B1(n10166), .B2(n10578), .ZN(
        P2_U3396) );
  INV_X1 U11261 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U11262 ( .A1(n10580), .A2(n10169), .B1(n10168), .B2(n10578), .ZN(
        P2_U3399) );
  INV_X1 U11263 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U11264 ( .A1(n10580), .A2(n10171), .B1(n10170), .B2(n10578), .ZN(
        P2_U3402) );
  INV_X1 U11265 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U11266 ( .A1(n10580), .A2(n10173), .B1(n10172), .B2(n10578), .ZN(
        P2_U3405) );
  INV_X1 U11267 ( .A(n10174), .ZN(n10175) );
  AOI22_X1 U11268 ( .A1(n10580), .A2(n10175), .B1(n5269), .B2(n10578), .ZN(
        P2_U3408) );
  AOI22_X1 U11269 ( .A1(n10580), .A2(n10176), .B1(n5297), .B2(n10578), .ZN(
        P2_U3411) );
  AOI22_X1 U11270 ( .A1(n10580), .A2(n10177), .B1(n5314), .B2(n10578), .ZN(
        P2_U3414) );
  INV_X1 U11271 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U11272 ( .A1(n10580), .A2(n10179), .B1(n10178), .B2(n10578), .ZN(
        P2_U3417) );
  AOI22_X1 U11273 ( .A1(n10580), .A2(n10180), .B1(n5362), .B2(n10578), .ZN(
        P2_U3420) );
  INV_X1 U11274 ( .A(n10181), .ZN(n10184) );
  AOI21_X1 U11275 ( .B1(n10186), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n10185), .ZN(
        n10183) );
  OAI22_X1 U11276 ( .A1(n10185), .A2(n10184), .B1(n10183), .B2(n10182), .ZN(
        ADD_1068_U5) );
  AOI21_X1 U11277 ( .B1(n10366), .B2(n10187), .A(n10186), .ZN(ADD_1068_U46) );
  NOR2_X1 U11278 ( .A1(n10189), .A2(n10188), .ZN(n10191) );
  XNOR2_X1 U11279 ( .A(n10191), .B(n10190), .ZN(ADD_1068_U55) );
  XNOR2_X1 U11280 ( .A(n10193), .B(n10192), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11281 ( .A(n10195), .B(n10194), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11282 ( .A(n10197), .B(n10196), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11283 ( .A(n10199), .B(n10198), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11284 ( .A(n10201), .B(n10200), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11285 ( .A(n10203), .B(n10202), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11286 ( .A(n10205), .B(n10204), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11287 ( .A(n10207), .B(n10206), .ZN(ADD_1068_U63) );
  AOI22_X1 U11288 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(keyinput225), .B1(
        P2_ADDR_REG_9__SCAN_IN), .B2(keyinput171), .ZN(n10208) );
  OAI221_X1 U11289 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(keyinput225), .C1(
        P2_ADDR_REG_9__SCAN_IN), .C2(keyinput171), .A(n10208), .ZN(n10215) );
  AOI22_X1 U11290 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput206), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(keyinput238), .ZN(n10209) );
  OAI221_X1 U11291 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput206), .C1(
        P2_DATAO_REG_3__SCAN_IN), .C2(keyinput238), .A(n10209), .ZN(n10214) );
  AOI22_X1 U11292 ( .A1(P1_REG0_REG_30__SCAN_IN), .A2(keyinput243), .B1(
        P1_REG3_REG_28__SCAN_IN), .B2(keyinput244), .ZN(n10210) );
  OAI221_X1 U11293 ( .B1(P1_REG0_REG_30__SCAN_IN), .B2(keyinput243), .C1(
        P1_REG3_REG_28__SCAN_IN), .C2(keyinput244), .A(n10210), .ZN(n10213) );
  AOI22_X1 U11294 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(keyinput241), .B1(
        P1_REG2_REG_23__SCAN_IN), .B2(keyinput164), .ZN(n10211) );
  OAI221_X1 U11295 ( .B1(P1_REG0_REG_11__SCAN_IN), .B2(keyinput241), .C1(
        P1_REG2_REG_23__SCAN_IN), .C2(keyinput164), .A(n10211), .ZN(n10212) );
  NOR4_X1 U11296 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n10243) );
  AOI22_X1 U11297 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(keyinput186), .B1(
        P2_REG1_REG_21__SCAN_IN), .B2(keyinput191), .ZN(n10216) );
  OAI221_X1 U11298 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(keyinput186), .C1(
        P2_REG1_REG_21__SCAN_IN), .C2(keyinput191), .A(n10216), .ZN(n10223) );
  AOI22_X1 U11299 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput234), .B1(
        P2_REG0_REG_28__SCAN_IN), .B2(keyinput220), .ZN(n10217) );
  OAI221_X1 U11300 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput234), .C1(
        P2_REG0_REG_28__SCAN_IN), .C2(keyinput220), .A(n10217), .ZN(n10222) );
  AOI22_X1 U11301 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(keyinput166), .B1(
        P2_REG1_REG_6__SCAN_IN), .B2(keyinput203), .ZN(n10218) );
  OAI221_X1 U11302 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(keyinput166), .C1(
        P2_REG1_REG_6__SCAN_IN), .C2(keyinput203), .A(n10218), .ZN(n10221) );
  AOI22_X1 U11303 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(keyinput219), .B1(
        P1_REG1_REG_13__SCAN_IN), .B2(keyinput231), .ZN(n10219) );
  OAI221_X1 U11304 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(keyinput219), .C1(
        P1_REG1_REG_13__SCAN_IN), .C2(keyinput231), .A(n10219), .ZN(n10220) );
  NOR4_X1 U11305 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10242) );
  AOI22_X1 U11306 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(keyinput170), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput139), .ZN(n10224) );
  OAI221_X1 U11307 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(keyinput170), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput139), .A(n10224), .ZN(n10231)
         );
  AOI22_X1 U11308 ( .A1(SI_31_), .A2(keyinput180), .B1(P2_IR_REG_31__SCAN_IN), 
        .B2(keyinput146), .ZN(n10225) );
  OAI221_X1 U11309 ( .B1(SI_31_), .B2(keyinput180), .C1(P2_IR_REG_31__SCAN_IN), 
        .C2(keyinput146), .A(n10225), .ZN(n10230) );
  AOI22_X1 U11310 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(keyinput128), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(keyinput224), .ZN(n10226) );
  OAI221_X1 U11311 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(keyinput128), .C1(
        P1_DATAO_REG_6__SCAN_IN), .C2(keyinput224), .A(n10226), .ZN(n10229) );
  AOI22_X1 U11312 ( .A1(SI_17_), .A2(keyinput187), .B1(P2_IR_REG_2__SCAN_IN), 
        .B2(keyinput245), .ZN(n10227) );
  OAI221_X1 U11313 ( .B1(SI_17_), .B2(keyinput187), .C1(P2_IR_REG_2__SCAN_IN), 
        .C2(keyinput245), .A(n10227), .ZN(n10228) );
  NOR4_X1 U11314 ( .A1(n10231), .A2(n10230), .A3(n10229), .A4(n10228), .ZN(
        n10241) );
  AOI22_X1 U11315 ( .A1(P2_REG0_REG_7__SCAN_IN), .A2(keyinput177), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput137), .ZN(n10232) );
  OAI221_X1 U11316 ( .B1(P2_REG0_REG_7__SCAN_IN), .B2(keyinput177), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput137), .A(n10232), .ZN(n10239) );
  AOI22_X1 U11317 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(keyinput173), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput182), .ZN(n10233) );
  OAI221_X1 U11318 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(keyinput173), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput182), .A(n10233), .ZN(n10238)
         );
  AOI22_X1 U11319 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(keyinput222), .B1(SI_29_), 
        .B2(keyinput210), .ZN(n10234) );
  OAI221_X1 U11320 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(keyinput222), .C1(SI_29_), .C2(keyinput210), .A(n10234), .ZN(n10237) );
  AOI22_X1 U11321 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(keyinput212), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(keyinput140), .ZN(n10235) );
  OAI221_X1 U11322 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(keyinput212), .C1(
        P1_DATAO_REG_5__SCAN_IN), .C2(keyinput140), .A(n10235), .ZN(n10236) );
  NOR4_X1 U11323 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10240) );
  NAND4_X1 U11324 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n10384) );
  AOI22_X1 U11325 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput235), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(keyinput211), .ZN(n10244) );
  OAI221_X1 U11326 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput235), .C1(
        P1_DATAO_REG_7__SCAN_IN), .C2(keyinput211), .A(n10244), .ZN(n10251) );
  AOI22_X1 U11327 ( .A1(P1_REG0_REG_15__SCAN_IN), .A2(keyinput174), .B1(
        P2_D_REG_30__SCAN_IN), .B2(keyinput154), .ZN(n10245) );
  OAI221_X1 U11328 ( .B1(P1_REG0_REG_15__SCAN_IN), .B2(keyinput174), .C1(
        P2_D_REG_30__SCAN_IN), .C2(keyinput154), .A(n10245), .ZN(n10250) );
  AOI22_X1 U11329 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(keyinput147), .B1(
        P1_REG3_REG_6__SCAN_IN), .B2(keyinput131), .ZN(n10246) );
  OAI221_X1 U11330 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(keyinput147), .C1(
        P1_REG3_REG_6__SCAN_IN), .C2(keyinput131), .A(n10246), .ZN(n10249) );
  AOI22_X1 U11331 ( .A1(P1_REG0_REG_23__SCAN_IN), .A2(keyinput253), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput167), .ZN(n10247) );
  OAI221_X1 U11332 ( .B1(P1_REG0_REG_23__SCAN_IN), .B2(keyinput253), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput167), .A(n10247), .ZN(n10248) );
  NOR4_X1 U11333 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10280) );
  AOI22_X1 U11334 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(keyinput240), .B1(
        P2_REG1_REG_27__SCAN_IN), .B2(keyinput216), .ZN(n10252) );
  OAI221_X1 U11335 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(keyinput240), .C1(
        P2_REG1_REG_27__SCAN_IN), .C2(keyinput216), .A(n10252), .ZN(n10259) );
  AOI22_X1 U11336 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(keyinput188), .B1(
        P2_IR_REG_28__SCAN_IN), .B2(keyinput178), .ZN(n10253) );
  OAI221_X1 U11337 ( .B1(P1_REG0_REG_10__SCAN_IN), .B2(keyinput188), .C1(
        P2_IR_REG_28__SCAN_IN), .C2(keyinput178), .A(n10253), .ZN(n10258) );
  AOI22_X1 U11338 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(keyinput202), .B1(
        P2_REG1_REG_13__SCAN_IN), .B2(keyinput141), .ZN(n10254) );
  OAI221_X1 U11339 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(keyinput202), .C1(
        P2_REG1_REG_13__SCAN_IN), .C2(keyinput141), .A(n10254), .ZN(n10257) );
  AOI22_X1 U11340 ( .A1(P1_REG2_REG_22__SCAN_IN), .A2(keyinput181), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput248), .ZN(n10255) );
  OAI221_X1 U11341 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(keyinput181), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput248), .A(n10255), .ZN(n10256) );
  NOR4_X1 U11342 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10279) );
  AOI22_X1 U11343 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(keyinput247), .B1(
        P2_D_REG_0__SCAN_IN), .B2(keyinput197), .ZN(n10260) );
  OAI221_X1 U11344 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(keyinput247), .C1(
        P2_D_REG_0__SCAN_IN), .C2(keyinput197), .A(n10260), .ZN(n10267) );
  AOI22_X1 U11345 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(keyinput189), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput160), .ZN(n10261) );
  OAI221_X1 U11346 ( .B1(P2_IR_REG_23__SCAN_IN), .B2(keyinput189), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput160), .A(n10261), .ZN(n10266) );
  AOI22_X1 U11347 ( .A1(P1_D_REG_22__SCAN_IN), .A2(keyinput249), .B1(
        P2_REG0_REG_30__SCAN_IN), .B2(keyinput208), .ZN(n10262) );
  OAI221_X1 U11348 ( .B1(P1_D_REG_22__SCAN_IN), .B2(keyinput249), .C1(
        P2_REG0_REG_30__SCAN_IN), .C2(keyinput208), .A(n10262), .ZN(n10265) );
  AOI22_X1 U11349 ( .A1(P1_D_REG_28__SCAN_IN), .A2(keyinput169), .B1(SI_4_), 
        .B2(keyinput129), .ZN(n10263) );
  OAI221_X1 U11350 ( .B1(P1_D_REG_28__SCAN_IN), .B2(keyinput169), .C1(SI_4_), 
        .C2(keyinput129), .A(n10263), .ZN(n10264) );
  NOR4_X1 U11351 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10278) );
  AOI22_X1 U11352 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput165), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput230), .ZN(n10268) );
  OAI221_X1 U11353 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput165), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput230), .A(n10268), .ZN(n10276) );
  AOI22_X1 U11354 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(keyinput215), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput255), .ZN(n10269) );
  OAI221_X1 U11355 ( .B1(P1_REG1_REG_28__SCAN_IN), .B2(keyinput215), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput255), .A(n10269), .ZN(n10275) );
  AOI22_X1 U11356 ( .A1(P1_REG0_REG_24__SCAN_IN), .A2(keyinput134), .B1(
        P2_D_REG_29__SCAN_IN), .B2(keyinput175), .ZN(n10270) );
  OAI221_X1 U11357 ( .B1(P1_REG0_REG_24__SCAN_IN), .B2(keyinput134), .C1(
        P2_D_REG_29__SCAN_IN), .C2(keyinput175), .A(n10270), .ZN(n10274) );
  AOI22_X1 U11358 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput144), .B1(n10272), 
        .B2(keyinput138), .ZN(n10271) );
  OAI221_X1 U11359 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput144), .C1(n10272), .C2(keyinput138), .A(n10271), .ZN(n10273) );
  NOR4_X1 U11360 ( .A1(n10276), .A2(n10275), .A3(n10274), .A4(n10273), .ZN(
        n10277) );
  NAND4_X1 U11361 ( .A1(n10280), .A2(n10279), .A3(n10278), .A4(n10277), .ZN(
        n10383) );
  INV_X1 U11362 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10422) );
  AOI22_X1 U11363 ( .A1(n10400), .A2(keyinput196), .B1(keyinput190), .B2(
        n10422), .ZN(n10281) );
  OAI221_X1 U11364 ( .B1(n10400), .B2(keyinput196), .C1(n10422), .C2(
        keyinput190), .A(n10281), .ZN(n10291) );
  INV_X1 U11365 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U11366 ( .A1(n6046), .A2(keyinput193), .B1(keyinput226), .B2(n10283), .ZN(n10282) );
  OAI221_X1 U11367 ( .B1(n6046), .B2(keyinput193), .C1(n10283), .C2(
        keyinput226), .A(n10282), .ZN(n10290) );
  AOI22_X1 U11368 ( .A1(n10285), .A2(keyinput213), .B1(n8088), .B2(keyinput184), .ZN(n10284) );
  OAI221_X1 U11369 ( .B1(n10285), .B2(keyinput213), .C1(n8088), .C2(
        keyinput184), .A(n10284), .ZN(n10289) );
  XNOR2_X1 U11370 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput198), .ZN(n10287)
         );
  XNOR2_X1 U11371 ( .A(keyinput136), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n10286)
         );
  NAND2_X1 U11372 ( .A1(n10287), .A2(n10286), .ZN(n10288) );
  NOR4_X1 U11373 ( .A1(n10291), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10328) );
  AOI22_X1 U11374 ( .A1(n10458), .A2(keyinput221), .B1(keyinput223), .B2(
        n10293), .ZN(n10292) );
  OAI221_X1 U11375 ( .B1(n10458), .B2(keyinput221), .C1(n10293), .C2(
        keyinput223), .A(n10292), .ZN(n10298) );
  AOI22_X1 U11376 ( .A1(n10295), .A2(keyinput172), .B1(n10469), .B2(
        keyinput233), .ZN(n10294) );
  OAI221_X1 U11377 ( .B1(n10295), .B2(keyinput172), .C1(n10469), .C2(
        keyinput233), .A(n10294), .ZN(n10297) );
  XOR2_X1 U11378 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput183), .Z(n10296) );
  OR3_X1 U11379 ( .A1(n10298), .A2(n10297), .A3(n10296), .ZN(n10303) );
  AOI22_X1 U11380 ( .A1(n10300), .A2(keyinput161), .B1(keyinput239), .B2(
        n10414), .ZN(n10299) );
  OAI221_X1 U11381 ( .B1(n10300), .B2(keyinput161), .C1(n10414), .C2(
        keyinput239), .A(n10299), .ZN(n10302) );
  XNOR2_X1 U11382 ( .A(n10396), .B(keyinput130), .ZN(n10301) );
  NOR3_X1 U11383 ( .A1(n10303), .A2(n10302), .A3(n10301), .ZN(n10327) );
  INV_X1 U11384 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U11385 ( .A1(n10470), .A2(keyinput155), .B1(keyinput168), .B2(
        n10305), .ZN(n10304) );
  OAI221_X1 U11386 ( .B1(n10470), .B2(keyinput155), .C1(n10305), .C2(
        keyinput168), .A(n10304), .ZN(n10314) );
  INV_X1 U11387 ( .A(SI_12_), .ZN(n10440) );
  AOI22_X1 U11388 ( .A1(n10307), .A2(keyinput135), .B1(n10440), .B2(
        keyinput252), .ZN(n10306) );
  OAI221_X1 U11389 ( .B1(n10307), .B2(keyinput135), .C1(n10440), .C2(
        keyinput252), .A(n10306), .ZN(n10313) );
  XNOR2_X1 U11390 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(keyinput201), .ZN(n10311)
         );
  XNOR2_X1 U11391 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput242), .ZN(n10310)
         );
  XNOR2_X1 U11392 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput209), .ZN(n10309)
         );
  XNOR2_X1 U11393 ( .A(P1_REG0_REG_18__SCAN_IN), .B(keyinput185), .ZN(n10308)
         );
  NAND4_X1 U11394 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10312) );
  NOR3_X1 U11395 ( .A1(n10314), .A2(n10313), .A3(n10312), .ZN(n10326) );
  AOI22_X1 U11396 ( .A1(n5362), .A2(keyinput227), .B1(keyinput163), .B2(n10316), .ZN(n10315) );
  OAI221_X1 U11397 ( .B1(n5362), .B2(keyinput227), .C1(n10316), .C2(
        keyinput163), .A(n10315), .ZN(n10324) );
  AOI22_X1 U11398 ( .A1(n10454), .A2(keyinput179), .B1(n7389), .B2(keyinput217), .ZN(n10317) );
  OAI221_X1 U11399 ( .B1(n10454), .B2(keyinput179), .C1(n7389), .C2(
        keyinput217), .A(n10317), .ZN(n10323) );
  AOI22_X1 U11400 ( .A1(n10319), .A2(keyinput254), .B1(keyinput194), .B2(
        n10489), .ZN(n10318) );
  OAI221_X1 U11401 ( .B1(n10319), .B2(keyinput254), .C1(n10489), .C2(
        keyinput194), .A(n10318), .ZN(n10322) );
  AOI22_X1 U11402 ( .A1(n7087), .A2(keyinput145), .B1(n8053), .B2(keyinput158), 
        .ZN(n10320) );
  OAI221_X1 U11403 ( .B1(n7087), .B2(keyinput145), .C1(n8053), .C2(keyinput158), .A(n10320), .ZN(n10321) );
  NOR4_X1 U11404 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10325) );
  NAND4_X1 U11405 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10382) );
  AOI22_X1 U11406 ( .A1(n8812), .A2(keyinput246), .B1(n10330), .B2(keyinput200), .ZN(n10329) );
  OAI221_X1 U11407 ( .B1(n8812), .B2(keyinput246), .C1(n10330), .C2(
        keyinput200), .A(n10329), .ZN(n10333) );
  XOR2_X1 U11408 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput204), .Z(n10332) );
  XNOR2_X1 U11409 ( .A(n10411), .B(keyinput205), .ZN(n10331) );
  OR3_X1 U11410 ( .A1(n10333), .A2(n10332), .A3(n10331), .ZN(n10341) );
  AOI22_X1 U11411 ( .A1(n8639), .A2(keyinput195), .B1(keyinput142), .B2(n10335), .ZN(n10334) );
  OAI221_X1 U11412 ( .B1(n8639), .B2(keyinput195), .C1(n10335), .C2(
        keyinput142), .A(n10334), .ZN(n10340) );
  INV_X1 U11413 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U11414 ( .A1(n10338), .A2(keyinput143), .B1(keyinput237), .B2(
        n10337), .ZN(n10336) );
  OAI221_X1 U11415 ( .B1(n10338), .B2(keyinput143), .C1(n10337), .C2(
        keyinput237), .A(n10336), .ZN(n10339) );
  NOR3_X1 U11416 ( .A1(n10341), .A2(n10340), .A3(n10339), .ZN(n10380) );
  AOI22_X1 U11417 ( .A1(n10408), .A2(keyinput236), .B1(n10438), .B2(
        keyinput156), .ZN(n10342) );
  OAI221_X1 U11418 ( .B1(n10408), .B2(keyinput236), .C1(n10438), .C2(
        keyinput156), .A(n10342), .ZN(n10352) );
  AOI22_X1 U11419 ( .A1(n10344), .A2(keyinput162), .B1(keyinput148), .B2(
        n10415), .ZN(n10343) );
  OAI221_X1 U11420 ( .B1(n10344), .B2(keyinput162), .C1(n10415), .C2(
        keyinput148), .A(n10343), .ZN(n10351) );
  AOI22_X1 U11421 ( .A1(n10347), .A2(keyinput192), .B1(keyinput132), .B2(
        n10346), .ZN(n10345) );
  OAI221_X1 U11422 ( .B1(n10347), .B2(keyinput192), .C1(n10346), .C2(
        keyinput132), .A(n10345), .ZN(n10350) );
  INV_X1 U11423 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10476) );
  AOI22_X1 U11424 ( .A1(n10476), .A2(keyinput232), .B1(n5864), .B2(keyinput149), .ZN(n10348) );
  OAI221_X1 U11425 ( .B1(n10476), .B2(keyinput232), .C1(n5864), .C2(
        keyinput149), .A(n10348), .ZN(n10349) );
  NOR4_X1 U11426 ( .A1(n10352), .A2(n10351), .A3(n10350), .A4(n10349), .ZN(
        n10379) );
  INV_X1 U11427 ( .A(SI_13_), .ZN(n10425) );
  AOI22_X1 U11428 ( .A1(n10354), .A2(keyinput251), .B1(keyinput207), .B2(
        n10425), .ZN(n10353) );
  OAI221_X1 U11429 ( .B1(n10354), .B2(keyinput251), .C1(n10425), .C2(
        keyinput207), .A(n10353), .ZN(n10364) );
  AOI22_X1 U11430 ( .A1(n10357), .A2(keyinput157), .B1(n10356), .B2(
        keyinput199), .ZN(n10355) );
  OAI221_X1 U11431 ( .B1(n10357), .B2(keyinput157), .C1(n10356), .C2(
        keyinput199), .A(n10355), .ZN(n10363) );
  XNOR2_X1 U11432 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput250), .ZN(n10361)
         );
  XNOR2_X1 U11433 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput151), .ZN(n10360) );
  XNOR2_X1 U11434 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput150), .ZN(n10359) );
  XNOR2_X1 U11435 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput153), .ZN(n10358)
         );
  NAND4_X1 U11436 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10362) );
  NOR3_X1 U11437 ( .A1(n10364), .A2(n10363), .A3(n10362), .ZN(n10378) );
  INV_X1 U11438 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U11439 ( .A1(n10367), .A2(keyinput133), .B1(keyinput152), .B2(
        n10366), .ZN(n10365) );
  OAI221_X1 U11440 ( .B1(n10367), .B2(keyinput133), .C1(n10366), .C2(
        keyinput152), .A(n10365), .ZN(n10376) );
  AOI22_X1 U11441 ( .A1(n10466), .A2(keyinput176), .B1(n10369), .B2(
        keyinput159), .ZN(n10368) );
  OAI221_X1 U11442 ( .B1(n10466), .B2(keyinput176), .C1(n10369), .C2(
        keyinput159), .A(n10368), .ZN(n10375) );
  AOI22_X1 U11443 ( .A1(n5299), .A2(keyinput218), .B1(n10421), .B2(keyinput229), .ZN(n10370) );
  OAI221_X1 U11444 ( .B1(n5299), .B2(keyinput218), .C1(n10421), .C2(
        keyinput229), .A(n10370), .ZN(n10374) );
  AOI22_X1 U11445 ( .A1(n10372), .A2(keyinput228), .B1(n10473), .B2(
        keyinput214), .ZN(n10371) );
  OAI221_X1 U11446 ( .B1(n10372), .B2(keyinput228), .C1(n10473), .C2(
        keyinput214), .A(n10371), .ZN(n10373) );
  NOR4_X1 U11447 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10377) );
  NAND4_X1 U11448 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10381) );
  NOR4_X1 U11449 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10577) );
  AOI22_X1 U11450 ( .A1(P1_D_REG_19__SCAN_IN), .A2(keyinput10), .B1(
        P2_REG1_REG_13__SCAN_IN), .B2(keyinput13), .ZN(n10385) );
  OAI221_X1 U11451 ( .B1(P1_D_REG_19__SCAN_IN), .B2(keyinput10), .C1(
        P2_REG1_REG_13__SCAN_IN), .C2(keyinput13), .A(n10385), .ZN(n10393) );
  AOI22_X1 U11452 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(keyinput19), .B1(SI_17_), 
        .B2(keyinput59), .ZN(n10386) );
  OAI221_X1 U11453 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(keyinput19), .C1(SI_17_), 
        .C2(keyinput59), .A(n10386), .ZN(n10392) );
  AOI22_X1 U11454 ( .A1(P1_D_REG_30__SCAN_IN), .A2(keyinput14), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput122), .ZN(n10387) );
  OAI221_X1 U11455 ( .B1(P1_D_REG_30__SCAN_IN), .B2(keyinput14), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput122), .A(n10387), .ZN(n10391)
         );
  AOI22_X1 U11456 ( .A1(n8005), .A2(keyinput52), .B1(n10389), .B2(keyinput102), 
        .ZN(n10388) );
  OAI221_X1 U11457 ( .B1(n8005), .B2(keyinput52), .C1(n10389), .C2(keyinput102), .A(n10388), .ZN(n10390) );
  NOR4_X1 U11458 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n10436) );
  AOI22_X1 U11459 ( .A1(n5189), .A2(keyinput117), .B1(keyinput84), .B2(n5954), 
        .ZN(n10394) );
  OAI221_X1 U11460 ( .B1(n5189), .B2(keyinput117), .C1(n5954), .C2(keyinput84), 
        .A(n10394), .ZN(n10406) );
  AOI22_X1 U11461 ( .A1(n10397), .A2(keyinput80), .B1(n10396), .B2(keyinput2), 
        .ZN(n10395) );
  OAI221_X1 U11462 ( .B1(n10397), .B2(keyinput80), .C1(n10396), .C2(keyinput2), 
        .A(n10395), .ZN(n10405) );
  AOI22_X1 U11463 ( .A1(n10400), .A2(keyinput68), .B1(n10399), .B2(keyinput88), 
        .ZN(n10398) );
  OAI221_X1 U11464 ( .B1(n10400), .B2(keyinput68), .C1(n10399), .C2(keyinput88), .A(n10398), .ZN(n10404) );
  XNOR2_X1 U11465 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput23), .ZN(n10402) );
  XNOR2_X1 U11466 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput16), .ZN(n10401) );
  NAND2_X1 U11467 ( .A1(n10402), .A2(n10401), .ZN(n10403) );
  NOR4_X1 U11468 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n10435) );
  AOI22_X1 U11469 ( .A1(n10409), .A2(keyinput125), .B1(n10408), .B2(
        keyinput108), .ZN(n10407) );
  OAI221_X1 U11470 ( .B1(n10409), .B2(keyinput125), .C1(n10408), .C2(
        keyinput108), .A(n10407), .ZN(n10419) );
  AOI22_X1 U11471 ( .A1(n8088), .A2(keyinput56), .B1(keyinput77), .B2(n10411), 
        .ZN(n10410) );
  OAI221_X1 U11472 ( .B1(n8088), .B2(keyinput56), .C1(n10411), .C2(keyinput77), 
        .A(n10410), .ZN(n10418) );
  AOI22_X1 U11473 ( .A1(n8812), .A2(keyinput118), .B1(n5813), .B2(keyinput69), 
        .ZN(n10412) );
  OAI221_X1 U11474 ( .B1(n8812), .B2(keyinput118), .C1(n5813), .C2(keyinput69), 
        .A(n10412), .ZN(n10417) );
  AOI22_X1 U11475 ( .A1(n10415), .A2(keyinput20), .B1(keyinput111), .B2(n10414), .ZN(n10413) );
  OAI221_X1 U11476 ( .B1(n10415), .B2(keyinput20), .C1(n10414), .C2(
        keyinput111), .A(n10413), .ZN(n10416) );
  NOR4_X1 U11477 ( .A1(n10419), .A2(n10418), .A3(n10417), .A4(n10416), .ZN(
        n10434) );
  AOI22_X1 U11478 ( .A1(n10422), .A2(keyinput62), .B1(n10421), .B2(keyinput101), .ZN(n10420) );
  OAI221_X1 U11479 ( .B1(n10422), .B2(keyinput62), .C1(n10421), .C2(
        keyinput101), .A(n10420), .ZN(n10432) );
  AOI22_X1 U11480 ( .A1(n10425), .A2(keyinput79), .B1(keyinput46), .B2(n10424), 
        .ZN(n10423) );
  OAI221_X1 U11481 ( .B1(n10425), .B2(keyinput79), .C1(n10424), .C2(keyinput46), .A(n10423), .ZN(n10431) );
  XNOR2_X1 U11482 ( .A(SI_4_), .B(keyinput1), .ZN(n10429) );
  XNOR2_X1 U11483 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput127), .ZN(n10428) );
  XNOR2_X1 U11484 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput50), .ZN(n10427) );
  XNOR2_X1 U11485 ( .A(keyinput91), .B(P1_REG2_REG_0__SCAN_IN), .ZN(n10426) );
  NAND4_X1 U11486 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10430) );
  NOR3_X1 U11487 ( .A1(n10432), .A2(n10431), .A3(n10430), .ZN(n10433) );
  NAND4_X1 U11488 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .ZN(
        n10576) );
  AOI22_X1 U11489 ( .A1(n10438), .A2(keyinput28), .B1(keyinput3), .B2(n6008), 
        .ZN(n10437) );
  OAI221_X1 U11490 ( .B1(n10438), .B2(keyinput28), .C1(n6008), .C2(keyinput3), 
        .A(n10437), .ZN(n10448) );
  XNOR2_X1 U11491 ( .A(n10439), .B(keyinput70), .ZN(n10447) );
  XNOR2_X1 U11492 ( .A(keyinput124), .B(n10440), .ZN(n10446) );
  XNOR2_X1 U11493 ( .A(P2_REG0_REG_28__SCAN_IN), .B(keyinput92), .ZN(n10444)
         );
  XNOR2_X1 U11494 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput81), .ZN(n10443) );
  XNOR2_X1 U11495 ( .A(P1_REG1_REG_28__SCAN_IN), .B(keyinput87), .ZN(n10442)
         );
  XNOR2_X1 U11496 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput78), .ZN(n10441) );
  NAND4_X1 U11497 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        n10445) );
  NOR4_X1 U11498 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10499) );
  AOI22_X1 U11499 ( .A1(n10451), .A2(keyinput106), .B1(keyinput74), .B2(n10450), .ZN(n10449) );
  OAI221_X1 U11500 ( .B1(n10451), .B2(keyinput106), .C1(n10450), .C2(
        keyinput74), .A(n10449), .ZN(n10464) );
  AOI22_X1 U11501 ( .A1(n10454), .A2(keyinput51), .B1(n10453), .B2(keyinput25), 
        .ZN(n10452) );
  OAI221_X1 U11502 ( .B1(n10454), .B2(keyinput51), .C1(n10453), .C2(keyinput25), .A(n10452), .ZN(n10463) );
  AOI22_X1 U11503 ( .A1(n10457), .A2(keyinput57), .B1(n10456), .B2(keyinput39), 
        .ZN(n10455) );
  OAI221_X1 U11504 ( .B1(n10457), .B2(keyinput57), .C1(n10456), .C2(keyinput39), .A(n10455), .ZN(n10462) );
  XOR2_X1 U11505 ( .A(n10458), .B(keyinput93), .Z(n10460) );
  XNOR2_X1 U11506 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput107), .ZN(n10459) );
  NAND2_X1 U11507 ( .A1(n10460), .A2(n10459), .ZN(n10461) );
  NOR4_X1 U11508 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10498) );
  AOI22_X1 U11509 ( .A1(n10467), .A2(keyinput6), .B1(n10466), .B2(keyinput48), 
        .ZN(n10465) );
  OAI221_X1 U11510 ( .B1(n10467), .B2(keyinput6), .C1(n10466), .C2(keyinput48), 
        .A(n10465), .ZN(n10480) );
  AOI22_X1 U11511 ( .A1(n10470), .A2(keyinput27), .B1(n10469), .B2(keyinput105), .ZN(n10468) );
  OAI221_X1 U11512 ( .B1(n10470), .B2(keyinput27), .C1(n10469), .C2(
        keyinput105), .A(n10468), .ZN(n10479) );
  AOI22_X1 U11513 ( .A1(n10473), .A2(keyinput86), .B1(keyinput0), .B2(n10472), 
        .ZN(n10471) );
  OAI221_X1 U11514 ( .B1(n10473), .B2(keyinput86), .C1(n10472), .C2(keyinput0), 
        .A(n10471), .ZN(n10478) );
  AOI22_X1 U11515 ( .A1(n10476), .A2(keyinput104), .B1(n10475), .B2(
        keyinput121), .ZN(n10474) );
  OAI221_X1 U11516 ( .B1(n10476), .B2(keyinput104), .C1(n10475), .C2(
        keyinput121), .A(n10474), .ZN(n10477) );
  NOR4_X1 U11517 ( .A1(n10480), .A2(n10479), .A3(n10478), .A4(n10477), .ZN(
        n10497) );
  AOI22_X1 U11518 ( .A1(n10483), .A2(keyinput110), .B1(keyinput43), .B2(n10482), .ZN(n10481) );
  OAI221_X1 U11519 ( .B1(n10483), .B2(keyinput110), .C1(n10482), .C2(
        keyinput43), .A(n10481), .ZN(n10495) );
  AOI22_X1 U11520 ( .A1(n10486), .A2(keyinput47), .B1(keyinput42), .B2(n10485), 
        .ZN(n10484) );
  OAI221_X1 U11521 ( .B1(n10486), .B2(keyinput47), .C1(n10485), .C2(keyinput42), .A(n10484), .ZN(n10494) );
  INV_X1 U11522 ( .A(SI_29_), .ZN(n10488) );
  AOI22_X1 U11523 ( .A1(n10489), .A2(keyinput66), .B1(n10488), .B2(keyinput82), 
        .ZN(n10487) );
  OAI221_X1 U11524 ( .B1(n10489), .B2(keyinput66), .C1(n10488), .C2(keyinput82), .A(n10487), .ZN(n10493) );
  XNOR2_X1 U11525 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput114), .ZN(n10491)
         );
  XNOR2_X1 U11526 ( .A(SI_25_), .B(keyinput71), .ZN(n10490) );
  NAND2_X1 U11527 ( .A1(n10491), .A2(n10490), .ZN(n10492) );
  NOR4_X1 U11528 ( .A1(n10495), .A2(n10494), .A3(n10493), .A4(n10492), .ZN(
        n10496) );
  NAND4_X1 U11529 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10575) );
  OAI22_X1 U11530 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(keyinput31), .B1(
        keyinput36), .B2(P1_REG2_REG_23__SCAN_IN), .ZN(n10500) );
  AOI221_X1 U11531 ( .B1(P1_DATAO_REG_21__SCAN_IN), .B2(keyinput31), .C1(
        P1_REG2_REG_23__SCAN_IN), .C2(keyinput36), .A(n10500), .ZN(n10507) );
  OAI22_X1 U11532 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput54), .B1(
        keyinput89), .B2(P2_REG2_REG_8__SCAN_IN), .ZN(n10501) );
  AOI221_X1 U11533 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput54), .C1(
        P2_REG2_REG_8__SCAN_IN), .C2(keyinput89), .A(n10501), .ZN(n10506) );
  OAI22_X1 U11534 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput76), .B1(
        P2_ADDR_REG_0__SCAN_IN), .B2(keyinput24), .ZN(n10502) );
  AOI221_X1 U11535 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput76), .C1(
        keyinput24), .C2(P2_ADDR_REG_0__SCAN_IN), .A(n10502), .ZN(n10505) );
  OAI22_X1 U11536 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput9), .B1(
        P2_REG1_REG_24__SCAN_IN), .B2(keyinput44), .ZN(n10503) );
  AOI221_X1 U11537 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput9), .C1(
        keyinput44), .C2(P2_REG1_REG_24__SCAN_IN), .A(n10503), .ZN(n10504) );
  NAND4_X1 U11538 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10504), .ZN(
        n10535) );
  OAI22_X1 U11539 ( .A1(P2_D_REG_30__SCAN_IN), .A2(keyinput26), .B1(
        P2_ADDR_REG_10__SCAN_IN), .B2(keyinput95), .ZN(n10508) );
  AOI221_X1 U11540 ( .B1(P2_D_REG_30__SCAN_IN), .B2(keyinput26), .C1(
        keyinput95), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n10508), .ZN(n10515) );
  OAI22_X1 U11541 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(keyinput96), .B1(
        keyinput103), .B2(P1_REG1_REG_13__SCAN_IN), .ZN(n10509) );
  AOI221_X1 U11542 ( .B1(P1_DATAO_REG_6__SCAN_IN), .B2(keyinput96), .C1(
        P1_REG1_REG_13__SCAN_IN), .C2(keyinput103), .A(n10509), .ZN(n10514) );
  OAI22_X1 U11543 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput85), .B1(
        keyinput7), .B2(P1_REG1_REG_17__SCAN_IN), .ZN(n10510) );
  AOI221_X1 U11544 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput85), .C1(
        P1_REG1_REG_17__SCAN_IN), .C2(keyinput7), .A(n10510), .ZN(n10513) );
  OAI22_X1 U11545 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(keyinput61), .B1(
        P2_REG2_REG_2__SCAN_IN), .B2(keyinput94), .ZN(n10511) );
  AOI221_X1 U11546 ( .B1(P2_IR_REG_23__SCAN_IN), .B2(keyinput61), .C1(
        keyinput94), .C2(P2_REG2_REG_2__SCAN_IN), .A(n10511), .ZN(n10512) );
  NAND4_X1 U11547 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10534) );
  OAI22_X1 U11548 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput11), .B1(
        P1_REG0_REG_2__SCAN_IN), .B2(keyinput109), .ZN(n10516) );
  AOI221_X1 U11549 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput11), .C1(
        keyinput109), .C2(P1_REG0_REG_2__SCAN_IN), .A(n10516), .ZN(n10523) );
  OAI22_X1 U11550 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(keyinput60), .B1(
        P2_ADDR_REG_17__SCAN_IN), .B2(keyinput40), .ZN(n10517) );
  AOI221_X1 U11551 ( .B1(P1_REG0_REG_10__SCAN_IN), .B2(keyinput60), .C1(
        keyinput40), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n10517), .ZN(n10522) );
  OAI22_X1 U11552 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(keyinput12), .B1(
        keyinput116), .B2(P1_REG3_REG_28__SCAN_IN), .ZN(n10518) );
  AOI221_X1 U11553 ( .B1(P1_DATAO_REG_5__SCAN_IN), .B2(keyinput12), .C1(
        P1_REG3_REG_28__SCAN_IN), .C2(keyinput116), .A(n10518), .ZN(n10521) );
  OAI22_X1 U11554 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput72), .B1(
        keyinput17), .B2(P1_REG2_REG_5__SCAN_IN), .ZN(n10519) );
  AOI221_X1 U11555 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput72), .C1(
        P1_REG2_REG_5__SCAN_IN), .C2(keyinput17), .A(n10519), .ZN(n10520) );
  NAND4_X1 U11556 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n10533) );
  OAI22_X1 U11557 ( .A1(P2_REG1_REG_21__SCAN_IN), .A2(keyinput63), .B1(
        keyinput65), .B2(P1_REG3_REG_8__SCAN_IN), .ZN(n10524) );
  AOI221_X1 U11558 ( .B1(P2_REG1_REG_21__SCAN_IN), .B2(keyinput63), .C1(
        P1_REG3_REG_8__SCAN_IN), .C2(keyinput65), .A(n10524), .ZN(n10531) );
  OAI22_X1 U11559 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(keyinput45), .B1(
        P1_REG0_REG_11__SCAN_IN), .B2(keyinput113), .ZN(n10525) );
  AOI221_X1 U11560 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(keyinput45), .C1(
        keyinput113), .C2(P1_REG0_REG_11__SCAN_IN), .A(n10525), .ZN(n10530) );
  OAI22_X1 U11561 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(keyinput55), .B1(
        P2_REG0_REG_10__SCAN_IN), .B2(keyinput99), .ZN(n10526) );
  AOI221_X1 U11562 ( .B1(P1_DATAO_REG_1__SCAN_IN), .B2(keyinput55), .C1(
        keyinput99), .C2(P2_REG0_REG_10__SCAN_IN), .A(n10526), .ZN(n10529) );
  OAI22_X1 U11563 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(keyinput123), .B1(
        P1_REG0_REG_30__SCAN_IN), .B2(keyinput115), .ZN(n10527) );
  AOI221_X1 U11564 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(keyinput123), .C1(
        keyinput115), .C2(P1_REG0_REG_30__SCAN_IN), .A(n10527), .ZN(n10528) );
  NAND4_X1 U11565 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10532) );
  NOR4_X1 U11566 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n10573) );
  OAI22_X1 U11567 ( .A1(P2_D_REG_20__SCAN_IN), .A2(keyinput33), .B1(
        keyinput126), .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n10536) );
  AOI221_X1 U11568 ( .B1(P2_D_REG_20__SCAN_IN), .B2(keyinput33), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput126), .A(n10536), .ZN(n10543)
         );
  OAI22_X1 U11569 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(keyinput34), .B1(
        P1_ADDR_REG_6__SCAN_IN), .B2(keyinput112), .ZN(n10537) );
  AOI221_X1 U11570 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(keyinput34), .C1(
        keyinput112), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n10537), .ZN(n10542) );
  OAI22_X1 U11571 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput30), .B1(
        P1_REG3_REG_19__SCAN_IN), .B2(keyinput29), .ZN(n10538) );
  AOI221_X1 U11572 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput30), .C1(
        keyinput29), .C2(P1_REG3_REG_19__SCAN_IN), .A(n10538), .ZN(n10541) );
  OAI22_X1 U11573 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput120), .B1(
        keyinput119), .B2(P1_REG1_REG_3__SCAN_IN), .ZN(n10539) );
  AOI221_X1 U11574 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput120), .C1(
        P1_REG1_REG_3__SCAN_IN), .C2(keyinput119), .A(n10539), .ZN(n10540) );
  NAND4_X1 U11575 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10571) );
  OAI22_X1 U11576 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput100), .B1(
        P2_REG1_REG_6__SCAN_IN), .B2(keyinput75), .ZN(n10544) );
  AOI221_X1 U11577 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput100), .C1(
        keyinput75), .C2(P2_REG1_REG_6__SCAN_IN), .A(n10544), .ZN(n10551) );
  OAI22_X1 U11578 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(keyinput73), .B1(
        P2_REG0_REG_7__SCAN_IN), .B2(keyinput49), .ZN(n10545) );
  AOI221_X1 U11579 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(keyinput73), .C1(
        keyinput49), .C2(P2_REG0_REG_7__SCAN_IN), .A(n10545), .ZN(n10550) );
  OAI22_X1 U11580 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput18), .B1(
        keyinput53), .B2(P1_REG2_REG_22__SCAN_IN), .ZN(n10546) );
  AOI221_X1 U11581 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput18), .C1(
        P1_REG2_REG_22__SCAN_IN), .C2(keyinput53), .A(n10546), .ZN(n10549) );
  OAI22_X1 U11582 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(keyinput90), .B1(
        P1_REG2_REG_18__SCAN_IN), .B2(keyinput98), .ZN(n10547) );
  AOI221_X1 U11583 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(keyinput90), .C1(
        keyinput98), .C2(P1_REG2_REG_18__SCAN_IN), .A(n10547), .ZN(n10548) );
  NAND4_X1 U11584 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .ZN(
        n10570) );
  OAI22_X1 U11585 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput15), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput21), .ZN(n10552) );
  AOI221_X1 U11586 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput15), .C1(
        keyinput21), .C2(P1_IR_REG_19__SCAN_IN), .A(n10552), .ZN(n10559) );
  OAI22_X1 U11587 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(keyinput83), .B1(
        keyinput35), .B2(P1_D_REG_27__SCAN_IN), .ZN(n10553) );
  AOI221_X1 U11588 ( .B1(P1_DATAO_REG_7__SCAN_IN), .B2(keyinput83), .C1(
        P1_D_REG_27__SCAN_IN), .C2(keyinput35), .A(n10553), .ZN(n10558) );
  OAI22_X1 U11589 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(keyinput5), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput22), .ZN(n10554) );
  AOI221_X1 U11590 ( .B1(P2_REG0_REG_22__SCAN_IN), .B2(keyinput5), .C1(
        keyinput22), .C2(P1_IR_REG_2__SCAN_IN), .A(n10554), .ZN(n10557) );
  OAI22_X1 U11591 ( .A1(P2_D_REG_3__SCAN_IN), .A2(keyinput64), .B1(keyinput8), 
        .B2(P1_REG2_REG_11__SCAN_IN), .ZN(n10555) );
  AOI221_X1 U11592 ( .B1(P2_D_REG_3__SCAN_IN), .B2(keyinput64), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(keyinput8), .A(n10555), .ZN(n10556) );
  NAND4_X1 U11593 ( .A1(n10559), .A2(n10558), .A3(n10557), .A4(n10556), .ZN(
        n10569) );
  OAI22_X1 U11594 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput37), .B1(
        P1_D_REG_28__SCAN_IN), .B2(keyinput41), .ZN(n10560) );
  AOI221_X1 U11595 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput37), .C1(
        keyinput41), .C2(P1_D_REG_28__SCAN_IN), .A(n10560), .ZN(n10567) );
  OAI22_X1 U11596 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(keyinput4), .B1(
        keyinput58), .B2(P1_REG3_REG_0__SCAN_IN), .ZN(n10561) );
  AOI221_X1 U11597 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(keyinput4), .C1(
        P1_REG3_REG_0__SCAN_IN), .C2(keyinput58), .A(n10561), .ZN(n10566) );
  OAI22_X1 U11598 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(keyinput67), .B1(
        P2_ADDR_REG_14__SCAN_IN), .B2(keyinput97), .ZN(n10562) );
  AOI221_X1 U11599 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(keyinput67), .C1(
        keyinput97), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n10562), .ZN(n10565) );
  OAI22_X1 U11600 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput32), .B1(
        P1_REG2_REG_10__SCAN_IN), .B2(keyinput38), .ZN(n10563) );
  AOI221_X1 U11601 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput32), .C1(
        keyinput38), .C2(P1_REG2_REG_10__SCAN_IN), .A(n10563), .ZN(n10564) );
  NAND4_X1 U11602 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(
        n10568) );
  NOR4_X1 U11603 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n10572) );
  NAND2_X1 U11604 ( .A1(n10573), .A2(n10572), .ZN(n10574) );
  NOR4_X1 U11605 ( .A1(n10577), .A2(n10576), .A3(n10575), .A4(n10574), .ZN(
        n10582) );
  AOI22_X1 U11606 ( .A1(n10580), .A2(n10579), .B1(P2_REG0_REG_11__SCAN_IN), 
        .B2(n10578), .ZN(n10581) );
  XNOR2_X1 U11607 ( .A(n10582), .B(n10581), .ZN(P2_U3423) );
  XNOR2_X1 U11608 ( .A(n10584), .B(n10583), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11609 ( .A(n10586), .B(n10585), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11610 ( .A(n10588), .B(n10587), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11611 ( .A(n10590), .B(n10589), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11612 ( .A(n10592), .B(n10591), .ZN(ADD_1068_U48) );
  XOR2_X1 U11613 ( .A(n10594), .B(n10593), .Z(ADD_1068_U54) );
  XOR2_X1 U11614 ( .A(n10596), .B(n10595), .Z(ADD_1068_U53) );
  XNOR2_X1 U11615 ( .A(n10598), .B(n10597), .ZN(ADD_1068_U52) );
  INV_X1 U7512 ( .A(n6284), .ZN(n6265) );
  CLKBUF_X1 U5035 ( .A(n5947), .Z(n5935) );
  CLKBUF_X1 U5101 ( .A(n5918), .Z(n6481) );
  INV_X1 U6495 ( .A(n5949), .ZN(n6522) );
endmodule

