

module b14_C_SARLock_k_64_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2028, n2029, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718;

  AOI211_X1 U2271 ( .C1(n2899), .C2(n4683), .A(n4682), .B(n4681), .ZN(n4710)
         );
  NAND2_X1 U2272 ( .A1(n2860), .A2(n3686), .ZN(n3175) );
  NAND2_X1 U2273 ( .A1(n3157), .A2(n2371), .ZN(n3164) );
  NAND2_X1 U2274 ( .A1(n3155), .A2(n3158), .ZN(n3157) );
  OR2_X2 U2275 ( .A1(n2805), .A2(n3088), .ZN(n3657) );
  CLKBUF_X3 U2276 ( .A(n2273), .Z(n3720) );
  OAI21_X2 U2277 ( .B1(n2363), .B2(n2279), .A(n2278), .ZN(n3124) );
  XNOR2_X1 U2278 ( .A(n2297), .B(n2296), .ZN(n3844) );
  XNOR2_X1 U2279 ( .A(n2260), .B(n2261), .ZN(n3905) );
  CLKBUF_X2 U2280 ( .A(IR_REG_0__SCAN_IN), .Z(n4488) );
  NOR2_X1 U2282 ( .A1(n2193), .A2(n2209), .ZN(n2192) );
  INV_X1 U2283 ( .A(n2675), .ZN(n2773) );
  CLKBUF_X2 U2284 ( .A(n2272), .Z(n2780) );
  NOR2_X2 U2285 ( .A1(n4470), .A2(n2949), .ZN(n2272) );
  AOI21_X2 U2288 ( .B1(n3016), .B2(REG1_REG_6__SCAN_IN), .A(n3015), .ZN(n3855)
         );
  NAND2_X2 U2289 ( .A1(n4318), .A2(n4319), .ZN(n4317) );
  NAND2_X2 U2290 ( .A1(n2869), .A2(n3700), .ZN(n4318) );
  AOI22_X1 U2291 ( .A1(n3120), .A2(n3121), .B1(n2286), .B2(n2691), .ZN(n3065)
         );
  OAI21_X2 U2292 ( .B1(n4123), .B2(n3784), .A(n3788), .ZN(n2882) );
  NAND2_X2 U2293 ( .A1(n2873), .A2(n3783), .ZN(n4123) );
  AOI21_X1 U2294 ( .B1(n3175), .B2(n3669), .A(n3673), .ZN(n3301) );
  OAI21_X2 U2295 ( .B1(n3983), .B2(n3791), .A(n3753), .ZN(n3967) );
  AND3_X2 U2296 ( .A1(n2882), .A2(n3712), .A3(n3793), .ZN(n3983) );
  NAND2_X1 U2297 ( .A1(n2161), .A2(n2164), .ZN(n3539) );
  NAND2_X1 U2298 ( .A1(n3521), .A2(n2618), .ZN(n3529) );
  NAND2_X1 U2299 ( .A1(n2151), .A2(n2152), .ZN(n2570) );
  NAND2_X1 U2300 ( .A1(n3349), .A2(n2466), .ZN(n3371) );
  NAND2_X1 U2301 ( .A1(n2863), .A2(n3678), .ZN(n3333) );
  NOR2_X1 U2302 ( .A1(n3393), .A2(n2180), .ZN(n2179) );
  INV_X1 U2303 ( .A(n2182), .ZN(n2180) );
  NAND2_X1 U2304 ( .A1(n2285), .A2(n2284), .ZN(n3121) );
  OAI21_X1 U2305 ( .B1(n2792), .B2(n4148), .A(n4332), .ZN(n3632) );
  INV_X4 U2306 ( .A(n2691), .ZN(n2735) );
  AND2_X2 U2307 ( .A1(n2853), .A2(n2771), .ZN(n2691) );
  NAND2_X1 U2308 ( .A1(n3661), .A2(n3664), .ZN(n3103) );
  AND2_X1 U2309 ( .A1(n3666), .A2(n3663), .ZN(n3771) );
  INV_X2 U2310 ( .A(n3825), .ZN(U4043) );
  NAND2_X1 U2311 ( .A1(n2254), .A2(n2253), .ZN(n2319) );
  NAND3_X1 U2312 ( .A1(n2740), .A2(n4471), .A3(n2936), .ZN(n2256) );
  NAND2_X1 U2313 ( .A1(n2949), .A2(n4470), .ZN(n2309) );
  OR2_X1 U2314 ( .A1(n2217), .A2(n2775), .ZN(n2215) );
  AND2_X1 U2315 ( .A1(n2244), .A2(n2104), .ZN(n2217) );
  INV_X1 U2316 ( .A(n2315), .ZN(n2210) );
  INV_X1 U2317 ( .A(IR_REG_2__SCAN_IN), .ZN(n2296) );
  INV_X1 U2318 ( .A(IR_REG_8__SCAN_IN), .ZN(n2206) );
  INV_X1 U2319 ( .A(IR_REG_7__SCAN_IN), .ZN(n2204) );
  NOR2_X1 U2320 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2063)
         );
  NOR2_X1 U2321 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2208)
         );
  NOR2_X1 U2322 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2062)
         );
  INV_X1 U2323 ( .A(IR_REG_14__SCAN_IN), .ZN(n2525) );
  INV_X1 U2324 ( .A(IR_REG_13__SCAN_IN), .ZN(n4235) );
  INV_X1 U2325 ( .A(IR_REG_6__SCAN_IN), .ZN(n2227) );
  NAND2_X1 U2326 ( .A1(n2131), .A2(n2212), .ZN(n2250) );
  OR3_X1 U2327 ( .A1(n4123), .A2(n4078), .A3(n4000), .ZN(n4058) );
  AND2_X2 U2328 ( .A1(n2190), .A2(n2210), .ZN(n2359) );
  AOI21_X2 U2329 ( .B1(n3539), .B2(n3541), .A(n3540), .ZN(n3623) );
  NAND2_X1 U2331 ( .A1(n2259), .A2(n2256), .ZN(n2732) );
  OR2_X4 U2332 ( .A1(n2259), .A2(n2283), .ZN(n2325) );
  AND2_X1 U2333 ( .A1(n2269), .A2(n2268), .ZN(n2028) );
  AND2_X1 U2334 ( .A1(n2269), .A2(n2268), .ZN(n2029) );
  AND2_X4 U2335 ( .A1(n2269), .A2(n2268), .ZN(n2324) );
  CLKBUF_X1 U2336 ( .A(n2732), .Z(n2031) );
  OAI21_X2 U2337 ( .B1(n2855), .B2(n3657), .A(n2856), .ZN(n3106) );
  NAND2_X2 U2338 ( .A1(n2502), .A2(n3392), .ZN(n3459) );
  NOR2_X2 U2339 ( .A1(n2523), .A2(n2230), .ZN(n2584) );
  NAND2_X2 U2340 ( .A1(n2234), .A2(IR_REG_31__SCAN_IN), .ZN(n2260) );
  NAND2_X2 U2341 ( .A1(n2266), .A2(n2267), .ZN(n2259) );
  INV_X2 U2342 ( .A(n2899), .ZN(n2269) );
  AOI21_X2 U2343 ( .B1(n3565), .B2(n2051), .A(n2167), .ZN(n3519) );
  AOI21_X2 U2344 ( .B1(n2576), .B2(n2575), .A(n2574), .ZN(n3565) );
  AOI21_X1 U2345 ( .B1(n2265), .B2(n2028), .A(n2270), .ZN(n2287) );
  BUF_X2 U2346 ( .A(n2267), .Z(n2760) );
  INV_X4 U2347 ( .A(n2325), .ZN(n2657) );
  XNOR2_X2 U2348 ( .A(n2237), .B(n2236), .ZN(n2266) );
  AND2_X1 U2349 ( .A1(n2210), .A2(n2188), .ZN(n2187) );
  INV_X1 U2350 ( .A(IR_REG_22__SCAN_IN), .ZN(n2188) );
  NOR2_X1 U2351 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2211)
         );
  XNOR2_X1 U2352 ( .A(n2988), .B(n4497), .ZN(n4493) );
  AND2_X1 U2353 ( .A1(n2170), .A2(n2177), .ZN(n2169) );
  INV_X1 U2354 ( .A(n3613), .ZN(n2177) );
  NAND2_X1 U2355 ( .A1(n2175), .A2(n2171), .ZN(n2170) );
  OR2_X1 U2356 ( .A1(n4555), .A2(n3864), .ZN(n3865) );
  INV_X1 U2357 ( .A(IR_REG_25__SCAN_IN), .ZN(n2212) );
  INV_X1 U2358 ( .A(IR_REG_10__SCAN_IN), .ZN(n2207) );
  AND2_X1 U2359 ( .A1(n3508), .A2(n3509), .ZN(n2666) );
  NAND2_X1 U2360 ( .A1(n2962), .A2(n2777), .ZN(n2251) );
  OR2_X1 U2361 ( .A1(n3032), .A2(n2992), .ZN(n3014) );
  NAND2_X1 U2362 ( .A1(n2143), .A2(n3891), .ZN(n2141) );
  INV_X1 U2363 ( .A(n3865), .ZN(n2143) );
  NOR2_X1 U2364 ( .A1(n4582), .A2(n3868), .ZN(n3870) );
  NAND2_X1 U2365 ( .A1(n4603), .A2(n3873), .ZN(n4617) );
  AND2_X1 U2366 ( .A1(n2684), .A2(REG3_REG_25__SCAN_IN), .ZN(n2712) );
  AOI21_X1 U2367 ( .B1(n2084), .B2(n2083), .A(n2082), .ZN(n4101) );
  NOR2_X1 U2368 ( .A1(n2087), .A2(n2035), .ZN(n2083) );
  OAI21_X1 U2369 ( .B1(n2085), .B2(n2035), .A(n2057), .ZN(n2082) );
  NOR2_X1 U2370 ( .A1(n2194), .A2(n2105), .ZN(n2104) );
  INV_X1 U2371 ( .A(n2211), .ZN(n2105) );
  NAND2_X1 U2372 ( .A1(n2195), .A2(n2777), .ZN(n2194) );
  INV_X1 U2373 ( .A(IR_REG_28__SCAN_IN), .ZN(n2777) );
  OAI21_X2 U2374 ( .B1(n2250), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2962) );
  INV_X1 U2375 ( .A(IR_REG_20__SCAN_IN), .ZN(n2236) );
  NAND2_X1 U2376 ( .A1(n2730), .A2(n2729), .ZN(n3942) );
  NAND2_X1 U2377 ( .A1(n4604), .A2(n4605), .ZN(n4603) );
  XNOR2_X1 U2378 ( .A(n3925), .B(n3924), .ZN(n3490) );
  INV_X1 U2379 ( .A(n3498), .ZN(n2155) );
  XNOR2_X1 U2380 ( .A(n2343), .B(n2691), .ZN(n2348) );
  NOR2_X1 U2381 ( .A1(n4535), .A2(n2059), .ZN(n3862) );
  AND2_X1 U2382 ( .A1(n2122), .A2(n2121), .ZN(n3897) );
  NAND2_X1 U2383 ( .A1(n3896), .A2(REG2_REG_15__SCAN_IN), .ZN(n2121) );
  INV_X1 U2384 ( .A(n3736), .ZN(n2066) );
  AOI21_X1 U2385 ( .B1(n2070), .B2(n2841), .A(n2081), .ZN(n2069) );
  INV_X1 U2386 ( .A(n2072), .ZN(n2070) );
  INV_X1 U2387 ( .A(n2074), .ZN(n2071) );
  AND2_X1 U2388 ( .A1(n3616), .A2(n4093), .ZN(n2839) );
  AOI21_X1 U2389 ( .B1(n3767), .B2(n2827), .A(n2045), .ZN(n2103) );
  INV_X1 U2390 ( .A(n2827), .ZN(n2101) );
  OR2_X1 U2391 ( .A1(n3222), .A2(n3253), .ZN(n3667) );
  NAND2_X1 U2392 ( .A1(n3222), .A2(n3253), .ZN(n3672) );
  AND2_X1 U2393 ( .A1(n2760), .A2(n2932), .ZN(n2958) );
  NAND2_X1 U2394 ( .A1(n4113), .A2(n4069), .ZN(n2130) );
  AOI21_X1 U2395 ( .B1(n2831), .B2(n2830), .A(n2829), .ZN(n4312) );
  AND2_X1 U2396 ( .A1(n3500), .A2(n3464), .ZN(n2829) );
  NAND2_X1 U2397 ( .A1(n4328), .A2(n3421), .ZN(n2830) );
  INV_X1 U2398 ( .A(n3410), .ZN(n2831) );
  OR2_X1 U2399 ( .A1(n2244), .A2(n2775), .ZN(n2758) );
  INV_X1 U2400 ( .A(IR_REG_23__SCAN_IN), .ZN(n2757) );
  INV_X1 U2401 ( .A(IR_REG_5__SCAN_IN), .ZN(n2191) );
  INV_X1 U2402 ( .A(IR_REG_15__SCAN_IN), .ZN(n2546) );
  OR2_X1 U2403 ( .A1(n2474), .A2(n2775), .ZN(n2490) );
  NAND2_X1 U2404 ( .A1(n2210), .A2(n2197), .ZN(n2357) );
  CLKBUF_X1 U2405 ( .A(n2359), .Z(n2360) );
  NAND2_X1 U2406 ( .A1(n2160), .A2(n2515), .ZN(n2154) );
  XNOR2_X1 U2407 ( .A(n2322), .B(n2735), .ZN(n2327) );
  NAND2_X1 U2408 ( .A1(n2321), .A2(n2320), .ZN(n2322) );
  INV_X1 U2409 ( .A(n2168), .ZN(n2167) );
  AOI22_X1 U2410 ( .A1(n2169), .A2(n2172), .B1(n2173), .B2(n3567), .ZN(n2168)
         );
  INV_X1 U2411 ( .A(n2666), .ZN(n2162) );
  NOR2_X1 U2412 ( .A1(n2683), .A2(n2678), .ZN(n2166) );
  NOR2_X1 U2413 ( .A1(n2678), .A2(n2679), .ZN(n2681) );
  NAND2_X1 U2414 ( .A1(n3372), .A2(n3373), .ZN(n2182) );
  NAND2_X1 U2415 ( .A1(n3371), .A2(n2183), .ZN(n2181) );
  NAND2_X1 U2416 ( .A1(n2185), .A2(n2184), .ZN(n2183) );
  INV_X1 U2417 ( .A(n3372), .ZN(n2185) );
  INV_X1 U2418 ( .A(n3373), .ZN(n2184) );
  OR2_X1 U2419 ( .A1(n3937), .A2(n2786), .ZN(n2718) );
  NAND2_X1 U2420 ( .A1(n2273), .A2(REG1_REG_0__SCAN_IN), .ZN(n2275) );
  AND2_X1 U2421 ( .A1(n2113), .A2(n2112), .ZN(n3020) );
  NAND2_X1 U2422 ( .A1(n3031), .A2(REG2_REG_5__SCAN_IN), .ZN(n2112) );
  XNOR2_X1 U2423 ( .A(n3862), .B(n4655), .ZN(n4546) );
  OR2_X1 U2424 ( .A1(n4546), .A2(n4547), .ZN(n2144) );
  NOR2_X1 U2425 ( .A1(n3892), .A2(n3891), .ZN(n3895) );
  AND3_X1 U2426 ( .A1(n2141), .A2(n3866), .A3(REG1_REG_14__SCAN_IN), .ZN(n4568) );
  XNOR2_X1 U2427 ( .A(n3870), .B(n3869), .ZN(n4593) );
  INV_X1 U2428 ( .A(n2120), .ZN(n2118) );
  NOR2_X1 U2429 ( .A1(n3929), .A2(n3930), .ZN(n4345) );
  OR2_X1 U2430 ( .A1(n2723), .A2(n4208), .ZN(n3910) );
  OR2_X1 U2431 ( .A1(n3800), .A2(n3718), .ZN(n3940) );
  OR2_X1 U2432 ( .A1(n2848), .A2(n2199), .ZN(n2095) );
  NOR2_X1 U2433 ( .A1(n2099), .A2(n2042), .ZN(n2098) );
  INV_X1 U2434 ( .A(n2845), .ZN(n2099) );
  INV_X1 U2435 ( .A(n3546), .ZN(n4008) );
  NOR2_X1 U2436 ( .A1(n2839), .A2(n2080), .ZN(n2079) );
  INV_X1 U2437 ( .A(n2838), .ZN(n2080) );
  AOI21_X1 U2438 ( .B1(n2088), .B2(n2086), .A(n2053), .ZN(n2085) );
  INV_X1 U2439 ( .A(n2834), .ZN(n2086) );
  INV_X1 U2440 ( .A(n2088), .ZN(n2087) );
  AND2_X1 U2441 ( .A1(n4142), .A2(n2054), .ZN(n2088) );
  NAND2_X1 U2442 ( .A1(n4310), .A2(n2833), .ZN(n3428) );
  NAND2_X1 U2443 ( .A1(n4308), .A2(n2832), .ZN(n2833) );
  OAI21_X1 U2444 ( .B1(n3337), .B2(n2826), .A(n2825), .ZN(n3443) );
  OR2_X1 U2445 ( .A1(n2200), .A2(n2823), .ZN(n3278) );
  AND2_X1 U2446 ( .A1(n3675), .A2(n3685), .ZN(n3762) );
  AND2_X1 U2447 ( .A1(n2887), .A2(n2886), .ZN(n4129) );
  AND2_X1 U2448 ( .A1(n4012), .A2(n2038), .ZN(n3935) );
  NAND2_X1 U2449 ( .A1(n3935), .A2(n2898), .ZN(n3929) );
  NOR2_X1 U2450 ( .A1(n2033), .A2(n4033), .ZN(n4380) );
  INV_X1 U2451 ( .A(IR_REG_29__SCAN_IN), .ZN(n2216) );
  NAND2_X1 U2452 ( .A1(n2046), .A2(n2212), .ZN(n2196) );
  INV_X1 U2453 ( .A(IR_REG_26__SCAN_IN), .ZN(n2214) );
  INV_X1 U2454 ( .A(n2246), .ZN(n2131) );
  NAND2_X1 U2455 ( .A1(n2758), .A2(n2757), .ZN(n2756) );
  OAI21_X1 U2456 ( .B1(n2758), .B2(n2757), .A(n2756), .ZN(n2960) );
  AND2_X1 U2457 ( .A1(n2063), .A2(n2062), .ZN(n2189) );
  INV_X1 U2458 ( .A(IR_REG_19__SCAN_IN), .ZN(n2261) );
  INV_X1 U2459 ( .A(IR_REG_18__SCAN_IN), .ZN(n2232) );
  INV_X1 U2460 ( .A(IR_REG_16__SCAN_IN), .ZN(n2561) );
  OR2_X1 U2461 ( .A1(n2788), .A2(n2787), .ZN(n3630) );
  INV_X1 U2462 ( .A(n2932), .ZN(n3816) );
  NAND2_X1 U2463 ( .A1(n2702), .A2(n2701), .ZN(n3970) );
  OR2_X1 U2464 ( .A1(n2656), .A2(n2655), .ZN(n4034) );
  OAI22_X1 U2465 ( .A1(n4493), .A2(n2147), .B1(n2989), .B2(n2146), .ZN(n3032)
         );
  INV_X1 U2466 ( .A(n2991), .ZN(n2146) );
  NAND2_X1 U2467 ( .A1(n2991), .A2(REG1_REG_4__SCAN_IN), .ZN(n2147) );
  XNOR2_X1 U2468 ( .A(n3014), .B(n2999), .ZN(n3016) );
  NAND2_X1 U2469 ( .A1(n4551), .A2(n3889), .ZN(n4562) );
  NOR2_X1 U2470 ( .A1(n4583), .A2(n4569), .ZN(n2140) );
  NAND2_X1 U2471 ( .A1(n4619), .A2(n4607), .ZN(n4623) );
  NOR2_X1 U2472 ( .A1(n4617), .A2(n4616), .ZN(n4624) );
  NAND2_X1 U2473 ( .A1(n4600), .A2(n2120), .ZN(n4614) );
  NOR2_X1 U2474 ( .A1(n3922), .A2(n2898), .ZN(n3923) );
  INV_X1 U2475 ( .A(n3942), .ZN(n3922) );
  NAND2_X1 U2476 ( .A1(n4076), .A2(n3183), .ZN(n3928) );
  OAI21_X1 U2477 ( .B1(n3490), .B2(n4685), .A(n2892), .ZN(n2904) );
  OR2_X1 U2478 ( .A1(n3359), .A2(n2866), .ZN(n2869) );
  INV_X1 U2479 ( .A(n2324), .ZN(n2719) );
  INV_X1 U2480 ( .A(n2175), .ZN(n2172) );
  NOR2_X1 U2481 ( .A1(n3612), .A2(n2171), .ZN(n2173) );
  OR2_X1 U2482 ( .A1(n2962), .A2(n2213), .ZN(n2252) );
  AOI21_X1 U2483 ( .B1(n2153), .B2(n2159), .A(n2058), .ZN(n2152) );
  NOR2_X1 U2484 ( .A1(n2199), .A2(n2097), .ZN(n2096) );
  INV_X1 U2485 ( .A(n2098), .ZN(n2097) );
  NOR2_X1 U2486 ( .A1(n2670), .A2(n3580), .ZN(n2684) );
  NAND2_X1 U2487 ( .A1(n3667), .A2(n3672), .ZN(n3242) );
  NOR2_X1 U2488 ( .A1(n3545), .A2(n3582), .ZN(n2132) );
  NOR2_X1 U2489 ( .A1(n3464), .A2(n2135), .ZN(n2134) );
  NOR2_X1 U2490 ( .A1(n2034), .A2(n3267), .ZN(n2125) );
  INV_X1 U2491 ( .A(n3226), .ZN(n2124) );
  INV_X1 U2492 ( .A(n2196), .ZN(n2195) );
  INV_X1 U2493 ( .A(IR_REG_17__SCAN_IN), .ZN(n2231) );
  NAND2_X1 U2494 ( .A1(n2229), .A2(n4235), .ZN(n2523) );
  INV_X1 U2495 ( .A(n2509), .ZN(n2229) );
  NAND2_X1 U2497 ( .A1(n2516), .A2(REG3_REG_14__SCAN_IN), .ZN(n2538) );
  AND2_X1 U2498 ( .A1(n2533), .A2(n2534), .ZN(n3498) );
  NAND2_X1 U2499 ( .A1(n3322), .A2(n3323), .ZN(n2178) );
  INV_X1 U2500 ( .A(n3974), .ZN(n3545) );
  INV_X1 U2501 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2553) );
  OR2_X1 U2502 ( .A1(n2538), .A2(n3644), .ZN(n2554) );
  OAI21_X1 U2503 ( .B1(n2568), .B2(n2567), .A(n2573), .ZN(n3557) );
  NAND2_X1 U2504 ( .A1(n2331), .A2(n2330), .ZN(n3194) );
  NAND2_X1 U2505 ( .A1(n3231), .A2(n3232), .ZN(n2186) );
  OR2_X1 U2506 ( .A1(n2636), .A2(n2635), .ZN(n3593) );
  AND2_X1 U2507 ( .A1(n2636), .A2(n2635), .ZN(n3591) );
  INV_X1 U2508 ( .A(n3421), .ZN(n3464) );
  NAND2_X1 U2509 ( .A1(n2477), .A2(n2476), .ZN(n3373) );
  XNOR2_X1 U2510 ( .A(n2480), .B(n2735), .ZN(n3372) );
  XNOR2_X1 U2511 ( .A(n2602), .B(n2735), .ZN(n3613) );
  XNOR2_X1 U2512 ( .A(n2387), .B(n2735), .ZN(n3165) );
  NAND2_X1 U2513 ( .A1(n2384), .A2(n2383), .ZN(n3166) );
  NOR2_X1 U2514 ( .A1(n2695), .A2(n2694), .ZN(n3540) );
  INV_X1 U2515 ( .A(n3648), .ZN(n3627) );
  OR2_X1 U2516 ( .A1(n2788), .A2(n2791), .ZN(n2792) );
  OR2_X1 U2517 ( .A1(n2786), .A2(REG3_REG_3__SCAN_IN), .ZN(n2312) );
  NAND2_X1 U2518 ( .A1(n3006), .A2(n2969), .ZN(n3846) );
  NAND2_X1 U2519 ( .A1(n2136), .A2(n2967), .ZN(n2983) );
  XNOR2_X1 U2520 ( .A(n2994), .B(n2981), .ZN(n2993) );
  NAND3_X1 U2521 ( .A1(n2108), .A2(n2107), .A3(n2109), .ZN(n2113) );
  INV_X1 U2522 ( .A(n3035), .ZN(n2109) );
  NAND2_X1 U2523 ( .A1(n2039), .A2(n2111), .ZN(n2107) );
  INV_X1 U2524 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U2525 ( .A1(n2150), .A2(REG1_REG_8__SCAN_IN), .ZN(n2149) );
  OAI21_X1 U2526 ( .B1(n2428), .B2(n4660), .A(n4520), .ZN(n3884) );
  AND2_X1 U2527 ( .A1(n2047), .A2(n2144), .ZN(n4557) );
  NAND2_X1 U2528 ( .A1(n4540), .A2(n3886), .ZN(n3888) );
  OR2_X1 U2529 ( .A1(n4579), .A2(n4578), .ZN(n2122) );
  XNOR2_X1 U2530 ( .A(n3897), .B(n3869), .ZN(n4590) );
  NAND2_X1 U2531 ( .A1(n4590), .A2(n2552), .ZN(n4589) );
  AND2_X1 U2532 ( .A1(n2959), .A2(n2363), .ZN(n2976) );
  NAND2_X1 U2533 ( .A1(n4647), .A2(n2579), .ZN(n2120) );
  NAND2_X1 U2534 ( .A1(n4620), .A2(REG2_REG_18__SCAN_IN), .ZN(n2119) );
  NAND2_X1 U2535 ( .A1(n2064), .A2(n2850), .ZN(n3925) );
  NOR2_X1 U2536 ( .A1(n2851), .A2(n2066), .ZN(n2065) );
  OAI21_X1 U2537 ( .B1(n3949), .B2(n3656), .A(n2884), .ZN(n3939) );
  INV_X1 U2538 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3512) );
  NAND2_X1 U2539 ( .A1(n2643), .A2(n2642), .ZN(n2651) );
  AND2_X1 U2540 ( .A1(n3725), .A2(DATAI_22_), .ZN(n4033) );
  AOI21_X1 U2541 ( .B1(n2068), .B2(n2041), .A(n2067), .ZN(n4023) );
  INV_X1 U2542 ( .A(n2069), .ZN(n2067) );
  NAND2_X1 U2543 ( .A1(n2073), .A2(n2032), .ZN(n2072) );
  INV_X1 U2544 ( .A(n2076), .ZN(n2073) );
  AOI21_X1 U2545 ( .B1(n2078), .B2(n2077), .A(n2040), .ZN(n2076) );
  INV_X1 U2546 ( .A(n2079), .ZN(n2077) );
  NAND2_X1 U2547 ( .A1(n2032), .A2(n2078), .ZN(n2074) );
  OR2_X1 U2548 ( .A1(n3749), .A2(n3748), .ZN(n4040) );
  INV_X1 U2549 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4211) );
  INV_X1 U2550 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2603) );
  INV_X1 U2551 ( .A(n4125), .ZN(n2837) );
  AND2_X1 U2552 ( .A1(n3755), .A2(n3754), .ZN(n4084) );
  OR2_X1 U2553 ( .A1(n2593), .A2(n4276), .ZN(n2604) );
  AOI21_X1 U2554 ( .B1(n2103), .B2(n2101), .A(n2055), .ZN(n2100) );
  INV_X1 U2555 ( .A(n2103), .ZN(n2102) );
  NOR2_X1 U2556 ( .A1(n2482), .A2(n2481), .ZN(n2503) );
  OR2_X1 U2557 ( .A1(n3443), .A2(n3767), .ZN(n3441) );
  OR2_X1 U2558 ( .A1(n2467), .A2(n3376), .ZN(n2482) );
  AND2_X1 U2559 ( .A1(n3358), .A2(n3698), .ZN(n3767) );
  NOR2_X1 U2560 ( .A1(n2429), .A2(n3325), .ZN(n2449) );
  OR2_X1 U2561 ( .A1(n3271), .A2(n3683), .ZN(n2863) );
  NAND2_X1 U2562 ( .A1(n2091), .A2(n2090), .ZN(n3337) );
  AOI21_X1 U2563 ( .B1(n2092), .B2(n2824), .A(n2056), .ZN(n2091) );
  INV_X1 U2564 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2407) );
  OR2_X1 U2565 ( .A1(n2408), .A2(n2407), .ZN(n2429) );
  INV_X1 U2566 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4251) );
  OR2_X1 U2567 ( .A1(n2390), .A2(n4251), .ZN(n2408) );
  INV_X1 U2568 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2350) );
  OR2_X1 U2569 ( .A1(n3246), .A2(n2858), .ZN(n2859) );
  NAND2_X1 U2570 ( .A1(n3241), .A2(n3242), .ZN(n3245) );
  INV_X1 U2571 ( .A(n3242), .ZN(n3772) );
  INV_X1 U2572 ( .A(n4086), .ZN(n4323) );
  INV_X1 U2573 ( .A(n4350), .ZN(n4148) );
  NOR2_X1 U2574 ( .A1(n3138), .A2(n3147), .ZN(n3254) );
  AND2_X1 U2575 ( .A1(n2908), .A2(n2807), .ZN(n3104) );
  INV_X1 U2576 ( .A(n4129), .ZN(n4320) );
  AND2_X1 U2577 ( .A1(n3086), .A2(n4472), .ZN(n4350) );
  NAND2_X1 U2578 ( .A1(n4012), .A2(n2037), .ZN(n3956) );
  NAND2_X1 U2579 ( .A1(n4012), .A2(n2132), .ZN(n3973) );
  NAND2_X1 U2580 ( .A1(n4012), .A2(n3992), .ZN(n3991) );
  INV_X1 U2581 ( .A(n3515), .ZN(n4014) );
  AND2_X1 U2582 ( .A1(n4380), .A2(n4014), .ZN(n4012) );
  NAND2_X1 U2583 ( .A1(n2129), .A2(n2128), .ZN(n2127) );
  INV_X1 U2584 ( .A(n2130), .ZN(n2129) );
  NOR2_X1 U2585 ( .A1(n3526), .A2(n4045), .ZN(n2128) );
  NAND2_X1 U2586 ( .A1(n3725), .A2(DATAI_20_), .ZN(n4069) );
  NOR3_X1 U2587 ( .A1(n4131), .A2(n3526), .A3(n3620), .ZN(n4091) );
  NOR2_X1 U2588 ( .A1(n4131), .A2(n3620), .ZN(n4103) );
  OR2_X1 U2589 ( .A1(n4404), .A2(n4124), .ZN(n4131) );
  AND2_X1 U2590 ( .A1(n3449), .A2(n2133), .ZN(n4154) );
  AND2_X1 U2591 ( .A1(n2036), .A2(n3434), .ZN(n2133) );
  NAND2_X1 U2592 ( .A1(n3449), .A2(n2036), .ZN(n4307) );
  NAND2_X1 U2593 ( .A1(n3449), .A2(n2134), .ZN(n4306) );
  AND2_X1 U2594 ( .A1(n3452), .A2(n3451), .ZN(n3449) );
  NAND2_X1 U2595 ( .A1(n3449), .A2(n3366), .ZN(n3420) );
  NAND2_X1 U2596 ( .A1(n2124), .A2(n2123), .ZN(n3338) );
  AND2_X1 U2597 ( .A1(n2125), .A2(n3275), .ZN(n2123) );
  NOR2_X1 U2598 ( .A1(n3338), .A2(n3354), .ZN(n3452) );
  NAND2_X1 U2599 ( .A1(n2124), .A2(n2125), .ZN(n3293) );
  NOR2_X1 U2600 ( .A1(n3226), .A2(n2034), .ZN(n3307) );
  OR2_X1 U2601 ( .A1(n3252), .A2(n3224), .ZN(n3226) );
  NOR2_X1 U2602 ( .A1(n3226), .A2(n3184), .ZN(n3306) );
  INV_X1 U2603 ( .A(n4692), .ZN(n4685) );
  OR2_X1 U2604 ( .A1(n3113), .A2(n3114), .ZN(n3138) );
  NOR2_X1 U2605 ( .A1(n2896), .A2(n2916), .ZN(n2903) );
  CLKBUF_X1 U2606 ( .A(n2761), .Z(n3086) );
  AND2_X1 U2607 ( .A1(n2256), .A2(n2759), .ZN(n2961) );
  NAND2_X1 U2608 ( .A1(n2741), .A2(n2740), .ZN(n2952) );
  AND2_X1 U2609 ( .A1(n2548), .A2(n2560), .ZN(n3896) );
  CLKBUF_X1 U2610 ( .A(n2523), .Z(n2524) );
  XNOR2_X1 U2611 ( .A(n2490), .B(IR_REG_11__SCAN_IN), .ZN(n3877) );
  AND2_X1 U2612 ( .A1(n2362), .A2(n2361), .ZN(n3031) );
  NOR2_X2 U2613 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2295)
         );
  XNOR2_X1 U2614 ( .A(n2403), .B(n2404), .ZN(n3232) );
  NAND2_X1 U2615 ( .A1(n2158), .A2(n2157), .ZN(n2156) );
  INV_X1 U2616 ( .A(n3459), .ZN(n2158) );
  AND2_X1 U2617 ( .A1(n3725), .A2(DATAI_23_), .ZN(n3515) );
  CLKBUF_X1 U2618 ( .A(n3519), .Z(n3520) );
  AND2_X1 U2619 ( .A1(n3725), .A2(DATAI_21_), .ZN(n4045) );
  AOI22_X1 U2620 ( .A1(n2683), .A2(n2165), .B1(n2678), .B2(n2679), .ZN(n2164)
         );
  INV_X1 U2621 ( .A(n2681), .ZN(n2165) );
  CLKBUF_X1 U2622 ( .A(n3155), .Z(n3156) );
  NAND2_X1 U2623 ( .A1(n2163), .A2(n2678), .ZN(n3576) );
  NAND2_X1 U2624 ( .A1(n3506), .A2(n2680), .ZN(n2163) );
  XNOR2_X1 U2625 ( .A(n2445), .B(n2446), .ZN(n3323) );
  INV_X1 U2626 ( .A(n4488), .ZN(n2279) );
  NAND2_X1 U2627 ( .A1(n2363), .A2(DATAI_0_), .ZN(n2278) );
  INV_X1 U2628 ( .A(n3560), .ZN(n3643) );
  INV_X1 U2629 ( .A(n3630), .ZN(n3645) );
  CLKBUF_X1 U2630 ( .A(n3601), .Z(n3602) );
  OAI21_X1 U2631 ( .B1(n2363), .B2(n2300), .A(n2299), .ZN(n3101) );
  NAND2_X1 U2632 ( .A1(n2363), .A2(n2298), .ZN(n2299) );
  INV_X1 U2633 ( .A(n3632), .ZN(n3560) );
  CLKBUF_X1 U2634 ( .A(n3095), .Z(n3096) );
  INV_X1 U2635 ( .A(n3653), .ZN(n3608) );
  OR2_X1 U2636 ( .A1(n3565), .A2(n3567), .ZN(n2174) );
  OR2_X1 U2637 ( .A1(n2774), .A2(n3069), .ZN(n3650) );
  INV_X1 U2638 ( .A(n3631), .ZN(n3952) );
  NAND4_X1 U2639 ( .A1(n2649), .A2(n2648), .A3(n2647), .A4(n2646), .ZN(n4046)
         );
  OR2_X1 U2640 ( .A1(n2256), .A2(n4644), .ZN(n3825) );
  NAND4_X1 U2641 ( .A1(n2336), .A2(n2335), .A3(n2334), .A4(n2333), .ZN(n3222)
         );
  OR2_X1 U2642 ( .A1(n2786), .A2(n3255), .ZN(n2333) );
  OR2_X1 U2643 ( .A1(n3724), .A2(n2111), .ZN(n2334) );
  OR2_X1 U2644 ( .A1(n2332), .A2(n2968), .ZN(n2291) );
  OR2_X1 U2645 ( .A1(n2309), .A2(n2290), .ZN(n2292) );
  CLKBUF_X1 U2646 ( .A(n2265), .Z(n3123) );
  NAND2_X1 U2647 ( .A1(n2272), .A2(REG0_REG_0__SCAN_IN), .ZN(n2276) );
  OR2_X1 U2648 ( .A1(n2309), .A2(n2271), .ZN(n2277) );
  INV_X1 U2649 ( .A(n3844), .ZN(n2300) );
  XNOR2_X1 U2650 ( .A(n2983), .B(n2981), .ZN(n2982) );
  OR2_X1 U2651 ( .A1(n4493), .A2(n2987), .ZN(n2145) );
  INV_X1 U2652 ( .A(n2110), .ZN(n3036) );
  NAND2_X1 U2653 ( .A1(n3026), .A2(n3025), .ZN(n3879) );
  INV_X1 U2654 ( .A(n3024), .ZN(n3025) );
  AND2_X1 U2655 ( .A1(n2149), .A2(n2148), .ZN(n4517) );
  XNOR2_X1 U2656 ( .A(n3884), .B(n4658), .ZN(n4532) );
  XNOR2_X1 U2657 ( .A(n3888), .B(n4655), .ZN(n4552) );
  NAND2_X1 U2658 ( .A1(n4552), .A2(REG2_REG_12__SCAN_IN), .ZN(n4551) );
  INV_X1 U2659 ( .A(n2144), .ZN(n4545) );
  NAND2_X1 U2660 ( .A1(n3894), .A2(n3893), .ZN(n4567) );
  NAND2_X1 U2661 ( .A1(n3892), .A2(n3891), .ZN(n3893) );
  NAND2_X1 U2662 ( .A1(n2141), .A2(n3866), .ZN(n4570) );
  INV_X1 U2663 ( .A(n4568), .ZN(n2138) );
  NAND2_X1 U2664 ( .A1(n4591), .A2(n3871), .ZN(n4604) );
  NAND2_X1 U2665 ( .A1(n2115), .A2(n2114), .ZN(n3902) );
  NAND2_X1 U2666 ( .A1(n2117), .A2(n2119), .ZN(n2114) );
  AND2_X1 U2667 ( .A1(n3910), .A2(n2724), .ZN(n3491) );
  NAND2_X1 U2668 ( .A1(n2849), .A2(n3736), .ZN(n3934) );
  NAND2_X1 U2669 ( .A1(n2846), .A2(n2098), .ZN(n3965) );
  NAND2_X1 U2670 ( .A1(n2846), .A2(n2845), .ZN(n3981) );
  NAND2_X1 U2671 ( .A1(n4099), .A2(n2079), .ZN(n2075) );
  OAI21_X1 U2672 ( .B1(n3428), .B2(n2087), .A(n2085), .ZN(n4121) );
  NAND2_X1 U2673 ( .A1(n4154), .A2(n4153), .ZN(n4404) );
  NAND2_X1 U2674 ( .A1(n2089), .A2(n2088), .ZN(n4140) );
  AND2_X1 U2675 ( .A1(n2089), .A2(n2054), .ZN(n4141) );
  NAND2_X1 U2676 ( .A1(n3428), .A2(n2834), .ZN(n2089) );
  INV_X1 U2677 ( .A(n3290), .ZN(n2093) );
  INV_X1 U2678 ( .A(n3905), .ZN(n4314) );
  AND2_X1 U2679 ( .A1(n4118), .A2(n2899), .ZN(n4633) );
  OR2_X1 U2680 ( .A1(n2893), .A2(n2791), .ZN(n4332) );
  INV_X1 U2681 ( .A(n3124), .ZN(n3088) );
  AND2_X1 U2682 ( .A1(n3657), .A2(n3658), .ZN(n3738) );
  CLKBUF_X1 U2683 ( .A(n2922), .Z(n4485) );
  INV_X1 U2684 ( .A(n4332), .ZN(n4631) );
  NAND2_X1 U2685 ( .A1(n4333), .A2(n2923), .ZN(n4076) );
  AND2_X2 U2686 ( .A1(n2903), .A2(n2902), .ZN(n4718) );
  INV_X1 U2687 ( .A(n4718), .ZN(n4715) );
  AOI21_X1 U2688 ( .B1(n2899), .B2(n4356), .A(n4355), .ZN(n4357) );
  NAND2_X1 U2689 ( .A1(n4706), .A2(n2899), .ZN(n4468) );
  AND2_X2 U2690 ( .A1(n2903), .A2(n2919), .ZN(n4706) );
  NAND2_X1 U2691 ( .A1(n2952), .A2(n2961), .ZN(n4641) );
  NAND2_X1 U2692 ( .A1(n2939), .A2(IR_REG_31__SCAN_IN), .ZN(n2218) );
  XNOR2_X1 U2693 ( .A(n2778), .B(n2777), .ZN(n4478) );
  CLKBUF_X1 U2694 ( .A(n2962), .Z(n2963) );
  XNOR2_X1 U2695 ( .A(n2248), .B(IR_REG_25__SCAN_IN), .ZN(n2936) );
  XNOR2_X1 U2697 ( .A(n2245), .B(IR_REG_24__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U2698 ( .A1(n2960), .A2(STATE_REG_SCAN_IN), .ZN(n4644) );
  XNOR2_X1 U2699 ( .A(n2263), .B(IR_REG_22__SCAN_IN), .ZN(n2932) );
  INV_X1 U2700 ( .A(IR_REG_21__SCAN_IN), .ZN(n2241) );
  INV_X1 U2701 ( .A(n4620), .ZN(n4646) );
  INV_X1 U2702 ( .A(n3877), .ZN(n4656) );
  INV_X1 U2703 ( .A(n3878), .ZN(n4660) );
  OAI21_X1 U2704 ( .B1(n2397), .B2(n2396), .A(n2414), .ZN(n4473) );
  INV_X1 U2705 ( .A(n2986), .ZN(n4497) );
  AND2_X1 U2706 ( .A1(n2337), .A2(n2318), .ZN(n4476) );
  NAND2_X1 U2707 ( .A1(n4488), .A2(IR_REG_31__SCAN_IN), .ZN(n2106) );
  NOR2_X1 U2708 ( .A1(n4626), .A2(n4625), .ZN(n4628) );
  OAI21_X1 U2709 ( .B1(n4624), .B2(n4623), .A(n4622), .ZN(n4625) );
  OR2_X1 U2710 ( .A1(n3493), .A2(n4417), .ZN(n2900) );
  OR2_X1 U2711 ( .A1(n4087), .A2(n4069), .ZN(n2032) );
  INV_X1 U2712 ( .A(n2159), .ZN(n2157) );
  NOR2_X1 U2713 ( .A1(n2515), .A2(n2160), .ZN(n2159) );
  OR2_X1 U2714 ( .A1(n4131), .A2(n2127), .ZN(n2033) );
  OR2_X1 U2715 ( .A1(n3184), .A2(n3233), .ZN(n2034) );
  AND2_X1 U2716 ( .A1(n2836), .A2(n4132), .ZN(n2035) );
  AND2_X1 U2717 ( .A1(n2134), .A2(n4308), .ZN(n2036) );
  XNOR2_X1 U2718 ( .A(n2513), .B(n2691), .ZN(n3461) );
  AOI22_X1 U2719 ( .A1(n4125), .A2(n2324), .B1(n2657), .B2(n3620), .ZN(n3612)
         );
  AND2_X1 U2720 ( .A1(n2132), .A2(n3957), .ZN(n2037) );
  INV_X1 U2721 ( .A(n4583), .ZN(n2142) );
  AND2_X1 U2722 ( .A1(n2037), .A2(n2720), .ZN(n2038) );
  INV_X1 U2723 ( .A(n3366), .ZN(n2135) );
  NAND4_X2 U2724 ( .A1(n2294), .A2(n2293), .A3(n2292), .A4(n2291), .ZN(n2809)
         );
  INV_X1 U2725 ( .A(n2780), .ZN(n2674) );
  NAND2_X1 U2726 ( .A1(n2997), .A2(n4497), .ZN(n2039) );
  NAND2_X1 U2727 ( .A1(n2174), .A2(n3566), .ZN(n3611) );
  NAND2_X1 U2728 ( .A1(n2949), .A2(n2222), .ZN(n2332) );
  MUX2_X1 U2729 ( .A(n4476), .B(DATAI_3_), .S(n2363), .Z(n3147) );
  XNOR2_X1 U2730 ( .A(n2215), .B(n2216), .ZN(n2222) );
  INV_X1 U2731 ( .A(n2222), .ZN(n4470) );
  NAND2_X1 U2732 ( .A1(n3506), .A2(n2681), .ZN(n3577) );
  AND2_X1 U2733 ( .A1(n4087), .A2(n4069), .ZN(n2040) );
  AND2_X1 U2734 ( .A1(n2071), .A2(n2841), .ZN(n2041) );
  NOR2_X1 U2735 ( .A1(n4008), .A2(n3992), .ZN(n2042) );
  AND2_X1 U2736 ( .A1(n2138), .A2(n3866), .ZN(n2043) );
  INV_X1 U2737 ( .A(n2803), .ZN(n2806) );
  AND2_X1 U2738 ( .A1(n2461), .A2(n2448), .ZN(n2044) );
  OR2_X1 U2739 ( .A1(n2839), .A2(n2840), .ZN(n2078) );
  NOR2_X1 U2740 ( .A1(n2828), .A2(n3366), .ZN(n2045) );
  XNOR2_X1 U2741 ( .A(n2304), .B(n2735), .ZN(n2305) );
  AND2_X1 U2742 ( .A1(n2214), .A2(n2213), .ZN(n2046) );
  OR2_X1 U2743 ( .A1(n3862), .A2(n4655), .ZN(n2047) );
  NAND2_X1 U2744 ( .A1(n3829), .A2(n3324), .ZN(n2048) );
  AND2_X1 U2745 ( .A1(n4600), .A2(n2116), .ZN(n2049) );
  NOR2_X1 U2746 ( .A1(n2166), .A2(n2162), .ZN(n2050) );
  NAND4_X1 U2747 ( .A1(n2277), .A2(n2276), .A3(n2275), .A4(n2274), .ZN(n2805)
         );
  OR2_X1 U2748 ( .A1(n2169), .A2(n2173), .ZN(n2051) );
  AND2_X1 U2749 ( .A1(n2406), .A2(n2422), .ZN(n2052) );
  NAND2_X1 U2750 ( .A1(n4099), .A2(n2838), .ZN(n4077) );
  NAND2_X1 U2751 ( .A1(n2075), .A2(n2078), .ZN(n4056) );
  OAI21_X1 U2752 ( .B1(n4099), .B2(n2074), .A(n2072), .ZN(n4039) );
  NAND2_X1 U2753 ( .A1(n2181), .A2(n2182), .ZN(n3391) );
  NAND2_X1 U2754 ( .A1(n2156), .A2(n2154), .ZN(n3497) );
  AND2_X1 U2755 ( .A1(n4126), .A2(n2835), .ZN(n2053) );
  NAND2_X1 U2756 ( .A1(n2178), .A2(n2448), .ZN(n3347) );
  NAND2_X1 U2757 ( .A1(n3559), .A2(n3434), .ZN(n2054) );
  INV_X1 U2758 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2111) );
  XOR2_X1 U2759 ( .A(n2765), .B(n2766), .Z(n3480) );
  AND2_X1 U2760 ( .A1(n2828), .A2(n3366), .ZN(n2055) );
  NOR2_X1 U2761 ( .A1(n3829), .A2(n3324), .ZN(n2056) );
  NAND2_X1 U2762 ( .A1(n4145), .A2(n4124), .ZN(n2057) );
  INV_X1 U2763 ( .A(n3460), .ZN(n2160) );
  AOI21_X1 U2764 ( .B1(n3500), .B2(n2324), .A(n2514), .ZN(n3460) );
  AND2_X1 U2765 ( .A1(n2155), .A2(n2154), .ZN(n2153) );
  BUF_X1 U2766 ( .A(n2259), .Z(n2853) );
  INV_X1 U2767 ( .A(n3526), .ZN(n4093) );
  INV_X1 U2768 ( .A(n3887), .ZN(n4655) );
  XNOR2_X1 U2769 ( .A(n2243), .B(IR_REG_26__SCAN_IN), .ZN(n2740) );
  INV_X1 U2770 ( .A(n3566), .ZN(n2171) );
  NAND2_X1 U2771 ( .A1(n3441), .A2(n2827), .ZN(n3364) );
  NAND2_X1 U2772 ( .A1(n2186), .A2(n2406), .ZN(n3259) );
  NAND2_X1 U2773 ( .A1(n3725), .A2(DATAI_24_), .ZN(n3992) );
  AND2_X1 U2774 ( .A1(n2536), .A2(n2535), .ZN(n2058) );
  AND2_X1 U2775 ( .A1(n3877), .A2(REG1_REG_11__SCAN_IN), .ZN(n2059) );
  NAND2_X1 U2776 ( .A1(n2178), .A2(n2044), .ZN(n3349) );
  INV_X1 U2777 ( .A(n2126), .ZN(n4068) );
  NOR3_X1 U2778 ( .A1(n4131), .A2(n2130), .A3(n3526), .ZN(n2126) );
  NAND2_X1 U2779 ( .A1(n2346), .A2(n2345), .ZN(n3195) );
  OAI21_X1 U2780 ( .B1(n3182), .B2(n2820), .A(n2819), .ZN(n3290) );
  INV_X1 U2781 ( .A(n2265), .ZN(n2804) );
  NOR2_X1 U2782 ( .A1(n3858), .A2(n4662), .ZN(n3859) );
  INV_X1 U2783 ( .A(n3859), .ZN(n2148) );
  NAND2_X1 U2784 ( .A1(n2286), .A2(n2198), .ZN(n3120) );
  AND2_X1 U2785 ( .A1(n3725), .A2(DATAI_27_), .ZN(n3941) );
  NAND2_X1 U2786 ( .A1(n3725), .A2(DATAI_26_), .ZN(n3957) );
  AND2_X1 U2787 ( .A1(n2145), .A2(n2989), .ZN(n2060) );
  AND2_X1 U2788 ( .A1(n4602), .A2(n2119), .ZN(n2061) );
  INV_X1 U2789 ( .A(n2117), .ZN(n2116) );
  OR2_X1 U2790 ( .A1(n4615), .A2(n2118), .ZN(n2117) );
  NAND2_X1 U2791 ( .A1(n2217), .A2(n2216), .ZN(n2939) );
  NAND2_X1 U2792 ( .A1(n3106), .A2(n3770), .ZN(n3105) );
  OAI21_X2 U2793 ( .B1(n3939), .B2(n3940), .A(n2885), .ZN(n3913) );
  OAI21_X2 U2794 ( .B1(n3967), .B2(n2883), .A(n3742), .ZN(n3949) );
  AOI21_X1 U2795 ( .B1(n3913), .B2(n3912), .A(n3911), .ZN(n3914) );
  NAND2_X1 U2796 ( .A1(n2857), .A2(n3666), .ZN(n3246) );
  NAND2_X1 U2797 ( .A1(n2864), .A2(n3692), .ZN(n3444) );
  OR2_X2 U2798 ( .A1(n3218), .A2(n3215), .ZN(n2860) );
  NAND2_X1 U2799 ( .A1(n2849), .A2(n2065), .ZN(n2064) );
  INV_X1 U2800 ( .A(n4099), .ZN(n2068) );
  AND2_X1 U2801 ( .A1(n4063), .A2(n4049), .ZN(n2081) );
  INV_X1 U2802 ( .A(n3428), .ZN(n2084) );
  NAND2_X1 U2803 ( .A1(n3290), .A2(n2824), .ZN(n2090) );
  INV_X1 U2804 ( .A(n2821), .ZN(n2092) );
  NAND2_X1 U2805 ( .A1(n2093), .A2(n2821), .ZN(n3279) );
  NAND2_X1 U2806 ( .A1(n2846), .A2(n2096), .ZN(n2094) );
  NAND2_X1 U2807 ( .A1(n2094), .A2(n2095), .ZN(n3948) );
  OAI21_X1 U2808 ( .B1(n3443), .B2(n2102), .A(n2100), .ZN(n3410) );
  NAND2_X1 U2809 ( .A1(n2244), .A2(n2211), .ZN(n2246) );
  MUX2_X1 U2810 ( .A(n2970), .B(REG2_REG_1__SCAN_IN), .S(n3013), .Z(n3006) );
  XNOR2_X2 U2811 ( .A(n2106), .B(n2249), .ZN(n3013) );
  NAND2_X1 U2812 ( .A1(n4495), .A2(n2039), .ZN(n2108) );
  OAI21_X1 U2813 ( .B1(n4495), .B2(n2111), .A(n2039), .ZN(n2110) );
  INV_X1 U2814 ( .A(n2113), .ZN(n3034) );
  NAND2_X1 U2815 ( .A1(n4601), .A2(n2061), .ZN(n2115) );
  NAND2_X1 U2816 ( .A1(n4601), .A2(n4602), .ZN(n4600) );
  INV_X1 U2817 ( .A(n2122), .ZN(n4577) );
  NOR2_X1 U2818 ( .A1(n4566), .A2(n3895), .ZN(n4579) );
  NAND2_X1 U2819 ( .A1(n2982), .A2(REG1_REG_3__SCAN_IN), .ZN(n2985) );
  NAND2_X1 U2820 ( .A1(n2966), .A2(n3841), .ZN(n2136) );
  NAND2_X1 U2821 ( .A1(n3867), .A2(n2142), .ZN(n2137) );
  NAND2_X1 U2822 ( .A1(n2139), .A2(n2137), .ZN(n4582) );
  NAND3_X1 U2823 ( .A1(n2141), .A2(n3866), .A3(n2140), .ZN(n2139) );
  NOR2_X1 U2824 ( .A1(n3859), .A2(n2149), .ZN(n4505) );
  NAND2_X1 U2825 ( .A1(n2148), .A2(n2150), .ZN(n4506) );
  NAND2_X1 U2826 ( .A1(n3858), .A2(n4662), .ZN(n2150) );
  INV_X1 U2827 ( .A(n3194), .ZN(n2346) );
  NAND2_X1 U2828 ( .A1(n3459), .A2(n2153), .ZN(n2151) );
  NAND2_X1 U2829 ( .A1(n3507), .A2(n2666), .ZN(n3506) );
  NAND2_X1 U2830 ( .A1(n3507), .A2(n2050), .ZN(n2161) );
  AOI21_X1 U2831 ( .B1(n3567), .B2(n3566), .A(n2176), .ZN(n2175) );
  INV_X1 U2832 ( .A(n3612), .ZN(n2176) );
  NAND2_X1 U2833 ( .A1(n2181), .A2(n2179), .ZN(n2502) );
  NAND2_X1 U2834 ( .A1(n2186), .A2(n2052), .ZN(n2427) );
  AND2_X2 U2835 ( .A1(n2197), .A2(n2191), .ZN(n2190) );
  AND4_X2 U2836 ( .A1(n2192), .A2(n2228), .A3(n2190), .A4(n2187), .ZN(n2244)
         );
  NAND3_X1 U2837 ( .A1(n2359), .A2(n2192), .A3(n2228), .ZN(n2262) );
  NAND2_X1 U2838 ( .A1(n2189), .A2(n2227), .ZN(n2193) );
  AND2_X2 U2839 ( .A1(n2473), .A2(n2208), .ZN(n2228) );
  NOR2_X1 U2840 ( .A1(n2246), .A2(n2196), .ZN(n2776) );
  XNOR2_X1 U2841 ( .A(n2264), .B(n2691), .ZN(n2288) );
  NAND2_X1 U2842 ( .A1(n2258), .A2(n2257), .ZN(n2264) );
  INV_X1 U2843 ( .A(n3641), .ZN(n2832) );
  INV_X1 U2844 ( .A(IR_REG_27__SCAN_IN), .ZN(n2213) );
  AND2_X1 U2845 ( .A1(n2316), .A2(n2338), .ZN(n2197) );
  OR2_X1 U2846 ( .A1(n2256), .A2(n2282), .ZN(n2198) );
  AND2_X1 U2847 ( .A1(n3988), .A2(n3545), .ZN(n2199) );
  INV_X1 U2848 ( .A(n3899), .ZN(n4647) );
  INV_X1 U2849 ( .A(n2732), .ZN(n2268) );
  INV_X1 U2850 ( .A(n4113), .ZN(n3620) );
  INV_X1 U2851 ( .A(IR_REG_30__SCAN_IN), .ZN(n2940) );
  AND2_X1 U2852 ( .A1(n2921), .A2(n4332), .ZN(n2922) );
  INV_X1 U2853 ( .A(n4649), .ZN(n3869) );
  NOR2_X1 U2854 ( .A1(n3272), .A2(n3267), .ZN(n2200) );
  INV_X1 U2855 ( .A(n3831), .ZN(n2818) );
  OR2_X1 U2856 ( .A1(n2288), .A2(n2287), .ZN(n2201) );
  OR2_X1 U2857 ( .A1(n4034), .A2(n3515), .ZN(n2202) );
  NOR2_X1 U2858 ( .A1(n4491), .A2(n4487), .ZN(n4607) );
  AND3_X1 U2859 ( .A1(n2796), .A2(n2795), .A3(n3608), .ZN(n2203) );
  INV_X1 U2860 ( .A(n3348), .ZN(n2461) );
  INV_X1 U2861 ( .A(n3198), .ZN(n2345) );
  NAND2_X1 U2862 ( .A1(n2303), .A2(n2302), .ZN(n2304) );
  INV_X1 U2863 ( .A(n3579), .ZN(n2683) );
  INV_X1 U2864 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3872) );
  NAND2_X1 U2865 ( .A1(n2808), .A2(n3133), .ZN(n2810) );
  AND2_X1 U2866 ( .A1(n3896), .A2(REG1_REG_15__SCAN_IN), .ZN(n3868) );
  NAND2_X1 U2867 ( .A1(n2837), .A2(n4113), .ZN(n2838) );
  INV_X1 U2868 ( .A(n4153), .ZN(n2835) );
  INV_X1 U2869 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2481) );
  NOR2_X1 U2870 ( .A1(n3762), .A2(n2200), .ZN(n2821) );
  INV_X1 U2871 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4276) );
  NAND2_X1 U2872 ( .A1(n2577), .A2(REG3_REG_17__SCAN_IN), .ZN(n2593) );
  OR2_X1 U2873 ( .A1(n3911), .A2(n2852), .ZN(n3924) );
  OR2_X1 U2874 ( .A1(n3970), .A2(n3951), .ZN(n3736) );
  OR2_X1 U2875 ( .A1(n2651), .A2(n3512), .ZN(n2670) );
  INV_X1 U2876 ( .A(n4046), .ZN(n2842) );
  AND2_X1 U2877 ( .A1(n2503), .A2(REG3_REG_13__SCAN_IN), .ZN(n2516) );
  INV_X1 U2878 ( .A(n3827), .ZN(n2828) );
  OR2_X1 U2879 ( .A1(n3830), .A2(n3305), .ZN(n3675) );
  NAND2_X1 U2880 ( .A1(n2708), .A2(n3624), .ZN(n3481) );
  NOR2_X1 U2881 ( .A1(n2619), .A2(n4211), .ZN(n2643) );
  OR2_X1 U2882 ( .A1(n2788), .A2(n2779), .ZN(n3648) );
  INV_X1 U2883 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3376) );
  INV_X1 U2884 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3644) );
  INV_X1 U2885 ( .A(n4478), .ZN(n3834) );
  AND2_X1 U2886 ( .A1(n3631), .A2(n3941), .ZN(n3800) );
  INV_X1 U2887 ( .A(n3826), .ZN(n4087) );
  OR2_X1 U2888 ( .A1(n4478), .A2(n2888), .ZN(n4327) );
  INV_X1 U2889 ( .A(n4327), .ZN(n4144) );
  INV_X1 U2890 ( .A(n2961), .ZN(n2791) );
  AND2_X1 U2891 ( .A1(n2752), .A2(n2953), .ZN(n2753) );
  INV_X1 U2892 ( .A(n3957), .ZN(n3951) );
  INV_X1 U2893 ( .A(n4132), .ZN(n4124) );
  OR2_X1 U2894 ( .A1(n2895), .A2(n3068), .ZN(n2916) );
  INV_X1 U2895 ( .A(IR_REG_7__SCAN_IN), .ZN(n2396) );
  INV_X1 U2896 ( .A(n4308), .ZN(n4322) );
  OR2_X1 U2897 ( .A1(n2604), .A2(n2603), .ZN(n2619) );
  NOR2_X1 U2898 ( .A1(n2554), .A2(n2553), .ZN(n2577) );
  OR2_X1 U2899 ( .A1(n4478), .A2(n3833), .ZN(n3837) );
  AND2_X1 U2900 ( .A1(n2718), .A2(n2717), .ZN(n3631) );
  AND4_X1 U2901 ( .A1(n2633), .A2(n2632), .A3(n2631), .A4(n2630), .ZN(n4063)
         );
  NAND2_X1 U2902 ( .A1(n4532), .A2(REG2_REG_10__SCAN_IN), .ZN(n4531) );
  NOR2_X1 U2903 ( .A1(n4491), .A2(n3834), .ZN(n4621) );
  AND2_X1 U2904 ( .A1(n3670), .A2(n3686), .ZN(n3768) );
  INV_X1 U2905 ( .A(n4633), .ZN(n4136) );
  AOI21_X1 U2906 ( .B1(n2754), .B2(n2954), .A(n2753), .ZN(n2902) );
  NAND2_X1 U2907 ( .A1(n3725), .A2(DATAI_25_), .ZN(n3974) );
  INV_X1 U2908 ( .A(n3267), .ZN(n3294) );
  NAND2_X1 U2909 ( .A1(n4067), .A2(n4700), .ZN(n4692) );
  AND2_X1 U2910 ( .A1(n2266), .A2(n2789), .ZN(n4676) );
  NAND2_X1 U2911 ( .A1(n2756), .A2(IR_REG_31__SCAN_IN), .ZN(n2245) );
  AND2_X1 U2912 ( .A1(n2440), .A2(n2455), .ZN(n3878) );
  AND2_X1 U2913 ( .A1(n2978), .A2(n2977), .ZN(n4599) );
  INV_X1 U2914 ( .A(n3650), .ZN(n3617) );
  OR2_X1 U2915 ( .A1(n2792), .A2(n2763), .ZN(n3653) );
  INV_X1 U2916 ( .A(n4621), .ZN(n4612) );
  INV_X1 U2917 ( .A(n4607), .ZN(n4618) );
  INV_X1 U2918 ( .A(n3928), .ZN(n4159) );
  NAND2_X1 U2919 ( .A1(n4718), .A2(n2899), .ZN(n4417) );
  OR2_X1 U2920 ( .A1(n3493), .A2(n4468), .ZN(n2906) );
  AND3_X1 U2921 ( .A1(n4697), .A2(n4696), .A3(n4695), .ZN(n4714) );
  INV_X1 U2922 ( .A(n4706), .ZN(n4704) );
  INV_X1 U2923 ( .A(n4471), .ZN(n2953) );
  INV_X1 U2924 ( .A(n3890), .ZN(n4653) );
  INV_X1 U2925 ( .A(n2999), .ZN(n4475) );
  INV_X2 U2926 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2927 ( .A(IR_REG_9__SCAN_IN), .ZN(n2205) );
  AND3_X2 U2928 ( .A1(n2206), .A2(n2205), .A3(n2204), .ZN(n2439) );
  AND2_X2 U2929 ( .A1(n2439), .A2(n2207), .ZN(n2473) );
  NOR2_X2 U2930 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2238)
         );
  NAND4_X1 U2931 ( .A1(n2238), .A2(n2231), .A3(n2525), .A4(n4235), .ZN(n2209)
         );
  NAND2_X1 U2932 ( .A1(n2295), .A2(n2296), .ZN(n2315) );
  INV_X2 U2933 ( .A(IR_REG_3__SCAN_IN), .ZN(n2316) );
  INV_X2 U2934 ( .A(IR_REG_4__SCAN_IN), .ZN(n2338) );
  XNOR2_X2 U2935 ( .A(n2218), .B(IR_REG_30__SCAN_IN), .ZN(n2949) );
  NAND2_X1 U2936 ( .A1(n2272), .A2(REG0_REG_1__SCAN_IN), .ZN(n2220) );
  NOR2_X1 U2937 ( .A1(n2949), .A2(n2222), .ZN(n2273) );
  NAND2_X1 U2938 ( .A1(n2273), .A2(REG1_REG_1__SCAN_IN), .ZN(n2219) );
  AND2_X1 U2939 ( .A1(n2220), .A2(n2219), .ZN(n2226) );
  INV_X1 U2940 ( .A(n2332), .ZN(n2221) );
  NAND2_X1 U2941 ( .A1(n2221), .A2(REG2_REG_1__SCAN_IN), .ZN(n2225) );
  INV_X1 U2942 ( .A(n2309), .ZN(n2223) );
  NAND2_X1 U2943 ( .A1(n2223), .A2(REG3_REG_1__SCAN_IN), .ZN(n2224) );
  NAND3_X1 U2944 ( .A1(n2226), .A2(n2225), .A3(n2224), .ZN(n2265) );
  AND2_X2 U2945 ( .A1(n2359), .A2(n2227), .ZN(n2380) );
  NAND2_X1 U2946 ( .A1(n2380), .A2(n2228), .ZN(n2509) );
  NAND3_X1 U2947 ( .A1(n2546), .A2(n2525), .A3(n2561), .ZN(n2230) );
  NAND2_X1 U2948 ( .A1(n2584), .A2(n2231), .ZN(n2599) );
  INV_X1 U2949 ( .A(n2599), .ZN(n2233) );
  NAND2_X1 U2950 ( .A1(n2233), .A2(n2232), .ZN(n2234) );
  NAND2_X1 U2951 ( .A1(n2260), .A2(n2261), .ZN(n2235) );
  INV_X1 U2952 ( .A(n2238), .ZN(n2239) );
  NAND2_X1 U2953 ( .A1(n2239), .A2(IR_REG_31__SCAN_IN), .ZN(n2240) );
  NAND2_X1 U2954 ( .A1(n2260), .A2(n2240), .ZN(n2242) );
  XNOR2_X2 U2955 ( .A(n2242), .B(n2241), .ZN(n2267) );
  NAND2_X1 U2956 ( .A1(n2250), .A2(IR_REG_31__SCAN_IN), .ZN(n2243) );
  NAND2_X1 U2957 ( .A1(n2246), .A2(IR_REG_31__SCAN_IN), .ZN(n2248) );
  INV_X1 U2958 ( .A(n2256), .ZN(n2283) );
  NAND2_X1 U2959 ( .A1(n2265), .A2(n2657), .ZN(n2258) );
  INV_X1 U2960 ( .A(IR_REG_1__SCAN_IN), .ZN(n2249) );
  INV_X1 U2961 ( .A(DATAI_1_), .ZN(n2255) );
  NAND2_X1 U2962 ( .A1(n2252), .A2(n2251), .ZN(n2254) );
  NAND2_X1 U2963 ( .A1(n2777), .A2(IR_REG_27__SCAN_IN), .ZN(n2253) );
  MUX2_X1 U2964 ( .A(n3013), .B(n2255), .S(n2319), .Z(n2803) );
  OR2_X1 U2965 ( .A1(n2803), .A2(n2732), .ZN(n2257) );
  NAND2_X1 U2966 ( .A1(n2262), .A2(IR_REG_31__SCAN_IN), .ZN(n2263) );
  NAND2_X1 U2967 ( .A1(n3905), .A2(n2932), .ZN(n2771) );
  INV_X1 U2968 ( .A(n2760), .ZN(n2790) );
  AND2_X2 U2969 ( .A1(n2790), .A2(n3816), .ZN(n2761) );
  AND2_X4 U2970 ( .A1(n2266), .A2(n2761), .ZN(n2899) );
  NOR2_X1 U2971 ( .A1(n2803), .A2(n2325), .ZN(n2270) );
  XNOR2_X1 U2972 ( .A(n2288), .B(n2287), .ZN(n3064) );
  INV_X1 U2973 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2271) );
  NAND2_X1 U2974 ( .A1(n2221), .A2(REG2_REG_0__SCAN_IN), .ZN(n2274) );
  NAND2_X1 U2975 ( .A1(n2805), .A2(n2657), .ZN(n2281) );
  BUF_X4 U2976 ( .A(n2319), .Z(n2363) );
  NAND2_X1 U2977 ( .A1(n3124), .A2(n2268), .ZN(n2280) );
  AND2_X1 U2978 ( .A1(n2281), .A2(n2280), .ZN(n2286) );
  INV_X1 U2979 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2282) );
  NAND2_X1 U2980 ( .A1(n2805), .A2(n2029), .ZN(n2285) );
  AOI22_X1 U2981 ( .A1(n3124), .A2(n2657), .B1(n2283), .B2(n4488), .ZN(n2284)
         );
  OAI21_X1 U2982 ( .B1(n3064), .B2(n3065), .A(n2201), .ZN(n2289) );
  INV_X1 U2983 ( .A(n2289), .ZN(n3094) );
  NAND2_X1 U2984 ( .A1(n2272), .A2(REG0_REG_2__SCAN_IN), .ZN(n2294) );
  NAND2_X1 U2985 ( .A1(n2273), .A2(REG1_REG_2__SCAN_IN), .ZN(n2293) );
  INV_X1 U2986 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2290) );
  INV_X1 U2987 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2968) );
  OR2_X1 U2988 ( .A1(n2295), .A2(n2775), .ZN(n2297) );
  INV_X1 U2989 ( .A(DATAI_2_), .ZN(n2298) );
  NOR2_X1 U2990 ( .A1(n3101), .A2(n2325), .ZN(n2301) );
  AOI21_X1 U2991 ( .B1(n2809), .B2(n2324), .A(n2301), .ZN(n2306) );
  NAND2_X1 U2992 ( .A1(n2809), .A2(n2657), .ZN(n2303) );
  OR2_X1 U2993 ( .A1(n3101), .A2(n2732), .ZN(n2302) );
  XNOR2_X1 U2994 ( .A(n2306), .B(n2305), .ZN(n3093) );
  NAND2_X1 U2995 ( .A1(n3094), .A2(n3093), .ZN(n3095) );
  INV_X1 U2996 ( .A(n2305), .ZN(n2307) );
  NAND2_X1 U2997 ( .A1(n2307), .A2(n2306), .ZN(n2308) );
  NAND2_X1 U2998 ( .A1(n3095), .A2(n2308), .ZN(n3145) );
  NAND2_X1 U2999 ( .A1(n3720), .A2(REG1_REG_3__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U3000 ( .A1(n2272), .A2(REG0_REG_3__SCAN_IN), .ZN(n2313) );
  INV_X1 U3002 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2310) );
  OR2_X1 U3003 ( .A1(n2332), .A2(n2310), .ZN(n2311) );
  NAND4_X2 U3004 ( .A1(n2314), .A2(n2313), .A3(n2312), .A4(n2311), .ZN(n2323)
         );
  NAND2_X1 U3005 ( .A1(n2323), .A2(n2657), .ZN(n2321) );
  NAND2_X1 U3006 ( .A1(n2315), .A2(IR_REG_31__SCAN_IN), .ZN(n2317) );
  NAND2_X1 U3007 ( .A1(n2317), .A2(n2316), .ZN(n2337) );
  OR2_X1 U3008 ( .A1(n2317), .A2(n2316), .ZN(n2318) );
  NAND2_X1 U3009 ( .A1(n3147), .A2(n2268), .ZN(n2320) );
  AND2_X1 U3010 ( .A1(n3147), .A2(n2657), .ZN(n2326) );
  AOI21_X1 U3011 ( .B1(n2323), .B2(n2324), .A(n2326), .ZN(n2328) );
  XNOR2_X1 U3012 ( .A(n2327), .B(n2328), .ZN(n3146) );
  NAND2_X1 U3013 ( .A1(n3145), .A2(n3146), .ZN(n2331) );
  INV_X1 U3014 ( .A(n2327), .ZN(n2329) );
  NAND2_X1 U3015 ( .A1(n2329), .A2(n2328), .ZN(n2330) );
  NAND2_X1 U3016 ( .A1(n3720), .A2(REG1_REG_4__SCAN_IN), .ZN(n2336) );
  NAND2_X1 U3017 ( .A1(n2780), .A2(REG0_REG_4__SCAN_IN), .ZN(n2335) );
  INV_X2 U3018 ( .A(n2221), .ZN(n3724) );
  NAND2_X1 U3019 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2351) );
  OAI21_X1 U3020 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2351), .ZN(n3255) );
  INV_X1 U3021 ( .A(n2325), .ZN(n2675) );
  NAND2_X1 U3022 ( .A1(n3222), .A2(n2675), .ZN(n2342) );
  NAND2_X1 U3023 ( .A1(n2337), .A2(IR_REG_31__SCAN_IN), .ZN(n2339) );
  XNOR2_X1 U3024 ( .A(n2339), .B(n2338), .ZN(n2986) );
  INV_X1 U3025 ( .A(DATAI_4_), .ZN(n2340) );
  MUX2_X1 U3026 ( .A(n2986), .B(n2340), .S(n2363), .Z(n3253) );
  OR2_X1 U3027 ( .A1(n3253), .A2(n2031), .ZN(n2341) );
  NAND2_X1 U3028 ( .A1(n2342), .A2(n2341), .ZN(n2343) );
  NOR2_X1 U3029 ( .A1(n3253), .A2(n2773), .ZN(n2344) );
  AOI21_X1 U3030 ( .B1(n3222), .B2(n2324), .A(n2344), .ZN(n2347) );
  XNOR2_X1 U3031 ( .A(n2348), .B(n2347), .ZN(n3198) );
  OR2_X1 U3032 ( .A1(n2348), .A2(n2347), .ZN(n2349) );
  NAND2_X1 U3033 ( .A1(n3195), .A2(n2349), .ZN(n3155) );
  NAND2_X1 U3034 ( .A1(n3720), .A2(REG1_REG_5__SCAN_IN), .ZN(n2356) );
  NAND2_X1 U3035 ( .A1(n2780), .A2(REG0_REG_5__SCAN_IN), .ZN(n2355) );
  AND2_X1 U3036 ( .A1(n2351), .A2(n2350), .ZN(n2352) );
  NOR2_X1 U3037 ( .A1(n2351), .A2(n2350), .ZN(n2373) );
  OR2_X1 U3038 ( .A1(n2352), .A2(n2373), .ZN(n3227) );
  OR2_X1 U3039 ( .A1(n2786), .A2(n3227), .ZN(n2354) );
  INV_X1 U3040 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3223) );
  OR2_X1 U3041 ( .A1(n3724), .A2(n3223), .ZN(n2353) );
  NAND4_X1 U3042 ( .A1(n2356), .A2(n2355), .A3(n2354), .A4(n2353), .ZN(n3832)
         );
  INV_X1 U3043 ( .A(n2325), .ZN(n2731) );
  NAND2_X1 U3044 ( .A1(n3832), .A2(n2731), .ZN(n2365) );
  NAND2_X1 U3045 ( .A1(n2357), .A2(IR_REG_31__SCAN_IN), .ZN(n2358) );
  MUX2_X1 U3046 ( .A(IR_REG_31__SCAN_IN), .B(n2358), .S(IR_REG_5__SCAN_IN), 
        .Z(n2362) );
  INV_X1 U3047 ( .A(n2360), .ZN(n2361) );
  MUX2_X1 U3048 ( .A(n3031), .B(DATAI_5_), .S(n3725), .Z(n3224) );
  NAND2_X1 U3049 ( .A1(n3224), .A2(n2268), .ZN(n2364) );
  NAND2_X1 U3050 ( .A1(n2365), .A2(n2364), .ZN(n2366) );
  XNOR2_X1 U3051 ( .A(n2366), .B(n2735), .ZN(n2370) );
  AND2_X1 U3052 ( .A1(n3224), .A2(n2731), .ZN(n2367) );
  AOI21_X1 U3053 ( .B1(n3832), .B2(n2324), .A(n2367), .ZN(n2368) );
  XNOR2_X1 U3054 ( .A(n2370), .B(n2368), .ZN(n3158) );
  INV_X1 U3055 ( .A(n2368), .ZN(n2369) );
  NAND2_X1 U3056 ( .A1(n2370), .A2(n2369), .ZN(n2371) );
  NAND2_X1 U3057 ( .A1(n3720), .A2(REG1_REG_6__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U3058 ( .A1(n2780), .A2(REG0_REG_6__SCAN_IN), .ZN(n2377) );
  INV_X1 U3059 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2372) );
  OR2_X1 U3060 ( .A1(n3724), .A2(n2372), .ZN(n2376) );
  NAND2_X1 U3061 ( .A1(n2373), .A2(REG3_REG_6__SCAN_IN), .ZN(n2390) );
  OR2_X1 U3062 ( .A1(n2373), .A2(REG3_REG_6__SCAN_IN), .ZN(n2374) );
  NAND2_X1 U3063 ( .A1(n2390), .A2(n2374), .ZN(n3168) );
  OR2_X1 U3064 ( .A1(n2786), .A2(n3168), .ZN(n2375) );
  NAND4_X1 U3065 ( .A1(n2378), .A2(n2377), .A3(n2376), .A4(n2375), .ZN(n3831)
         );
  NAND2_X1 U3066 ( .A1(n3831), .A2(n2324), .ZN(n2384) );
  NOR2_X1 U3067 ( .A1(n2360), .A2(n2775), .ZN(n2379) );
  MUX2_X1 U3068 ( .A(n2775), .B(n2379), .S(IR_REG_6__SCAN_IN), .Z(n2382) );
  OR2_X1 U3069 ( .A1(n2382), .A2(n2381), .ZN(n2999) );
  MUX2_X1 U3070 ( .A(n4475), .B(DATAI_6_), .S(n3725), .Z(n3184) );
  NAND2_X1 U3071 ( .A1(n3184), .A2(n2731), .ZN(n2383) );
  NAND2_X1 U3072 ( .A1(n3831), .A2(n2731), .ZN(n2386) );
  NAND2_X1 U3073 ( .A1(n3184), .A2(n2268), .ZN(n2385) );
  NAND2_X1 U3074 ( .A1(n2386), .A2(n2385), .ZN(n2387) );
  OAI21_X2 U3075 ( .B1(n3164), .B2(n3166), .A(n3165), .ZN(n2389) );
  NAND2_X1 U3076 ( .A1(n3164), .A2(n3166), .ZN(n2388) );
  NAND2_X1 U3077 ( .A1(n2389), .A2(n2388), .ZN(n3231) );
  NAND2_X1 U3078 ( .A1(n3720), .A2(REG1_REG_7__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3079 ( .A1(n2780), .A2(REG0_REG_7__SCAN_IN), .ZN(n2394) );
  INV_X1 U3080 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3019) );
  OR2_X1 U3081 ( .A1(n3724), .A2(n3019), .ZN(n2393) );
  NAND2_X1 U3082 ( .A1(n2390), .A2(n4251), .ZN(n2391) );
  NAND2_X1 U3083 ( .A1(n2408), .A2(n2391), .ZN(n3309) );
  OR2_X1 U3084 ( .A1(n2786), .A2(n3309), .ZN(n2392) );
  NAND4_X1 U3085 ( .A1(n2395), .A2(n2394), .A3(n2393), .A4(n2392), .ZN(n3830)
         );
  NAND2_X1 U3086 ( .A1(n3830), .A2(n2731), .ZN(n2400) );
  OR2_X1 U3087 ( .A1(n2381), .A2(n2775), .ZN(n2397) );
  NAND2_X1 U3088 ( .A1(n2397), .A2(n2396), .ZN(n2414) );
  INV_X1 U3089 ( .A(DATAI_7_), .ZN(n2398) );
  MUX2_X1 U3090 ( .A(n4473), .B(n2398), .S(n3725), .Z(n3305) );
  OR2_X1 U3091 ( .A1(n3305), .A2(n2732), .ZN(n2399) );
  NAND2_X1 U3092 ( .A1(n2400), .A2(n2399), .ZN(n2401) );
  XNOR2_X1 U3093 ( .A(n2401), .B(n2735), .ZN(n2403) );
  NOR2_X1 U3094 ( .A1(n3305), .A2(n2773), .ZN(n2402) );
  AOI21_X1 U3095 ( .B1(n3830), .B2(n2324), .A(n2402), .ZN(n2404) );
  INV_X1 U3096 ( .A(n2403), .ZN(n2405) );
  OR2_X1 U3097 ( .A1(n2405), .A2(n2404), .ZN(n2406) );
  NAND2_X1 U3098 ( .A1(n3720), .A2(REG1_REG_8__SCAN_IN), .ZN(n2413) );
  NAND2_X1 U3099 ( .A1(n2780), .A2(REG0_REG_8__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3100 ( .A1(n2408), .A2(n2407), .ZN(n2409) );
  NAND2_X1 U3101 ( .A1(n2429), .A2(n2409), .ZN(n3295) );
  OR2_X1 U3102 ( .A1(n2786), .A2(n3295), .ZN(n2411) );
  INV_X1 U3103 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3296) );
  OR2_X1 U3104 ( .A1(n3724), .A2(n3296), .ZN(n2410) );
  NAND4_X1 U3105 ( .A1(n2413), .A2(n2412), .A3(n2411), .A4(n2410), .ZN(n3272)
         );
  NAND2_X1 U3106 ( .A1(n3272), .A2(n2731), .ZN(n2418) );
  NAND2_X1 U3107 ( .A1(n2414), .A2(IR_REG_31__SCAN_IN), .ZN(n2416) );
  INV_X1 U3108 ( .A(IR_REG_8__SCAN_IN), .ZN(n2415) );
  XNOR2_X1 U3109 ( .A(n2416), .B(n2415), .ZN(n4662) );
  INV_X1 U3110 ( .A(n4662), .ZN(n3880) );
  MUX2_X1 U3111 ( .A(n3880), .B(DATAI_8_), .S(n3725), .Z(n3267) );
  NAND2_X1 U3112 ( .A1(n3267), .A2(n2268), .ZN(n2417) );
  NAND2_X1 U3113 ( .A1(n2418), .A2(n2417), .ZN(n2419) );
  XNOR2_X1 U3114 ( .A(n2419), .B(n2735), .ZN(n2423) );
  NAND2_X1 U3115 ( .A1(n3272), .A2(n2324), .ZN(n2421) );
  NAND2_X1 U3116 ( .A1(n3267), .A2(n2731), .ZN(n2420) );
  NAND2_X1 U3117 ( .A1(n2421), .A2(n2420), .ZN(n2424) );
  AND2_X1 U3118 ( .A1(n2423), .A2(n2424), .ZN(n3261) );
  INV_X1 U3119 ( .A(n3261), .ZN(n2422) );
  INV_X1 U3120 ( .A(n2423), .ZN(n2426) );
  INV_X1 U3121 ( .A(n2424), .ZN(n2425) );
  NAND2_X1 U3122 ( .A1(n2426), .A2(n2425), .ZN(n3260) );
  NAND2_X1 U3123 ( .A1(n2427), .A2(n3260), .ZN(n3322) );
  NAND2_X1 U3124 ( .A1(n3720), .A2(REG1_REG_9__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U3125 ( .A1(n2780), .A2(REG0_REG_9__SCAN_IN), .ZN(n2434) );
  INV_X1 U3126 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2428) );
  OR2_X1 U3127 ( .A1(n3724), .A2(n2428), .ZN(n2433) );
  INV_X1 U3128 ( .A(n2449), .ZN(n2431) );
  NAND2_X1 U3129 ( .A1(n2429), .A2(n3325), .ZN(n2430) );
  NAND2_X1 U3130 ( .A1(n2431), .A2(n2430), .ZN(n3282) );
  OR2_X1 U3131 ( .A1(n2786), .A2(n3282), .ZN(n2432) );
  NAND4_X1 U3132 ( .A1(n2435), .A2(n2434), .A3(n2433), .A4(n2432), .ZN(n3829)
         );
  NAND2_X1 U3133 ( .A1(n3829), .A2(n2731), .ZN(n2442) );
  NOR2_X1 U3134 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2436)
         );
  NAND2_X1 U3135 ( .A1(n2381), .A2(n2436), .ZN(n2437) );
  NAND2_X1 U3136 ( .A1(n2437), .A2(IR_REG_31__SCAN_IN), .ZN(n2438) );
  MUX2_X1 U3137 ( .A(IR_REG_31__SCAN_IN), .B(n2438), .S(IR_REG_9__SCAN_IN), 
        .Z(n2440) );
  NAND2_X1 U3138 ( .A1(n2381), .A2(n2439), .ZN(n2455) );
  MUX2_X1 U3139 ( .A(n3878), .B(DATAI_9_), .S(n3725), .Z(n3324) );
  NAND2_X1 U3140 ( .A1(n3324), .A2(n2268), .ZN(n2441) );
  NAND2_X1 U3141 ( .A1(n2442), .A2(n2441), .ZN(n2443) );
  XNOR2_X1 U3142 ( .A(n2443), .B(n2735), .ZN(n2445) );
  AND2_X1 U3143 ( .A1(n3324), .A2(n2675), .ZN(n2444) );
  AOI21_X1 U3144 ( .B1(n3829), .B2(n2324), .A(n2444), .ZN(n2446) );
  INV_X1 U3145 ( .A(n2445), .ZN(n2447) );
  NAND2_X1 U3146 ( .A1(n2447), .A2(n2446), .ZN(n2448) );
  NAND2_X1 U3147 ( .A1(n3720), .A2(REG1_REG_10__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U31480 ( .A1(n2780), .A2(REG0_REG_10__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U31490 ( .A1(n2449), .A2(REG3_REG_10__SCAN_IN), .ZN(n2467) );
  OR2_X1 U3150 ( .A1(n2449), .A2(REG3_REG_10__SCAN_IN), .ZN(n2450) );
  NAND2_X1 U3151 ( .A1(n2467), .A2(n2450), .ZN(n3357) );
  OR2_X1 U3152 ( .A1(n2786), .A2(n3357), .ZN(n2452) );
  INV_X1 U3153 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3342) );
  OR2_X1 U3154 ( .A1(n3724), .A2(n3342), .ZN(n2451) );
  NAND4_X1 U3155 ( .A1(n2454), .A2(n2453), .A3(n2452), .A4(n2451), .ZN(n3828)
         );
  NAND2_X1 U3156 ( .A1(n3828), .A2(n2675), .ZN(n2458) );
  NAND2_X1 U3157 ( .A1(n2455), .A2(IR_REG_31__SCAN_IN), .ZN(n2456) );
  XNOR2_X1 U3158 ( .A(n2456), .B(IR_REG_10__SCAN_IN), .ZN(n3883) );
  MUX2_X1 U3159 ( .A(n3883), .B(DATAI_10_), .S(n3725), .Z(n3354) );
  NAND2_X1 U3160 ( .A1(n3354), .A2(n2268), .ZN(n2457) );
  NAND2_X1 U3161 ( .A1(n2458), .A2(n2457), .ZN(n2459) );
  XNOR2_X1 U3162 ( .A(n2459), .B(n2691), .ZN(n2462) );
  AND2_X1 U3163 ( .A1(n3354), .A2(n2675), .ZN(n2460) );
  AOI21_X1 U3164 ( .B1(n3828), .B2(n2324), .A(n2460), .ZN(n2463) );
  XNOR2_X1 U3165 ( .A(n2462), .B(n2463), .ZN(n3348) );
  INV_X1 U3166 ( .A(n2462), .ZN(n2465) );
  INV_X1 U3167 ( .A(n2463), .ZN(n2464) );
  NAND2_X1 U3168 ( .A1(n2465), .A2(n2464), .ZN(n2466) );
  NAND2_X1 U3169 ( .A1(n3720), .A2(REG1_REG_11__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U3170 ( .A1(n2780), .A2(REG0_REG_11__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U3171 ( .A1(n2467), .A2(n3376), .ZN(n2468) );
  NAND2_X1 U3172 ( .A1(n2482), .A2(n2468), .ZN(n3453) );
  OR2_X1 U3173 ( .A1(n2786), .A2(n3453), .ZN(n2470) );
  INV_X1 U3174 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3454) );
  OR2_X1 U3175 ( .A1(n3724), .A2(n3454), .ZN(n2469) );
  NAND4_X1 U3176 ( .A1(n2472), .A2(n2471), .A3(n2470), .A4(n2469), .ZN(n3396)
         );
  NAND2_X1 U3177 ( .A1(n3396), .A2(n2324), .ZN(n2477) );
  AND2_X1 U3178 ( .A1(n2473), .A2(n2381), .ZN(n2474) );
  INV_X1 U3179 ( .A(DATAI_11_), .ZN(n2475) );
  MUX2_X1 U3180 ( .A(n4656), .B(n2475), .S(n3725), .Z(n3451) );
  OR2_X1 U3181 ( .A1(n3451), .A2(n2773), .ZN(n2476) );
  NAND2_X1 U3182 ( .A1(n3396), .A2(n2657), .ZN(n2479) );
  OR2_X1 U3183 ( .A1(n3451), .A2(n2031), .ZN(n2478) );
  NAND2_X1 U3184 ( .A1(n2479), .A2(n2478), .ZN(n2480) );
  NAND2_X1 U3185 ( .A1(n3720), .A2(REG1_REG_12__SCAN_IN), .ZN(n2488) );
  NAND2_X1 U3186 ( .A1(n2780), .A2(REG0_REG_12__SCAN_IN), .ZN(n2487) );
  INV_X1 U3187 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3367) );
  OR2_X1 U3188 ( .A1(n3724), .A2(n3367), .ZN(n2486) );
  INV_X1 U3189 ( .A(n2503), .ZN(n2484) );
  NAND2_X1 U3190 ( .A1(n2482), .A2(n2481), .ZN(n2483) );
  NAND2_X1 U3191 ( .A1(n2484), .A2(n2483), .ZN(n3398) );
  OR2_X1 U3192 ( .A1(n2786), .A2(n3398), .ZN(n2485) );
  NAND4_X1 U3193 ( .A1(n2488), .A2(n2487), .A3(n2486), .A4(n2485), .ZN(n3827)
         );
  NAND2_X1 U3194 ( .A1(n3827), .A2(n2675), .ZN(n2494) );
  INV_X1 U3195 ( .A(IR_REG_11__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U3196 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  NAND2_X1 U3197 ( .A1(n2491), .A2(IR_REG_31__SCAN_IN), .ZN(n2492) );
  XNOR2_X1 U3198 ( .A(n2492), .B(IR_REG_12__SCAN_IN), .ZN(n3887) );
  INV_X1 U3199 ( .A(DATAI_12_), .ZN(n4654) );
  MUX2_X1 U3200 ( .A(n4655), .B(n4654), .S(n3725), .Z(n3366) );
  OR2_X1 U3201 ( .A1(n3366), .A2(n2031), .ZN(n2493) );
  NAND2_X1 U3202 ( .A1(n2494), .A2(n2493), .ZN(n2495) );
  XNOR2_X1 U3203 ( .A(n2495), .B(n2735), .ZN(n2498) );
  NAND2_X1 U3204 ( .A1(n3827), .A2(n2324), .ZN(n2497) );
  OR2_X1 U3205 ( .A1(n3366), .A2(n2773), .ZN(n2496) );
  NAND2_X1 U3206 ( .A1(n2497), .A2(n2496), .ZN(n2499) );
  AND2_X1 U3207 ( .A1(n2498), .A2(n2499), .ZN(n3393) );
  INV_X1 U3208 ( .A(n2498), .ZN(n2501) );
  INV_X1 U3209 ( .A(n2499), .ZN(n2500) );
  NAND2_X1 U32100 ( .A1(n2501), .A2(n2500), .ZN(n3392) );
  NAND2_X1 U32110 ( .A1(n3720), .A2(REG1_REG_13__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U32120 ( .A1(n2780), .A2(REG0_REG_13__SCAN_IN), .ZN(n2507) );
  INV_X1 U32130 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3423) );
  OR2_X1 U32140 ( .A1(n3724), .A2(n3423), .ZN(n2506) );
  NOR2_X1 U32150 ( .A1(n2503), .A2(REG3_REG_13__SCAN_IN), .ZN(n2504) );
  OR2_X1 U32160 ( .A1(n2516), .A2(n2504), .ZN(n3463) );
  OR2_X1 U32170 ( .A1(n2786), .A2(n3463), .ZN(n2505) );
  NAND4_X1 U32180 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n3500)
         );
  NAND2_X1 U32190 ( .A1(n3500), .A2(n2675), .ZN(n2512) );
  NAND2_X1 U32200 ( .A1(n2509), .A2(IR_REG_31__SCAN_IN), .ZN(n2510) );
  XNOR2_X1 U32210 ( .A(n2510), .B(IR_REG_13__SCAN_IN), .ZN(n3890) );
  INV_X1 U32220 ( .A(DATAI_13_), .ZN(n4652) );
  MUX2_X1 U32230 ( .A(n4653), .B(n4652), .S(n2363), .Z(n3421) );
  OR2_X1 U32240 ( .A1(n3421), .A2(n2031), .ZN(n2511) );
  NAND2_X1 U32250 ( .A1(n2512), .A2(n2511), .ZN(n2513) );
  NOR2_X1 U32260 ( .A1(n3421), .A2(n2773), .ZN(n2514) );
  INV_X1 U32270 ( .A(n3461), .ZN(n2515) );
  NAND2_X1 U32280 ( .A1(n3720), .A2(REG1_REG_14__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32290 ( .A1(n2780), .A2(REG0_REG_14__SCAN_IN), .ZN(n2521) );
  OR2_X1 U32300 ( .A1(n2516), .A2(REG3_REG_14__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32310 ( .A1(n2538), .A2(n2517), .ZN(n4331) );
  OR2_X1 U32320 ( .A1(n2786), .A2(n4331), .ZN(n2520) );
  INV_X1 U32330 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2518) );
  OR2_X1 U32340 ( .A1(n3724), .A2(n2518), .ZN(n2519) );
  NAND4_X1 U32350 ( .A1(n2522), .A2(n2521), .A3(n2520), .A4(n2519), .ZN(n3641)
         );
  NAND2_X1 U32360 ( .A1(n3641), .A2(n2731), .ZN(n2529) );
  NAND2_X1 U32370 ( .A1(n2524), .A2(IR_REG_31__SCAN_IN), .ZN(n2526) );
  XNOR2_X1 U32380 ( .A(n2526), .B(n2525), .ZN(n3891) );
  INV_X1 U32390 ( .A(DATAI_14_), .ZN(n2527) );
  MUX2_X1 U32400 ( .A(n3891), .B(n2527), .S(n3725), .Z(n4308) );
  OR2_X1 U32410 ( .A1(n4308), .A2(n2031), .ZN(n2528) );
  NAND2_X1 U32420 ( .A1(n2529), .A2(n2528), .ZN(n2530) );
  XNOR2_X1 U32430 ( .A(n2530), .B(n2735), .ZN(n2533) );
  NAND2_X1 U32440 ( .A1(n3641), .A2(n2324), .ZN(n2532) );
  OR2_X1 U32450 ( .A1(n4308), .A2(n2773), .ZN(n2531) );
  NAND2_X1 U32460 ( .A1(n2532), .A2(n2531), .ZN(n2534) );
  INV_X1 U32470 ( .A(n2533), .ZN(n2536) );
  INV_X1 U32480 ( .A(n2534), .ZN(n2535) );
  NAND2_X1 U32490 ( .A1(n3720), .A2(REG1_REG_15__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U32500 ( .A1(n2780), .A2(REG0_REG_15__SCAN_IN), .ZN(n2542) );
  INV_X1 U32510 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2537) );
  OR2_X1 U32520 ( .A1(n3724), .A2(n2537), .ZN(n2541) );
  NAND2_X1 U32530 ( .A1(n2538), .A2(n3644), .ZN(n2539) );
  NAND2_X1 U32540 ( .A1(n2554), .A2(n2539), .ZN(n3436) );
  OR2_X1 U32550 ( .A1(n2786), .A2(n3436), .ZN(n2540) );
  NAND4_X1 U32560 ( .A1(n2543), .A2(n2542), .A3(n2541), .A4(n2540), .ZN(n4324)
         );
  NAND2_X1 U32570 ( .A1(n4324), .A2(n2731), .ZN(n2550) );
  OR2_X1 U32580 ( .A1(n2524), .A2(IR_REG_14__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U32590 ( .A1(n2544), .A2(IR_REG_31__SCAN_IN), .ZN(n2547) );
  INV_X1 U32600 ( .A(n2547), .ZN(n2545) );
  NAND2_X1 U32610 ( .A1(n2545), .A2(IR_REG_15__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32620 ( .A1(n2547), .A2(n2546), .ZN(n2560) );
  MUX2_X1 U32630 ( .A(n3896), .B(DATAI_15_), .S(n2363), .Z(n3642) );
  NAND2_X1 U32640 ( .A1(n3642), .A2(n2268), .ZN(n2549) );
  NAND2_X1 U32650 ( .A1(n2550), .A2(n2549), .ZN(n2551) );
  XNOR2_X1 U32660 ( .A(n2551), .B(n2691), .ZN(n2569) );
  NOR2_X1 U32670 ( .A1(n2570), .A2(n2569), .ZN(n3554) );
  NAND2_X1 U32680 ( .A1(n3720), .A2(REG1_REG_16__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U32690 ( .A1(n2780), .A2(REG0_REG_16__SCAN_IN), .ZN(n2558) );
  INV_X1 U32700 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2552) );
  OR2_X1 U32710 ( .A1(n3724), .A2(n2552), .ZN(n2557) );
  AND2_X1 U32720 ( .A1(n2554), .A2(n2553), .ZN(n2555) );
  OR2_X1 U32730 ( .A1(n2555), .A2(n2577), .ZN(n4151) );
  OR2_X1 U32740 ( .A1(n2786), .A2(n4151), .ZN(n2556) );
  NAND4_X1 U32750 ( .A1(n2559), .A2(n2558), .A3(n2557), .A4(n2556), .ZN(n4126)
         );
  NAND2_X1 U32760 ( .A1(n4126), .A2(n2731), .ZN(n2564) );
  NAND2_X1 U32770 ( .A1(n2560), .A2(IR_REG_31__SCAN_IN), .ZN(n2562) );
  XNOR2_X1 U32780 ( .A(n2562), .B(n2561), .ZN(n4649) );
  INV_X1 U32790 ( .A(DATAI_16_), .ZN(n4648) );
  MUX2_X1 U32800 ( .A(n4649), .B(n4648), .S(n2363), .Z(n4153) );
  OR2_X1 U32810 ( .A1(n4153), .A2(n2031), .ZN(n2563) );
  NAND2_X1 U32820 ( .A1(n2564), .A2(n2563), .ZN(n2565) );
  XNOR2_X1 U32830 ( .A(n2565), .B(n2691), .ZN(n2568) );
  NOR2_X1 U32840 ( .A1(n4153), .A2(n2773), .ZN(n2566) );
  AOI21_X1 U32850 ( .B1(n4126), .B2(n2324), .A(n2566), .ZN(n2567) );
  NAND2_X1 U32860 ( .A1(n2568), .A2(n2567), .ZN(n2573) );
  NOR2_X2 U32870 ( .A1(n3554), .A2(n3557), .ZN(n2576) );
  NAND2_X1 U32880 ( .A1(n2570), .A2(n2569), .ZN(n3555) );
  NAND2_X1 U32890 ( .A1(n4324), .A2(n2324), .ZN(n2572) );
  NAND2_X1 U32900 ( .A1(n3642), .A2(n2675), .ZN(n2571) );
  NAND2_X1 U32910 ( .A1(n2572), .A2(n2571), .ZN(n3639) );
  NAND2_X1 U32920 ( .A1(n3555), .A2(n3639), .ZN(n2575) );
  INV_X1 U32930 ( .A(n2573), .ZN(n2574) );
  NAND2_X1 U32940 ( .A1(n3720), .A2(REG1_REG_17__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U32950 ( .A1(n2780), .A2(REG0_REG_17__SCAN_IN), .ZN(n2582) );
  OR2_X1 U32960 ( .A1(n2577), .A2(REG3_REG_17__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U32970 ( .A1(n2593), .A2(n2578), .ZN(n3569) );
  OR2_X1 U32980 ( .A1(n2786), .A2(n3569), .ZN(n2581) );
  INV_X1 U32990 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2579) );
  OR2_X1 U33000 ( .A1(n3724), .A2(n2579), .ZN(n2580) );
  NAND4_X1 U33010 ( .A1(n2583), .A2(n2582), .A3(n2581), .A4(n2580), .ZN(n4145)
         );
  NAND2_X1 U33020 ( .A1(n4145), .A2(n2731), .ZN(n2588) );
  OR2_X1 U33030 ( .A1(n2584), .A2(n2775), .ZN(n2585) );
  XNOR2_X1 U33040 ( .A(n2585), .B(IR_REG_17__SCAN_IN), .ZN(n3899) );
  INV_X1 U33050 ( .A(DATAI_17_), .ZN(n2586) );
  MUX2_X1 U33060 ( .A(n4647), .B(n2586), .S(n3725), .Z(n4132) );
  OR2_X1 U33070 ( .A1(n4132), .A2(n2031), .ZN(n2587) );
  NAND2_X1 U33080 ( .A1(n2588), .A2(n2587), .ZN(n2589) );
  XNOR2_X1 U33090 ( .A(n2589), .B(n2691), .ZN(n2592) );
  NOR2_X1 U33100 ( .A1(n4132), .A2(n2773), .ZN(n2590) );
  AOI21_X1 U33110 ( .B1(n4145), .B2(n2324), .A(n2590), .ZN(n2591) );
  NOR2_X1 U33120 ( .A1(n2592), .A2(n2591), .ZN(n3567) );
  NAND2_X1 U33130 ( .A1(n2592), .A2(n2591), .ZN(n3566) );
  NAND2_X1 U33140 ( .A1(n3720), .A2(REG1_REG_18__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U33150 ( .A1(n2780), .A2(REG0_REG_18__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U33160 ( .A1(n2593), .A2(n4276), .ZN(n2594) );
  NAND2_X1 U33170 ( .A1(n2604), .A2(n2594), .ZN(n4106) );
  OR2_X1 U33180 ( .A1(n2786), .A2(n4106), .ZN(n2596) );
  INV_X1 U33190 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4107) );
  OR2_X1 U33200 ( .A1(n3724), .A2(n4107), .ZN(n2595) );
  NAND4_X1 U33210 ( .A1(n2598), .A2(n2597), .A3(n2596), .A4(n2595), .ZN(n4125)
         );
  NAND2_X1 U33220 ( .A1(n2599), .A2(IR_REG_31__SCAN_IN), .ZN(n2600) );
  XNOR2_X1 U33230 ( .A(n2600), .B(IR_REG_18__SCAN_IN), .ZN(n4620) );
  INV_X1 U33240 ( .A(DATAI_18_), .ZN(n2601) );
  MUX2_X1 U33250 ( .A(n4646), .B(n2601), .S(n2363), .Z(n4113) );
  AOI22_X1 U33260 ( .A1(n4125), .A2(n2731), .B1(n2268), .B2(n3620), .ZN(n2602)
         );
  NAND2_X1 U33270 ( .A1(n3720), .A2(REG1_REG_19__SCAN_IN), .ZN(n2609) );
  NAND2_X1 U33280 ( .A1(n2780), .A2(REG0_REG_19__SCAN_IN), .ZN(n2608) );
  OR2_X1 U33290 ( .A1(n3724), .A2(n3900), .ZN(n2607) );
  NAND2_X1 U33300 ( .A1(n2604), .A2(n2603), .ZN(n2605) );
  NAND2_X1 U33310 ( .A1(n2619), .A2(n2605), .ZN(n4094) );
  OR2_X1 U33320 ( .A1(n2786), .A2(n4094), .ZN(n2606) );
  NAND4_X1 U33330 ( .A1(n2609), .A2(n2608), .A3(n2607), .A4(n2606), .ZN(n4110)
         );
  NAND2_X1 U33340 ( .A1(n4110), .A2(n2731), .ZN(n2611) );
  MUX2_X1 U33350 ( .A(n4314), .B(DATAI_19_), .S(n2363), .Z(n3526) );
  NAND2_X1 U33360 ( .A1(n3526), .A2(n2268), .ZN(n2610) );
  NAND2_X1 U33370 ( .A1(n2611), .A2(n2610), .ZN(n2612) );
  XNOR2_X1 U33380 ( .A(n2612), .B(n2735), .ZN(n2616) );
  NAND2_X1 U33390 ( .A1(n4110), .A2(n2324), .ZN(n2614) );
  NAND2_X1 U33400 ( .A1(n3526), .A2(n2675), .ZN(n2613) );
  NAND2_X1 U33410 ( .A1(n2614), .A2(n2613), .ZN(n2615) );
  NOR2_X1 U33420 ( .A1(n2616), .A2(n2615), .ZN(n2617) );
  AOI21_X1 U33430 ( .B1(n2616), .B2(n2615), .A(n2617), .ZN(n3522) );
  NAND2_X1 U33440 ( .A1(n3519), .A2(n3522), .ZN(n3521) );
  INV_X1 U33450 ( .A(n2617), .ZN(n2618) );
  NAND2_X1 U33460 ( .A1(n3720), .A2(REG1_REG_20__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U33470 ( .A1(n2780), .A2(REG0_REG_20__SCAN_IN), .ZN(n2624) );
  INV_X1 U33480 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4071) );
  OR2_X1 U33490 ( .A1(n3724), .A2(n4071), .ZN(n2623) );
  INV_X1 U33500 ( .A(n2643), .ZN(n2621) );
  NAND2_X1 U33510 ( .A1(n2619), .A2(n4211), .ZN(n2620) );
  NAND2_X1 U33520 ( .A1(n2621), .A2(n2620), .ZN(n4070) );
  OR2_X1 U3353 ( .A1(n2786), .A2(n4070), .ZN(n2622) );
  NAND4_X1 U33540 ( .A1(n2625), .A2(n2624), .A3(n2623), .A4(n2622), .ZN(n3826)
         );
  NAND2_X1 U3355 ( .A1(n3826), .A2(n2731), .ZN(n2627) );
  OR2_X1 U3356 ( .A1(n4069), .A2(n2031), .ZN(n2626) );
  NAND2_X1 U3357 ( .A1(n2627), .A2(n2626), .ZN(n2628) );
  XNOR2_X1 U3358 ( .A(n2628), .B(n2691), .ZN(n2636) );
  NOR2_X1 U3359 ( .A1(n2773), .A2(n4069), .ZN(n2629) );
  AOI21_X1 U3360 ( .B1(n3826), .B2(n2324), .A(n2629), .ZN(n2635) );
  NAND2_X1 U3361 ( .A1(n3529), .A2(n3593), .ZN(n3590) );
  NAND2_X1 U3362 ( .A1(n3720), .A2(REG1_REG_21__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3363 ( .A1(n2780), .A2(REG0_REG_21__SCAN_IN), .ZN(n2632) );
  XNOR2_X1 U3364 ( .A(n2643), .B(REG3_REG_21__SCAN_IN), .ZN(n4050) );
  OR2_X1 U3365 ( .A1(n2786), .A2(n4050), .ZN(n2631) );
  INV_X1 U3366 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4051) );
  OR2_X1 U3367 ( .A1(n3724), .A2(n4051), .ZN(n2630) );
  INV_X1 U3368 ( .A(n4045), .ZN(n4049) );
  OAI22_X1 U3369 ( .A1(n4063), .A2(n2773), .B1(n2031), .B2(n4049), .ZN(n2634)
         );
  XNOR2_X1 U3370 ( .A(n2634), .B(n2735), .ZN(n2638) );
  OAI22_X1 U3371 ( .A1(n4063), .A2(n2719), .B1(n2773), .B2(n4049), .ZN(n2637)
         );
  NOR2_X1 U3372 ( .A1(n2638), .A2(n2637), .ZN(n3531) );
  NOR2_X1 U3373 ( .A1(n3531), .A2(n3591), .ZN(n2639) );
  AND2_X1 U3374 ( .A1(n2638), .A2(n2637), .ZN(n3530) );
  AOI21_X2 U3375 ( .B1(n3590), .B2(n2639), .A(n3530), .ZN(n3601) );
  NAND2_X1 U3376 ( .A1(n3720), .A2(REG1_REG_22__SCAN_IN), .ZN(n2649) );
  NAND2_X1 U3377 ( .A1(n2780), .A2(REG0_REG_22__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U3378 ( .A1(n2643), .A2(REG3_REG_21__SCAN_IN), .ZN(n2641) );
  INV_X1 U3379 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U3380 ( .A1(n2641), .A2(n2640), .ZN(n2644) );
  AND2_X1 U3381 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2642) );
  NAND2_X1 U3382 ( .A1(n2644), .A2(n2651), .ZN(n4025) );
  OR2_X1 U3383 ( .A1(n2786), .A2(n4025), .ZN(n2647) );
  INV_X1 U3384 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2645) );
  OR2_X1 U3385 ( .A1(n3724), .A2(n2645), .ZN(n2646) );
  INV_X1 U3386 ( .A(n4033), .ZN(n2843) );
  OAI22_X1 U3387 ( .A1(n2842), .A2(n2719), .B1(n2773), .B2(n2843), .ZN(n2663)
         );
  OAI22_X1 U3388 ( .A1(n2842), .A2(n2773), .B1(n2031), .B2(n2843), .ZN(n2650)
         );
  XNOR2_X1 U3389 ( .A(n2650), .B(n2735), .ZN(n2662) );
  XOR2_X1 U3390 ( .A(n2663), .B(n2662), .Z(n3603) );
  NAND2_X1 U3391 ( .A1(n3601), .A2(n3603), .ZN(n3507) );
  NAND2_X1 U3392 ( .A1(n2651), .A2(n3512), .ZN(n2652) );
  NAND2_X1 U3393 ( .A1(n2670), .A2(n2652), .ZN(n4015) );
  INV_X1 U3394 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4016) );
  OAI22_X1 U3395 ( .A1(n4015), .A2(n2786), .B1(n3724), .B2(n4016), .ZN(n2656)
         );
  NAND2_X1 U3396 ( .A1(n3720), .A2(REG1_REG_23__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3397 ( .A1(n2780), .A2(REG0_REG_23__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U3398 ( .A1(n2654), .A2(n2653), .ZN(n2655) );
  NAND2_X1 U3399 ( .A1(n4034), .A2(n2657), .ZN(n2659) );
  NAND2_X1 U3400 ( .A1(n3515), .A2(n2268), .ZN(n2658) );
  NAND2_X1 U3401 ( .A1(n2659), .A2(n2658), .ZN(n2660) );
  XNOR2_X1 U3402 ( .A(n2660), .B(n2735), .ZN(n2667) );
  AND2_X1 U3403 ( .A1(n2731), .A2(n3515), .ZN(n2661) );
  AOI21_X1 U3404 ( .B1(n4034), .B2(n2324), .A(n2661), .ZN(n2668) );
  XNOR2_X1 U3405 ( .A(n2667), .B(n2668), .ZN(n3508) );
  INV_X1 U3406 ( .A(n2662), .ZN(n2665) );
  INV_X1 U3407 ( .A(n2663), .ZN(n2664) );
  NAND2_X1 U3408 ( .A1(n2665), .A2(n2664), .ZN(n3509) );
  INV_X1 U3409 ( .A(n2667), .ZN(n2669) );
  NOR2_X1 U3410 ( .A1(n2669), .A2(n2668), .ZN(n2679) );
  INV_X1 U3411 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4435) );
  INV_X1 U3412 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3580) );
  AND2_X1 U3413 ( .A1(n2670), .A2(n3580), .ZN(n2671) );
  NOR2_X1 U3414 ( .A1(n2684), .A2(n2671), .ZN(n3993) );
  NAND2_X1 U3415 ( .A1(n3993), .A2(n2223), .ZN(n2673) );
  AOI22_X1 U3416 ( .A1(n2221), .A2(REG2_REG_24__SCAN_IN), .B1(n3720), .B2(
        REG1_REG_24__SCAN_IN), .ZN(n2672) );
  OAI211_X1 U3417 ( .C1(n2674), .C2(n4435), .A(n2673), .B(n2672), .ZN(n3546)
         );
  NAND2_X1 U3418 ( .A1(n3546), .A2(n2324), .ZN(n2677) );
  INV_X1 U3419 ( .A(n3992), .ZN(n3582) );
  NAND2_X1 U3420 ( .A1(n2675), .A2(n3582), .ZN(n2676) );
  NAND2_X1 U3421 ( .A1(n2677), .A2(n2676), .ZN(n2678) );
  INV_X1 U3422 ( .A(n2679), .ZN(n2680) );
  OAI22_X1 U3423 ( .A1(n4008), .A2(n2773), .B1(n2031), .B2(n3992), .ZN(n2682)
         );
  XOR2_X1 U3424 ( .A(n2735), .B(n2682), .Z(n3579) );
  NOR2_X1 U3425 ( .A1(n2684), .A2(REG3_REG_25__SCAN_IN), .ZN(n2685) );
  OR2_X1 U3426 ( .A1(n2712), .A2(n2685), .ZN(n3544) );
  AOI22_X1 U3427 ( .A1(n3720), .A2(REG1_REG_25__SCAN_IN), .B1(n2780), .B2(
        REG0_REG_25__SCAN_IN), .ZN(n2688) );
  INV_X1 U3428 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2686) );
  OR2_X1 U3429 ( .A1(n3724), .A2(n2686), .ZN(n2687) );
  OAI211_X1 U3430 ( .C1(n3544), .C2(n2786), .A(n2688), .B(n2687), .ZN(n3988)
         );
  NAND2_X1 U3431 ( .A1(n3988), .A2(n2731), .ZN(n2690) );
  OR2_X1 U3432 ( .A1(n3974), .A2(n2031), .ZN(n2689) );
  NAND2_X1 U3433 ( .A1(n2690), .A2(n2689), .ZN(n2692) );
  XNOR2_X1 U3434 ( .A(n2692), .B(n2691), .ZN(n2695) );
  NOR2_X1 U3435 ( .A1(n2773), .A2(n3974), .ZN(n2693) );
  AOI21_X1 U3436 ( .B1(n3988), .B2(n2324), .A(n2693), .ZN(n2694) );
  NAND2_X1 U3437 ( .A1(n2695), .A2(n2694), .ZN(n3541) );
  INV_X1 U3438 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2696) );
  XNOR2_X1 U3439 ( .A(n2712), .B(n2696), .ZN(n3959) );
  NAND2_X1 U3440 ( .A1(n3959), .A2(n2223), .ZN(n2702) );
  INV_X1 U3441 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2699) );
  NAND2_X1 U3442 ( .A1(n3720), .A2(REG1_REG_26__SCAN_IN), .ZN(n2698) );
  NAND2_X1 U3443 ( .A1(n2780), .A2(REG0_REG_26__SCAN_IN), .ZN(n2697) );
  OAI211_X1 U3444 ( .C1(n2699), .C2(n3724), .A(n2698), .B(n2697), .ZN(n2700)
         );
  INV_X1 U3445 ( .A(n2700), .ZN(n2701) );
  NOR2_X1 U3446 ( .A1(n3957), .A2(n2031), .ZN(n2703) );
  AOI21_X1 U3447 ( .B1(n3970), .B2(n2731), .A(n2703), .ZN(n2704) );
  XNOR2_X1 U3448 ( .A(n2704), .B(n2735), .ZN(n2707) );
  NOR2_X1 U3449 ( .A1(n2773), .A2(n3957), .ZN(n2705) );
  AOI21_X1 U3450 ( .B1(n3970), .B2(n2324), .A(n2705), .ZN(n2706) );
  OR2_X1 U3451 ( .A1(n2707), .A2(n2706), .ZN(n3625) );
  NAND2_X1 U3452 ( .A1(n3623), .A2(n3625), .ZN(n2708) );
  NAND2_X1 U3453 ( .A1(n2707), .A2(n2706), .ZN(n3624) );
  INV_X1 U3454 ( .A(n3481), .ZN(n2722) );
  NAND2_X1 U3455 ( .A1(n2712), .A2(REG3_REG_26__SCAN_IN), .ZN(n2710) );
  INV_X1 U3456 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2709) );
  NAND2_X1 U3457 ( .A1(n2710), .A2(n2709), .ZN(n2713) );
  AND2_X1 U34580 ( .A1(REG3_REG_26__SCAN_IN), .A2(REG3_REG_27__SCAN_IN), .ZN(
        n2711) );
  NAND2_X1 U34590 ( .A1(n2712), .A2(n2711), .ZN(n2723) );
  NAND2_X1 U3460 ( .A1(n2713), .A2(n2723), .ZN(n3937) );
  INV_X1 U3461 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3936) );
  NAND2_X1 U3462 ( .A1(n3720), .A2(REG1_REG_27__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U3463 ( .A1(n2780), .A2(REG0_REG_27__SCAN_IN), .ZN(n2714) );
  OAI211_X1 U3464 ( .C1(n3936), .C2(n3724), .A(n2715), .B(n2714), .ZN(n2716)
         );
  INV_X1 U3465 ( .A(n2716), .ZN(n2717) );
  INV_X1 U3466 ( .A(n3941), .ZN(n2720) );
  OAI22_X1 U34670 ( .A1(n3631), .A2(n2719), .B1(n2720), .B2(n2773), .ZN(n2765)
         );
  OAI22_X1 U3468 ( .A1(n3631), .A2(n2773), .B1(n2720), .B2(n2031), .ZN(n2721)
         );
  XNOR2_X1 U34690 ( .A(n2721), .B(n2735), .ZN(n2766) );
  NAND2_X1 U3470 ( .A1(n2722), .A2(n3480), .ZN(n2802) );
  INV_X1 U34710 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4208) );
  NAND2_X1 U3472 ( .A1(n2723), .A2(n4208), .ZN(n2724) );
  NAND2_X1 U34730 ( .A1(n3491), .A2(n2223), .ZN(n2730) );
  INV_X1 U3474 ( .A(REG2_REG_28__SCAN_IN), .ZN(n2727) );
  NAND2_X1 U34750 ( .A1(n3720), .A2(REG1_REG_28__SCAN_IN), .ZN(n2726) );
  NAND2_X1 U3476 ( .A1(n2780), .A2(REG0_REG_28__SCAN_IN), .ZN(n2725) );
  OAI211_X1 U34770 ( .C1(n2727), .C2(n3724), .A(n2726), .B(n2725), .ZN(n2728)
         );
  INV_X1 U3478 ( .A(n2728), .ZN(n2729) );
  NAND2_X1 U34790 ( .A1(n3942), .A2(n2731), .ZN(n2734) );
  NAND2_X1 U3480 ( .A1(n3725), .A2(DATAI_28_), .ZN(n2898) );
  OR2_X1 U34810 ( .A1(n2898), .A2(n2031), .ZN(n2733) );
  NAND2_X1 U3482 ( .A1(n2734), .A2(n2733), .ZN(n2736) );
  XNOR2_X1 U34830 ( .A(n2736), .B(n2735), .ZN(n2738) );
  INV_X1 U3484 ( .A(n2898), .ZN(n3921) );
  AOI22_X1 U34850 ( .A1(n3942), .A2(n2324), .B1(n2675), .B2(n3921), .ZN(n2737)
         );
  XNOR2_X1 U3486 ( .A(n2738), .B(n2737), .ZN(n2796) );
  INV_X1 U34870 ( .A(n2796), .ZN(n2764) );
  INV_X1 U3488 ( .A(n2936), .ZN(n2955) );
  NAND2_X1 U34890 ( .A1(n2953), .A2(n2955), .ZN(n2739) );
  MUX2_X1 U3490 ( .A(n2953), .B(n2739), .S(B_REG_SCAN_IN), .Z(n2741) );
  OAI22_X1 U34910 ( .A1(n2952), .A2(D_REG_1__SCAN_IN), .B1(n2740), .B2(n2936), 
        .ZN(n2917) );
  NOR4_X1 U3492 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2750) );
  NOR4_X1 U34930 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2749) );
  OR4_X1 U3494 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2747) );
  NOR4_X1 U34950 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2745) );
  NOR4_X1 U3496 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2744) );
  NOR4_X1 U34970 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2743) );
  NOR4_X1 U3498 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2742) );
  NAND4_X1 U34990 ( .A1(n2745), .A2(n2744), .A3(n2743), .A4(n2742), .ZN(n2746)
         );
  NOR4_X1 U3500 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(n2747), 
        .A4(n2746), .ZN(n2748) );
  AND3_X1 U35010 ( .A1(n2750), .A2(n2749), .A3(n2748), .ZN(n2751) );
  NOR2_X1 U3502 ( .A1(n2952), .A2(n2751), .ZN(n2895) );
  NOR2_X1 U35030 ( .A1(n2917), .A2(n2895), .ZN(n2755) );
  INV_X1 U3504 ( .A(n2952), .ZN(n2754) );
  INV_X1 U35050 ( .A(D_REG_0__SCAN_IN), .ZN(n2954) );
  INV_X1 U35060 ( .A(n2740), .ZN(n2752) );
  NAND2_X1 U35070 ( .A1(n2755), .A2(n2902), .ZN(n2788) );
  INV_X1 U35080 ( .A(n4644), .ZN(n2759) );
  INV_X1 U35090 ( .A(n2958), .ZN(n2888) );
  NAND2_X1 U35100 ( .A1(n3086), .A2(n4314), .ZN(n2762) );
  NAND2_X1 U35110 ( .A1(n2888), .A2(n2762), .ZN(n2767) );
  INV_X1 U35120 ( .A(n2266), .ZN(n4472) );
  OR2_X1 U35130 ( .A1(n2767), .A2(n4350), .ZN(n2763) );
  NAND2_X1 U35140 ( .A1(n2764), .A2(n3608), .ZN(n2801) );
  NAND2_X1 U35150 ( .A1(n2766), .A2(n2765), .ZN(n2795) );
  NAND2_X1 U35160 ( .A1(n2802), .A2(n2203), .ZN(n2800) );
  NAND2_X1 U35170 ( .A1(n4148), .A2(n2767), .ZN(n2768) );
  NAND2_X1 U35180 ( .A1(n2788), .A2(n2768), .ZN(n3071) );
  NAND2_X1 U35190 ( .A1(n2266), .A2(n3905), .ZN(n2769) );
  NAND2_X1 U35200 ( .A1(n2958), .A2(n2769), .ZN(n2894) );
  AND3_X1 U35210 ( .A1(n2894), .A2(n2960), .A3(n2256), .ZN(n2770) );
  AOI21_X1 U35220 ( .B1(n3071), .B2(n2770), .A(U3149), .ZN(n2774) );
  OR2_X1 U35230 ( .A1(n2771), .A2(n4644), .ZN(n2772) );
  NOR2_X1 U35240 ( .A1(n2773), .A2(n2772), .ZN(n3815) );
  AND2_X1 U35250 ( .A1(n2788), .A2(n3815), .ZN(n3069) );
  OR2_X1 U35260 ( .A1(n2776), .A2(n2775), .ZN(n2778) );
  NAND2_X1 U35270 ( .A1(n3815), .A2(n3834), .ZN(n2779) );
  INV_X1 U35280 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2783) );
  NAND2_X1 U35290 ( .A1(n2780), .A2(REG0_REG_29__SCAN_IN), .ZN(n2782) );
  NAND2_X1 U35300 ( .A1(n3720), .A2(REG1_REG_29__SCAN_IN), .ZN(n2781) );
  OAI211_X1 U35310 ( .C1(n3724), .C2(n2783), .A(n2782), .B(n2781), .ZN(n2784)
         );
  INV_X1 U35320 ( .A(n2784), .ZN(n2785) );
  OAI21_X1 U35330 ( .B1(n3910), .B2(n2786), .A(n2785), .ZN(n3823) );
  NAND2_X1 U35340 ( .A1(n3815), .A2(n4478), .ZN(n2787) );
  AOI22_X1 U35350 ( .A1(n3823), .A2(n3645), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2794) );
  AND2_X1 U35360 ( .A1(n4314), .A2(n3816), .ZN(n2789) );
  NAND2_X1 U35370 ( .A1(n4676), .A2(n2790), .ZN(n2893) );
  NAND2_X1 U35380 ( .A1(n3643), .A2(n3921), .ZN(n2793) );
  OAI211_X1 U35390 ( .C1(n3631), .C2(n3648), .A(n2794), .B(n2793), .ZN(n2798)
         );
  NOR3_X1 U35400 ( .A1(n2796), .A2(n3653), .A3(n2795), .ZN(n2797) );
  AOI211_X1 U35410 ( .C1(n3491), .C2(n3650), .A(n2798), .B(n2797), .ZN(n2799)
         );
  OAI211_X1 U35420 ( .C1(n2802), .C2(n2801), .A(n2800), .B(n2799), .ZN(U3217)
         );
  NAND2_X1 U35430 ( .A1(n2265), .A2(n2803), .ZN(n3659) );
  NAND2_X1 U35440 ( .A1(n2804), .A2(n2806), .ZN(n2856) );
  AND2_X1 U35450 ( .A1(n2805), .A2(n3124), .ZN(n2909) );
  NAND2_X1 U35460 ( .A1(n2855), .A2(n2909), .ZN(n2908) );
  NAND2_X1 U35470 ( .A1(n3123), .A2(n2806), .ZN(n2807) );
  OR2_X1 U35480 ( .A1(n2809), .A2(n3101), .ZN(n3661) );
  NAND2_X1 U35490 ( .A1(n2809), .A2(n3101), .ZN(n3664) );
  NAND2_X1 U35500 ( .A1(n3104), .A2(n3103), .ZN(n3102) );
  INV_X1 U35510 ( .A(n2323), .ZN(n2808) );
  INV_X1 U35520 ( .A(n3101), .ZN(n3114) );
  OR2_X1 U35530 ( .A1(n2809), .A2(n3114), .ZN(n3127) );
  AND2_X1 U35540 ( .A1(n2810), .A2(n3127), .ZN(n2811) );
  NAND2_X1 U35550 ( .A1(n3102), .A2(n2811), .ZN(n2813) );
  NAND2_X1 U35560 ( .A1(n2323), .A2(n3147), .ZN(n2812) );
  NAND2_X1 U35570 ( .A1(n2813), .A2(n2812), .ZN(n3241) );
  INV_X1 U35580 ( .A(n3253), .ZN(n3191) );
  NAND2_X1 U35590 ( .A1(n3222), .A2(n3191), .ZN(n2814) );
  NAND2_X1 U35600 ( .A1(n3245), .A2(n2814), .ZN(n3216) );
  OR2_X1 U35610 ( .A1(n3832), .A2(n3224), .ZN(n2815) );
  NAND2_X1 U35620 ( .A1(n3216), .A2(n2815), .ZN(n2817) );
  NAND2_X1 U35630 ( .A1(n3832), .A2(n3224), .ZN(n2816) );
  NAND2_X1 U35640 ( .A1(n2817), .A2(n2816), .ZN(n3182) );
  AND2_X1 U35650 ( .A1(n3831), .A2(n3184), .ZN(n2820) );
  NAND2_X1 U35660 ( .A1(n2818), .A2(n3176), .ZN(n2819) );
  NAND2_X1 U35670 ( .A1(n3830), .A2(n3305), .ZN(n3685) );
  INV_X1 U35680 ( .A(n3305), .ZN(n3233) );
  NAND2_X1 U35690 ( .A1(n3830), .A2(n3233), .ZN(n3291) );
  NAND2_X1 U35700 ( .A1(n3272), .A2(n3267), .ZN(n2822) );
  AND2_X1 U35710 ( .A1(n3291), .A2(n2822), .ZN(n2823) );
  AND2_X1 U35720 ( .A1(n2048), .A2(n3278), .ZN(n2824) );
  NOR2_X1 U35730 ( .A1(n3828), .A2(n3354), .ZN(n2826) );
  NAND2_X1 U35740 ( .A1(n3828), .A2(n3354), .ZN(n2825) );
  OR2_X1 U35750 ( .A1(n3396), .A2(n3451), .ZN(n3358) );
  NAND2_X1 U35760 ( .A1(n3396), .A2(n3451), .ZN(n3698) );
  INV_X1 U35770 ( .A(n3451), .ZN(n3375) );
  OR2_X1 U35780 ( .A1(n3396), .A2(n3375), .ZN(n2827) );
  INV_X1 U35790 ( .A(n3500), .ZN(n4328) );
  OR2_X1 U35800 ( .A1(n3641), .A2(n4308), .ZN(n3702) );
  NAND2_X1 U35810 ( .A1(n3641), .A2(n4308), .ZN(n3681) );
  NAND2_X1 U3582 ( .A1(n3702), .A2(n3681), .ZN(n4311) );
  NAND2_X1 U3583 ( .A1(n4312), .A2(n4311), .ZN(n4310) );
  NAND2_X1 U3584 ( .A1(n4324), .A2(n3642), .ZN(n2834) );
  INV_X1 U3585 ( .A(n4324), .ZN(n3559) );
  INV_X1 U3586 ( .A(n3642), .ZN(n3434) );
  OR2_X1 U3587 ( .A1(n4126), .A2(n4153), .ZN(n3786) );
  NAND2_X1 U3588 ( .A1(n4126), .A2(n4153), .ZN(n3783) );
  NAND2_X1 U3589 ( .A1(n3786), .A2(n3783), .ZN(n4142) );
  INV_X1 U3590 ( .A(n4126), .ZN(n3572) );
  INV_X1 U3591 ( .A(n4145), .ZN(n2836) );
  OR2_X1 U3592 ( .A1(n4125), .A2(n4113), .ZN(n4081) );
  NAND2_X1 U3593 ( .A1(n4125), .A2(n4113), .ZN(n4082) );
  NAND2_X1 U3594 ( .A1(n4081), .A2(n4082), .ZN(n4100) );
  NAND2_X1 U3595 ( .A1(n4101), .A2(n4100), .ZN(n4099) );
  NAND2_X1 U3596 ( .A1(n4110), .A2(n3526), .ZN(n2840) );
  INV_X1 U3597 ( .A(n4110), .ZN(n3616) );
  INV_X1 U3598 ( .A(n4063), .ZN(n3824) );
  NAND2_X1 U3599 ( .A1(n3824), .A2(n4045), .ZN(n2841) );
  NAND2_X1 U3600 ( .A1(n2842), .A2(n4033), .ZN(n4005) );
  NAND2_X1 U3601 ( .A1(n4046), .A2(n2843), .ZN(n2880) );
  NAND2_X1 U3602 ( .A1(n4005), .A2(n2880), .ZN(n4022) );
  NAND2_X1 U3603 ( .A1(n4023), .A2(n4022), .ZN(n4021) );
  NAND2_X1 U3604 ( .A1(n4046), .A2(n4033), .ZN(n2844) );
  NAND2_X1 U3605 ( .A1(n4021), .A2(n2844), .ZN(n3998) );
  NAND2_X1 U3606 ( .A1(n3998), .A2(n2202), .ZN(n2846) );
  NAND2_X1 U3607 ( .A1(n4034), .A2(n3515), .ZN(n2845) );
  OR2_X1 U3608 ( .A1(n3988), .A2(n3545), .ZN(n2847) );
  NAND2_X1 U3609 ( .A1(n4008), .A2(n3992), .ZN(n3964) );
  AND2_X1 U3610 ( .A1(n2847), .A2(n3964), .ZN(n2848) );
  NAND2_X1 U3611 ( .A1(n3970), .A2(n3951), .ZN(n3735) );
  NAND2_X1 U3612 ( .A1(n3948), .A2(n3735), .ZN(n2849) );
  NOR2_X1 U3613 ( .A1(n3952), .A2(n3941), .ZN(n2851) );
  NAND2_X1 U3614 ( .A1(n3952), .A2(n3941), .ZN(n2850) );
  NOR2_X1 U3615 ( .A1(n3942), .A2(n2898), .ZN(n3911) );
  NAND2_X1 U3616 ( .A1(n3942), .A2(n2898), .ZN(n3912) );
  INV_X1 U3617 ( .A(n3912), .ZN(n2852) );
  XNOR2_X1 U3618 ( .A(n2853), .B(n2932), .ZN(n2854) );
  NAND2_X1 U3619 ( .A1(n2854), .A2(n3905), .ZN(n4067) );
  INV_X1 U3620 ( .A(n4676), .ZN(n4700) );
  INV_X1 U3621 ( .A(n3103), .ZN(n3770) );
  NAND2_X1 U3622 ( .A1(n3105), .A2(n3661), .ZN(n3130) );
  INV_X1 U3623 ( .A(n3147), .ZN(n3133) );
  OR2_X1 U3624 ( .A1(n2323), .A2(n3133), .ZN(n3666) );
  NAND2_X1 U3625 ( .A1(n2323), .A2(n3133), .ZN(n3663) );
  NAND2_X1 U3626 ( .A1(n3130), .A2(n3771), .ZN(n2857) );
  INV_X1 U3627 ( .A(n3667), .ZN(n2858) );
  NAND2_X1 U3628 ( .A1(n2859), .A2(n3672), .ZN(n3218) );
  INV_X1 U3629 ( .A(n3224), .ZN(n3217) );
  AND2_X1 U3630 ( .A1(n3832), .A2(n3217), .ZN(n3215) );
  OR2_X1 U3631 ( .A1(n3832), .A2(n3217), .ZN(n3686) );
  INV_X1 U3632 ( .A(n3184), .ZN(n3176) );
  NAND2_X1 U3633 ( .A1(n3831), .A2(n3176), .ZN(n3669) );
  NOR2_X1 U3634 ( .A1(n3831), .A2(n3176), .ZN(n3673) );
  NAND2_X1 U3635 ( .A1(n3301), .A2(n3675), .ZN(n2861) );
  NAND2_X1 U3636 ( .A1(n2861), .A2(n3685), .ZN(n3286) );
  OR2_X1 U3637 ( .A1(n3272), .A2(n3294), .ZN(n3679) );
  NAND2_X1 U3638 ( .A1(n3286), .A2(n3679), .ZN(n2862) );
  NAND2_X1 U3639 ( .A1(n3272), .A2(n3294), .ZN(n3689) );
  NAND2_X1 U3640 ( .A1(n2862), .A2(n3689), .ZN(n3271) );
  INV_X1 U3641 ( .A(n3324), .ZN(n3275) );
  AND2_X1 U3642 ( .A1(n3829), .A2(n3275), .ZN(n3683) );
  OR2_X1 U3643 ( .A1(n3829), .A2(n3275), .ZN(n3678) );
  INV_X1 U3644 ( .A(n3354), .ZN(n3340) );
  NAND2_X1 U3645 ( .A1(n3828), .A2(n3340), .ZN(n3697) );
  NAND2_X1 U3646 ( .A1(n3333), .A2(n3697), .ZN(n2864) );
  OR2_X1 U3647 ( .A1(n3828), .A2(n3340), .ZN(n3692) );
  NAND2_X1 U3648 ( .A1(n3444), .A2(n3698), .ZN(n3359) );
  NAND2_X1 U3649 ( .A1(n3827), .A2(n3366), .ZN(n3412) );
  NAND2_X1 U3650 ( .A1(n3500), .A2(n3421), .ZN(n2865) );
  NAND2_X1 U3651 ( .A1(n3412), .A2(n2865), .ZN(n2866) );
  INV_X1 U3652 ( .A(n2866), .ZN(n3699) );
  OR2_X1 U3653 ( .A1(n3827), .A2(n3366), .ZN(n3411) );
  NAND2_X1 U3654 ( .A1(n3358), .A2(n3411), .ZN(n2868) );
  NOR2_X1 U3655 ( .A1(n3500), .A2(n3421), .ZN(n2867) );
  AOI21_X1 U3656 ( .B1(n3699), .B2(n2868), .A(n2867), .ZN(n3700) );
  INV_X1 U3657 ( .A(n4311), .ZN(n4319) );
  OR2_X1 U3658 ( .A1(n4324), .A2(n3434), .ZN(n3701) );
  NAND2_X1 U3659 ( .A1(n4324), .A2(n3434), .ZN(n3682) );
  NAND2_X1 U3660 ( .A1(n3701), .A2(n3682), .ZN(n3760) );
  INV_X1 U3661 ( .A(n3702), .ZN(n2870) );
  NOR2_X1 U3662 ( .A1(n3760), .A2(n2870), .ZN(n2871) );
  NAND2_X1 U3663 ( .A1(n4317), .A2(n2871), .ZN(n2872) );
  NAND2_X1 U3664 ( .A1(n2872), .A2(n3682), .ZN(n4143) );
  INV_X1 U3665 ( .A(n4142), .ZN(n3763) );
  NAND2_X1 U3666 ( .A1(n4143), .A2(n3763), .ZN(n2873) );
  NAND2_X1 U3667 ( .A1(n4145), .A2(n4132), .ZN(n3999) );
  AND2_X1 U3668 ( .A1(n3826), .A2(n4069), .ZN(n4003) );
  INV_X1 U3669 ( .A(n4003), .ZN(n2874) );
  NAND2_X1 U3670 ( .A1(n3999), .A2(n2874), .ZN(n2875) );
  NAND2_X1 U3671 ( .A1(n4110), .A2(n4093), .ZN(n3754) );
  AND2_X1 U3672 ( .A1(n4082), .A2(n3754), .ZN(n2877) );
  INV_X1 U3673 ( .A(n2877), .ZN(n4000) );
  OR2_X1 U3674 ( .A1(n2875), .A2(n4000), .ZN(n3784) );
  OR2_X1 U3675 ( .A1(n4145), .A2(n4132), .ZN(n4079) );
  NAND2_X1 U3676 ( .A1(n4081), .A2(n4079), .ZN(n2876) );
  NAND2_X1 U3677 ( .A1(n2877), .A2(n2876), .ZN(n2878) );
  OR2_X1 U3678 ( .A1(n4110), .A2(n4093), .ZN(n3755) );
  AND2_X1 U3679 ( .A1(n2878), .A2(n3755), .ZN(n4057) );
  INV_X1 U3680 ( .A(n4069), .ZN(n4061) );
  NAND2_X1 U3681 ( .A1(n4087), .A2(n4061), .ZN(n2879) );
  AOI21_X1 U3682 ( .B1(n4057), .B2(n2879), .A(n4003), .ZN(n4001) );
  NAND2_X1 U3683 ( .A1(n4063), .A2(n4045), .ZN(n4004) );
  NAND2_X1 U3684 ( .A1(n4004), .A2(n4005), .ZN(n3715) );
  NOR2_X1 U3685 ( .A1(n4001), .A2(n3715), .ZN(n3788) );
  INV_X1 U3686 ( .A(n4034), .ZN(n3986) );
  NOR2_X1 U3687 ( .A1(n3986), .A2(n3515), .ZN(n3751) );
  INV_X1 U3688 ( .A(n2880), .ZN(n2881) );
  NOR2_X1 U3689 ( .A1(n3751), .A2(n2881), .ZN(n3712) );
  NOR2_X1 U3690 ( .A1(n4063), .A2(n4045), .ZN(n3749) );
  NAND2_X1 U3691 ( .A1(n3749), .A2(n4005), .ZN(n3793) );
  OR2_X1 U3692 ( .A1(n3546), .A2(n3992), .ZN(n3752) );
  NAND2_X1 U3693 ( .A1(n3986), .A2(n3515), .ZN(n3750) );
  NAND2_X1 U3694 ( .A1(n3752), .A2(n3750), .ZN(n3791) );
  NAND2_X1 U3695 ( .A1(n3546), .A2(n3992), .ZN(n3753) );
  NAND2_X1 U3696 ( .A1(n3988), .A2(n3974), .ZN(n3743) );
  INV_X1 U3697 ( .A(n3743), .ZN(n2883) );
  OR2_X1 U3698 ( .A1(n3988), .A2(n3974), .ZN(n3742) );
  NOR2_X1 U3699 ( .A1(n3970), .A2(n3957), .ZN(n3656) );
  AND2_X1 U3700 ( .A1(n3970), .A2(n3957), .ZN(n3716) );
  INV_X1 U3701 ( .A(n3716), .ZN(n2884) );
  NOR2_X1 U3702 ( .A1(n3631), .A2(n3941), .ZN(n3718) );
  INV_X1 U3703 ( .A(n3800), .ZN(n2885) );
  XNOR2_X1 U3704 ( .A(n3913), .B(n3924), .ZN(n2891) );
  NAND2_X1 U3705 ( .A1(n4472), .A2(n2267), .ZN(n2887) );
  NAND2_X1 U3706 ( .A1(n4314), .A2(n2932), .ZN(n2886) );
  NAND2_X1 U3707 ( .A1(n2958), .A2(n4478), .ZN(n4086) );
  AOI22_X1 U3708 ( .A1(n3823), .A2(n4323), .B1(n4350), .B2(n3921), .ZN(n2890)
         );
  NAND2_X1 U3709 ( .A1(n3952), .A2(n4144), .ZN(n2889) );
  OAI211_X1 U3710 ( .C1(n2891), .C2(n4129), .A(n2890), .B(n2889), .ZN(n3495)
         );
  INV_X1 U3711 ( .A(n3495), .ZN(n2892) );
  NAND2_X1 U3712 ( .A1(n2917), .A2(n2893), .ZN(n2896) );
  NAND2_X1 U3713 ( .A1(n2894), .A2(n2961), .ZN(n3068) );
  MUX2_X1 U3714 ( .A(REG1_REG_28__SCAN_IN), .B(n2904), .S(n4718), .Z(n2897) );
  INV_X1 U3715 ( .A(n2897), .ZN(n2901) );
  NAND2_X1 U3716 ( .A1(n2803), .A2(n3088), .ZN(n3113) );
  NAND2_X1 U3717 ( .A1(n3254), .A2(n3253), .ZN(n3252) );
  OAI21_X1 U3718 ( .B1(n3935), .B2(n2898), .A(n3929), .ZN(n3493) );
  NAND2_X1 U3719 ( .A1(n2901), .A2(n2900), .ZN(U3546) );
  INV_X1 U3720 ( .A(n2902), .ZN(n2919) );
  MUX2_X1 U3721 ( .A(REG0_REG_28__SCAN_IN), .B(n2904), .S(n4706), .Z(n2905) );
  INV_X1 U3722 ( .A(n2905), .ZN(n2907) );
  NAND2_X1 U3723 ( .A1(n2907), .A2(n2906), .ZN(U3514) );
  OAI21_X1 U3724 ( .B1(n2855), .B2(n2909), .A(n2908), .ZN(n3078) );
  NAND2_X1 U3725 ( .A1(n2805), .A2(n4144), .ZN(n2911) );
  NAND2_X1 U3726 ( .A1(n2809), .A2(n4323), .ZN(n2910) );
  OAI211_X1 U3727 ( .C1(n2803), .C2(n4148), .A(n2911), .B(n2910), .ZN(n2912)
         );
  INV_X1 U3728 ( .A(n2912), .ZN(n2915) );
  XNOR2_X1 U3729 ( .A(n2855), .B(n3657), .ZN(n2913) );
  NAND2_X1 U3730 ( .A1(n2913), .A2(n4320), .ZN(n2914) );
  OAI211_X1 U3731 ( .C1(n3078), .C2(n4067), .A(n2915), .B(n2914), .ZN(n3080)
         );
  INV_X1 U3732 ( .A(n2916), .ZN(n2920) );
  INV_X1 U3733 ( .A(n2917), .ZN(n2918) );
  NAND3_X1 U3734 ( .A1(n2920), .A2(n2919), .A3(n2918), .ZN(n2921) );
  MUX2_X1 U3735 ( .A(n3080), .B(REG2_REG_1__SCAN_IN), .S(n4485), .Z(n2927) );
  NOR2_X1 U3736 ( .A1(n2922), .A2(n4314), .ZN(n4118) );
  OAI21_X1 U3737 ( .B1(n3088), .B2(n2803), .A(n3113), .ZN(n3077) );
  NOR2_X1 U3738 ( .A1(n4136), .A2(n3077), .ZN(n2926) );
  NOR2_X1 U3739 ( .A1(n2259), .A2(n3905), .ZN(n2923) );
  INV_X1 U3740 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2924) );
  OAI22_X1 U3741 ( .A1(n3078), .A2(n4076), .B1(n2924), .B2(n4332), .ZN(n2925)
         );
  OR3_X1 U3742 ( .A1(n2927), .A2(n2926), .A3(n2925), .ZN(U3289) );
  MUX2_X1 U3743 ( .A(n3844), .B(n2298), .S(U3149), .Z(n2928) );
  INV_X1 U3744 ( .A(n2928), .ZN(U3350) );
  INV_X1 U3745 ( .A(n3031), .ZN(n3038) );
  INV_X1 U3746 ( .A(DATAI_5_), .ZN(n2929) );
  MUX2_X1 U3747 ( .A(n3038), .B(n2929), .S(U3149), .Z(n2930) );
  INV_X1 U3748 ( .A(n2930), .ZN(U3347) );
  MUX2_X1 U3749 ( .A(n3013), .B(n2255), .S(U3149), .Z(n2931) );
  INV_X1 U3750 ( .A(n2931), .ZN(U3351) );
  INV_X1 U3751 ( .A(DATAI_22_), .ZN(n2934) );
  NAND2_X1 U3752 ( .A1(n2932), .A2(STATE_REG_SCAN_IN), .ZN(n2933) );
  OAI21_X1 U3753 ( .B1(STATE_REG_SCAN_IN), .B2(n2934), .A(n2933), .ZN(U3330)
         );
  MUX2_X1 U3754 ( .A(n2527), .B(n3891), .S(STATE_REG_SCAN_IN), .Z(n2935) );
  INV_X1 U3755 ( .A(n2935), .ZN(U3338) );
  INV_X1 U3756 ( .A(DATAI_25_), .ZN(n2938) );
  NAND2_X1 U3757 ( .A1(n2936), .A2(STATE_REG_SCAN_IN), .ZN(n2937) );
  OAI21_X1 U3758 ( .B1(STATE_REG_SCAN_IN), .B2(n2938), .A(n2937), .ZN(U3327)
         );
  NAND3_X1 U3759 ( .A1(n2940), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n2942) );
  INV_X1 U3760 ( .A(DATAI_31_), .ZN(n2941) );
  OAI22_X1 U3761 ( .A1(n2939), .A2(n2942), .B1(STATE_REG_SCAN_IN), .B2(n2941), 
        .ZN(U3321) );
  INV_X1 U3762 ( .A(DATAI_26_), .ZN(n2944) );
  NAND2_X1 U3763 ( .A1(n2740), .A2(STATE_REG_SCAN_IN), .ZN(n2943) );
  OAI21_X1 U3764 ( .B1(STATE_REG_SCAN_IN), .B2(n2944), .A(n2943), .ZN(U3326)
         );
  INV_X1 U3765 ( .A(DATAI_19_), .ZN(n2945) );
  MUX2_X1 U3766 ( .A(n2945), .B(n3905), .S(STATE_REG_SCAN_IN), .Z(n2946) );
  INV_X1 U3767 ( .A(n2946), .ZN(U3333) );
  INV_X1 U3768 ( .A(DATAI_21_), .ZN(n2948) );
  NAND2_X1 U3769 ( .A1(n2267), .A2(STATE_REG_SCAN_IN), .ZN(n2947) );
  OAI21_X1 U3770 ( .B1(STATE_REG_SCAN_IN), .B2(n2948), .A(n2947), .ZN(U3331)
         );
  INV_X1 U3771 ( .A(DATAI_30_), .ZN(n2951) );
  NAND2_X1 U3772 ( .A1(n2949), .A2(STATE_REG_SCAN_IN), .ZN(n2950) );
  OAI21_X1 U3773 ( .B1(STATE_REG_SCAN_IN), .B2(n2951), .A(n2950), .ZN(U3322)
         );
  NOR2_X1 U3774 ( .A1(n2740), .A2(n4644), .ZN(n2956) );
  AOI22_X1 U3775 ( .A1(n4641), .A2(n2954), .B1(n2956), .B2(n2953), .ZN(U3458)
         );
  INV_X1 U3776 ( .A(D_REG_1__SCAN_IN), .ZN(n2957) );
  AOI22_X1 U3777 ( .A1(n4641), .A2(n2957), .B1(n2956), .B2(n2955), .ZN(U3459)
         );
  INV_X1 U3778 ( .A(n4476), .ZN(n2981) );
  NAND2_X1 U3779 ( .A1(n2958), .A2(n2960), .ZN(n2959) );
  OR2_X1 U3780 ( .A1(n2960), .A2(U3149), .ZN(n3821) );
  INV_X1 U3781 ( .A(n3821), .ZN(n3817) );
  OR2_X1 U3782 ( .A1(n2961), .A2(n3817), .ZN(n2977) );
  NAND2_X1 U3783 ( .A1(n2976), .A2(n2977), .ZN(n4491) );
  XNOR2_X1 U3784 ( .A(n2963), .B(IR_REG_27__SCAN_IN), .ZN(n4487) );
  XNOR2_X1 U3785 ( .A(n3013), .B(REG1_REG_1__SCAN_IN), .ZN(n3004) );
  AND2_X1 U3786 ( .A1(n4488), .A2(REG1_REG_0__SCAN_IN), .ZN(n3005) );
  INV_X1 U3787 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2964) );
  NOR2_X1 U3788 ( .A1(n3013), .A2(n2964), .ZN(n2965) );
  AOI21_X1 U3789 ( .B1(n3004), .B2(n3005), .A(n2965), .ZN(n3842) );
  INV_X1 U3790 ( .A(n3842), .ZN(n2966) );
  XNOR2_X1 U3791 ( .A(n3844), .B(REG1_REG_2__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U3792 ( .A1(n2300), .A2(REG1_REG_2__SCAN_IN), .ZN(n2967) );
  XOR2_X1 U3793 ( .A(n2982), .B(REG1_REG_3__SCAN_IN), .Z(n2975) );
  INV_X1 U3794 ( .A(n4487), .ZN(n3833) );
  NOR2_X2 U3795 ( .A1(n4491), .A2(n3837), .ZN(n4609) );
  MUX2_X1 U3796 ( .A(n2968), .B(REG2_REG_2__SCAN_IN), .S(n3844), .Z(n2972) );
  INV_X1 U3797 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2970) );
  AND2_X1 U3798 ( .A1(n4488), .A2(REG2_REG_0__SCAN_IN), .ZN(n2969) );
  OR2_X1 U3799 ( .A1(n3013), .A2(n2970), .ZN(n3845) );
  NAND2_X1 U3800 ( .A1(n3846), .A2(n3845), .ZN(n2971) );
  NAND2_X1 U3801 ( .A1(n2972), .A2(n2971), .ZN(n3849) );
  NAND2_X1 U3802 ( .A1(n2300), .A2(REG2_REG_2__SCAN_IN), .ZN(n2973) );
  NAND2_X1 U3803 ( .A1(n3849), .A2(n2973), .ZN(n2994) );
  XOR2_X1 U3804 ( .A(n2993), .B(REG2_REG_3__SCAN_IN), .Z(n2974) );
  AOI22_X1 U3805 ( .A1(n4607), .A2(n2975), .B1(n4609), .B2(n2974), .ZN(n2980)
         );
  INV_X1 U3806 ( .A(n2976), .ZN(n2978) );
  INV_X1 U3807 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3140) );
  NOR2_X1 U3808 ( .A1(STATE_REG_SCAN_IN), .A2(n3140), .ZN(n3148) );
  AOI21_X1 U3809 ( .B1(n4599), .B2(ADDR_REG_3__SCAN_IN), .A(n3148), .ZN(n2979)
         );
  OAI211_X1 U3810 ( .C1(n2981), .C2(n4612), .A(n2980), .B(n2979), .ZN(U3243)
         );
  NOR2_X1 U3811 ( .A1(n4599), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U3812 ( .A1(n2983), .A2(n4476), .ZN(n2984) );
  NAND2_X1 U3813 ( .A1(n2985), .A2(n2984), .ZN(n2988) );
  INV_X1 U3814 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2987) );
  NAND2_X1 U3815 ( .A1(n2988), .A2(n4497), .ZN(n2989) );
  INV_X1 U3816 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2990) );
  MUX2_X1 U3817 ( .A(REG1_REG_5__SCAN_IN), .B(n2990), .S(n3031), .Z(n2991) );
  AND2_X1 U3818 ( .A1(n3031), .A2(REG1_REG_5__SCAN_IN), .ZN(n2992) );
  XNOR2_X1 U3819 ( .A(n3016), .B(REG1_REG_6__SCAN_IN), .ZN(n3003) );
  NAND2_X1 U3820 ( .A1(n2993), .A2(REG2_REG_3__SCAN_IN), .ZN(n2996) );
  NAND2_X1 U3821 ( .A1(n2994), .A2(n4476), .ZN(n2995) );
  NAND2_X1 U3822 ( .A1(n2996), .A2(n2995), .ZN(n2997) );
  XNOR2_X1 U3823 ( .A(n2997), .B(n4497), .ZN(n4495) );
  MUX2_X1 U3824 ( .A(n3223), .B(REG2_REG_5__SCAN_IN), .S(n3031), .Z(n3035) );
  XNOR2_X1 U3825 ( .A(n3020), .B(n4475), .ZN(n3022) );
  XOR2_X1 U3826 ( .A(REG2_REG_6__SCAN_IN), .B(n3022), .Z(n3001) );
  AND2_X1 U3827 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3169) );
  AOI21_X1 U3828 ( .B1(n4599), .B2(ADDR_REG_6__SCAN_IN), .A(n3169), .ZN(n2998)
         );
  OAI21_X1 U3829 ( .B1(n4612), .B2(n2999), .A(n2998), .ZN(n3000) );
  AOI21_X1 U3830 ( .B1(n4609), .B2(n3001), .A(n3000), .ZN(n3002) );
  OAI21_X1 U3831 ( .B1(n3003), .B2(n4618), .A(n3002), .ZN(U3246) );
  XOR2_X1 U3832 ( .A(n3005), .B(n3004), .Z(n3010) );
  INV_X1 U3833 ( .A(n4609), .ZN(n4613) );
  INV_X1 U3834 ( .A(n3846), .ZN(n3008) );
  AOI21_X1 U3835 ( .B1(n4488), .B2(REG2_REG_0__SCAN_IN), .A(n3006), .ZN(n3007)
         );
  NOR3_X1 U3836 ( .A1(n4613), .A2(n3008), .A3(n3007), .ZN(n3009) );
  AOI21_X1 U3837 ( .B1(n4607), .B2(n3010), .A(n3009), .ZN(n3012) );
  AOI22_X1 U3838 ( .A1(n4599), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3011) );
  OAI211_X1 U3839 ( .C1(n3013), .C2(n4612), .A(n3012), .B(n3011), .ZN(U3241)
         );
  AND2_X1 U3840 ( .A1(n3014), .A2(n4475), .ZN(n3015) );
  INV_X1 U3841 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4711) );
  XNOR2_X1 U3842 ( .A(n4473), .B(n4711), .ZN(n3017) );
  XNOR2_X1 U3843 ( .A(n3855), .B(n3017), .ZN(n3030) );
  NOR2_X1 U3844 ( .A1(STATE_REG_SCAN_IN), .A2(n4251), .ZN(n3234) );
  NOR2_X1 U3845 ( .A1(n4612), .A2(n4473), .ZN(n3018) );
  AOI211_X1 U3846 ( .C1(n4599), .C2(ADDR_REG_7__SCAN_IN), .A(n3234), .B(n3018), 
        .ZN(n3029) );
  MUX2_X1 U3847 ( .A(n3019), .B(REG2_REG_7__SCAN_IN), .S(n4473), .Z(n3027) );
  INV_X1 U3848 ( .A(n3020), .ZN(n3021) );
  AOI22_X1 U3849 ( .A1(n3022), .A2(REG2_REG_6__SCAN_IN), .B1(n4475), .B2(n3021), .ZN(n3023) );
  INV_X1 U3850 ( .A(n3023), .ZN(n3026) );
  MUX2_X1 U3851 ( .A(REG2_REG_7__SCAN_IN), .B(n3019), .S(n4473), .Z(n3024) );
  OAI211_X1 U3852 ( .C1(n3027), .C2(n3026), .A(n3879), .B(n4609), .ZN(n3028)
         );
  OAI211_X1 U3853 ( .C1(n3030), .C2(n4618), .A(n3029), .B(n3028), .ZN(U3247)
         );
  MUX2_X1 U3854 ( .A(n2990), .B(REG1_REG_5__SCAN_IN), .S(n3031), .Z(n3033) );
  AOI211_X1 U3855 ( .C1(n2060), .C2(n3033), .A(n3032), .B(n4618), .ZN(n3041)
         );
  AOI211_X1 U3856 ( .C1(n3036), .C2(n3035), .A(n3034), .B(n4613), .ZN(n3040)
         );
  NAND2_X1 U3857 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3159) );
  NAND2_X1 U3858 ( .A1(n4599), .A2(ADDR_REG_5__SCAN_IN), .ZN(n3037) );
  OAI211_X1 U3859 ( .C1(n4612), .C2(n3038), .A(n3159), .B(n3037), .ZN(n3039)
         );
  OR3_X1 U3860 ( .A1(n3041), .A2(n3040), .A3(n3039), .ZN(U3245) );
  INV_X1 U3861 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n3043) );
  NAND2_X1 U3862 ( .A1(n3222), .A2(U4043), .ZN(n3042) );
  OAI21_X1 U3863 ( .B1(U4043), .B2(n3043), .A(n3042), .ZN(U3554) );
  INV_X1 U3864 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n3045) );
  NAND2_X1 U3865 ( .A1(n3396), .A2(U4043), .ZN(n3044) );
  OAI21_X1 U3866 ( .B1(U4043), .B2(n3045), .A(n3044), .ZN(U3561) );
  INV_X1 U3867 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n3047) );
  NAND2_X1 U3868 ( .A1(n3272), .A2(U4043), .ZN(n3046) );
  OAI21_X1 U3869 ( .B1(U4043), .B2(n3047), .A(n3046), .ZN(U3558) );
  INV_X1 U3870 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n3049) );
  NAND2_X1 U3871 ( .A1(n4125), .A2(U4043), .ZN(n3048) );
  OAI21_X1 U3872 ( .B1(U4043), .B2(n3049), .A(n3048), .ZN(U3568) );
  INV_X1 U3873 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U3874 ( .A1(n3641), .A2(U4043), .ZN(n3050) );
  OAI21_X1 U3875 ( .B1(U4043), .B2(n3051), .A(n3050), .ZN(U3564) );
  INV_X1 U3876 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n3053) );
  NAND2_X1 U3877 ( .A1(n3500), .A2(U4043), .ZN(n3052) );
  OAI21_X1 U3878 ( .B1(U4043), .B2(n3053), .A(n3052), .ZN(U3563) );
  INV_X1 U3879 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n3058) );
  INV_X1 U3880 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3056) );
  NAND2_X1 U3881 ( .A1(n3720), .A2(REG1_REG_30__SCAN_IN), .ZN(n3055) );
  NAND2_X1 U3882 ( .A1(n2780), .A2(REG0_REG_30__SCAN_IN), .ZN(n3054) );
  OAI211_X1 U3883 ( .C1(n3724), .C2(n3056), .A(n3055), .B(n3054), .ZN(n3916)
         );
  NAND2_X1 U3884 ( .A1(n3916), .A2(U4043), .ZN(n3057) );
  OAI21_X1 U3885 ( .B1(U4043), .B2(n3058), .A(n3057), .ZN(U3580) );
  INV_X1 U3886 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n3060) );
  NAND2_X1 U3887 ( .A1(n3123), .A2(U4043), .ZN(n3059) );
  OAI21_X1 U3888 ( .B1(U4043), .B2(n3060), .A(n3059), .ZN(U3551) );
  NAND2_X1 U3889 ( .A1(n2805), .A2(n3088), .ZN(n3658) );
  NOR2_X1 U3890 ( .A1(n3738), .A2(n4700), .ZN(n3062) );
  INV_X1 U3891 ( .A(n4067), .ZN(n4330) );
  NOR2_X1 U3892 ( .A1(n4330), .A2(n4320), .ZN(n3061) );
  OAI22_X1 U3893 ( .A1(n3738), .A2(n3061), .B1(n2804), .B2(n4086), .ZN(n3090)
         );
  AOI211_X1 U3894 ( .C1(n3124), .C2(n3086), .A(n3062), .B(n3090), .ZN(n4664)
         );
  NAND2_X1 U3895 ( .A1(n4715), .A2(REG1_REG_0__SCAN_IN), .ZN(n3063) );
  OAI21_X1 U3896 ( .B1(n4664), .B2(n4715), .A(n3063), .ZN(U3518) );
  AOI21_X1 U3897 ( .B1(n3064), .B2(n3065), .A(n3653), .ZN(n3067) );
  OR2_X1 U3898 ( .A1(n3064), .A2(n3065), .ZN(n3066) );
  NAND2_X1 U3899 ( .A1(n3067), .A2(n3066), .ZN(n3076) );
  NOR2_X1 U3900 ( .A1(n3069), .A2(n3068), .ZN(n3070) );
  NAND2_X1 U3901 ( .A1(n3071), .A2(n3070), .ZN(n3122) );
  INV_X1 U3902 ( .A(n2805), .ZN(n3073) );
  INV_X1 U3903 ( .A(n2809), .ZN(n3072) );
  OAI22_X1 U3904 ( .A1(n3073), .A2(n3648), .B1(n3630), .B2(n3072), .ZN(n3074)
         );
  AOI21_X1 U3905 ( .B1(REG3_REG_1__SCAN_IN), .B2(n3122), .A(n3074), .ZN(n3075)
         );
  OAI211_X1 U3906 ( .C1(n3560), .C2(n2803), .A(n3076), .B(n3075), .ZN(U3219)
         );
  OAI22_X1 U3907 ( .A1(n3078), .A2(n4700), .B1(n2269), .B2(n3077), .ZN(n3079)
         );
  NOR2_X1 U3908 ( .A1(n3080), .A2(n3079), .ZN(n4666) );
  NAND2_X1 U3909 ( .A1(n4715), .A2(REG1_REG_1__SCAN_IN), .ZN(n3081) );
  OAI21_X1 U3910 ( .B1(n4666), .B2(n4715), .A(n3081), .ZN(U3519) );
  INV_X1 U3911 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n3083) );
  NAND2_X1 U3912 ( .A1(n3546), .A2(U4043), .ZN(n3082) );
  OAI21_X1 U3913 ( .B1(U4043), .B2(n3083), .A(n3082), .ZN(U3574) );
  INV_X1 U3914 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n3085) );
  NAND2_X1 U3915 ( .A1(n3988), .A2(U4043), .ZN(n3084) );
  OAI21_X1 U3916 ( .B1(U4043), .B2(n3085), .A(n3084), .ZN(U3575) );
  AOI21_X1 U3917 ( .B1(n3086), .B2(n3905), .A(n4350), .ZN(n3087) );
  NOR2_X1 U3918 ( .A1(n3088), .A2(n3087), .ZN(n3089) );
  INV_X2 U3919 ( .A(n2922), .ZN(n4333) );
  OAI21_X1 U3920 ( .B1(n3090), .B2(n3089), .A(n4333), .ZN(n3092) );
  AOI22_X1 U3921 ( .A1(n4485), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4631), .ZN(n3091) );
  OAI211_X1 U3922 ( .C1(n3738), .C2(n4076), .A(n3092), .B(n3091), .ZN(U3290)
         );
  OAI21_X1 U3923 ( .B1(n3093), .B2(n3094), .A(n3096), .ZN(n3097) );
  NAND2_X1 U3924 ( .A1(n3097), .A2(n3608), .ZN(n3100) );
  OAI22_X1 U3925 ( .A1(n2808), .A2(n3630), .B1(n3648), .B2(n2804), .ZN(n3098)
         );
  AOI21_X1 U3926 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3122), .A(n3098), .ZN(n3099)
         );
  OAI211_X1 U3927 ( .C1(n3560), .C2(n3101), .A(n3100), .B(n3099), .ZN(U3234)
         );
  OAI21_X1 U3928 ( .B1(n3104), .B2(n3103), .A(n3102), .ZN(n4635) );
  OAI21_X1 U3929 ( .B1(n3770), .B2(n3106), .A(n3105), .ZN(n3107) );
  NAND2_X1 U3930 ( .A1(n3107), .A2(n4320), .ZN(n3109) );
  AOI22_X1 U3931 ( .A1(n3123), .A2(n4144), .B1(n4350), .B2(n3114), .ZN(n3108)
         );
  OAI211_X1 U3932 ( .C1(n2808), .C2(n4086), .A(n3109), .B(n3108), .ZN(n3110)
         );
  AOI21_X1 U3933 ( .B1(n4330), .B2(n4635), .A(n3110), .ZN(n4638) );
  INV_X1 U3934 ( .A(n4638), .ZN(n3111) );
  AOI21_X1 U3935 ( .B1(n4676), .B2(n4635), .A(n3111), .ZN(n3119) );
  INV_X1 U3936 ( .A(n3138), .ZN(n3112) );
  AOI21_X1 U3937 ( .B1(n3114), .B2(n3113), .A(n3112), .ZN(n4632) );
  INV_X1 U3938 ( .A(n4468), .ZN(n3207) );
  INV_X1 U3939 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3115) );
  NOR2_X1 U3940 ( .A1(n4706), .A2(n3115), .ZN(n3116) );
  AOI21_X1 U3941 ( .B1(n4632), .B2(n3207), .A(n3116), .ZN(n3117) );
  OAI21_X1 U3942 ( .B1(n3119), .B2(n4704), .A(n3117), .ZN(U3471) );
  INV_X1 U3943 ( .A(n4417), .ZN(n3211) );
  AOI22_X1 U3944 ( .A1(n4632), .A2(n3211), .B1(REG1_REG_2__SCAN_IN), .B2(n4715), .ZN(n3118) );
  OAI21_X1 U3945 ( .B1(n3119), .B2(n4715), .A(n3118), .ZN(U3520) );
  XNOR2_X1 U3946 ( .A(n3120), .B(n3121), .ZN(n3835) );
  AOI22_X1 U3947 ( .A1(n3645), .A2(n3123), .B1(n3122), .B2(REG3_REG_0__SCAN_IN), .ZN(n3126) );
  NAND2_X1 U3948 ( .A1(n3643), .A2(n3124), .ZN(n3125) );
  OAI211_X1 U3949 ( .C1(n3835), .C2(n3653), .A(n3126), .B(n3125), .ZN(U3229)
         );
  NAND2_X1 U3950 ( .A1(n3102), .A2(n3127), .ZN(n3129) );
  INV_X1 U3951 ( .A(n3771), .ZN(n3128) );
  XNOR2_X1 U3952 ( .A(n3129), .B(n3128), .ZN(n4668) );
  NAND2_X1 U3953 ( .A1(n4668), .A2(n4330), .ZN(n3137) );
  XNOR2_X1 U3954 ( .A(n3130), .B(n3771), .ZN(n3135) );
  NAND2_X1 U3955 ( .A1(n2809), .A2(n4144), .ZN(n3132) );
  NAND2_X1 U3956 ( .A1(n3222), .A2(n4323), .ZN(n3131) );
  OAI211_X1 U3957 ( .C1(n3133), .C2(n4148), .A(n3132), .B(n3131), .ZN(n3134)
         );
  AOI21_X1 U3958 ( .B1(n3135), .B2(n4320), .A(n3134), .ZN(n3136) );
  AND2_X1 U3959 ( .A1(n3137), .A2(n3136), .ZN(n4670) );
  INV_X1 U3960 ( .A(n4076), .ZN(n4634) );
  AND2_X1 U3961 ( .A1(n3138), .A2(n3147), .ZN(n3139) );
  NOR2_X1 U3962 ( .A1(n3254), .A2(n3139), .ZN(n4667) );
  INV_X1 U3963 ( .A(n4667), .ZN(n3142) );
  AOI22_X1 U3964 ( .A1(n2922), .A2(REG2_REG_3__SCAN_IN), .B1(n4631), .B2(n3140), .ZN(n3141) );
  OAI21_X1 U3965 ( .B1(n4136), .B2(n3142), .A(n3141), .ZN(n3143) );
  AOI21_X1 U3966 ( .B1(n4668), .B2(n4634), .A(n3143), .ZN(n3144) );
  OAI21_X1 U3967 ( .B1(n4670), .B2(n4485), .A(n3144), .ZN(U3287) );
  XOR2_X1 U3968 ( .A(n3146), .B(n3145), .Z(n3154) );
  INV_X1 U3969 ( .A(n3222), .ZN(n3151) );
  NAND2_X1 U3970 ( .A1(n3643), .A2(n3147), .ZN(n3150) );
  AOI21_X1 U3971 ( .B1(n3627), .B2(n2809), .A(n3148), .ZN(n3149) );
  OAI211_X1 U3972 ( .C1(n3151), .C2(n3630), .A(n3150), .B(n3149), .ZN(n3152)
         );
  AOI21_X1 U3973 ( .B1(n3140), .B2(n3650), .A(n3152), .ZN(n3153) );
  OAI21_X1 U3974 ( .B1(n3154), .B2(n3653), .A(n3153), .ZN(U3215) );
  OAI211_X1 U3975 ( .C1(n3156), .C2(n3158), .A(n3157), .B(n3608), .ZN(n3163)
         );
  NAND2_X1 U3976 ( .A1(n3627), .A2(n3222), .ZN(n3160) );
  OAI211_X1 U3977 ( .C1(n2818), .C2(n3630), .A(n3160), .B(n3159), .ZN(n3161)
         );
  AOI21_X1 U3978 ( .B1(n3224), .B2(n3643), .A(n3161), .ZN(n3162) );
  OAI211_X1 U3979 ( .C1(n3617), .C2(n3227), .A(n3163), .B(n3162), .ZN(U3224)
         );
  XOR2_X1 U3980 ( .A(n3166), .B(n3165), .Z(n3167) );
  XNOR2_X1 U3981 ( .A(n3164), .B(n3167), .ZN(n3174) );
  INV_X1 U3982 ( .A(n3168), .ZN(n3185) );
  INV_X1 U3983 ( .A(n3830), .ZN(n3177) );
  NAND2_X1 U3984 ( .A1(n3632), .A2(n3184), .ZN(n3171) );
  AOI21_X1 U3985 ( .B1(n3627), .B2(n3832), .A(n3169), .ZN(n3170) );
  OAI211_X1 U3986 ( .C1(n3177), .C2(n3630), .A(n3171), .B(n3170), .ZN(n3172)
         );
  AOI21_X1 U3987 ( .B1(n3185), .B2(n3650), .A(n3172), .ZN(n3173) );
  OAI21_X1 U3988 ( .B1(n3174), .B2(n3653), .A(n3173), .ZN(U3236) );
  INV_X1 U3989 ( .A(n3669), .ZN(n3687) );
  OR2_X1 U3990 ( .A1(n3673), .A2(n3687), .ZN(n3181) );
  XNOR2_X1 U3991 ( .A(n3175), .B(n3181), .ZN(n3180) );
  OAI22_X1 U3992 ( .A1(n3177), .A2(n4086), .B1(n4148), .B2(n3176), .ZN(n3178)
         );
  AOI21_X1 U3993 ( .B1(n4144), .B2(n3832), .A(n3178), .ZN(n3179) );
  OAI21_X1 U3994 ( .B1(n3180), .B2(n4129), .A(n3179), .ZN(n3203) );
  INV_X1 U3995 ( .A(n3203), .ZN(n3190) );
  INV_X1 U3996 ( .A(n3181), .ZN(n3759) );
  XNOR2_X1 U3997 ( .A(n3182), .B(n3759), .ZN(n3204) );
  NAND2_X1 U3998 ( .A1(n4333), .A2(n4330), .ZN(n3183) );
  AOI21_X1 U3999 ( .B1(n3184), .B2(n3226), .A(n3306), .ZN(n3212) );
  INV_X1 U4000 ( .A(n3212), .ZN(n3187) );
  AOI22_X1 U4001 ( .A1(n4485), .A2(REG2_REG_6__SCAN_IN), .B1(n3185), .B2(n4631), .ZN(n3186) );
  OAI21_X1 U4002 ( .B1(n3187), .B2(n4136), .A(n3186), .ZN(n3188) );
  AOI21_X1 U4003 ( .B1(n3204), .B2(n3928), .A(n3188), .ZN(n3189) );
  OAI21_X1 U4004 ( .B1(n3190), .B2(n4485), .A(n3189), .ZN(U3284) );
  INV_X1 U4005 ( .A(n3255), .ZN(n3201) );
  NAND2_X1 U4006 ( .A1(n3643), .A2(n3191), .ZN(n3193) );
  INV_X1 U4007 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4255) );
  NOR2_X1 U4008 ( .A1(STATE_REG_SCAN_IN), .A2(n4255), .ZN(n4498) );
  AOI21_X1 U4009 ( .B1(n3645), .B2(n3832), .A(n4498), .ZN(n3192) );
  OAI211_X1 U4010 ( .C1(n2808), .C2(n3648), .A(n3193), .B(n3192), .ZN(n3200)
         );
  CLKBUF_X1 U4011 ( .A(n3194), .Z(n3197) );
  INV_X1 U4012 ( .A(n3195), .ZN(n3196) );
  AOI211_X1 U4013 ( .C1(n3198), .C2(n3197), .A(n3653), .B(n3196), .ZN(n3199)
         );
  AOI211_X1 U4014 ( .C1(n3201), .C2(n3650), .A(n3200), .B(n3199), .ZN(n3202)
         );
  INV_X1 U4015 ( .A(n3202), .ZN(U3227) );
  AOI21_X1 U4016 ( .B1(n3204), .B2(n4692), .A(n3203), .ZN(n3214) );
  INV_X1 U4017 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3205) );
  NOR2_X1 U4018 ( .A1(n4706), .A2(n3205), .ZN(n3206) );
  AOI21_X1 U4019 ( .B1(n3212), .B2(n3207), .A(n3206), .ZN(n3208) );
  OAI21_X1 U4020 ( .B1(n3214), .B2(n4704), .A(n3208), .ZN(U3479) );
  INV_X1 U4021 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3209) );
  NOR2_X1 U4022 ( .A1(n4718), .A2(n3209), .ZN(n3210) );
  AOI21_X1 U4023 ( .B1(n3212), .B2(n3211), .A(n3210), .ZN(n3213) );
  OAI21_X1 U4024 ( .B1(n3214), .B2(n4715), .A(n3213), .ZN(U3524) );
  INV_X1 U4025 ( .A(n3215), .ZN(n3670) );
  XOR2_X1 U4026 ( .A(n3216), .B(n3768), .Z(n4679) );
  OAI22_X1 U4027 ( .A1(n2818), .A2(n4086), .B1(n4148), .B2(n3217), .ZN(n3221)
         );
  XNOR2_X1 U4028 ( .A(n3218), .B(n3768), .ZN(n3219) );
  NOR2_X1 U4029 ( .A1(n3219), .A2(n4129), .ZN(n3220) );
  AOI211_X1 U4030 ( .C1(n4144), .C2(n3222), .A(n3221), .B(n3220), .ZN(n4680)
         );
  MUX2_X1 U4031 ( .A(n3223), .B(n4680), .S(n4333), .Z(n3230) );
  NAND2_X1 U4032 ( .A1(n3252), .A2(n3224), .ZN(n3225) );
  AND2_X1 U4033 ( .A1(n3226), .A2(n3225), .ZN(n4683) );
  INV_X1 U4034 ( .A(n3227), .ZN(n3228) );
  AOI22_X1 U4035 ( .A1(n4683), .A2(n4633), .B1(n3228), .B2(n4631), .ZN(n3229)
         );
  OAI211_X1 U4036 ( .C1(n4159), .C2(n4679), .A(n3230), .B(n3229), .ZN(U3285)
         );
  XNOR2_X1 U4037 ( .A(n3231), .B(n3232), .ZN(n3240) );
  INV_X1 U4038 ( .A(n3309), .ZN(n3238) );
  INV_X1 U4039 ( .A(n3272), .ZN(n3328) );
  NAND2_X1 U4040 ( .A1(n3632), .A2(n3233), .ZN(n3236) );
  AOI21_X1 U4041 ( .B1(n3627), .B2(n3831), .A(n3234), .ZN(n3235) );
  OAI211_X1 U4042 ( .C1(n3328), .C2(n3630), .A(n3236), .B(n3235), .ZN(n3237)
         );
  AOI21_X1 U40430 ( .B1(n3238), .B2(n3650), .A(n3237), .ZN(n3239) );
  OAI21_X1 U4044 ( .B1(n3240), .B2(n3653), .A(n3239), .ZN(U3210) );
  INV_X1 U4045 ( .A(n3241), .ZN(n3243) );
  NAND2_X1 U4046 ( .A1(n3243), .A2(n3772), .ZN(n3244) );
  NAND2_X1 U4047 ( .A1(n3245), .A2(n3244), .ZN(n4672) );
  XOR2_X1 U4048 ( .A(n3772), .B(n3246), .Z(n3251) );
  NAND2_X1 U4049 ( .A1(n2323), .A2(n4144), .ZN(n3247) );
  OAI21_X1 U4050 ( .B1(n3253), .B2(n4148), .A(n3247), .ZN(n3249) );
  NOR2_X1 U4051 ( .A1(n4672), .A2(n4067), .ZN(n3248) );
  AOI211_X1 U4052 ( .C1(n4323), .C2(n3832), .A(n3249), .B(n3248), .ZN(n3250)
         );
  OAI21_X1 U4053 ( .B1(n4129), .B2(n3251), .A(n3250), .ZN(n4674) );
  OAI211_X1 U4054 ( .C1(n3254), .C2(n3253), .A(n3252), .B(n2899), .ZN(n4673)
         );
  OAI22_X1 U4055 ( .A1(n4673), .A2(n4314), .B1(n4332), .B2(n3255), .ZN(n3256)
         );
  OAI21_X1 U4056 ( .B1(n4674), .B2(n3256), .A(n4333), .ZN(n3258) );
  NAND2_X1 U4057 ( .A1(n4485), .A2(REG2_REG_4__SCAN_IN), .ZN(n3257) );
  OAI211_X1 U4058 ( .C1(n4672), .C2(n4076), .A(n3258), .B(n3257), .ZN(U3286)
         );
  INV_X1 U4059 ( .A(n3260), .ZN(n3262) );
  NOR2_X1 U4060 ( .A1(n3262), .A2(n3261), .ZN(n3263) );
  XNOR2_X1 U4061 ( .A(n3259), .B(n3263), .ZN(n3269) );
  INV_X1 U4062 ( .A(n3829), .ZN(n3352) );
  NAND2_X1 U4063 ( .A1(n3627), .A2(n3830), .ZN(n3264) );
  NAND2_X1 U4064 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4508) );
  OAI211_X1 U4065 ( .C1(n3352), .C2(n3630), .A(n3264), .B(n4508), .ZN(n3266)
         );
  NOR2_X1 U4066 ( .A1(n3617), .A2(n3295), .ZN(n3265) );
  AOI211_X1 U4067 ( .C1(n3267), .C2(n3632), .A(n3266), .B(n3265), .ZN(n3268)
         );
  OAI21_X1 U4068 ( .B1(n3269), .B2(n3653), .A(n3268), .ZN(U3218) );
  INV_X1 U4069 ( .A(n3683), .ZN(n3690) );
  AND2_X1 U4070 ( .A1(n3690), .A2(n3678), .ZN(n3758) );
  INV_X1 U4071 ( .A(n3758), .ZN(n3270) );
  XNOR2_X1 U4072 ( .A(n3271), .B(n3270), .ZN(n3277) );
  NAND2_X1 U4073 ( .A1(n3272), .A2(n4144), .ZN(n3274) );
  NAND2_X1 U4074 ( .A1(n3828), .A2(n4323), .ZN(n3273) );
  OAI211_X1 U4075 ( .C1(n3275), .C2(n4148), .A(n3274), .B(n3273), .ZN(n3276)
         );
  AOI21_X1 U4076 ( .B1(n3277), .B2(n4320), .A(n3276), .ZN(n4697) );
  NAND2_X1 U4077 ( .A1(n3279), .A2(n3278), .ZN(n3280) );
  XNOR2_X1 U4078 ( .A(n3280), .B(n3758), .ZN(n4693) );
  NAND2_X1 U4079 ( .A1(n3293), .A2(n3324), .ZN(n3281) );
  NAND2_X1 U4080 ( .A1(n3338), .A2(n3281), .ZN(n4694) );
  INV_X1 U4081 ( .A(n3282), .ZN(n3330) );
  AOI22_X1 U4082 ( .A1(n2922), .A2(REG2_REG_9__SCAN_IN), .B1(n3330), .B2(n4631), .ZN(n3283) );
  OAI21_X1 U4083 ( .B1(n4694), .B2(n4136), .A(n3283), .ZN(n3284) );
  AOI21_X1 U4084 ( .B1(n4693), .B2(n3928), .A(n3284), .ZN(n3285) );
  OAI21_X1 U4085 ( .B1(n4697), .B2(n2922), .A(n3285), .ZN(U3281) );
  AND2_X1 U4086 ( .A1(n3679), .A2(n3689), .ZN(n3757) );
  XNOR2_X1 U4087 ( .A(n3286), .B(n3757), .ZN(n3289) );
  OAI22_X1 U4088 ( .A1(n3352), .A2(n4086), .B1(n4148), .B2(n3294), .ZN(n3287)
         );
  AOI21_X1 U4089 ( .B1(n4144), .B2(n3830), .A(n3287), .ZN(n3288) );
  OAI21_X1 U4090 ( .B1(n3289), .B2(n4129), .A(n3288), .ZN(n3315) );
  INV_X1 U4091 ( .A(n3315), .ZN(n3300) );
  OR2_X1 U4092 ( .A1(n3290), .A2(n3762), .ZN(n4689) );
  NAND2_X1 U4093 ( .A1(n4689), .A2(n3291), .ZN(n3292) );
  XNOR2_X1 U4094 ( .A(n3292), .B(n3757), .ZN(n3316) );
  OAI21_X1 U4095 ( .B1(n3307), .B2(n3294), .A(n3293), .ZN(n3321) );
  NOR2_X1 U4096 ( .A1(n3321), .A2(n4136), .ZN(n3298) );
  OAI22_X1 U4097 ( .A1(n4333), .A2(n3296), .B1(n3295), .B2(n4332), .ZN(n3297)
         );
  AOI211_X1 U4098 ( .C1(n3316), .C2(n3928), .A(n3298), .B(n3297), .ZN(n3299)
         );
  OAI21_X1 U4099 ( .B1(n3300), .B2(n4485), .A(n3299), .ZN(U3282) );
  XNOR2_X1 U4100 ( .A(n3301), .B(n3762), .ZN(n3304) );
  OAI22_X1 U4101 ( .A1(n3328), .A2(n4086), .B1(n4148), .B2(n3305), .ZN(n3302)
         );
  AOI21_X1 U4102 ( .B1(n4144), .B2(n3831), .A(n3302), .ZN(n3303) );
  OAI21_X1 U4103 ( .B1(n3304), .B2(n4129), .A(n3303), .ZN(n4687) );
  INV_X1 U4104 ( .A(n4687), .ZN(n3314) );
  OAI21_X1 U4105 ( .B1(n3306), .B2(n3305), .A(n2899), .ZN(n3308) );
  NOR2_X1 U4106 ( .A1(n3308), .A2(n3307), .ZN(n4688) );
  OAI22_X1 U4107 ( .A1(n4333), .A2(n3019), .B1(n3309), .B2(n4332), .ZN(n3312)
         );
  INV_X1 U4108 ( .A(n4689), .ZN(n3310) );
  AND2_X1 U4109 ( .A1(n3290), .A2(n3762), .ZN(n4686) );
  NOR3_X1 U4110 ( .A1(n3310), .A2(n4686), .A3(n4159), .ZN(n3311) );
  AOI211_X1 U4111 ( .C1(n4118), .C2(n4688), .A(n3312), .B(n3311), .ZN(n3313)
         );
  OAI21_X1 U4112 ( .B1(n4485), .B2(n3314), .A(n3313), .ZN(U3283) );
  INV_X1 U4113 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4507) );
  AOI21_X1 U4114 ( .B1(n3316), .B2(n4692), .A(n3315), .ZN(n3318) );
  MUX2_X1 U4115 ( .A(n4507), .B(n3318), .S(n4718), .Z(n3317) );
  OAI21_X1 U4116 ( .B1(n3321), .B2(n4417), .A(n3317), .ZN(U3526) );
  INV_X1 U4117 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3319) );
  MUX2_X1 U4118 ( .A(n3319), .B(n3318), .S(n4706), .Z(n3320) );
  OAI21_X1 U4119 ( .B1(n3321), .B2(n4468), .A(n3320), .ZN(U3483) );
  XOR2_X1 U4120 ( .A(n3322), .B(n3323), .Z(n3332) );
  NAND2_X1 U4121 ( .A1(n3643), .A2(n3324), .ZN(n3327) );
  NOR2_X1 U4122 ( .A1(STATE_REG_SCAN_IN), .A2(n3325), .ZN(n4519) );
  AOI21_X1 U4123 ( .B1(n3645), .B2(n3828), .A(n4519), .ZN(n3326) );
  OAI211_X1 U4124 ( .C1(n3328), .C2(n3648), .A(n3327), .B(n3326), .ZN(n3329)
         );
  AOI21_X1 U4125 ( .B1(n3330), .B2(n3650), .A(n3329), .ZN(n3331) );
  OAI21_X1 U4126 ( .B1(n3332), .B2(n3653), .A(n3331), .ZN(U3228) );
  AND2_X1 U4127 ( .A1(n3692), .A2(n3697), .ZN(n3766) );
  XNOR2_X1 U4128 ( .A(n3333), .B(n3766), .ZN(n3334) );
  NAND2_X1 U4129 ( .A1(n3334), .A2(n4320), .ZN(n3336) );
  AOI22_X1 U4130 ( .A1(n3396), .A2(n4323), .B1(n4350), .B2(n3354), .ZN(n3335)
         );
  OAI211_X1 U4131 ( .C1(n3352), .C2(n4327), .A(n3336), .B(n3335), .ZN(n3384)
         );
  INV_X1 U4132 ( .A(n3384), .ZN(n3346) );
  XOR2_X1 U4133 ( .A(n3337), .B(n3766), .Z(n3385) );
  INV_X1 U4134 ( .A(n3338), .ZN(n3341) );
  INV_X1 U4135 ( .A(n3452), .ZN(n3339) );
  OAI21_X1 U4136 ( .B1(n3341), .B2(n3340), .A(n3339), .ZN(n3390) );
  NOR2_X1 U4137 ( .A1(n3390), .A2(n4136), .ZN(n3344) );
  OAI22_X1 U4138 ( .A1(n4333), .A2(n3342), .B1(n3357), .B2(n4332), .ZN(n3343)
         );
  AOI211_X1 U4139 ( .C1(n3385), .C2(n3928), .A(n3344), .B(n3343), .ZN(n3345)
         );
  OAI21_X1 U4140 ( .B1(n4485), .B2(n3346), .A(n3345), .ZN(U3280) );
  AOI21_X1 U4141 ( .B1(n3347), .B2(n3348), .A(n3653), .ZN(n3350) );
  NAND2_X1 U4142 ( .A1(n3350), .A2(n3349), .ZN(n3356) );
  NAND2_X1 U4143 ( .A1(n3645), .A2(n3396), .ZN(n3351) );
  NAND2_X1 U4144 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4528) );
  OAI211_X1 U4145 ( .C1(n3352), .C2(n3648), .A(n3351), .B(n4528), .ZN(n3353)
         );
  AOI21_X1 U4146 ( .B1(n3354), .B2(n3643), .A(n3353), .ZN(n3355) );
  OAI211_X1 U4147 ( .C1(n3617), .C2(n3357), .A(n3356), .B(n3355), .ZN(U3214)
         );
  NAND2_X1 U4148 ( .A1(n3359), .A2(n3358), .ZN(n3414) );
  AND2_X1 U4149 ( .A1(n3411), .A2(n3412), .ZN(n3745) );
  XNOR2_X1 U4150 ( .A(n3414), .B(n3745), .ZN(n3363) );
  NAND2_X1 U4151 ( .A1(n3396), .A2(n4144), .ZN(n3361) );
  NAND2_X1 U4152 ( .A1(n3500), .A2(n4323), .ZN(n3360) );
  OAI211_X1 U4153 ( .C1(n3366), .C2(n4148), .A(n3361), .B(n3360), .ZN(n3362)
         );
  AOI21_X1 U4154 ( .B1(n3363), .B2(n4320), .A(n3362), .ZN(n3404) );
  INV_X1 U4155 ( .A(n3745), .ZN(n3365) );
  XNOR2_X1 U4156 ( .A(n3364), .B(n3365), .ZN(n3403) );
  OAI21_X1 U4157 ( .B1(n3449), .B2(n3366), .A(n3420), .ZN(n3409) );
  NOR2_X1 U4158 ( .A1(n3409), .A2(n4136), .ZN(n3369) );
  OAI22_X1 U4159 ( .A1(n4333), .A2(n3367), .B1(n3398), .B2(n4332), .ZN(n3368)
         );
  AOI211_X1 U4160 ( .C1(n3403), .C2(n3928), .A(n3369), .B(n3368), .ZN(n3370)
         );
  OAI21_X1 U4161 ( .B1(n4485), .B2(n3404), .A(n3370), .ZN(U3278) );
  XOR2_X1 U4162 ( .A(n3373), .B(n3372), .Z(n3374) );
  XNOR2_X1 U4163 ( .A(n3371), .B(n3374), .ZN(n3383) );
  INV_X1 U4164 ( .A(n3453), .ZN(n3381) );
  INV_X1 U4165 ( .A(n3828), .ZN(n3379) );
  NAND2_X1 U4166 ( .A1(n3632), .A2(n3375), .ZN(n3378) );
  NOR2_X1 U4167 ( .A1(STATE_REG_SCAN_IN), .A2(n3376), .ZN(n4538) );
  AOI21_X1 U4168 ( .B1(n3645), .B2(n3827), .A(n4538), .ZN(n3377) );
  OAI211_X1 U4169 ( .C1(n3379), .C2(n3648), .A(n3378), .B(n3377), .ZN(n3380)
         );
  AOI21_X1 U4170 ( .B1(n3381), .B2(n3650), .A(n3380), .ZN(n3382) );
  OAI21_X1 U4171 ( .B1(n3383), .B2(n3653), .A(n3382), .ZN(U3233) );
  INV_X1 U4172 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4527) );
  AOI21_X1 U4173 ( .B1(n3385), .B2(n4692), .A(n3384), .ZN(n3387) );
  MUX2_X1 U4174 ( .A(n4527), .B(n3387), .S(n4718), .Z(n3386) );
  OAI21_X1 U4175 ( .B1(n3390), .B2(n4417), .A(n3386), .ZN(U3528) );
  INV_X1 U4176 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3388) );
  MUX2_X1 U4177 ( .A(n3388), .B(n3387), .S(n4706), .Z(n3389) );
  OAI21_X1 U4178 ( .B1(n3390), .B2(n4468), .A(n3389), .ZN(U3487) );
  INV_X1 U4179 ( .A(n3392), .ZN(n3394) );
  NOR2_X1 U4180 ( .A1(n3394), .A2(n3393), .ZN(n3395) );
  XNOR2_X1 U4181 ( .A(n3391), .B(n3395), .ZN(n3402) );
  NAND2_X1 U4182 ( .A1(n3627), .A2(n3396), .ZN(n3397) );
  NAND2_X1 U4183 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4548) );
  OAI211_X1 U4184 ( .C1(n4328), .C2(n3630), .A(n3397), .B(n4548), .ZN(n3400)
         );
  NOR2_X1 U4185 ( .A1(n3617), .A2(n3398), .ZN(n3399) );
  AOI211_X1 U4186 ( .C1(n2135), .C2(n3632), .A(n3400), .B(n3399), .ZN(n3401)
         );
  OAI21_X1 U4187 ( .B1(n3402), .B2(n3653), .A(n3401), .ZN(U3221) );
  NAND2_X1 U4188 ( .A1(n3403), .A2(n4692), .ZN(n3405) );
  AND2_X1 U4189 ( .A1(n3405), .A2(n3404), .ZN(n3407) );
  INV_X1 U4190 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4236) );
  MUX2_X1 U4191 ( .A(n3407), .B(n4236), .S(n4704), .Z(n3406) );
  OAI21_X1 U4192 ( .B1(n3409), .B2(n4468), .A(n3406), .ZN(U3491) );
  INV_X1 U4193 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4547) );
  MUX2_X1 U4194 ( .A(n4547), .B(n3407), .S(n4718), .Z(n3408) );
  OAI21_X1 U4195 ( .B1(n4417), .B2(n3409), .A(n3408), .ZN(U3530) );
  XNOR2_X1 U4196 ( .A(n3500), .B(n3421), .ZN(n3747) );
  XOR2_X1 U4197 ( .A(n3747), .B(n3410), .Z(n3472) );
  INV_X1 U4198 ( .A(n3411), .ZN(n3413) );
  OAI21_X1 U4199 ( .B1(n3414), .B2(n3413), .A(n3412), .ZN(n3415) );
  XNOR2_X1 U4200 ( .A(n3415), .B(n3747), .ZN(n3418) );
  AOI22_X1 U4201 ( .A1(n3641), .A2(n4323), .B1(n4350), .B2(n3464), .ZN(n3416)
         );
  OAI21_X1 U4202 ( .B1(n2828), .B2(n4327), .A(n3416), .ZN(n3417) );
  AOI21_X1 U4203 ( .B1(n3418), .B2(n4320), .A(n3417), .ZN(n3419) );
  OAI21_X1 U4204 ( .B1(n3472), .B2(n4067), .A(n3419), .ZN(n3473) );
  NAND2_X1 U4205 ( .A1(n3473), .A2(n4333), .ZN(n3427) );
  INV_X1 U4206 ( .A(n3420), .ZN(n3422) );
  OAI21_X1 U4207 ( .B1(n3422), .B2(n3421), .A(n4306), .ZN(n3479) );
  INV_X1 U4208 ( .A(n3479), .ZN(n3425) );
  OAI22_X1 U4209 ( .A1(n4333), .A2(n3423), .B1(n3463), .B2(n4332), .ZN(n3424)
         );
  AOI21_X1 U4210 ( .B1(n3425), .B2(n4633), .A(n3424), .ZN(n3426) );
  OAI211_X1 U4211 ( .C1(n3472), .C2(n4076), .A(n3427), .B(n3426), .ZN(U3277)
         );
  XNOR2_X1 U4212 ( .A(n3428), .B(n3760), .ZN(n4410) );
  INV_X1 U4213 ( .A(n4410), .ZN(n3440) );
  NAND2_X1 U4214 ( .A1(n4317), .A2(n3702), .ZN(n3429) );
  XNOR2_X1 U4215 ( .A(n3429), .B(n3760), .ZN(n3432) );
  OAI22_X1 U4216 ( .A1(n3572), .A2(n4086), .B1(n4148), .B2(n3434), .ZN(n3430)
         );
  AOI21_X1 U4217 ( .B1(n4144), .B2(n3641), .A(n3430), .ZN(n3431) );
  OAI21_X1 U4218 ( .B1(n3432), .B2(n4129), .A(n3431), .ZN(n4409) );
  INV_X1 U4219 ( .A(n4307), .ZN(n3435) );
  INV_X1 U4220 ( .A(n4154), .ZN(n3433) );
  OAI21_X1 U4221 ( .B1(n3435), .B2(n3434), .A(n3433), .ZN(n4464) );
  INV_X1 U4222 ( .A(n3436), .ZN(n3651) );
  AOI22_X1 U4223 ( .A1(n4485), .A2(REG2_REG_15__SCAN_IN), .B1(n3651), .B2(
        n4631), .ZN(n3437) );
  OAI21_X1 U4224 ( .B1(n4464), .B2(n4136), .A(n3437), .ZN(n3438) );
  AOI21_X1 U4225 ( .B1(n4409), .B2(n4333), .A(n3438), .ZN(n3439) );
  OAI21_X1 U4226 ( .B1(n3440), .B2(n4159), .A(n3439), .ZN(U3275) );
  INV_X1 U4227 ( .A(n3441), .ZN(n3442) );
  AOI21_X1 U4228 ( .B1(n3767), .B2(n3443), .A(n3442), .ZN(n4701) );
  XOR2_X1 U4229 ( .A(n3767), .B(n3444), .Z(n3448) );
  OAI22_X1 U4230 ( .A1(n2828), .A2(n4086), .B1(n4148), .B2(n3451), .ZN(n3446)
         );
  NOR2_X1 U4231 ( .A1(n4701), .A2(n4067), .ZN(n3445) );
  AOI211_X1 U4232 ( .C1(n4144), .C2(n3828), .A(n3446), .B(n3445), .ZN(n3447)
         );
  OAI21_X1 U4233 ( .B1(n4129), .B2(n3448), .A(n3447), .ZN(n4703) );
  NAND2_X1 U4234 ( .A1(n4703), .A2(n4333), .ZN(n3458) );
  INV_X1 U4235 ( .A(n3449), .ZN(n3450) );
  OAI21_X1 U4236 ( .B1(n3452), .B2(n3451), .A(n3450), .ZN(n4699) );
  INV_X1 U4237 ( .A(n4699), .ZN(n3456) );
  OAI22_X1 U4238 ( .A1(n4333), .A2(n3454), .B1(n3453), .B2(n4332), .ZN(n3455)
         );
  AOI21_X1 U4239 ( .B1(n3456), .B2(n4633), .A(n3455), .ZN(n3457) );
  OAI211_X1 U4240 ( .C1(n4701), .C2(n4076), .A(n3458), .B(n3457), .ZN(U3279)
         );
  XNOR2_X1 U4241 ( .A(n3461), .B(n3460), .ZN(n3462) );
  XNOR2_X1 U4242 ( .A(n3459), .B(n3462), .ZN(n3471) );
  INV_X1 U4243 ( .A(n3463), .ZN(n3469) );
  NAND2_X1 U4244 ( .A1(n3632), .A2(n3464), .ZN(n3467) );
  INV_X1 U4245 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3465) );
  NOR2_X1 U4246 ( .A1(STATE_REG_SCAN_IN), .A2(n3465), .ZN(n4559) );
  AOI21_X1 U4247 ( .B1(n3645), .B2(n3641), .A(n4559), .ZN(n3466) );
  OAI211_X1 U4248 ( .C1(n2828), .C2(n3648), .A(n3467), .B(n3466), .ZN(n3468)
         );
  AOI21_X1 U4249 ( .B1(n3469), .B2(n3650), .A(n3468), .ZN(n3470) );
  OAI21_X1 U4250 ( .B1(n3471), .B2(n3653), .A(n3470), .ZN(U3231) );
  INV_X1 U4251 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3475) );
  INV_X1 U4252 ( .A(n3472), .ZN(n3474) );
  AOI21_X1 U4253 ( .B1(n4676), .B2(n3474), .A(n3473), .ZN(n3477) );
  MUX2_X1 U4254 ( .A(n3475), .B(n3477), .S(n4706), .Z(n3476) );
  OAI21_X1 U4255 ( .B1(n3479), .B2(n4468), .A(n3476), .ZN(U3493) );
  INV_X1 U4256 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3863) );
  MUX2_X1 U4257 ( .A(n3863), .B(n3477), .S(n4718), .Z(n3478) );
  OAI21_X1 U4258 ( .B1(n4417), .B2(n3479), .A(n3478), .ZN(U3531) );
  XNOR2_X1 U4259 ( .A(n3481), .B(n3480), .ZN(n3482) );
  NAND2_X1 U4260 ( .A1(n3482), .A2(n3608), .ZN(n3489) );
  AOI22_X1 U4261 ( .A1(n3942), .A2(n3645), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3487) );
  INV_X1 U4262 ( .A(n3937), .ZN(n3483) );
  NAND2_X1 U4263 ( .A1(n3483), .A2(n3650), .ZN(n3486) );
  NAND2_X1 U4264 ( .A1(n3643), .A2(n3941), .ZN(n3485) );
  NAND2_X1 U4265 ( .A1(n3970), .A2(n3627), .ZN(n3484) );
  AND4_X1 U4266 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(n3488)
         );
  NAND2_X1 U4267 ( .A1(n3489), .A2(n3488), .ZN(U3211) );
  AOI22_X1 U4268 ( .A1(n3491), .A2(n4631), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4485), .ZN(n3492) );
  OAI21_X1 U4269 ( .B1(n3493), .B2(n4136), .A(n3492), .ZN(n3494) );
  AOI21_X1 U4270 ( .B1(n3495), .B2(n4333), .A(n3494), .ZN(n3496) );
  OAI21_X1 U4271 ( .B1(n3490), .B2(n4159), .A(n3496), .ZN(U3262) );
  NOR2_X1 U4272 ( .A1(n2058), .A2(n3498), .ZN(n3499) );
  XNOR2_X1 U4273 ( .A(n3497), .B(n3499), .ZN(n3505) );
  NAND2_X1 U4274 ( .A1(n3627), .A2(n3500), .ZN(n3501) );
  NAND2_X1 U4275 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4574) );
  OAI211_X1 U4276 ( .C1(n3559), .C2(n3630), .A(n3501), .B(n4574), .ZN(n3503)
         );
  NOR2_X1 U4277 ( .A1(n3617), .A2(n4331), .ZN(n3502) );
  AOI211_X1 U4278 ( .C1(n4322), .C2(n3643), .A(n3503), .B(n3502), .ZN(n3504)
         );
  OAI21_X1 U4279 ( .B1(n3505), .B2(n3653), .A(n3504), .ZN(U3212) );
  NAND2_X1 U4280 ( .A1(n3506), .A2(n3608), .ZN(n3518) );
  AOI21_X1 U4281 ( .B1(n3507), .B2(n3509), .A(n3508), .ZN(n3517) );
  NAND2_X1 U4282 ( .A1(n3546), .A2(n3645), .ZN(n3511) );
  NAND2_X1 U4283 ( .A1(n3627), .A2(n4046), .ZN(n3510) );
  OAI211_X1 U4284 ( .C1(STATE_REG_SCAN_IN), .C2(n3512), .A(n3511), .B(n3510), 
        .ZN(n3514) );
  NOR2_X1 U4285 ( .A1(n3617), .A2(n4015), .ZN(n3513) );
  AOI211_X1 U4286 ( .C1(n3515), .C2(n3632), .A(n3514), .B(n3513), .ZN(n3516)
         );
  OAI21_X1 U4287 ( .B1(n3518), .B2(n3517), .A(n3516), .ZN(U3213) );
  OAI21_X1 U4288 ( .B1(n3522), .B2(n3520), .A(n3521), .ZN(n3523) );
  NAND2_X1 U4289 ( .A1(n3523), .A2(n3608), .ZN(n3528) );
  NAND2_X1 U4290 ( .A1(n3627), .A2(n4125), .ZN(n3524) );
  NAND2_X1 U4291 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3904) );
  OAI211_X1 U4292 ( .C1(n4087), .C2(n3630), .A(n3524), .B(n3904), .ZN(n3525)
         );
  AOI21_X1 U4293 ( .B1(n3526), .B2(n3643), .A(n3525), .ZN(n3527) );
  OAI211_X1 U4294 ( .C1(n3617), .C2(n4094), .A(n3528), .B(n3527), .ZN(U3216)
         );
  OAI21_X1 U4295 ( .B1(n3529), .B2(n3591), .A(n3593), .ZN(n3533) );
  NOR2_X1 U4296 ( .A1(n3531), .A2(n3530), .ZN(n3532) );
  XNOR2_X1 U4297 ( .A(n3533), .B(n3532), .ZN(n3538) );
  AOI22_X1 U4298 ( .A1(n3645), .A2(n4046), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3534) );
  OAI21_X1 U4299 ( .B1(n4087), .B2(n3648), .A(n3534), .ZN(n3536) );
  NOR2_X1 U4300 ( .A1(n3617), .A2(n4050), .ZN(n3535) );
  AOI211_X1 U4301 ( .C1(n4045), .C2(n3632), .A(n3536), .B(n3535), .ZN(n3537)
         );
  OAI21_X1 U4302 ( .B1(n3538), .B2(n3653), .A(n3537), .ZN(U3220) );
  INV_X1 U4303 ( .A(n3540), .ZN(n3542) );
  NAND2_X1 U4304 ( .A1(n3542), .A2(n3541), .ZN(n3543) );
  XNOR2_X1 U4305 ( .A(n3539), .B(n3543), .ZN(n3552) );
  AOI22_X1 U4306 ( .A1(n3970), .A2(n3645), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3550) );
  INV_X1 U4307 ( .A(n3544), .ZN(n3976) );
  NAND2_X1 U4308 ( .A1(n3650), .A2(n3976), .ZN(n3549) );
  NAND2_X1 U4309 ( .A1(n3643), .A2(n3545), .ZN(n3548) );
  NAND2_X1 U4310 ( .A1(n3546), .A2(n3627), .ZN(n3547) );
  NAND4_X1 U4311 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(n3551)
         );
  AOI21_X1 U4312 ( .B1(n3552), .B2(n3608), .A(n3551), .ZN(n3553) );
  INV_X1 U4313 ( .A(n3553), .ZN(U3222) );
  OAI21_X1 U4314 ( .B1(n3554), .B2(n3639), .A(n3555), .ZN(n3556) );
  XOR2_X1 U4315 ( .A(n3557), .B(n3556), .Z(n3558) );
  NAND2_X1 U4316 ( .A1(n3558), .A2(n3608), .ZN(n3564) );
  NAND2_X1 U4317 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4587) );
  OAI21_X1 U4318 ( .B1(n3648), .B2(n3559), .A(n4587), .ZN(n3562) );
  NOR2_X1 U4319 ( .A1(n3560), .A2(n4153), .ZN(n3561) );
  AOI211_X1 U4320 ( .C1(n3645), .C2(n4145), .A(n3562), .B(n3561), .ZN(n3563)
         );
  OAI211_X1 U4321 ( .C1(n3617), .C2(n4151), .A(n3564), .B(n3563), .ZN(U3223)
         );
  NOR2_X1 U4322 ( .A1(n3567), .A2(n2171), .ZN(n3568) );
  XNOR2_X1 U4323 ( .A(n3565), .B(n3568), .ZN(n3575) );
  INV_X1 U4324 ( .A(n3569), .ZN(n4134) );
  NAND2_X1 U4325 ( .A1(n3643), .A2(n4124), .ZN(n3571) );
  AND2_X1 U4326 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4598) );
  AOI21_X1 U4327 ( .B1(n3645), .B2(n4125), .A(n4598), .ZN(n3570) );
  OAI211_X1 U4328 ( .C1(n3572), .C2(n3648), .A(n3571), .B(n3570), .ZN(n3573)
         );
  AOI21_X1 U4329 ( .B1(n4134), .B2(n3650), .A(n3573), .ZN(n3574) );
  OAI21_X1 U4330 ( .B1(n3575), .B2(n3653), .A(n3574), .ZN(U3225) );
  NAND2_X1 U4331 ( .A1(n3576), .A2(n3577), .ZN(n3578) );
  XOR2_X1 U4332 ( .A(n3579), .B(n3578), .Z(n3588) );
  NOR2_X1 U4333 ( .A1(n3580), .A2(STATE_REG_SCAN_IN), .ZN(n3581) );
  AOI21_X1 U4334 ( .B1(n3988), .B2(n3645), .A(n3581), .ZN(n3586) );
  NAND2_X1 U4335 ( .A1(n3650), .A2(n3993), .ZN(n3585) );
  NAND2_X1 U4336 ( .A1(n3643), .A2(n3582), .ZN(n3584) );
  NAND2_X1 U4337 ( .A1(n3627), .A2(n4034), .ZN(n3583) );
  NAND4_X1 U4338 ( .A1(n3586), .A2(n3585), .A3(n3584), .A4(n3583), .ZN(n3587)
         );
  AOI21_X1 U4339 ( .B1(n3588), .B2(n3608), .A(n3587), .ZN(n3589) );
  INV_X1 U4340 ( .A(n3589), .ZN(U3226) );
  NOR2_X1 U4341 ( .A1(n3590), .A2(n3591), .ZN(n3595) );
  INV_X1 U4342 ( .A(n3591), .ZN(n3592) );
  AOI21_X1 U4343 ( .B1(n3593), .B2(n3592), .A(n3529), .ZN(n3594) );
  OAI21_X1 U4344 ( .B1(n3595), .B2(n3594), .A(n3608), .ZN(n3600) );
  OR2_X1 U4345 ( .A1(n3648), .A2(n3616), .ZN(n3597) );
  NAND2_X1 U4346 ( .A1(U3149), .A2(REG3_REG_20__SCAN_IN), .ZN(n3596) );
  OAI211_X1 U4347 ( .C1(n4063), .C2(n3630), .A(n3597), .B(n3596), .ZN(n3598)
         );
  AOI21_X1 U4348 ( .B1(n4061), .B2(n3632), .A(n3598), .ZN(n3599) );
  OAI211_X1 U4349 ( .C1(n3617), .C2(n4070), .A(n3600), .B(n3599), .ZN(U3230)
         );
  OAI21_X1 U4350 ( .B1(n3603), .B2(n3602), .A(n3507), .ZN(n3609) );
  NOR2_X1 U4351 ( .A1(n3617), .A2(n4025), .ZN(n3607) );
  NAND2_X1 U4352 ( .A1(n3643), .A2(n4033), .ZN(n3605) );
  AOI22_X1 U4353 ( .A1(n3645), .A2(n4034), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3604) );
  OAI211_X1 U4354 ( .C1(n4063), .C2(n3648), .A(n3605), .B(n3604), .ZN(n3606)
         );
  AOI211_X1 U4355 ( .C1(n3609), .C2(n3608), .A(n3607), .B(n3606), .ZN(n3610)
         );
  INV_X1 U4356 ( .A(n3610), .ZN(U3232) );
  XNOR2_X1 U4357 ( .A(n3613), .B(n3612), .ZN(n3614) );
  XNOR2_X1 U4358 ( .A(n3611), .B(n3614), .ZN(n3622) );
  NAND2_X1 U4359 ( .A1(n3627), .A2(n4145), .ZN(n3615) );
  NAND2_X1 U4360 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4627) );
  OAI211_X1 U4361 ( .C1(n3616), .C2(n3630), .A(n3615), .B(n4627), .ZN(n3619)
         );
  NOR2_X1 U4362 ( .A1(n3617), .A2(n4106), .ZN(n3618) );
  AOI211_X1 U4363 ( .C1(n3620), .C2(n3632), .A(n3619), .B(n3618), .ZN(n3621)
         );
  OAI21_X1 U4364 ( .B1(n3622), .B2(n3653), .A(n3621), .ZN(U3235) );
  NAND2_X1 U4365 ( .A1(n3625), .A2(n3624), .ZN(n3626) );
  XNOR2_X1 U4366 ( .A(n3623), .B(n3626), .ZN(n3637) );
  NAND2_X1 U4367 ( .A1(U3149), .A2(REG3_REG_26__SCAN_IN), .ZN(n3629) );
  NAND2_X1 U4368 ( .A1(n3988), .A2(n3627), .ZN(n3628) );
  OAI211_X1 U4369 ( .C1(n3631), .C2(n3630), .A(n3629), .B(n3628), .ZN(n3634)
         );
  AND2_X1 U4370 ( .A1(n3632), .A2(n3951), .ZN(n3633) );
  NOR2_X1 U4371 ( .A1(n3634), .A2(n3633), .ZN(n3636) );
  NAND2_X1 U4372 ( .A1(n3650), .A2(n3959), .ZN(n3635) );
  OAI211_X1 U4373 ( .C1(n3637), .C2(n3653), .A(n3636), .B(n3635), .ZN(U3237)
         );
  INV_X1 U4374 ( .A(n3555), .ZN(n3638) );
  NOR2_X1 U4375 ( .A1(n3554), .A2(n3638), .ZN(n3640) );
  XNOR2_X1 U4376 ( .A(n3640), .B(n3639), .ZN(n3654) );
  NAND2_X1 U4377 ( .A1(n3643), .A2(n3642), .ZN(n3647) );
  NOR2_X1 U4378 ( .A1(STATE_REG_SCAN_IN), .A2(n3644), .ZN(n4581) );
  AOI21_X1 U4379 ( .B1(n3645), .B2(n4126), .A(n4581), .ZN(n3646) );
  OAI211_X1 U4380 ( .C1(n2832), .C2(n3648), .A(n3647), .B(n3646), .ZN(n3649)
         );
  AOI21_X1 U4381 ( .B1(n3651), .B2(n3650), .A(n3649), .ZN(n3652) );
  OAI21_X1 U4382 ( .B1(n3654), .B2(n3653), .A(n3652), .ZN(U3238) );
  INV_X1 U4383 ( .A(n3742), .ZN(n3655) );
  NOR2_X1 U4384 ( .A1(n3656), .A2(n3655), .ZN(n3795) );
  INV_X1 U4385 ( .A(n3657), .ZN(n3660) );
  OAI211_X1 U4386 ( .C1(n3660), .C2(n2760), .A(n3659), .B(n3658), .ZN(n3662)
         );
  NAND3_X1 U4387 ( .A1(n3662), .A2(n3661), .A3(n2856), .ZN(n3665) );
  NAND3_X1 U4388 ( .A1(n3665), .A2(n3664), .A3(n3663), .ZN(n3668) );
  NAND3_X1 U4389 ( .A1(n3668), .A2(n3667), .A3(n3666), .ZN(n3671) );
  NAND4_X1 U4390 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3676)
         );
  INV_X1 U4391 ( .A(n3673), .ZN(n3674) );
  NAND3_X1 U4392 ( .A1(n3676), .A2(n3675), .A3(n3674), .ZN(n3677) );
  NAND3_X1 U4393 ( .A1(n3677), .A2(n3685), .A3(n3689), .ZN(n3680) );
  NAND3_X1 U4394 ( .A1(n3680), .A2(n3679), .A3(n3678), .ZN(n3696) );
  NAND2_X1 U4395 ( .A1(n3682), .A2(n3681), .ZN(n3684) );
  NOR2_X1 U4396 ( .A1(n3684), .A2(n3683), .ZN(n3695) );
  NAND2_X1 U4397 ( .A1(n3684), .A2(n3701), .ZN(n3781) );
  INV_X1 U4398 ( .A(n3685), .ZN(n3688) );
  NOR3_X1 U4399 ( .A1(n3688), .A2(n3687), .A3(n3686), .ZN(n3691) );
  NAND3_X1 U4400 ( .A1(n3691), .A2(n3690), .A3(n3689), .ZN(n3693) );
  NAND2_X1 U4401 ( .A1(n3693), .A2(n3692), .ZN(n3694) );
  AOI22_X1 U4402 ( .A1(n3696), .A2(n3695), .B1(n3781), .B2(n3694), .ZN(n3706)
         );
  NAND3_X1 U4403 ( .A1(n3699), .A2(n3698), .A3(n3697), .ZN(n3705) );
  INV_X1 U4404 ( .A(n3700), .ZN(n3703) );
  NAND2_X1 U4405 ( .A1(n3702), .A2(n3701), .ZN(n3782) );
  OAI21_X1 U4406 ( .B1(n3703), .B2(n3782), .A(n3781), .ZN(n3704) );
  OAI21_X1 U4407 ( .B1(n3706), .B2(n3705), .A(n3704), .ZN(n3707) );
  NAND2_X1 U4408 ( .A1(n3707), .A2(n3783), .ZN(n3708) );
  AOI21_X1 U4409 ( .B1(n3708), .B2(n3786), .A(n3784), .ZN(n3709) );
  NOR2_X1 U4410 ( .A1(n3709), .A2(n4001), .ZN(n3711) );
  INV_X1 U4411 ( .A(n3791), .ZN(n3710) );
  OAI21_X1 U4412 ( .B1(n3711), .B2(n3749), .A(n3710), .ZN(n3714) );
  OAI211_X1 U4413 ( .C1(n3712), .C2(n3791), .A(n3743), .B(n3753), .ZN(n3796)
         );
  INV_X1 U4414 ( .A(n3796), .ZN(n3713) );
  OAI21_X1 U4415 ( .B1(n3715), .B2(n3714), .A(n3713), .ZN(n3719) );
  NAND2_X1 U4416 ( .A1(n3725), .A2(DATAI_29_), .ZN(n3915) );
  NAND2_X1 U4417 ( .A1(n3823), .A2(n3915), .ZN(n3737) );
  NAND2_X1 U4418 ( .A1(n3737), .A2(n3912), .ZN(n3727) );
  NOR2_X1 U4419 ( .A1(n3716), .A2(n3727), .ZN(n3803) );
  INV_X1 U4420 ( .A(n3803), .ZN(n3717) );
  AOI211_X1 U4421 ( .C1(n3795), .C2(n3719), .A(n3718), .B(n3717), .ZN(n3729)
         );
  NOR2_X1 U4422 ( .A1(n3911), .A2(n3800), .ZN(n3728) );
  INV_X1 U4423 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3723) );
  NAND2_X1 U4424 ( .A1(n3720), .A2(REG1_REG_31__SCAN_IN), .ZN(n3722) );
  NAND2_X1 U4425 ( .A1(n2780), .A2(REG0_REG_31__SCAN_IN), .ZN(n3721) );
  OAI211_X1 U4426 ( .C1(n3724), .C2(n3723), .A(n3722), .B(n3721), .ZN(n4341)
         );
  NAND2_X1 U4427 ( .A1(n3725), .A2(DATAI_31_), .ZN(n4339) );
  NAND2_X1 U4428 ( .A1(n4341), .A2(n4339), .ZN(n3731) );
  NAND2_X1 U4429 ( .A1(n3725), .A2(DATAI_30_), .ZN(n4338) );
  OR2_X1 U4430 ( .A1(n3916), .A2(n4338), .ZN(n3726) );
  AND2_X1 U4431 ( .A1(n3731), .A2(n3726), .ZN(n3798) );
  OR2_X1 U4432 ( .A1(n3823), .A2(n3915), .ZN(n3794) );
  OAI211_X1 U4433 ( .C1(n3728), .C2(n3727), .A(n3798), .B(n3794), .ZN(n3802)
         );
  OR2_X1 U4434 ( .A1(n3729), .A2(n3802), .ZN(n3734) );
  NAND2_X1 U4435 ( .A1(n3916), .A2(n4338), .ZN(n3805) );
  OR2_X1 U4436 ( .A1(n4341), .A2(n4339), .ZN(n3730) );
  AND2_X1 U4437 ( .A1(n3805), .A2(n3730), .ZN(n3744) );
  INV_X1 U4438 ( .A(n3744), .ZN(n3732) );
  NAND2_X1 U4439 ( .A1(n3732), .A2(n3731), .ZN(n3733) );
  NAND2_X1 U4440 ( .A1(n3734), .A2(n3733), .ZN(n3813) );
  NAND2_X1 U4441 ( .A1(n3736), .A2(n3735), .ZN(n3950) );
  INV_X1 U4442 ( .A(n3950), .ZN(n3741) );
  NAND2_X1 U4443 ( .A1(n3794), .A2(n3737), .ZN(n3926) );
  NAND2_X1 U4444 ( .A1(n3738), .A2(n3798), .ZN(n3739) );
  OR2_X1 U4445 ( .A1(n3926), .A2(n3739), .ZN(n3740) );
  NOR3_X1 U4446 ( .A1(n3924), .A2(n3741), .A3(n3740), .ZN(n3780) );
  NAND2_X1 U4447 ( .A1(n3743), .A2(n3742), .ZN(n3968) );
  NAND2_X1 U4448 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  NOR4_X1 U4449 ( .A1(n3940), .A2(n3968), .A3(n3747), .A4(n3746), .ZN(n3779)
         );
  INV_X1 U4450 ( .A(n4004), .ZN(n3748) );
  INV_X1 U4451 ( .A(n3750), .ZN(n3982) );
  NOR2_X1 U4452 ( .A1(n3751), .A2(n3982), .ZN(n4007) );
  AND2_X1 U4453 ( .A1(n3753), .A2(n3752), .ZN(n3984) );
  XNOR2_X1 U4454 ( .A(n3826), .B(n4061), .ZN(n4059) );
  NAND4_X1 U4455 ( .A1(n4007), .A2(n3984), .A3(n4084), .A4(n4059), .ZN(n3756)
         );
  NOR3_X1 U4456 ( .A1(n4022), .A2(n4040), .A3(n3756), .ZN(n3778) );
  AND2_X1 U4457 ( .A1(n4079), .A2(n3999), .ZN(n4122) );
  NAND4_X1 U4458 ( .A1(n3759), .A2(n3758), .A3(n4122), .A4(n3757), .ZN(n3765)
         );
  INV_X1 U4459 ( .A(n3760), .ZN(n3761) );
  NAND4_X1 U4460 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n4319), .ZN(n3764)
         );
  NOR2_X1 U4461 ( .A1(n3765), .A2(n3764), .ZN(n3776) );
  INV_X1 U4462 ( .A(n4100), .ZN(n4108) );
  NAND4_X1 U4463 ( .A1(n3768), .A2(n4108), .A3(n3767), .A4(n3766), .ZN(n3774)
         );
  INV_X1 U4464 ( .A(n2855), .ZN(n3769) );
  NAND4_X1 U4465 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3773)
         );
  NOR2_X1 U4466 ( .A1(n3774), .A2(n3773), .ZN(n3775) );
  AND2_X1 U4467 ( .A1(n3776), .A2(n3775), .ZN(n3777) );
  NAND4_X1 U4468 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3811)
         );
  INV_X1 U4469 ( .A(n4338), .ZN(n4351) );
  OAI21_X1 U4470 ( .B1(n4318), .B2(n3782), .A(n3781), .ZN(n3787) );
  INV_X1 U4471 ( .A(n3783), .ZN(n3785) );
  AOI211_X1 U4472 ( .C1(n3787), .C2(n3786), .A(n3785), .B(n3784), .ZN(n3790)
         );
  INV_X1 U4473 ( .A(n3788), .ZN(n3789) );
  OR2_X1 U4474 ( .A1(n3790), .A2(n3789), .ZN(n3792) );
  AOI21_X1 U4475 ( .B1(n3793), .B2(n3792), .A(n3791), .ZN(n3797) );
  OAI211_X1 U4476 ( .C1(n3797), .C2(n3796), .A(n3795), .B(n3794), .ZN(n3801)
         );
  INV_X1 U4477 ( .A(n3798), .ZN(n3799) );
  NOR4_X1 U4478 ( .A1(n3801), .A2(n3911), .A3(n3800), .A4(n3799), .ZN(n3808)
         );
  INV_X1 U4479 ( .A(n3940), .ZN(n3804) );
  AOI21_X1 U4480 ( .B1(n3804), .B2(n3803), .A(n3802), .ZN(n3807) );
  AOI21_X1 U4481 ( .B1(n3805), .B2(n4341), .A(n4339), .ZN(n3806) );
  NOR3_X1 U4482 ( .A1(n3808), .A2(n3807), .A3(n3806), .ZN(n3809) );
  AOI21_X1 U4483 ( .B1(n4351), .B2(n4339), .A(n3809), .ZN(n3810) );
  MUX2_X1 U4484 ( .A(n3811), .B(n3810), .S(n2267), .Z(n3812) );
  MUX2_X1 U4485 ( .A(n3813), .B(n3812), .S(n4472), .Z(n3814) );
  XNOR2_X1 U4486 ( .A(n3814), .B(n3905), .ZN(n3822) );
  INV_X1 U4487 ( .A(n3815), .ZN(n3819) );
  NAND2_X1 U4488 ( .A1(n3817), .A2(n3816), .ZN(n3818) );
  OAI211_X1 U4489 ( .C1(n3819), .C2(n3837), .A(B_REG_SCAN_IN), .B(n3818), .ZN(
        n3820) );
  OAI21_X1 U4490 ( .B1(n3822), .B2(n3821), .A(n3820), .ZN(U3239) );
  MUX2_X1 U4491 ( .A(n4341), .B(DATAO_REG_31__SCAN_IN), .S(n3825), .Z(U3581)
         );
  MUX2_X1 U4492 ( .A(n3823), .B(DATAO_REG_29__SCAN_IN), .S(n3825), .Z(U3579)
         );
  MUX2_X1 U4493 ( .A(DATAO_REG_28__SCAN_IN), .B(n3942), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4494 ( .A(DATAO_REG_27__SCAN_IN), .B(n3952), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4495 ( .A(DATAO_REG_26__SCAN_IN), .B(n3970), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4496 ( .A(n4034), .B(DATAO_REG_23__SCAN_IN), .S(n3825), .Z(U3573)
         );
  MUX2_X1 U4497 ( .A(n4046), .B(DATAO_REG_22__SCAN_IN), .S(n3825), .Z(U3572)
         );
  MUX2_X1 U4498 ( .A(DATAO_REG_21__SCAN_IN), .B(n3824), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4499 ( .A(n3826), .B(DATAO_REG_20__SCAN_IN), .S(n3825), .Z(U3570)
         );
  MUX2_X1 U4500 ( .A(DATAO_REG_19__SCAN_IN), .B(n4110), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4501 ( .A(DATAO_REG_17__SCAN_IN), .B(n4145), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4502 ( .A(DATAO_REG_16__SCAN_IN), .B(n4126), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4503 ( .A(DATAO_REG_15__SCAN_IN), .B(n4324), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4504 ( .A(DATAO_REG_12__SCAN_IN), .B(n3827), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4505 ( .A(DATAO_REG_10__SCAN_IN), .B(n3828), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4506 ( .A(DATAO_REG_9__SCAN_IN), .B(n3829), .S(U4043), .Z(U3559) );
  MUX2_X1 U4507 ( .A(DATAO_REG_7__SCAN_IN), .B(n3830), .S(U4043), .Z(U3557) );
  MUX2_X1 U4508 ( .A(DATAO_REG_6__SCAN_IN), .B(n3831), .S(U4043), .Z(U3556) );
  MUX2_X1 U4509 ( .A(DATAO_REG_5__SCAN_IN), .B(n3832), .S(U4043), .Z(U3555) );
  MUX2_X1 U4510 ( .A(DATAO_REG_3__SCAN_IN), .B(n2323), .S(U4043), .Z(U3553) );
  MUX2_X1 U4511 ( .A(DATAO_REG_2__SCAN_IN), .B(n2809), .S(U4043), .Z(U3552) );
  MUX2_X1 U4512 ( .A(DATAO_REG_0__SCAN_IN), .B(n2805), .S(U4043), .Z(U3550) );
  NAND3_X1 U4513 ( .A1(n3835), .A2(n3834), .A3(n3833), .ZN(n3840) );
  INV_X1 U4514 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3836) );
  AOI21_X1 U4515 ( .B1(n4487), .B2(n3836), .A(n4478), .ZN(n4486) );
  OR2_X1 U4516 ( .A1(n3837), .A2(n3836), .ZN(n3838) );
  MUX2_X1 U4517 ( .A(n4486), .B(n3838), .S(n4488), .Z(n3839) );
  NAND3_X1 U4518 ( .A1(n3840), .A2(U4043), .A3(n3839), .ZN(n4503) );
  AOI22_X1 U4519 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4599), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3852) );
  XNOR2_X1 U4520 ( .A(n3842), .B(n3841), .ZN(n3843) );
  AOI22_X1 U4521 ( .A1(n2300), .A2(n4621), .B1(n4607), .B2(n3843), .ZN(n3851)
         );
  MUX2_X1 U4522 ( .A(REG2_REG_2__SCAN_IN), .B(n2968), .S(n3844), .Z(n3847) );
  NAND3_X1 U4523 ( .A1(n3847), .A2(n3846), .A3(n3845), .ZN(n3848) );
  NAND3_X1 U4524 ( .A1(n4609), .A2(n3849), .A3(n3848), .ZN(n3850) );
  NAND4_X1 U4525 ( .A1(n4503), .A2(n3852), .A3(n3851), .A4(n3850), .ZN(U3242)
         );
  INV_X1 U4526 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4527 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4646), .B1(n4620), .B2(
        n3853), .ZN(n4616) );
  OR2_X1 U4528 ( .A1(n4473), .A2(n4711), .ZN(n3854) );
  NAND2_X1 U4529 ( .A1(n3855), .A2(n3854), .ZN(n3857) );
  NAND2_X1 U4530 ( .A1(n4473), .A2(n4711), .ZN(n3856) );
  NAND2_X1 U4531 ( .A1(n3857), .A2(n3856), .ZN(n3858) );
  INV_X1 U4532 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U4533 ( .A1(n3878), .A2(n4713), .B1(REG1_REG_9__SCAN_IN), .B2(n4660), .ZN(n4516) );
  NOR2_X1 U4534 ( .A1(n4517), .A2(n4516), .ZN(n4515) );
  AOI21_X1 U4535 ( .B1(REG1_REG_9__SCAN_IN), .B2(n3878), .A(n4515), .ZN(n3860)
         );
  INV_X1 U4536 ( .A(n3883), .ZN(n4658) );
  NOR2_X1 U4537 ( .A1(n3860), .A2(n4658), .ZN(n3861) );
  XOR2_X1 U4538 ( .A(n3883), .B(n3860), .Z(n4526) );
  NOR2_X1 U4539 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  NOR2_X1 U4540 ( .A1(n3861), .A2(n4525), .ZN(n4537) );
  INV_X1 U4541 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4716) );
  AOI22_X1 U4542 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4656), .B1(n3877), .B2(
        n4716), .ZN(n4536) );
  NOR2_X1 U4543 ( .A1(n4537), .A2(n4536), .ZN(n4535) );
  AOI22_X1 U4544 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4653), .B1(n3890), .B2(
        n3863), .ZN(n4556) );
  NOR2_X1 U4545 ( .A1(n4557), .A2(n4556), .ZN(n4555) );
  AND2_X1 U4546 ( .A1(n3890), .A2(REG1_REG_13__SCAN_IN), .ZN(n3864) );
  INV_X1 U4547 ( .A(n3891), .ZN(n4573) );
  NAND2_X1 U4548 ( .A1(n3865), .A2(n4573), .ZN(n3866) );
  INV_X1 U4549 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4569) );
  INV_X1 U4550 ( .A(n3866), .ZN(n3867) );
  INV_X1 U4551 ( .A(n3896), .ZN(n4651) );
  INV_X1 U4552 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U4553 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4651), .B1(n3896), .B2(
        n4411), .ZN(n4583) );
  NAND2_X1 U4554 ( .A1(n3870), .A2(n4649), .ZN(n3871) );
  INV_X1 U4555 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U4556 ( .A1(n4593), .A2(n4592), .ZN(n4591) );
  AOI22_X1 U4557 ( .A1(n3899), .A2(REG1_REG_17__SCAN_IN), .B1(n3872), .B2(
        n4647), .ZN(n4605) );
  NAND2_X1 U4558 ( .A1(n4647), .A2(n3872), .ZN(n3873) );
  AOI21_X1 U4559 ( .B1(n4620), .B2(REG1_REG_18__SCAN_IN), .A(n4624), .ZN(n3875) );
  XNOR2_X1 U4560 ( .A(n4314), .B(REG1_REG_19__SCAN_IN), .ZN(n3874) );
  XNOR2_X1 U4561 ( .A(n3875), .B(n3874), .ZN(n3909) );
  AOI22_X1 U4562 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4646), .B1(n4620), .B2(
        n4107), .ZN(n4615) );
  NOR2_X1 U4563 ( .A1(n3899), .A2(REG2_REG_17__SCAN_IN), .ZN(n3876) );
  AOI21_X1 U4564 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3899), .A(n3876), .ZN(n4602) );
  NAND2_X1 U4565 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3877), .ZN(n3886) );
  AOI22_X1 U4566 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3877), .B1(n4656), .B2(
        n3454), .ZN(n4542) );
  AOI22_X1 U4567 ( .A1(n3878), .A2(REG2_REG_9__SCAN_IN), .B1(n2428), .B2(n4660), .ZN(n4522) );
  OAI21_X1 U4568 ( .B1(n3019), .B2(n4473), .A(n3879), .ZN(n3881) );
  NAND2_X1 U4569 ( .A1(n3881), .A2(n3880), .ZN(n3882) );
  XNOR2_X1 U4570 ( .A(n3881), .B(n4662), .ZN(n4512) );
  NAND2_X1 U4571 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4512), .ZN(n4511) );
  NAND2_X1 U4572 ( .A1(n3882), .A2(n4511), .ZN(n4521) );
  NAND2_X1 U4573 ( .A1(n4522), .A2(n4521), .ZN(n4520) );
  NAND2_X1 U4574 ( .A1(n3883), .A2(n3884), .ZN(n3885) );
  NAND2_X1 U4575 ( .A1(n3885), .A2(n4531), .ZN(n4541) );
  NAND2_X1 U4576 ( .A1(n4542), .A2(n4541), .ZN(n4540) );
  NAND2_X1 U4577 ( .A1(n3887), .A2(n3888), .ZN(n3889) );
  NOR2_X1 U4578 ( .A1(n3423), .A2(n4653), .ZN(n4560) );
  OAI22_X1 U4579 ( .A1(n4562), .A2(n4560), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3890), .ZN(n3892) );
  INV_X1 U4580 ( .A(n3895), .ZN(n3894) );
  NOR2_X1 U4581 ( .A1(n2518), .A2(n4567), .ZN(n4566) );
  AOI22_X1 U4582 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4651), .B1(n3896), .B2(
        n2537), .ZN(n4578) );
  NAND2_X1 U4583 ( .A1(n3897), .A2(n4649), .ZN(n3898) );
  NAND2_X1 U4584 ( .A1(n3898), .A2(n4589), .ZN(n4601) );
  INV_X1 U4585 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3900) );
  MUX2_X1 U4586 ( .A(n3900), .B(REG2_REG_19__SCAN_IN), .S(n3905), .Z(n3901) );
  XNOR2_X1 U4587 ( .A(n3902), .B(n3901), .ZN(n3907) );
  NAND2_X1 U4588 ( .A1(n4599), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3903) );
  OAI211_X1 U4589 ( .C1(n4612), .C2(n3905), .A(n3904), .B(n3903), .ZN(n3906)
         );
  AOI21_X1 U4590 ( .B1(n3907), .B2(n4609), .A(n3906), .ZN(n3908) );
  OAI21_X1 U4591 ( .B1(n3909), .B2(n4618), .A(n3908), .ZN(U3259) );
  INV_X1 U4592 ( .A(n3910), .ZN(n3920) );
  XOR2_X1 U4593 ( .A(n3926), .B(n3914), .Z(n3919) );
  AOI21_X1 U4594 ( .B1(n4487), .B2(B_REG_SCAN_IN), .A(n4086), .ZN(n4340) );
  INV_X1 U4595 ( .A(n3915), .ZN(n3930) );
  AOI22_X1 U4596 ( .A1(n3916), .A2(n4340), .B1(n4350), .B2(n3930), .ZN(n3918)
         );
  NAND2_X1 U4597 ( .A1(n3942), .A2(n4144), .ZN(n3917) );
  OAI211_X1 U4598 ( .C1(n3919), .C2(n4129), .A(n3918), .B(n3917), .ZN(n4355)
         );
  AOI21_X1 U4599 ( .B1(n4631), .B2(n3920), .A(n4355), .ZN(n3933) );
  AOI21_X1 U4600 ( .B1(n3925), .B2(n3924), .A(n3923), .ZN(n3927) );
  XNOR2_X1 U4601 ( .A(n3927), .B(n3926), .ZN(n4354) );
  NAND2_X1 U4602 ( .A1(n4354), .A2(n3928), .ZN(n3932) );
  AOI21_X1 U4603 ( .B1(n3930), .B2(n3929), .A(n4345), .ZN(n4356) );
  AOI22_X1 U4604 ( .A1(n4356), .A2(n4633), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4485), .ZN(n3931) );
  OAI211_X1 U4605 ( .C1(n4485), .C2(n3933), .A(n3932), .B(n3931), .ZN(U3354)
         );
  XOR2_X1 U4606 ( .A(n3940), .B(n3934), .Z(n4362) );
  AOI21_X1 U4607 ( .B1(n3941), .B2(n3956), .A(n3935), .ZN(n4360) );
  OAI22_X1 U4608 ( .A1(n3937), .A2(n4332), .B1(n4333), .B2(n3936), .ZN(n3938)
         );
  AOI21_X1 U4609 ( .B1(n4360), .B2(n4633), .A(n3938), .ZN(n3947) );
  XOR2_X1 U4610 ( .A(n3940), .B(n3939), .Z(n3945) );
  AOI22_X1 U4611 ( .A1(n3942), .A2(n4323), .B1(n4350), .B2(n3941), .ZN(n3944)
         );
  NAND2_X1 U4612 ( .A1(n3970), .A2(n4144), .ZN(n3943) );
  OAI211_X1 U4613 ( .C1(n3945), .C2(n4129), .A(n3944), .B(n3943), .ZN(n4359)
         );
  NAND2_X1 U4614 ( .A1(n4359), .A2(n4333), .ZN(n3946) );
  OAI211_X1 U4615 ( .C1(n4362), .C2(n4159), .A(n3947), .B(n3946), .ZN(U3263)
         );
  XOR2_X1 U4616 ( .A(n3950), .B(n3948), .Z(n4364) );
  INV_X1 U4617 ( .A(n4364), .ZN(n3963) );
  XOR2_X1 U4618 ( .A(n3950), .B(n3949), .Z(n3955) );
  AOI22_X1 U4619 ( .A1(n3988), .A2(n4144), .B1(n4350), .B2(n3951), .ZN(n3954)
         );
  NAND2_X1 U4620 ( .A1(n3952), .A2(n4323), .ZN(n3953) );
  OAI211_X1 U4621 ( .C1(n3955), .C2(n4129), .A(n3954), .B(n3953), .ZN(n4363)
         );
  INV_X1 U4622 ( .A(n3973), .ZN(n3958) );
  OAI21_X1 U4623 ( .B1(n3958), .B2(n3957), .A(n3956), .ZN(n4429) );
  AOI22_X1 U4624 ( .A1(n3959), .A2(n4631), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4485), .ZN(n3960) );
  OAI21_X1 U4625 ( .B1(n4429), .B2(n4136), .A(n3960), .ZN(n3961) );
  AOI21_X1 U4626 ( .B1(n4363), .B2(n4333), .A(n3961), .ZN(n3962) );
  OAI21_X1 U4627 ( .B1(n3963), .B2(n4159), .A(n3962), .ZN(U3264) );
  NAND2_X1 U4628 ( .A1(n3965), .A2(n3964), .ZN(n3966) );
  XNOR2_X1 U4629 ( .A(n3966), .B(n3968), .ZN(n4368) );
  INV_X1 U4630 ( .A(n4368), .ZN(n3980) );
  XOR2_X1 U4631 ( .A(n3968), .B(n3967), .Z(n3972) );
  OAI22_X1 U4632 ( .A1(n4008), .A2(n4327), .B1(n4148), .B2(n3974), .ZN(n3969)
         );
  AOI21_X1 U4633 ( .B1(n4323), .B2(n3970), .A(n3969), .ZN(n3971) );
  OAI21_X1 U4634 ( .B1(n3972), .B2(n4129), .A(n3971), .ZN(n4367) );
  INV_X1 U4635 ( .A(n3991), .ZN(n3975) );
  OAI21_X1 U4636 ( .B1(n3975), .B2(n3974), .A(n3973), .ZN(n4433) );
  AOI22_X1 U4637 ( .A1(n3976), .A2(n4631), .B1(n4485), .B2(
        REG2_REG_25__SCAN_IN), .ZN(n3977) );
  OAI21_X1 U4638 ( .B1(n4433), .B2(n4136), .A(n3977), .ZN(n3978) );
  AOI21_X1 U4639 ( .B1(n4367), .B2(n4333), .A(n3978), .ZN(n3979) );
  OAI21_X1 U4640 ( .B1(n3980), .B2(n4159), .A(n3979), .ZN(U3265) );
  XNOR2_X1 U4641 ( .A(n3981), .B(n3984), .ZN(n4372) );
  INV_X1 U4642 ( .A(n4372), .ZN(n3997) );
  NOR2_X1 U4643 ( .A1(n3983), .A2(n3982), .ZN(n3985) );
  XNOR2_X1 U4644 ( .A(n3985), .B(n3984), .ZN(n3990) );
  OAI22_X1 U4645 ( .A1(n3986), .A2(n4327), .B1(n4148), .B2(n3992), .ZN(n3987)
         );
  AOI21_X1 U4646 ( .B1(n3988), .B2(n4323), .A(n3987), .ZN(n3989) );
  OAI21_X1 U4647 ( .B1(n3990), .B2(n4129), .A(n3989), .ZN(n4371) );
  OAI21_X1 U4648 ( .B1(n4012), .B2(n3992), .A(n3991), .ZN(n4437) );
  AOI22_X1 U4649 ( .A1(n2922), .A2(REG2_REG_24__SCAN_IN), .B1(n3993), .B2(
        n4631), .ZN(n3994) );
  OAI21_X1 U4650 ( .B1(n4437), .B2(n4136), .A(n3994), .ZN(n3995) );
  AOI21_X1 U4651 ( .B1(n4371), .B2(n4333), .A(n3995), .ZN(n3996) );
  OAI21_X1 U4652 ( .B1(n3997), .B2(n4159), .A(n3996), .ZN(U3266) );
  XNOR2_X1 U4653 ( .A(n3998), .B(n4007), .ZN(n4376) );
  INV_X1 U4654 ( .A(n4376), .ZN(n4020) );
  INV_X1 U4655 ( .A(n3999), .ZN(n4078) );
  INV_X1 U4656 ( .A(n4001), .ZN(n4002) );
  OAI21_X1 U4657 ( .B1(n4058), .B2(n4003), .A(n4002), .ZN(n4042) );
  INV_X1 U4658 ( .A(n4040), .ZN(n4043) );
  NAND2_X1 U4659 ( .A1(n4042), .A2(n4043), .ZN(n4041) );
  NAND2_X1 U4660 ( .A1(n4041), .A2(n4004), .ZN(n4030) );
  INV_X1 U4661 ( .A(n4022), .ZN(n4031) );
  NAND2_X1 U4662 ( .A1(n4030), .A2(n4031), .ZN(n4029) );
  NAND2_X1 U4663 ( .A1(n4029), .A2(n4005), .ZN(n4006) );
  XOR2_X1 U4664 ( .A(n4007), .B(n4006), .Z(n4011) );
  OAI22_X1 U4665 ( .A1(n4008), .A2(n4086), .B1(n4148), .B2(n4014), .ZN(n4009)
         );
  AOI21_X1 U4666 ( .B1(n4144), .B2(n4046), .A(n4009), .ZN(n4010) );
  OAI21_X1 U4667 ( .B1(n4011), .B2(n4129), .A(n4010), .ZN(n4375) );
  INV_X1 U4668 ( .A(n4012), .ZN(n4013) );
  OAI21_X1 U4669 ( .B1(n4380), .B2(n4014), .A(n4013), .ZN(n4441) );
  NOR2_X1 U4670 ( .A1(n4441), .A2(n4136), .ZN(n4018) );
  OAI22_X1 U4671 ( .A1(n4333), .A2(n4016), .B1(n4015), .B2(n4332), .ZN(n4017)
         );
  AOI211_X1 U4672 ( .C1(n4375), .C2(n4333), .A(n4018), .B(n4017), .ZN(n4019)
         );
  OAI21_X1 U4673 ( .B1(n4020), .B2(n4159), .A(n4019), .ZN(U3267) );
  OAI21_X1 U4674 ( .B1(n4023), .B2(n4022), .A(n4021), .ZN(n4384) );
  INV_X1 U4675 ( .A(n4380), .ZN(n4028) );
  AND2_X1 U4676 ( .A1(n2033), .A2(n4033), .ZN(n4379) );
  NOR2_X1 U4677 ( .A1(n4379), .A2(n4136), .ZN(n4027) );
  NAND2_X1 U4678 ( .A1(n4485), .A2(REG2_REG_22__SCAN_IN), .ZN(n4024) );
  OAI21_X1 U4679 ( .B1(n4332), .B2(n4025), .A(n4024), .ZN(n4026) );
  AOI21_X1 U4680 ( .B1(n4028), .B2(n4027), .A(n4026), .ZN(n4038) );
  OAI21_X1 U4681 ( .B1(n4031), .B2(n4030), .A(n4029), .ZN(n4032) );
  NAND2_X1 U4682 ( .A1(n4032), .A2(n4320), .ZN(n4036) );
  AOI22_X1 U4683 ( .A1(n4034), .A2(n4323), .B1(n4350), .B2(n4033), .ZN(n4035)
         );
  OAI211_X1 U4684 ( .C1(n4063), .C2(n4327), .A(n4036), .B(n4035), .ZN(n4382)
         );
  NAND2_X1 U4685 ( .A1(n4382), .A2(n4333), .ZN(n4037) );
  OAI211_X1 U4686 ( .C1(n4384), .C2(n4159), .A(n4038), .B(n4037), .ZN(U3268)
         );
  XNOR2_X1 U4687 ( .A(n4039), .B(n4040), .ZN(n4386) );
  INV_X1 U4688 ( .A(n4386), .ZN(n4055) );
  OAI21_X1 U4689 ( .B1(n4043), .B2(n4042), .A(n4041), .ZN(n4044) );
  NAND2_X1 U4690 ( .A1(n4044), .A2(n4320), .ZN(n4048) );
  AOI22_X1 U4691 ( .A1(n4046), .A2(n4323), .B1(n4350), .B2(n4045), .ZN(n4047)
         );
  OAI211_X1 U4692 ( .C1(n4087), .C2(n4327), .A(n4048), .B(n4047), .ZN(n4385)
         );
  OAI21_X1 U4693 ( .B1(n2126), .B2(n4049), .A(n2033), .ZN(n4446) );
  NOR2_X1 U4694 ( .A1(n4446), .A2(n4136), .ZN(n4053) );
  OAI22_X1 U4695 ( .A1(n4333), .A2(n4051), .B1(n4050), .B2(n4332), .ZN(n4052)
         );
  AOI211_X1 U4696 ( .C1(n4385), .C2(n4333), .A(n4053), .B(n4052), .ZN(n4054)
         );
  OAI21_X1 U4697 ( .B1(n4055), .B2(n4159), .A(n4054), .ZN(U3269) );
  XOR2_X1 U4698 ( .A(n4059), .B(n4056), .Z(n4389) );
  NAND2_X1 U4699 ( .A1(n4058), .A2(n4057), .ZN(n4060) );
  XNOR2_X1 U4700 ( .A(n4060), .B(n4059), .ZN(n4065) );
  AOI22_X1 U4701 ( .A1(n4110), .A2(n4144), .B1(n4350), .B2(n4061), .ZN(n4062)
         );
  OAI21_X1 U4702 ( .B1(n4063), .B2(n4086), .A(n4062), .ZN(n4064) );
  AOI21_X1 U4703 ( .B1(n4065), .B2(n4320), .A(n4064), .ZN(n4066) );
  OAI21_X1 U4704 ( .B1(n4389), .B2(n4067), .A(n4066), .ZN(n4390) );
  NAND2_X1 U4705 ( .A1(n4390), .A2(n4333), .ZN(n4075) );
  OAI21_X1 U4706 ( .B1(n4091), .B2(n4069), .A(n4068), .ZN(n4450) );
  INV_X1 U4707 ( .A(n4450), .ZN(n4073) );
  OAI22_X1 U4708 ( .A1(n4333), .A2(n4071), .B1(n4070), .B2(n4332), .ZN(n4072)
         );
  AOI21_X1 U4709 ( .B1(n4073), .B2(n4633), .A(n4072), .ZN(n4074) );
  OAI211_X1 U4710 ( .C1(n4389), .C2(n4076), .A(n4075), .B(n4074), .ZN(U3270)
         );
  XOR2_X1 U4711 ( .A(n4084), .B(n4077), .Z(n4395) );
  INV_X1 U4712 ( .A(n4395), .ZN(n4098) );
  OR2_X1 U4713 ( .A1(n4123), .A2(n4078), .ZN(n4080) );
  NAND2_X1 U4714 ( .A1(n4080), .A2(n4079), .ZN(n4109) );
  INV_X1 U4715 ( .A(n4081), .ZN(n4083) );
  OAI21_X1 U4716 ( .B1(n4109), .B2(n4083), .A(n4082), .ZN(n4085) );
  XNOR2_X1 U4717 ( .A(n4085), .B(n4084), .ZN(n4090) );
  OAI22_X1 U4718 ( .A1(n4087), .A2(n4086), .B1(n4148), .B2(n4093), .ZN(n4088)
         );
  AOI21_X1 U4719 ( .B1(n4144), .B2(n4125), .A(n4088), .ZN(n4089) );
  OAI21_X1 U4720 ( .B1(n4090), .B2(n4129), .A(n4089), .ZN(n4394) );
  INV_X1 U4721 ( .A(n4091), .ZN(n4092) );
  OAI21_X1 U4722 ( .B1(n4103), .B2(n4093), .A(n4092), .ZN(n4454) );
  NOR2_X1 U4723 ( .A1(n4454), .A2(n4136), .ZN(n4096) );
  OAI22_X1 U4724 ( .A1(n4333), .A2(n3900), .B1(n4094), .B2(n4332), .ZN(n4095)
         );
  AOI211_X1 U4725 ( .C1(n4394), .C2(n4333), .A(n4096), .B(n4095), .ZN(n4097)
         );
  OAI21_X1 U4726 ( .B1(n4098), .B2(n4159), .A(n4097), .ZN(U3271) );
  OAI21_X1 U4727 ( .B1(n4101), .B2(n4100), .A(n4099), .ZN(n4102) );
  INV_X1 U4728 ( .A(n4102), .ZN(n4400) );
  INV_X1 U4729 ( .A(n4131), .ZN(n4105) );
  INV_X1 U4730 ( .A(n4103), .ZN(n4104) );
  OAI211_X1 U4731 ( .C1(n4105), .C2(n4113), .A(n4104), .B(n2899), .ZN(n4398)
         );
  INV_X1 U4732 ( .A(n4398), .ZN(n4119) );
  OAI22_X1 U4733 ( .A1(n4333), .A2(n4107), .B1(n4106), .B2(n4332), .ZN(n4117)
         );
  XNOR2_X1 U4734 ( .A(n4109), .B(n4108), .ZN(n4115) );
  NAND2_X1 U4735 ( .A1(n4145), .A2(n4144), .ZN(n4112) );
  NAND2_X1 U4736 ( .A1(n4110), .A2(n4323), .ZN(n4111) );
  OAI211_X1 U4737 ( .C1(n4113), .C2(n4148), .A(n4112), .B(n4111), .ZN(n4114)
         );
  AOI21_X1 U4738 ( .B1(n4115), .B2(n4320), .A(n4114), .ZN(n4399) );
  NOR2_X1 U4739 ( .A1(n4399), .A2(n4485), .ZN(n4116) );
  AOI211_X1 U4740 ( .C1(n4119), .C2(n4118), .A(n4117), .B(n4116), .ZN(n4120)
         );
  OAI21_X1 U4741 ( .B1(n4400), .B2(n4159), .A(n4120), .ZN(U3272) );
  XNOR2_X1 U4742 ( .A(n4121), .B(n4122), .ZN(n4402) );
  INV_X1 U4743 ( .A(n4402), .ZN(n4139) );
  XNOR2_X1 U4744 ( .A(n4123), .B(n4122), .ZN(n4130) );
  AOI22_X1 U4745 ( .A1(n4125), .A2(n4323), .B1(n4350), .B2(n4124), .ZN(n4128)
         );
  NAND2_X1 U4746 ( .A1(n4126), .A2(n4144), .ZN(n4127) );
  OAI211_X1 U4747 ( .C1(n4130), .C2(n4129), .A(n4128), .B(n4127), .ZN(n4401)
         );
  INV_X1 U4748 ( .A(n4404), .ZN(n4133) );
  OAI21_X1 U4749 ( .B1(n4133), .B2(n4132), .A(n4131), .ZN(n4459) );
  AOI22_X1 U4750 ( .A1(n2922), .A2(REG2_REG_17__SCAN_IN), .B1(n4134), .B2(
        n4631), .ZN(n4135) );
  OAI21_X1 U4751 ( .B1(n4459), .B2(n4136), .A(n4135), .ZN(n4137) );
  AOI21_X1 U4752 ( .B1(n4401), .B2(n4333), .A(n4137), .ZN(n4138) );
  OAI21_X1 U4753 ( .B1(n4139), .B2(n4159), .A(n4138), .ZN(U3273) );
  OAI21_X1 U4754 ( .B1(n4141), .B2(n4142), .A(n4140), .ZN(n4408) );
  XNOR2_X1 U4755 ( .A(n4143), .B(n4142), .ZN(n4150) );
  NAND2_X1 U4756 ( .A1(n4324), .A2(n4144), .ZN(n4147) );
  NAND2_X1 U4757 ( .A1(n4145), .A2(n4323), .ZN(n4146) );
  OAI211_X1 U4758 ( .C1(n4153), .C2(n4148), .A(n4147), .B(n4146), .ZN(n4149)
         );
  AOI21_X1 U4759 ( .B1(n4150), .B2(n4320), .A(n4149), .ZN(n4407) );
  NOR2_X1 U4760 ( .A1(n4332), .A2(n4151), .ZN(n4152) );
  AOI21_X1 U4761 ( .B1(n4485), .B2(REG2_REG_16__SCAN_IN), .A(n4152), .ZN(n4156) );
  OR2_X1 U4762 ( .A1(n4154), .A2(n4153), .ZN(n4405) );
  NAND3_X1 U4763 ( .A1(n4404), .A2(n4405), .A3(n4633), .ZN(n4155) );
  OAI211_X1 U4764 ( .C1(n4407), .C2(n4485), .A(n4156), .B(n4155), .ZN(n4157)
         );
  INV_X1 U4765 ( .A(n4157), .ZN(n4158) );
  OAI21_X1 U4766 ( .B1(n4408), .B2(n4159), .A(n4158), .ZN(U3274) );
  NOR3_X1 U4767 ( .A1(keyinput6), .A2(keyinput2), .A3(keyinput4), .ZN(n4173)
         );
  NAND2_X1 U4768 ( .A1(keyinput18), .A2(keyinput45), .ZN(n4163) );
  NOR2_X1 U4769 ( .A1(keyinput30), .A2(keyinput53), .ZN(n4161) );
  NOR4_X1 U4770 ( .A1(keyinput43), .A2(keyinput31), .A3(keyinput5), .A4(
        keyinput60), .ZN(n4160) );
  NAND4_X1 U4771 ( .A1(keyinput50), .A2(keyinput17), .A3(n4161), .A4(n4160), 
        .ZN(n4162) );
  NOR4_X1 U4772 ( .A1(keyinput54), .A2(keyinput59), .A3(n4163), .A4(n4162), 
        .ZN(n4172) );
  NAND3_X1 U4773 ( .A1(keyinput42), .A2(keyinput8), .A3(keyinput46), .ZN(n4170) );
  NOR2_X1 U4774 ( .A1(keyinput58), .A2(keyinput15), .ZN(n4164) );
  NAND3_X1 U4775 ( .A1(keyinput26), .A2(keyinput27), .A3(n4164), .ZN(n4169) );
  NOR3_X1 U4776 ( .A1(keyinput39), .A2(keyinput41), .A3(keyinput33), .ZN(n4167) );
  INV_X1 U4777 ( .A(keyinput29), .ZN(n4165) );
  NOR3_X1 U4778 ( .A1(keyinput52), .A2(keyinput20), .A3(n4165), .ZN(n4166) );
  NAND4_X1 U4779 ( .A1(keyinput49), .A2(n4167), .A3(keyinput24), .A4(n4166), 
        .ZN(n4168) );
  NOR4_X1 U4780 ( .A1(keyinput37), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(
        n4171) );
  NAND4_X1 U4781 ( .A1(keyinput36), .A2(n4173), .A3(n4172), .A4(n4171), .ZN(
        n4188) );
  NOR4_X1 U4782 ( .A1(keyinput10), .A2(keyinput19), .A3(keyinput63), .A4(
        keyinput32), .ZN(n4186) );
  NAND2_X1 U4783 ( .A1(keyinput55), .A2(keyinput51), .ZN(n4174) );
  NOR3_X1 U4784 ( .A1(keyinput47), .A2(keyinput11), .A3(n4174), .ZN(n4185) );
  INV_X1 U4785 ( .A(keyinput0), .ZN(n4175) );
  NAND4_X1 U4786 ( .A1(keyinput25), .A2(keyinput22), .A3(keyinput57), .A4(
        n4175), .ZN(n4176) );
  NOR4_X1 U4787 ( .A1(keyinput23), .A2(keyinput38), .A3(keyinput9), .A4(n4176), 
        .ZN(n4184) );
  NAND3_X1 U4788 ( .A1(keyinput34), .A2(keyinput56), .A3(keyinput40), .ZN(
        n4182) );
  NOR2_X1 U4789 ( .A1(keyinput48), .A2(keyinput14), .ZN(n4177) );
  NAND3_X1 U4790 ( .A1(keyinput12), .A2(keyinput16), .A3(n4177), .ZN(n4181) );
  NOR3_X1 U4791 ( .A1(keyinput35), .A2(keyinput21), .A3(keyinput7), .ZN(n4179)
         );
  NOR3_X1 U4792 ( .A1(keyinput3), .A2(keyinput28), .A3(keyinput62), .ZN(n4178)
         );
  NAND4_X1 U4793 ( .A1(keyinput61), .A2(n4179), .A3(keyinput44), .A4(n4178), 
        .ZN(n4180) );
  NOR4_X1 U4794 ( .A1(keyinput1), .A2(n4182), .A3(n4181), .A4(n4180), .ZN(
        n4183) );
  NAND4_X1 U4795 ( .A1(n4186), .A2(n4185), .A3(n4184), .A4(n4183), .ZN(n4187)
         );
  OAI21_X1 U4796 ( .B1(n4188), .B2(n4187), .A(keyinput13), .ZN(n4189) );
  NAND2_X1 U4797 ( .A1(n4189), .A2(REG3_REG_18__SCAN_IN), .ZN(n4305) );
  INV_X1 U4798 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4457) );
  INV_X1 U4799 ( .A(keyinput3), .ZN(n4191) );
  AOI22_X1 U4800 ( .A1(n4457), .A2(keyinput28), .B1(DATAO_REG_16__SCAN_IN), 
        .B2(n4191), .ZN(n4190) );
  OAI221_X1 U4801 ( .B1(n4457), .B2(keyinput28), .C1(n4191), .C2(
        DATAO_REG_16__SCAN_IN), .A(n4190), .ZN(n4202) );
  INV_X1 U4802 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4194) );
  INV_X1 U4803 ( .A(keyinput62), .ZN(n4193) );
  AOI22_X1 U4804 ( .A1(n4194), .A2(keyinput12), .B1(DATAO_REG_18__SCAN_IN), 
        .B2(n4193), .ZN(n4192) );
  OAI221_X1 U4805 ( .B1(n4194), .B2(keyinput12), .C1(n4193), .C2(
        DATAO_REG_18__SCAN_IN), .A(n4192), .ZN(n4201) );
  INV_X1 U4806 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4377) );
  INV_X1 U4807 ( .A(keyinput16), .ZN(n4196) );
  AOI22_X1 U4808 ( .A1(n4377), .A2(keyinput48), .B1(DATAO_REG_24__SCAN_IN), 
        .B2(n4196), .ZN(n4195) );
  OAI221_X1 U4809 ( .B1(n4377), .B2(keyinput48), .C1(n4196), .C2(
        DATAO_REG_24__SCAN_IN), .A(n4195), .ZN(n4200) );
  INV_X1 U4810 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4373) );
  INV_X1 U4811 ( .A(keyinput54), .ZN(n4198) );
  AOI22_X1 U4812 ( .A1(n4373), .A2(keyinput14), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(n4198), .ZN(n4197) );
  OAI221_X1 U4813 ( .B1(n4373), .B2(keyinput14), .C1(n4198), .C2(
        DATAO_REG_25__SCAN_IN), .A(n4197), .ZN(n4199) );
  NOR4_X1 U4814 ( .A1(n4202), .A2(n4201), .A3(n4200), .A4(n4199), .ZN(n4275)
         );
  INV_X1 U4815 ( .A(keyinput19), .ZN(n4205) );
  INV_X1 U4816 ( .A(keyinput63), .ZN(n4204) );
  AOI22_X1 U4817 ( .A1(n4205), .A2(DATAO_REG_11__SCAN_IN), .B1(
        DATAO_REG_13__SCAN_IN), .B2(n4204), .ZN(n4203) );
  OAI221_X1 U4818 ( .B1(n4205), .B2(DATAO_REG_11__SCAN_IN), .C1(n4204), .C2(
        DATAO_REG_13__SCAN_IN), .A(n4203), .ZN(n4217) );
  INV_X1 U4819 ( .A(keyinput32), .ZN(n4207) );
  AOI22_X1 U4820 ( .A1(n4208), .A2(keyinput51), .B1(DATAO_REG_14__SCAN_IN), 
        .B2(n4207), .ZN(n4206) );
  OAI221_X1 U4821 ( .B1(n4208), .B2(keyinput51), .C1(n4207), .C2(
        DATAO_REG_14__SCAN_IN), .A(n4206), .ZN(n4216) );
  INV_X1 U4822 ( .A(DATAI_24_), .ZN(n4210) );
  AOI22_X1 U4823 ( .A1(n4211), .A2(keyinput47), .B1(keyinput55), .B2(n4210), 
        .ZN(n4209) );
  OAI221_X1 U4824 ( .B1(n4211), .B2(keyinput47), .C1(n4210), .C2(keyinput55), 
        .A(n4209), .ZN(n4215) );
  INV_X1 U4825 ( .A(keyinput11), .ZN(n4213) );
  AOI22_X1 U4826 ( .A1(n3296), .A2(keyinput34), .B1(ADDR_REG_6__SCAN_IN), .B2(
        n4213), .ZN(n4212) );
  OAI221_X1 U4827 ( .B1(n3296), .B2(keyinput34), .C1(n4213), .C2(
        ADDR_REG_6__SCAN_IN), .A(n4212), .ZN(n4214) );
  NOR4_X1 U4828 ( .A1(n4217), .A2(n4216), .A3(n4215), .A4(n4214), .ZN(n4274)
         );
  INV_X1 U4829 ( .A(keyinput21), .ZN(n4219) );
  AOI22_X1 U4830 ( .A1(n3423), .A2(keyinput7), .B1(ADDR_REG_18__SCAN_IN), .B2(
        n4219), .ZN(n4218) );
  OAI221_X1 U4831 ( .B1(n3423), .B2(keyinput7), .C1(n4219), .C2(
        ADDR_REG_18__SCAN_IN), .A(n4218), .ZN(n4223) );
  INV_X1 U4832 ( .A(keyinput1), .ZN(n4221) );
  AOI22_X1 U4833 ( .A1(n4716), .A2(keyinput35), .B1(ADDR_REG_16__SCAN_IN), 
        .B2(n4221), .ZN(n4220) );
  OAI221_X1 U4834 ( .B1(n4716), .B2(keyinput35), .C1(n4221), .C2(
        ADDR_REG_16__SCAN_IN), .A(n4220), .ZN(n4222) );
  NOR2_X1 U4835 ( .A1(n4223), .A2(n4222), .ZN(n4246) );
  INV_X1 U4836 ( .A(D_REG_5__SCAN_IN), .ZN(n4640) );
  INV_X1 U4837 ( .A(D_REG_17__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U4838 ( .A1(n4640), .A2(keyinput49), .B1(keyinput41), .B2(n4639), 
        .ZN(n4224) );
  OAI221_X1 U4839 ( .B1(n4640), .B2(keyinput49), .C1(n4639), .C2(keyinput41), 
        .A(n4224), .ZN(n4229) );
  INV_X1 U4840 ( .A(keyinput56), .ZN(n4227) );
  INV_X1 U4841 ( .A(keyinput40), .ZN(n4226) );
  AOI22_X1 U4842 ( .A1(n4227), .A2(ADDR_REG_9__SCAN_IN), .B1(
        ADDR_REG_14__SCAN_IN), .B2(n4226), .ZN(n4225) );
  OAI221_X1 U4843 ( .B1(n4227), .B2(ADDR_REG_9__SCAN_IN), .C1(n4226), .C2(
        ADDR_REG_14__SCAN_IN), .A(n4225), .ZN(n4228) );
  NOR2_X1 U4844 ( .A1(n4229), .A2(n4228), .ZN(n4245) );
  INV_X1 U4845 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4684) );
  INV_X1 U4846 ( .A(DATAI_8_), .ZN(n4661) );
  AOI22_X1 U4847 ( .A1(n4684), .A2(keyinput42), .B1(n4661), .B2(keyinput8), 
        .ZN(n4230) );
  OAI221_X1 U4848 ( .B1(n4684), .B2(keyinput42), .C1(n4661), .C2(keyinput8), 
        .A(n4230), .ZN(n4233) );
  INV_X1 U4849 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4665) );
  INV_X1 U4850 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U4851 ( .A1(n4665), .A2(keyinput4), .B1(n4678), .B2(keyinput37), 
        .ZN(n4231) );
  OAI221_X1 U4852 ( .B1(n4665), .B2(keyinput4), .C1(n4678), .C2(keyinput37), 
        .A(n4231), .ZN(n4232) );
  NOR2_X1 U4853 ( .A1(n4233), .A2(n4232), .ZN(n4244) );
  AOI22_X1 U4854 ( .A1(n4236), .A2(keyinput60), .B1(n4235), .B2(keyinput6), 
        .ZN(n4234) );
  OAI221_X1 U4855 ( .B1(n4236), .B2(keyinput60), .C1(n4235), .C2(keyinput6), 
        .A(n4234), .ZN(n4242) );
  XNOR2_X1 U4856 ( .A(REG0_REG_13__SCAN_IN), .B(keyinput39), .ZN(n4240) );
  XNOR2_X1 U4857 ( .A(IR_REG_25__SCAN_IN), .B(keyinput24), .ZN(n4239) );
  XNOR2_X1 U4858 ( .A(IR_REG_31__SCAN_IN), .B(keyinput61), .ZN(n4238) );
  XNOR2_X1 U4859 ( .A(IR_REG_17__SCAN_IN), .B(keyinput44), .ZN(n4237) );
  NAND4_X1 U4860 ( .A1(n4240), .A2(n4239), .A3(n4238), .A4(n4237), .ZN(n4241)
         );
  NOR2_X1 U4861 ( .A1(n4242), .A2(n4241), .ZN(n4243) );
  NAND4_X1 U4862 ( .A1(n4246), .A2(n4245), .A3(n4244), .A4(n4243), .ZN(n4272)
         );
  INV_X1 U4863 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4691) );
  INV_X1 U4864 ( .A(DATAI_6_), .ZN(n4248) );
  AOI22_X1 U4865 ( .A1(n4691), .A2(keyinput2), .B1(keyinput36), .B2(n4248), 
        .ZN(n4247) );
  OAI221_X1 U4866 ( .B1(n4691), .B2(keyinput2), .C1(n4248), .C2(keyinput36), 
        .A(n4247), .ZN(n4253) );
  INV_X1 U4867 ( .A(DATAI_20_), .ZN(n4250) );
  AOI22_X1 U4868 ( .A1(n4251), .A2(keyinput26), .B1(keyinput27), .B2(n4250), 
        .ZN(n4249) );
  OAI221_X1 U4869 ( .B1(n4251), .B2(keyinput26), .C1(n4250), .C2(keyinput27), 
        .A(n4249), .ZN(n4252) );
  NOR2_X1 U4870 ( .A1(n4253), .A2(n4252), .ZN(n4270) );
  INV_X1 U4871 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4418) );
  AOI22_X1 U4872 ( .A1(n4255), .A2(keyinput15), .B1(keyinput52), .B2(n4418), 
        .ZN(n4254) );
  OAI221_X1 U4873 ( .B1(n4255), .B2(keyinput15), .C1(n4418), .C2(keyinput52), 
        .A(n4254), .ZN(n4256) );
  INV_X1 U4874 ( .A(n4256), .ZN(n4269) );
  INV_X1 U4875 ( .A(D_REG_2__SCAN_IN), .ZN(n4642) );
  INV_X1 U4876 ( .A(keyinput33), .ZN(n4257) );
  XNOR2_X1 U4877 ( .A(n4642), .B(n4257), .ZN(n4268) );
  XNOR2_X1 U4878 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput9), .ZN(n4261) );
  XNOR2_X1 U4879 ( .A(IR_REG_11__SCAN_IN), .B(keyinput5), .ZN(n4260) );
  XNOR2_X1 U4880 ( .A(IR_REG_22__SCAN_IN), .B(keyinput58), .ZN(n4259) );
  XNOR2_X1 U4881 ( .A(IR_REG_12__SCAN_IN), .B(keyinput31), .ZN(n4258) );
  NAND4_X1 U4882 ( .A1(n4261), .A2(n4260), .A3(n4259), .A4(n4258), .ZN(n4266)
         );
  XNOR2_X1 U4883 ( .A(DATAI_3_), .B(keyinput29), .ZN(n4264) );
  XNOR2_X1 U4884 ( .A(IR_REG_8__SCAN_IN), .B(keyinput46), .ZN(n4263) );
  XNOR2_X1 U4885 ( .A(keyinput20), .B(IR_REG_24__SCAN_IN), .ZN(n4262) );
  NAND3_X1 U4886 ( .A1(n4264), .A2(n4263), .A3(n4262), .ZN(n4265) );
  NOR2_X1 U4887 ( .A1(n4266), .A2(n4265), .ZN(n4267) );
  NAND4_X1 U4888 ( .A1(n4270), .A2(n4269), .A3(n4268), .A4(n4267), .ZN(n4271)
         );
  NOR2_X1 U4889 ( .A1(n4272), .A2(n4271), .ZN(n4273) );
  AND3_X1 U4890 ( .A1(n4275), .A2(n4274), .A3(n4273), .ZN(n4304) );
  AOI22_X1 U4891 ( .A1(keyinput23), .A2(n4107), .B1(keyinput13), .B2(n4276), 
        .ZN(n4277) );
  OAI21_X1 U4892 ( .B1(n4107), .B2(keyinput23), .A(n4277), .ZN(n4289) );
  INV_X1 U4893 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4280) );
  INV_X1 U4894 ( .A(keyinput38), .ZN(n4279) );
  AOI22_X1 U4895 ( .A1(n4280), .A2(keyinput25), .B1(ADDR_REG_19__SCAN_IN), 
        .B2(n4279), .ZN(n4278) );
  OAI221_X1 U4896 ( .B1(n4280), .B2(keyinput25), .C1(n4279), .C2(
        ADDR_REG_19__SCAN_IN), .A(n4278), .ZN(n4288) );
  INV_X1 U4897 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4707) );
  INV_X1 U4898 ( .A(keyinput22), .ZN(n4282) );
  AOI22_X1 U4899 ( .A1(n4707), .A2(keyinput0), .B1(DATAO_REG_4__SCAN_IN), .B2(
        n4282), .ZN(n4281) );
  OAI221_X1 U4900 ( .B1(n4707), .B2(keyinput0), .C1(n4282), .C2(
        DATAO_REG_4__SCAN_IN), .A(n4281), .ZN(n4287) );
  INV_X1 U4901 ( .A(keyinput57), .ZN(n4285) );
  INV_X1 U4902 ( .A(keyinput10), .ZN(n4284) );
  AOI22_X1 U4903 ( .A1(n4285), .A2(DATAO_REG_8__SCAN_IN), .B1(
        DATAO_REG_1__SCAN_IN), .B2(n4284), .ZN(n4283) );
  OAI221_X1 U4904 ( .B1(n4285), .B2(DATAO_REG_8__SCAN_IN), .C1(n4284), .C2(
        DATAO_REG_1__SCAN_IN), .A(n4283), .ZN(n4286) );
  NOR4_X1 U4905 ( .A1(n4289), .A2(n4288), .A3(n4287), .A4(n4286), .ZN(n4303)
         );
  INV_X1 U4906 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4292) );
  INV_X1 U4907 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4291) );
  AOI22_X1 U4908 ( .A1(n4292), .A2(keyinput45), .B1(n4291), .B2(keyinput50), 
        .ZN(n4290) );
  OAI221_X1 U4909 ( .B1(n4292), .B2(keyinput45), .C1(n4291), .C2(keyinput50), 
        .A(n4290), .ZN(n4301) );
  INV_X1 U4910 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4369) );
  INV_X1 U4911 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U4912 ( .A1(n4369), .A2(keyinput59), .B1(n4365), .B2(keyinput18), 
        .ZN(n4293) );
  OAI221_X1 U4913 ( .B1(n4369), .B2(keyinput59), .C1(n4365), .C2(keyinput18), 
        .A(n4293), .ZN(n4300) );
  INV_X1 U4914 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4421) );
  AOI22_X1 U4915 ( .A1(n4421), .A2(keyinput53), .B1(n2518), .B2(keyinput43), 
        .ZN(n4294) );
  OAI221_X1 U4916 ( .B1(n4421), .B2(keyinput53), .C1(n2518), .C2(keyinput43), 
        .A(n4294), .ZN(n4299) );
  INV_X1 U4917 ( .A(keyinput17), .ZN(n4297) );
  INV_X1 U4918 ( .A(keyinput30), .ZN(n4296) );
  AOI22_X1 U4919 ( .A1(n4297), .A2(DATAO_REG_29__SCAN_IN), .B1(
        DATAO_REG_30__SCAN_IN), .B2(n4296), .ZN(n4295) );
  OAI221_X1 U4920 ( .B1(n4297), .B2(DATAO_REG_29__SCAN_IN), .C1(n4296), .C2(
        DATAO_REG_30__SCAN_IN), .A(n4295), .ZN(n4298) );
  NOR4_X1 U4921 ( .A1(n4301), .A2(n4300), .A3(n4299), .A4(n4298), .ZN(n4302)
         );
  NAND4_X1 U4922 ( .A1(n4305), .A2(n4304), .A3(n4303), .A4(n4302), .ZN(n4337)
         );
  INV_X1 U4923 ( .A(n4306), .ZN(n4309) );
  OAI21_X1 U4924 ( .B1(n4309), .B2(n4308), .A(n4307), .ZN(n4469) );
  NOR2_X1 U4925 ( .A1(n4469), .A2(n2269), .ZN(n4316) );
  OAI21_X1 U4926 ( .B1(n4312), .B2(n4311), .A(n4310), .ZN(n4415) );
  INV_X1 U4927 ( .A(n4415), .ZN(n4313) );
  NOR2_X1 U4928 ( .A1(n4313), .A2(n2259), .ZN(n4315) );
  MUX2_X1 U4929 ( .A(n4316), .B(n4315), .S(n4314), .Z(n4335) );
  OAI21_X1 U4930 ( .B1(n4319), .B2(n4318), .A(n4317), .ZN(n4321) );
  NAND2_X1 U4931 ( .A1(n4321), .A2(n4320), .ZN(n4326) );
  AOI22_X1 U4932 ( .A1(n4324), .A2(n4323), .B1(n4350), .B2(n4322), .ZN(n4325)
         );
  OAI211_X1 U4933 ( .C1(n4328), .C2(n4327), .A(n4326), .B(n4325), .ZN(n4329)
         );
  AOI21_X1 U4934 ( .B1(n4415), .B2(n4330), .A(n4329), .ZN(n4413) );
  OAI211_X1 U4935 ( .C1(n4332), .C2(n4331), .A(n4413), .B(n4333), .ZN(n4334)
         );
  OAI22_X1 U4936 ( .A1(n4335), .A2(n4334), .B1(REG2_REG_14__SCAN_IN), .B2(
        n4333), .ZN(n4336) );
  XOR2_X1 U4937 ( .A(n4337), .B(n4336), .Z(U3276) );
  NAND2_X1 U4938 ( .A1(n4345), .A2(n4338), .ZN(n4346) );
  XNOR2_X1 U4939 ( .A(n4346), .B(n4339), .ZN(n4479) );
  INV_X1 U4940 ( .A(n4479), .ZN(n4420) );
  INV_X1 U4941 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4343) );
  INV_X1 U4942 ( .A(n4339), .ZN(n4342) );
  AND2_X1 U4943 ( .A1(n4341), .A2(n4340), .ZN(n4349) );
  AOI21_X1 U4944 ( .B1(n4342), .B2(n4350), .A(n4349), .ZN(n4481) );
  MUX2_X1 U4945 ( .A(n4343), .B(n4481), .S(n4718), .Z(n4344) );
  OAI21_X1 U4946 ( .B1(n4420), .B2(n4417), .A(n4344), .ZN(U3549) );
  INV_X1 U4947 ( .A(n4345), .ZN(n4348) );
  INV_X1 U4948 ( .A(n4346), .ZN(n4347) );
  AOI21_X1 U4949 ( .B1(n4351), .B2(n4348), .A(n4347), .ZN(n4482) );
  INV_X1 U4950 ( .A(n4482), .ZN(n4423) );
  INV_X1 U4951 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4352) );
  AOI21_X1 U4952 ( .B1(n4351), .B2(n4350), .A(n4349), .ZN(n4484) );
  MUX2_X1 U4953 ( .A(n4352), .B(n4484), .S(n4718), .Z(n4353) );
  OAI21_X1 U4954 ( .B1(n4423), .B2(n4417), .A(n4353), .ZN(U3548) );
  NAND2_X1 U4955 ( .A1(n4354), .A2(n4692), .ZN(n4358) );
  NAND2_X1 U4956 ( .A1(n4358), .A2(n4357), .ZN(n4424) );
  MUX2_X1 U4957 ( .A(REG1_REG_29__SCAN_IN), .B(n4424), .S(n4718), .Z(U3547) );
  AOI21_X1 U4958 ( .B1(n2899), .B2(n4360), .A(n4359), .ZN(n4361) );
  OAI21_X1 U4959 ( .B1(n4362), .B2(n4685), .A(n4361), .ZN(n4425) );
  MUX2_X1 U4960 ( .A(REG1_REG_27__SCAN_IN), .B(n4425), .S(n4718), .Z(U3545) );
  AOI21_X1 U4961 ( .B1(n4364), .B2(n4692), .A(n4363), .ZN(n4426) );
  MUX2_X1 U4962 ( .A(n4365), .B(n4426), .S(n4718), .Z(n4366) );
  OAI21_X1 U4963 ( .B1(n4417), .B2(n4429), .A(n4366), .ZN(U3544) );
  AOI21_X1 U4964 ( .B1(n4368), .B2(n4692), .A(n4367), .ZN(n4430) );
  MUX2_X1 U4965 ( .A(n4369), .B(n4430), .S(n4718), .Z(n4370) );
  OAI21_X1 U4966 ( .B1(n4417), .B2(n4433), .A(n4370), .ZN(U3543) );
  AOI21_X1 U4967 ( .B1(n4372), .B2(n4692), .A(n4371), .ZN(n4434) );
  MUX2_X1 U4968 ( .A(n4373), .B(n4434), .S(n4718), .Z(n4374) );
  OAI21_X1 U4969 ( .B1(n4417), .B2(n4437), .A(n4374), .ZN(U3542) );
  AOI21_X1 U4970 ( .B1(n4376), .B2(n4692), .A(n4375), .ZN(n4438) );
  MUX2_X1 U4971 ( .A(n4377), .B(n4438), .S(n4718), .Z(n4378) );
  OAI21_X1 U4972 ( .B1(n4417), .B2(n4441), .A(n4378), .ZN(U3541) );
  NOR3_X1 U4973 ( .A1(n4380), .A2(n4379), .A3(n2269), .ZN(n4381) );
  NOR2_X1 U4974 ( .A1(n4382), .A2(n4381), .ZN(n4383) );
  OAI21_X1 U4975 ( .B1(n4384), .B2(n4685), .A(n4383), .ZN(n4442) );
  MUX2_X1 U4976 ( .A(REG1_REG_22__SCAN_IN), .B(n4442), .S(n4718), .Z(U3540) );
  INV_X1 U4977 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4387) );
  AOI21_X1 U4978 ( .B1(n4386), .B2(n4692), .A(n4385), .ZN(n4443) );
  MUX2_X1 U4979 ( .A(n4387), .B(n4443), .S(n4718), .Z(n4388) );
  OAI21_X1 U4980 ( .B1(n4417), .B2(n4446), .A(n4388), .ZN(U3539) );
  INV_X1 U4981 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4392) );
  INV_X1 U4982 ( .A(n4389), .ZN(n4391) );
  AOI21_X1 U4983 ( .B1(n4676), .B2(n4391), .A(n4390), .ZN(n4447) );
  MUX2_X1 U4984 ( .A(n4392), .B(n4447), .S(n4718), .Z(n4393) );
  OAI21_X1 U4985 ( .B1(n4417), .B2(n4450), .A(n4393), .ZN(U3538) );
  INV_X1 U4986 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4396) );
  AOI21_X1 U4987 ( .B1(n4395), .B2(n4692), .A(n4394), .ZN(n4451) );
  MUX2_X1 U4988 ( .A(n4396), .B(n4451), .S(n4718), .Z(n4397) );
  OAI21_X1 U4989 ( .B1(n4417), .B2(n4454), .A(n4397), .ZN(U3537) );
  OAI211_X1 U4990 ( .C1(n4400), .C2(n4685), .A(n4399), .B(n4398), .ZN(n4455)
         );
  MUX2_X1 U4991 ( .A(REG1_REG_18__SCAN_IN), .B(n4455), .S(n4718), .Z(U3536) );
  AOI21_X1 U4992 ( .B1(n4402), .B2(n4692), .A(n4401), .ZN(n4456) );
  MUX2_X1 U4993 ( .A(n3872), .B(n4456), .S(n4718), .Z(n4403) );
  OAI21_X1 U4994 ( .B1(n4417), .B2(n4459), .A(n4403), .ZN(U3535) );
  NAND3_X1 U4995 ( .A1(n4405), .A2(n2899), .A3(n4404), .ZN(n4406) );
  OAI211_X1 U4996 ( .C1(n4408), .C2(n4685), .A(n4407), .B(n4406), .ZN(n4460)
         );
  MUX2_X1 U4997 ( .A(REG1_REG_16__SCAN_IN), .B(n4460), .S(n4718), .Z(U3534) );
  AOI21_X1 U4998 ( .B1(n4410), .B2(n4692), .A(n4409), .ZN(n4461) );
  MUX2_X1 U4999 ( .A(n4411), .B(n4461), .S(n4718), .Z(n4412) );
  OAI21_X1 U5000 ( .B1(n4417), .B2(n4464), .A(n4412), .ZN(U3533) );
  INV_X1 U5001 ( .A(n4413), .ZN(n4414) );
  AOI21_X1 U5002 ( .B1(n4676), .B2(n4415), .A(n4414), .ZN(n4465) );
  MUX2_X1 U5003 ( .A(n4569), .B(n4465), .S(n4718), .Z(n4416) );
  OAI21_X1 U5004 ( .B1(n4469), .B2(n4417), .A(n4416), .ZN(U3532) );
  MUX2_X1 U5005 ( .A(n4418), .B(n4481), .S(n4706), .Z(n4419) );
  OAI21_X1 U5006 ( .B1(n4420), .B2(n4468), .A(n4419), .ZN(U3517) );
  MUX2_X1 U5007 ( .A(n4421), .B(n4484), .S(n4706), .Z(n4422) );
  OAI21_X1 U5008 ( .B1(n4423), .B2(n4468), .A(n4422), .ZN(U3516) );
  MUX2_X1 U5009 ( .A(REG0_REG_29__SCAN_IN), .B(n4424), .S(n4706), .Z(U3515) );
  MUX2_X1 U5010 ( .A(REG0_REG_27__SCAN_IN), .B(n4425), .S(n4706), .Z(U3513) );
  INV_X1 U5011 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4427) );
  MUX2_X1 U5012 ( .A(n4427), .B(n4426), .S(n4706), .Z(n4428) );
  OAI21_X1 U5013 ( .B1(n4429), .B2(n4468), .A(n4428), .ZN(U3512) );
  INV_X1 U5014 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4431) );
  MUX2_X1 U5015 ( .A(n4431), .B(n4430), .S(n4706), .Z(n4432) );
  OAI21_X1 U5016 ( .B1(n4433), .B2(n4468), .A(n4432), .ZN(U3511) );
  MUX2_X1 U5017 ( .A(n4435), .B(n4434), .S(n4706), .Z(n4436) );
  OAI21_X1 U5018 ( .B1(n4437), .B2(n4468), .A(n4436), .ZN(U3510) );
  INV_X1 U5019 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4439) );
  MUX2_X1 U5020 ( .A(n4439), .B(n4438), .S(n4706), .Z(n4440) );
  OAI21_X1 U5021 ( .B1(n4441), .B2(n4468), .A(n4440), .ZN(U3509) );
  MUX2_X1 U5022 ( .A(REG0_REG_22__SCAN_IN), .B(n4442), .S(n4706), .Z(U3508) );
  INV_X1 U5023 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4444) );
  MUX2_X1 U5024 ( .A(n4444), .B(n4443), .S(n4706), .Z(n4445) );
  OAI21_X1 U5025 ( .B1(n4446), .B2(n4468), .A(n4445), .ZN(U3507) );
  INV_X1 U5026 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4448) );
  MUX2_X1 U5027 ( .A(n4448), .B(n4447), .S(n4706), .Z(n4449) );
  OAI21_X1 U5028 ( .B1(n4450), .B2(n4468), .A(n4449), .ZN(U3506) );
  INV_X1 U5029 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4452) );
  MUX2_X1 U5030 ( .A(n4452), .B(n4451), .S(n4706), .Z(n4453) );
  OAI21_X1 U5031 ( .B1(n4454), .B2(n4468), .A(n4453), .ZN(U3505) );
  MUX2_X1 U5032 ( .A(REG0_REG_18__SCAN_IN), .B(n4455), .S(n4706), .Z(U3503) );
  MUX2_X1 U5033 ( .A(n4457), .B(n4456), .S(n4706), .Z(n4458) );
  OAI21_X1 U5034 ( .B1(n4459), .B2(n4468), .A(n4458), .ZN(U3501) );
  MUX2_X1 U5035 ( .A(REG0_REG_16__SCAN_IN), .B(n4460), .S(n4706), .Z(U3499) );
  INV_X1 U5036 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4462) );
  MUX2_X1 U5037 ( .A(n4462), .B(n4461), .S(n4706), .Z(n4463) );
  OAI21_X1 U5038 ( .B1(n4464), .B2(n4468), .A(n4463), .ZN(U3497) );
  INV_X1 U5039 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4466) );
  MUX2_X1 U5040 ( .A(n4466), .B(n4465), .S(n4706), .Z(n4467) );
  OAI21_X1 U5041 ( .B1(n4469), .B2(n4468), .A(n4467), .ZN(U3495) );
  MUX2_X1 U5042 ( .A(DATAI_29_), .B(n4470), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U5043 ( .A(n4487), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5044 ( .A(n4471), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5045 ( .A(DATAI_20_), .B(n4472), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  INV_X1 U5046 ( .A(n4473), .ZN(n4474) );
  MUX2_X1 U5047 ( .A(DATAI_7_), .B(n4474), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5048 ( .A(n4475), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5049 ( .A(DATAI_4_), .B(n4497), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5050 ( .A(n4476), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5051 ( .A(DATAI_0_), .B(n4488), .S(STATE_REG_SCAN_IN), .Z(U3352) );
  INV_X1 U5052 ( .A(DATAI_28_), .ZN(n4477) );
  AOI22_X1 U5053 ( .A1(STATE_REG_SCAN_IN), .A2(n4478), .B1(n4477), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U5054 ( .A1(n4479), .A2(n4633), .B1(n4485), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4480) );
  OAI21_X1 U5055 ( .B1(n2922), .B2(n4481), .A(n4480), .ZN(U3260) );
  AOI22_X1 U5056 ( .A1(n4482), .A2(n4633), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4485), .ZN(n4483) );
  OAI21_X1 U5057 ( .B1(n4485), .B2(n4484), .A(n4483), .ZN(U3261) );
  OAI21_X1 U5058 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4487), .A(n4486), .ZN(n4489)
         );
  XOR2_X1 U5059 ( .A(n4489), .B(n4488), .Z(n4492) );
  AOI22_X1 U5060 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4599), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4490) );
  OAI21_X1 U5061 ( .B1(n4492), .B2(n4491), .A(n4490), .ZN(U3240) );
  XNOR2_X1 U5062 ( .A(n4493), .B(REG1_REG_4__SCAN_IN), .ZN(n4494) );
  NAND2_X1 U5063 ( .A1(n4607), .A2(n4494), .ZN(n4502) );
  XNOR2_X1 U5064 ( .A(n4495), .B(REG2_REG_4__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U5065 ( .A1(n4609), .A2(n4496), .ZN(n4501) );
  NAND2_X1 U5066 ( .A1(n4621), .A2(n4497), .ZN(n4500) );
  AOI21_X1 U5067 ( .B1(n4599), .B2(ADDR_REG_4__SCAN_IN), .A(n4498), .ZN(n4499)
         );
  AND4_X1 U5068 ( .A1(n4502), .A2(n4501), .A3(n4500), .A4(n4499), .ZN(n4504)
         );
  NAND2_X1 U5069 ( .A1(n4504), .A2(n4503), .ZN(U3244) );
  AOI211_X1 U5070 ( .C1(n4507), .C2(n4506), .A(n4505), .B(n4618), .ZN(n4510)
         );
  INV_X1 U5071 ( .A(n4508), .ZN(n4509) );
  AOI211_X1 U5072 ( .C1(n4599), .C2(ADDR_REG_8__SCAN_IN), .A(n4510), .B(n4509), 
        .ZN(n4514) );
  OAI211_X1 U5073 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4512), .A(n4609), .B(n4511), 
        .ZN(n4513) );
  OAI211_X1 U5074 ( .C1(n4612), .C2(n4662), .A(n4514), .B(n4513), .ZN(U3248)
         );
  AOI211_X1 U5075 ( .C1(n4517), .C2(n4516), .A(n4515), .B(n4618), .ZN(n4518)
         );
  AOI211_X1 U5076 ( .C1(n4599), .C2(ADDR_REG_9__SCAN_IN), .A(n4519), .B(n4518), 
        .ZN(n4524) );
  OAI211_X1 U5077 ( .C1(n4522), .C2(n4521), .A(n4609), .B(n4520), .ZN(n4523)
         );
  OAI211_X1 U5078 ( .C1(n4612), .C2(n4660), .A(n4524), .B(n4523), .ZN(U3249)
         );
  AOI211_X1 U5079 ( .C1(n4527), .C2(n4526), .A(n4525), .B(n4618), .ZN(n4530)
         );
  INV_X1 U5080 ( .A(n4528), .ZN(n4529) );
  AOI211_X1 U5081 ( .C1(n4599), .C2(ADDR_REG_10__SCAN_IN), .A(n4530), .B(n4529), .ZN(n4534) );
  OAI211_X1 U5082 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4532), .A(n4609), .B(n4531), .ZN(n4533) );
  OAI211_X1 U5083 ( .C1(n4612), .C2(n4658), .A(n4534), .B(n4533), .ZN(U3250)
         );
  AOI211_X1 U5084 ( .C1(n4537), .C2(n4536), .A(n4535), .B(n4618), .ZN(n4539)
         );
  AOI211_X1 U5085 ( .C1(n4599), .C2(ADDR_REG_11__SCAN_IN), .A(n4539), .B(n4538), .ZN(n4544) );
  OAI211_X1 U5086 ( .C1(n4542), .C2(n4541), .A(n4609), .B(n4540), .ZN(n4543)
         );
  OAI211_X1 U5087 ( .C1(n4612), .C2(n4656), .A(n4544), .B(n4543), .ZN(U3251)
         );
  AOI211_X1 U5088 ( .C1(n4547), .C2(n4546), .A(n4545), .B(n4618), .ZN(n4550)
         );
  INV_X1 U5089 ( .A(n4548), .ZN(n4549) );
  AOI211_X1 U5090 ( .C1(n4599), .C2(ADDR_REG_12__SCAN_IN), .A(n4550), .B(n4549), .ZN(n4554) );
  OAI211_X1 U5091 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4552), .A(n4609), .B(n4551), .ZN(n4553) );
  OAI211_X1 U5092 ( .C1(n4612), .C2(n4655), .A(n4554), .B(n4553), .ZN(U3252)
         );
  AOI211_X1 U5093 ( .C1(n4557), .C2(n4556), .A(n4555), .B(n4618), .ZN(n4558)
         );
  AOI211_X1 U5094 ( .C1(n4599), .C2(ADDR_REG_13__SCAN_IN), .A(n4559), .B(n4558), .ZN(n4565) );
  AOI21_X1 U5095 ( .B1(n3423), .B2(n4653), .A(n4560), .ZN(n4563) );
  AOI21_X1 U5096 ( .B1(n4563), .B2(n4562), .A(n4613), .ZN(n4561) );
  OAI21_X1 U5097 ( .B1(n4563), .B2(n4562), .A(n4561), .ZN(n4564) );
  OAI211_X1 U5098 ( .C1(n4612), .C2(n4653), .A(n4565), .B(n4564), .ZN(U3253)
         );
  INV_X1 U5099 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4576) );
  INV_X1 U5100 ( .A(n4599), .ZN(n4629) );
  AOI211_X1 U5101 ( .C1(n4567), .C2(n2518), .A(n4566), .B(n4613), .ZN(n4572)
         );
  AOI211_X1 U5102 ( .C1(n4570), .C2(n4569), .A(n4568), .B(n4618), .ZN(n4571)
         );
  AOI211_X1 U5103 ( .C1(n4621), .C2(n4573), .A(n4572), .B(n4571), .ZN(n4575)
         );
  OAI211_X1 U5104 ( .C1(n4576), .C2(n4629), .A(n4575), .B(n4574), .ZN(U3254)
         );
  AOI211_X1 U5105 ( .C1(n4579), .C2(n4578), .A(n4577), .B(n4613), .ZN(n4580)
         );
  AOI211_X1 U5106 ( .C1(n4599), .C2(ADDR_REG_15__SCAN_IN), .A(n4581), .B(n4580), .ZN(n4586) );
  AOI21_X1 U5107 ( .B1(n4583), .B2(n2043), .A(n4582), .ZN(n4584) );
  NAND2_X1 U5108 ( .A1(n4607), .A2(n4584), .ZN(n4585) );
  OAI211_X1 U5109 ( .C1(n4612), .C2(n4651), .A(n4586), .B(n4585), .ZN(U3255)
         );
  INV_X1 U5110 ( .A(n4587), .ZN(n4588) );
  AOI21_X1 U5111 ( .B1(ADDR_REG_16__SCAN_IN), .B2(n4599), .A(n4588), .ZN(n4597) );
  OAI21_X1 U5112 ( .B1(n4590), .B2(n2552), .A(n4589), .ZN(n4595) );
  OAI21_X1 U5113 ( .B1(n4593), .B2(n4592), .A(n4591), .ZN(n4594) );
  AOI22_X1 U5114 ( .A1(n4609), .A2(n4595), .B1(n4607), .B2(n4594), .ZN(n4596)
         );
  OAI211_X1 U5115 ( .C1(n4649), .C2(n4612), .A(n4597), .B(n4596), .ZN(U3256)
         );
  AOI21_X1 U5116 ( .B1(n4599), .B2(ADDR_REG_17__SCAN_IN), .A(n4598), .ZN(n4611) );
  OAI21_X1 U5117 ( .B1(n4602), .B2(n4601), .A(n4600), .ZN(n4608) );
  OAI21_X1 U5118 ( .B1(n4605), .B2(n4604), .A(n4603), .ZN(n4606) );
  AOI22_X1 U5119 ( .A1(n4609), .A2(n4608), .B1(n4607), .B2(n4606), .ZN(n4610)
         );
  OAI211_X1 U5120 ( .C1(n4647), .C2(n4612), .A(n4611), .B(n4610), .ZN(U3257)
         );
  INV_X1 U5121 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4630) );
  AOI211_X1 U5122 ( .C1(n4615), .C2(n4614), .A(n2049), .B(n4613), .ZN(n4626)
         );
  NAND2_X1 U5123 ( .A1(n4617), .A2(n4616), .ZN(n4619) );
  NAND2_X1 U5124 ( .A1(n4621), .A2(n4620), .ZN(n4622) );
  OAI211_X1 U5125 ( .C1(n4630), .C2(n4629), .A(n4628), .B(n4627), .ZN(U3258)
         );
  AOI22_X1 U5126 ( .A1(REG2_REG_2__SCAN_IN), .A2(n2922), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4631), .ZN(n4637) );
  AOI22_X1 U5127 ( .A1(n4635), .A2(n4634), .B1(n4633), .B2(n4632), .ZN(n4636)
         );
  OAI211_X1 U5128 ( .C1(n4485), .C2(n4638), .A(n4637), .B(n4636), .ZN(U3288)
         );
  AND2_X1 U5129 ( .A1(D_REG_31__SCAN_IN), .A2(n4641), .ZN(U3291) );
  AND2_X1 U5130 ( .A1(D_REG_30__SCAN_IN), .A2(n4641), .ZN(U3292) );
  AND2_X1 U5131 ( .A1(D_REG_29__SCAN_IN), .A2(n4641), .ZN(U3293) );
  AND2_X1 U5132 ( .A1(D_REG_28__SCAN_IN), .A2(n4641), .ZN(U3294) );
  AND2_X1 U5133 ( .A1(D_REG_27__SCAN_IN), .A2(n4641), .ZN(U3295) );
  AND2_X1 U5134 ( .A1(D_REG_26__SCAN_IN), .A2(n4641), .ZN(U3296) );
  AND2_X1 U5135 ( .A1(D_REG_25__SCAN_IN), .A2(n4641), .ZN(U3297) );
  AND2_X1 U5136 ( .A1(D_REG_24__SCAN_IN), .A2(n4641), .ZN(U3298) );
  AND2_X1 U5137 ( .A1(D_REG_23__SCAN_IN), .A2(n4641), .ZN(U3299) );
  AND2_X1 U5138 ( .A1(D_REG_22__SCAN_IN), .A2(n4641), .ZN(U3300) );
  AND2_X1 U5139 ( .A1(D_REG_21__SCAN_IN), .A2(n4641), .ZN(U3301) );
  AND2_X1 U5140 ( .A1(D_REG_20__SCAN_IN), .A2(n4641), .ZN(U3302) );
  AND2_X1 U5141 ( .A1(D_REG_19__SCAN_IN), .A2(n4641), .ZN(U3303) );
  AND2_X1 U5142 ( .A1(D_REG_18__SCAN_IN), .A2(n4641), .ZN(U3304) );
  INV_X1 U5143 ( .A(n4641), .ZN(n4643) );
  NOR2_X1 U5144 ( .A1(n4643), .A2(n4639), .ZN(U3305) );
  AND2_X1 U5145 ( .A1(D_REG_16__SCAN_IN), .A2(n4641), .ZN(U3306) );
  AND2_X1 U5146 ( .A1(D_REG_15__SCAN_IN), .A2(n4641), .ZN(U3307) );
  AND2_X1 U5147 ( .A1(D_REG_14__SCAN_IN), .A2(n4641), .ZN(U3308) );
  AND2_X1 U5148 ( .A1(D_REG_13__SCAN_IN), .A2(n4641), .ZN(U3309) );
  AND2_X1 U5149 ( .A1(D_REG_12__SCAN_IN), .A2(n4641), .ZN(U3310) );
  AND2_X1 U5150 ( .A1(D_REG_11__SCAN_IN), .A2(n4641), .ZN(U3311) );
  AND2_X1 U5151 ( .A1(D_REG_10__SCAN_IN), .A2(n4641), .ZN(U3312) );
  AND2_X1 U5152 ( .A1(D_REG_9__SCAN_IN), .A2(n4641), .ZN(U3313) );
  AND2_X1 U5153 ( .A1(D_REG_8__SCAN_IN), .A2(n4641), .ZN(U3314) );
  AND2_X1 U5154 ( .A1(D_REG_7__SCAN_IN), .A2(n4641), .ZN(U3315) );
  AND2_X1 U5155 ( .A1(D_REG_6__SCAN_IN), .A2(n4641), .ZN(U3316) );
  NOR2_X1 U5156 ( .A1(n4643), .A2(n4640), .ZN(U3317) );
  AND2_X1 U5157 ( .A1(D_REG_4__SCAN_IN), .A2(n4641), .ZN(U3318) );
  AND2_X1 U5158 ( .A1(D_REG_3__SCAN_IN), .A2(n4641), .ZN(U3319) );
  NOR2_X1 U5159 ( .A1(n4643), .A2(n4642), .ZN(U3320) );
  OAI21_X1 U5160 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4644), .ZN(
        n4645) );
  INV_X1 U5161 ( .A(n4645), .ZN(U3329) );
  AOI22_X1 U5162 ( .A1(STATE_REG_SCAN_IN), .A2(n4646), .B1(n2601), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5163 ( .A1(STATE_REG_SCAN_IN), .A2(n4647), .B1(n2586), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5164 ( .A1(STATE_REG_SCAN_IN), .A2(n4649), .B1(n4648), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5165 ( .A(DATAI_15_), .ZN(n4650) );
  AOI22_X1 U5166 ( .A1(STATE_REG_SCAN_IN), .A2(n4651), .B1(n4650), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5167 ( .A1(STATE_REG_SCAN_IN), .A2(n4653), .B1(n4652), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5168 ( .A1(STATE_REG_SCAN_IN), .A2(n4655), .B1(n4654), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5169 ( .A1(STATE_REG_SCAN_IN), .A2(n4656), .B1(n2475), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5170 ( .A(DATAI_10_), .ZN(n4657) );
  AOI22_X1 U5171 ( .A1(STATE_REG_SCAN_IN), .A2(n4658), .B1(n4657), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5172 ( .A(DATAI_9_), .ZN(n4659) );
  AOI22_X1 U5173 ( .A1(STATE_REG_SCAN_IN), .A2(n4660), .B1(n4659), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5174 ( .A1(STATE_REG_SCAN_IN), .A2(n4662), .B1(n4661), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5175 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4663) );
  AOI22_X1 U5176 ( .A1(n4706), .A2(n4664), .B1(n4663), .B2(n4704), .ZN(U3467)
         );
  AOI22_X1 U5177 ( .A1(n4706), .A2(n4666), .B1(n4665), .B2(n4704), .ZN(U3469)
         );
  AOI22_X1 U5178 ( .A1(n4668), .A2(n4676), .B1(n2899), .B2(n4667), .ZN(n4669)
         );
  AND2_X1 U5179 ( .A1(n4670), .A2(n4669), .ZN(n4708) );
  INV_X1 U5180 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4671) );
  AOI22_X1 U5181 ( .A1(n4706), .A2(n4708), .B1(n4671), .B2(n4704), .ZN(U3473)
         );
  INV_X1 U5182 ( .A(n4672), .ZN(n4677) );
  INV_X1 U5183 ( .A(n4673), .ZN(n4675) );
  AOI211_X1 U5184 ( .C1(n4677), .C2(n4676), .A(n4675), .B(n4674), .ZN(n4709)
         );
  AOI22_X1 U5185 ( .A1(n4706), .A2(n4709), .B1(n4678), .B2(n4704), .ZN(U3475)
         );
  NOR2_X1 U5186 ( .A1(n4679), .A2(n4685), .ZN(n4682) );
  INV_X1 U5187 ( .A(n4680), .ZN(n4681) );
  AOI22_X1 U5188 ( .A1(n4706), .A2(n4710), .B1(n4684), .B2(n4704), .ZN(U3477)
         );
  NOR2_X1 U5189 ( .A1(n4686), .A2(n4685), .ZN(n4690) );
  AOI211_X1 U5190 ( .C1(n4690), .C2(n4689), .A(n4688), .B(n4687), .ZN(n4712)
         );
  AOI22_X1 U5191 ( .A1(n4706), .A2(n4712), .B1(n4691), .B2(n4704), .ZN(U3481)
         );
  NAND2_X1 U5192 ( .A1(n4693), .A2(n4692), .ZN(n4696) );
  OR2_X1 U5193 ( .A1(n4694), .A2(n2269), .ZN(n4695) );
  INV_X1 U5194 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4698) );
  AOI22_X1 U5195 ( .A1(n4706), .A2(n4714), .B1(n4698), .B2(n4704), .ZN(U3485)
         );
  OAI22_X1 U5196 ( .A1(n4701), .A2(n4700), .B1(n2269), .B2(n4699), .ZN(n4702)
         );
  NOR2_X1 U5197 ( .A1(n4703), .A2(n4702), .ZN(n4717) );
  INV_X1 U5198 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5199 ( .A1(n4706), .A2(n4717), .B1(n4705), .B2(n4704), .ZN(U3489)
         );
  AOI22_X1 U5200 ( .A1(n4718), .A2(n4708), .B1(n4707), .B2(n4715), .ZN(U3521)
         );
  AOI22_X1 U5201 ( .A1(n4718), .A2(n4709), .B1(n2987), .B2(n4715), .ZN(U3522)
         );
  AOI22_X1 U5202 ( .A1(n4718), .A2(n4710), .B1(n2990), .B2(n4715), .ZN(U3523)
         );
  AOI22_X1 U5203 ( .A1(n4718), .A2(n4712), .B1(n4711), .B2(n4715), .ZN(U3525)
         );
  AOI22_X1 U5204 ( .A1(n4718), .A2(n4714), .B1(n4713), .B2(n4715), .ZN(U3527)
         );
  AOI22_X1 U5205 ( .A1(n4718), .A2(n4717), .B1(n4716), .B2(n4715), .ZN(U3529)
         );
  INV_X1 U2281 ( .A(IR_REG_31__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U2286 ( .A1(n3659), .A2(n2856), .ZN(n2855) );
  CLKBUF_X1 U2287 ( .A(n2363), .Z(n3725) );
  NAND2_X1 U2330 ( .A1(n2235), .A2(IR_REG_31__SCAN_IN), .ZN(n2237) );
  CLKBUF_X1 U2496 ( .A(n2380), .Z(n2381) );
  CLKBUF_X3 U2696 ( .A(n2309), .Z(n2786) );
endmodule

