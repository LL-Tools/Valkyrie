

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6427, n6428, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665;

  AND2_X1 U7175 ( .A1(n12592), .A2(n12591), .ZN(n15079) );
  INV_X1 U7176 ( .A(n15329), .ZN(n15057) );
  INV_X4 U7177 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U7178 ( .A1(n13770), .A2(n9080), .ZN(n13758) );
  NAND2_X1 U7179 ( .A1(n7485), .A2(n14844), .ZN(n14839) );
  NAND2_X1 U7180 ( .A1(n8456), .A2(n8455), .ZN(n13751) );
  INV_X1 U7181 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n15298) );
  NAND2_X1 U7182 ( .A1(n14322), .A2(n14321), .ZN(n14320) );
  INV_X1 U7183 ( .A(n14811), .ZN(n15087) );
  AND2_X1 U7184 ( .A1(n8332), .A2(n8331), .ZN(n14137) );
  AND2_X1 U7185 ( .A1(n8341), .A2(n8340), .ZN(n14133) );
  NAND2_X1 U7186 ( .A1(n7043), .A2(n15252), .ZN(n15030) );
  AND2_X1 U7187 ( .A1(n15191), .A2(n8843), .ZN(n15111) );
  NAND2_X1 U7188 ( .A1(n8909), .A2(n8908), .ZN(n15146) );
  BUF_X1 U7189 ( .A(n10632), .Z(n12569) );
  INV_X1 U7190 ( .A(n10720), .ZN(n9619) );
  INV_X2 U7191 ( .A(n12761), .ZN(n10074) );
  NAND2_X1 U7192 ( .A1(n14535), .A2(n14544), .ZN(n15365) );
  INV_X4 U7194 ( .A(n10632), .ZN(n13974) );
  AND2_X1 U7195 ( .A1(n12957), .A2(n12797), .ZN(n12930) );
  AND3_X1 U7196 ( .A1(n8850), .A2(n8849), .A3(n8848), .ZN(n11622) );
  INV_X1 U7197 ( .A(n9638), .ZN(n9288) );
  INV_X1 U7198 ( .A(n8843), .ZN(n10456) );
  NAND3_X1 U7199 ( .A1(n7913), .A2(n7912), .A3(n7911), .ZN(n12126) );
  NAND4_X2 U7200 ( .A1(n7924), .A2(n7923), .A3(n7922), .A4(n7921), .ZN(n13671)
         );
  INV_X1 U7201 ( .A(n9822), .ZN(n10165) );
  OR2_X1 U7202 ( .A1(n7967), .A2(n10415), .ZN(n7864) );
  CLKBUF_X2 U7203 ( .A(n7967), .Z(n8719) );
  INV_X1 U7204 ( .A(n8424), .ZN(n8282) );
  NAND2_X1 U7205 ( .A1(n9219), .A2(n11709), .ZN(n14387) );
  NAND2_X1 U7206 ( .A1(n10492), .A2(n7733), .ZN(n7967) );
  INV_X2 U7207 ( .A(n8018), .ZN(n7979) );
  NAND2_X1 U7208 ( .A1(n10492), .A2(n9755), .ZN(n7948) );
  NAND2_X1 U7209 ( .A1(n12404), .A2(n7879), .ZN(n8018) );
  NAND2_X1 U7210 ( .A1(n7842), .A2(n7843), .ZN(n7873) );
  INV_X1 U7211 ( .A(n15298), .ZN(n6427) );
  INV_X1 U7212 ( .A(n6427), .ZN(n6428) );
  INV_X1 U7213 ( .A(n6427), .ZN(P1_U3086) );
  INV_X2 U7214 ( .A(n8726), .ZN(n8770) );
  OAI21_X1 U7215 ( .B1(n13758), .B2(n7274), .A(n7273), .ZN(n13741) );
  INV_X1 U7216 ( .A(n10436), .ZN(n7733) );
  OAI21_X1 U7217 ( .B1(n7799), .B2(n6509), .A(n7189), .ZN(n13323) );
  INV_X1 U7218 ( .A(n12930), .ZN(n12946) );
  INV_X1 U7219 ( .A(n7019), .ZN(n6967) );
  NAND2_X1 U7220 ( .A1(n8493), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7870) );
  INV_X1 U7221 ( .A(n9648), .ZN(n9621) );
  INV_X1 U7222 ( .A(n9284), .ZN(n9644) );
  NOR2_X1 U7223 ( .A1(n14776), .A2(n14775), .ZN(n14777) );
  AND3_X1 U7224 ( .A1(n7236), .A2(n7235), .A3(n8844), .ZN(n8820) );
  INV_X1 U7225 ( .A(n14133), .ZN(n13831) );
  AND2_X1 U7226 ( .A1(n8199), .A2(n8198), .ZN(n13941) );
  BUF_X1 U7227 ( .A(n7956), .Z(n8279) );
  INV_X1 U7228 ( .A(n12038), .ZN(n11318) );
  OAI21_X1 U7229 ( .B1(n14320), .B2(n6704), .A(n6702), .ZN(n6705) );
  NOR2_X1 U7230 ( .A1(n7045), .A2(n9610), .ZN(n14363) );
  BUF_X1 U7231 ( .A(n9463), .Z(n6433) );
  AND2_X1 U7232 ( .A1(n8858), .A2(n8857), .ZN(n11635) );
  INV_X1 U7233 ( .A(n14958), .ZN(n14381) );
  INV_X1 U7234 ( .A(n11999), .ZN(n15552) );
  NAND2_X1 U7235 ( .A1(n8479), .A2(n8478), .ZN(n13720) );
  INV_X1 U7236 ( .A(n13901), .ZN(n14064) );
  CLKBUF_X3 U7237 ( .A(n7980), .Z(n8424) );
  INV_X1 U7238 ( .A(n13541), .ZN(n14129) );
  NAND2_X1 U7239 ( .A1(n8305), .A2(n8304), .ZN(n14140) );
  INV_X1 U7240 ( .A(n15365), .ZN(n15333) );
  INV_X1 U7241 ( .A(n9728), .ZN(n13507) );
  AND2_X1 U7242 ( .A1(n8074), .A2(n8073), .ZN(n12110) );
  NAND2_X1 U7243 ( .A1(n7947), .A2(n6488), .ZN(n13670) );
  INV_X2 U7244 ( .A(n13909), .ZN(n13987) );
  INV_X1 U7245 ( .A(n13955), .ZN(n7172) );
  NAND2_X1 U7246 ( .A1(n7851), .A2(n7852), .ZN(n14181) );
  NAND4_X1 U7247 ( .A1(n9280), .A2(n9279), .A3(n9278), .A4(n9277), .ZN(n14651)
         );
  XNOR2_X1 U7248 ( .A(n6982), .B(n14610), .ZN(n15073) );
  INV_X2 U7249 ( .A(n15049), .ZN(n15340) );
  AND2_X1 U7250 ( .A1(n9249), .A2(n9248), .ZN(n6430) );
  AND2_X2 U7251 ( .A1(n13761), .A2(n7407), .ZN(n6431) );
  NAND2_X2 U7252 ( .A1(n9119), .A2(n6943), .ZN(n9122) );
  NAND2_X2 U7253 ( .A1(n14738), .A2(n14737), .ZN(n14736) );
  INV_X2 U7254 ( .A(n14467), .ZN(n14541) );
  NAND2_X2 U7255 ( .A1(n13964), .A2(n9063), .ZN(n13948) );
  NAND2_X2 U7256 ( .A1(n6643), .A2(n7755), .ZN(n13964) );
  NAND2_X2 U7257 ( .A1(n6798), .A2(n11682), .ZN(n11926) );
  XNOR2_X2 U7258 ( .A(n12837), .B(n11767), .ZN(n12835) );
  OAI211_X2 U7259 ( .C1(n7059), .C2(n7058), .A(n6465), .B(n7057), .ZN(n11919)
         );
  BUF_X2 U7260 ( .A(n8582), .Z(n6432) );
  BUF_X2 U7261 ( .A(n9463), .Z(n6434) );
  NAND2_X1 U7262 ( .A1(n9220), .A2(n8965), .ZN(n9463) );
  OAI21_X4 U7263 ( .B1(n8830), .B2(n7297), .A(n7295), .ZN(n14654) );
  AND2_X4 U7264 ( .A1(n9634), .A2(n15365), .ZN(n9648) );
  AOI21_X2 U7265 ( .B1(n13981), .B2(n13982), .A(n6540), .ZN(n7812) );
  OAI21_X2 U7266 ( .B1(n12305), .B2(n9027), .A(n9026), .ZN(n13981) );
  INV_X8 U7267 ( .A(n7859), .ZN(n10436) );
  XNOR2_X2 U7268 ( .A(n7870), .B(n8494), .ZN(n9039) );
  NAND2_X1 U7269 ( .A1(n7068), .A2(n7072), .ZN(n7067) );
  AOI21_X2 U7270 ( .B1(n7805), .B2(n7804), .A(n6491), .ZN(n13210) );
  NAND2_X1 U7271 ( .A1(n8944), .A2(n8943), .ZN(n15077) );
  NAND2_X1 U7272 ( .A1(n9034), .A2(n9033), .ZN(n13852) );
  NAND2_X1 U7273 ( .A1(n8942), .A2(n8941), .ZN(n15082) );
  NAND2_X1 U7274 ( .A1(n14892), .A2(n14878), .ZN(n14855) );
  NAND2_X1 U7275 ( .A1(n8930), .A2(n8929), .ZN(n14889) );
  INV_X1 U7276 ( .A(n13742), .ZN(n13723) );
  OAI21_X1 U7277 ( .B1(n11760), .B2(n7712), .A(n7709), .ZN(n12150) );
  NAND2_X1 U7278 ( .A1(n8891), .A2(n8890), .ZN(n15230) );
  NAND2_X1 U7279 ( .A1(n6435), .A2(n12046), .ZN(n12041) );
  AND2_X1 U7280 ( .A1(n8040), .A2(n8039), .ZN(n11984) );
  XNOR2_X1 U7281 ( .A(n9893), .B(n12843), .ZN(n12139) );
  NAND2_X1 U7282 ( .A1(n9846), .A2(n9845), .ZN(n12842) );
  INV_X2 U7283 ( .A(n15583), .ZN(n9757) );
  AND3_X1 U7284 ( .A1(n9766), .A2(n9765), .A3(n9764), .ZN(n15573) );
  INV_X1 U7285 ( .A(n13668), .ZN(n11312) );
  NAND4_X2 U7286 ( .A1(n9294), .A2(n9293), .A3(n9292), .A4(n9291), .ZN(n14650)
         );
  INV_X1 U7287 ( .A(n11629), .ZN(n14399) );
  OR2_X1 U7288 ( .A1(n11370), .A2(n11453), .ZN(n15332) );
  BUF_X2 U7289 ( .A(n9903), .Z(n12758) );
  INV_X2 U7290 ( .A(n8571), .ZN(n12056) );
  AOI21_X1 U7291 ( .B1(n10074), .B2(SI_8_), .A(n6958), .ZN(n9845) );
  NAND2_X1 U7292 ( .A1(n6979), .A2(n7987), .ZN(n13669) );
  NAND2_X4 U7293 ( .A1(n10911), .A2(n10436), .ZN(n12761) );
  INV_X2 U7294 ( .A(n8965), .ZN(n15181) );
  INV_X2 U7295 ( .A(n7019), .ZN(n7920) );
  XNOR2_X1 U7296 ( .A(n7869), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8776) );
  AND4_X1 U7297 ( .A1(n8831), .A2(n6698), .A3(n6697), .A4(n6641), .ZN(n6442)
         );
  NAND2_X1 U7298 ( .A1(n6725), .A2(n7417), .ZN(n14551) );
  MUX2_X1 U7299 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15156), .S(n15420), .Z(
        P1_U3557) );
  NAND2_X1 U7300 ( .A1(n6897), .A2(n7356), .ZN(n8775) );
  OAI211_X1 U7301 ( .C1(n15325), .C2(n15073), .A(n7055), .B(n6796), .ZN(n15156) );
  AOI21_X1 U7302 ( .B1(n9217), .B2(n15561), .A(n9216), .ZN(n9218) );
  NAND2_X1 U7303 ( .A1(n13590), .A2(n8409), .ZN(n13565) );
  NOR3_X1 U7304 ( .A1(n14612), .A2(n14611), .A3(n14610), .ZN(n14613) );
  NAND2_X1 U7305 ( .A1(n7248), .A2(n6919), .ZN(n12588) );
  OAI21_X1 U7306 ( .B1(n8656), .B2(n7640), .A(n7638), .ZN(n8661) );
  NAND2_X1 U7307 ( .A1(n14812), .A2(n14830), .ZN(n15092) );
  NAND2_X1 U7308 ( .A1(n7067), .A2(n6536), .ZN(n12602) );
  NAND2_X1 U7309 ( .A1(n7074), .A2(n7752), .ZN(n14832) );
  NAND2_X1 U7310 ( .A1(n13801), .A2(n9037), .ZN(n13769) );
  AND2_X1 U7311 ( .A1(n7247), .A2(n14605), .ZN(n6919) );
  NOR2_X1 U7312 ( .A1(n7364), .A2(n10381), .ZN(n7363) );
  AND2_X1 U7313 ( .A1(n14753), .A2(n14754), .ZN(n14764) );
  NAND2_X1 U7314 ( .A1(n7662), .A2(n6534), .ZN(n13801) );
  NAND2_X1 U7315 ( .A1(n7420), .A2(n10162), .ZN(n7419) );
  XNOR2_X1 U7316 ( .A(n14016), .B(n13653), .ZN(n14011) );
  XNOR2_X1 U7317 ( .A(n14550), .B(n14548), .ZN(n14610) );
  NOR2_X1 U7318 ( .A1(n13720), .A2(n13751), .ZN(n7407) );
  NAND2_X1 U7319 ( .A1(n14869), .A2(n14880), .ZN(n14868) );
  NAND2_X1 U7320 ( .A1(n6473), .A2(n12353), .ZN(n14751) );
  AND2_X1 U7321 ( .A1(n13602), .A2(n13601), .ZN(n8358) );
  OAI21_X1 U7322 ( .B1(n12491), .B2(n12490), .A(n12492), .ZN(n12538) );
  CLKBUF_X1 U7323 ( .A(n13286), .Z(n6925) );
  XNOR2_X1 U7324 ( .A(n8683), .B(n8682), .ZN(n14176) );
  OAI21_X1 U7325 ( .B1(n10292), .B2(n10291), .A(n10293), .ZN(n12491) );
  CLKBUF_X1 U7326 ( .A(n13584), .Z(n6993) );
  NAND2_X1 U7327 ( .A1(n14954), .A2(n12415), .ZN(n7623) );
  AND2_X1 U7328 ( .A1(n6814), .A2(n6813), .ZN(n15279) );
  NAND2_X2 U7329 ( .A1(n8934), .A2(n8933), .ZN(n15104) );
  XNOR2_X1 U7330 ( .A(n8473), .B(n8454), .ZN(n14180) );
  NAND2_X1 U7331 ( .A1(n6877), .A2(n10267), .ZN(n10274) );
  AND2_X1 U7332 ( .A1(n12983), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U7333 ( .A1(n8936), .A2(n8935), .ZN(n14838) );
  NAND2_X1 U7334 ( .A1(n8398), .A2(n8397), .ZN(n14036) );
  NAND2_X1 U7335 ( .A1(n9595), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U7336 ( .A1(n8414), .A2(n6525), .ZN(n6831) );
  NAND2_X1 U7337 ( .A1(n6735), .A2(n8926), .ZN(n15128) );
  NAND2_X2 U7338 ( .A1(n8928), .A2(n8927), .ZN(n15122) );
  AND2_X1 U7339 ( .A1(n8261), .A2(n8260), .ZN(n13901) );
  NAND2_X1 U7340 ( .A1(n8922), .A2(n8921), .ZN(n15131) );
  NAND2_X1 U7341 ( .A1(n7373), .A2(n6501), .ZN(n12257) );
  NAND2_X1 U7342 ( .A1(n6915), .A2(n10143), .ZN(n10156) );
  XNOR2_X1 U7343 ( .A(n8389), .B(SI_22_), .ZN(n8931) );
  CLKBUF_X1 U7344 ( .A(n11760), .Z(n7014) );
  XNOR2_X1 U7345 ( .A(n15151), .B(n15026), .ZN(n15011) );
  INV_X1 U7346 ( .A(n13941), .ZN(n14074) );
  NAND2_X1 U7347 ( .A1(n7173), .A2(n8220), .ZN(n13955) );
  NAND2_X1 U7348 ( .A1(n7397), .A2(n14161), .ZN(n12281) );
  AND2_X1 U7349 ( .A1(n8126), .A2(n8125), .ZN(n12282) );
  INV_X1 U7350 ( .A(n11962), .ZN(n7397) );
  NAND2_X1 U7351 ( .A1(n8429), .A2(n8428), .ZN(n13795) );
  XNOR2_X1 U7352 ( .A(n8230), .B(n8229), .ZN(n11297) );
  AND2_X1 U7353 ( .A1(n11741), .A2(n6700), .ZN(n6699) );
  OAI21_X1 U7354 ( .B1(n10936), .B2(n6756), .A(n6754), .ZN(n11061) );
  NAND2_X1 U7355 ( .A1(n8887), .A2(n8886), .ZN(n14438) );
  NAND2_X1 U7356 ( .A1(n8252), .A2(n8251), .ZN(n8230) );
  NAND2_X1 U7357 ( .A1(n8145), .A2(n8144), .ZN(n8162) );
  NOR2_X1 U7358 ( .A1(n8540), .A2(n8777), .ZN(n13643) );
  OR2_X1 U7359 ( .A1(n8093), .A2(n8092), .ZN(n8115) );
  NAND2_X1 U7360 ( .A1(n15321), .A2(n11373), .ZN(n11633) );
  OAI21_X1 U7361 ( .B1(n9128), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9111), .ZN(
        n9156) );
  NAND2_X1 U7362 ( .A1(n8122), .A2(n8121), .ZN(n7187) );
  OAI21_X1 U7363 ( .B1(n14385), .B2(n14389), .A(n14391), .ZN(n15324) );
  AND2_X1 U7364 ( .A1(n8053), .A2(n8052), .ZN(n12015) );
  NAND2_X1 U7365 ( .A1(n8088), .A2(n8087), .ZN(n8122) );
  NAND2_X1 U7366 ( .A1(n8871), .A2(n8870), .ZN(n14424) );
  NOR2_X2 U7367 ( .A1(n12506), .A2(n14381), .ZN(n15235) );
  AND2_X1 U7368 ( .A1(n9286), .A2(n9285), .ZN(n11519) );
  INV_X1 U7369 ( .A(n12043), .ZN(n6435) );
  AOI21_X2 U7370 ( .B1(n10432), .B2(n7976), .A(n8017), .ZN(n11999) );
  INV_X2 U7371 ( .A(n12487), .ZN(n12496) );
  INV_X1 U7372 ( .A(n11635), .ZN(n15355) );
  NAND2_X1 U7373 ( .A1(n7170), .A2(n8071), .ZN(n8088) );
  NAND2_X1 U7374 ( .A1(n7978), .A2(n7977), .ZN(n12038) );
  AND2_X1 U7375 ( .A1(n9004), .A2(n11249), .ZN(n9005) );
  INV_X1 U7376 ( .A(n11336), .ZN(n6436) );
  INV_X1 U7377 ( .A(n12773), .ZN(n6437) );
  NAND4_X1 U7378 ( .A1(n9750), .A2(n9749), .A3(n9748), .A4(n9747), .ZN(n15596)
         );
  AND2_X1 U7379 ( .A1(n11248), .A2(n8791), .ZN(n11241) );
  NAND2_X2 U7380 ( .A1(n9834), .A2(n9833), .ZN(n12977) );
  AND3_X1 U7381 ( .A1(n9870), .A2(n9869), .A3(n9868), .ZN(n11767) );
  NAND2_X1 U7382 ( .A1(n7052), .A2(n7050), .ZN(n15330) );
  NAND2_X1 U7383 ( .A1(n6780), .A2(n9267), .ZN(n14652) );
  CLKBUF_X1 U7384 ( .A(n12269), .Z(n12101) );
  AND4_X1 U7385 ( .A1(n9234), .A2(n9233), .A3(n9232), .A4(n9231), .ZN(n11948)
         );
  NAND2_X1 U7386 ( .A1(n8007), .A2(n6964), .ZN(n13668) );
  OR2_X1 U7387 ( .A1(n11251), .A2(n12126), .ZN(n8791) );
  AND2_X1 U7388 ( .A1(n9831), .A2(n7825), .ZN(n9834) );
  AND2_X1 U7389 ( .A1(n8983), .A2(n8982), .ZN(n6710) );
  NAND4_X2 U7390 ( .A1(n9262), .A2(n9261), .A3(n9260), .A4(n9259), .ZN(n11381)
         );
  OAI211_X1 U7391 ( .C1(n8843), .C2(n10616), .A(n8842), .B(n8841), .ZN(n11629)
         );
  NAND2_X1 U7392 ( .A1(n7889), .A2(n7890), .ZN(n13673) );
  OAI21_X1 U7393 ( .B1(n7973), .B2(n7167), .A(n6551), .ZN(n6980) );
  AND4_X1 U7394 ( .A1(n8061), .A2(n8060), .A3(n8059), .A4(n8058), .ZN(n11702)
         );
  NAND2_X2 U7395 ( .A1(n14383), .A2(n14387), .ZN(n10720) );
  INV_X1 U7396 ( .A(n12797), .ZN(n6928) );
  BUF_X2 U7397 ( .A(n7976), .Z(n8718) );
  CLKBUF_X1 U7398 ( .A(n8949), .Z(n6952) );
  INV_X1 U7399 ( .A(n9723), .ZN(n10301) );
  AND4_X2 U7400 ( .A1(n7902), .A2(n6966), .A3(n7901), .A4(n7903), .ZN(n11251)
         );
  NAND2_X1 U7401 ( .A1(n8843), .A2(n7733), .ZN(n8859) );
  CLKBUF_X1 U7402 ( .A(n9826), .Z(n6957) );
  OAI21_X1 U7403 ( .B1(n8976), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8975) );
  NAND2_X1 U7404 ( .A1(n15190), .A2(n14958), .ZN(n14383) );
  AND2_X2 U7405 ( .A1(n13896), .A2(n8779), .ZN(n7940) );
  INV_X2 U7406 ( .A(n9826), .ZN(n12093) );
  NAND2_X1 U7407 ( .A1(n7920), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7922) );
  CLKBUF_X1 U7408 ( .A(n10911), .Z(n6924) );
  INV_X2 U7409 ( .A(n8002), .ZN(n8708) );
  INV_X1 U7410 ( .A(n14575), .ZN(n15190) );
  INV_X1 U7411 ( .A(n9725), .ZN(n7790) );
  CLKBUF_X2 U7412 ( .A(n8964), .Z(n12468) );
  NAND2_X1 U7413 ( .A1(n7880), .A2(n7879), .ZN(n7980) );
  NAND2_X1 U7414 ( .A1(n9687), .A2(n9689), .ZN(n10200) );
  AOI21_X1 U7415 ( .B1(n8046), .B2(n8037), .A(n8069), .ZN(n7340) );
  XNOR2_X1 U7416 ( .A(n9721), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9725) );
  INV_X1 U7417 ( .A(n13134), .ZN(n13517) );
  XNOR2_X1 U7418 ( .A(n8963), .B(n15173), .ZN(n8964) );
  NAND2_X1 U7419 ( .A1(n15172), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8963) );
  XNOR2_X1 U7420 ( .A(n8036), .B(SI_8_), .ZN(n8046) );
  NAND2_X1 U7421 ( .A1(n7244), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7243) );
  NAND2_X1 U7422 ( .A1(n7330), .A2(n8837), .ZN(n7934) );
  NAND2_X1 U7423 ( .A1(n9722), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7153) );
  XNOR2_X1 U7424 ( .A(n8957), .B(n8956), .ZN(n11709) );
  INV_X2 U7425 ( .A(n14175), .ZN(n6438) );
  AND2_X1 U7426 ( .A1(n6442), .A2(n6451), .ZN(n8954) );
  XNOR2_X1 U7427 ( .A(n7872), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13705) );
  NAND2_X1 U7428 ( .A1(n8923), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8924) );
  OR2_X1 U7429 ( .A1(n9734), .A2(n13502), .ZN(n6753) );
  OAI21_X1 U7430 ( .B1(n8958), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8959) );
  XNOR2_X1 U7431 ( .A(n9797), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10979) );
  AND3_X1 U7432 ( .A1(n6790), .A2(n7233), .A3(n6789), .ZN(n8828) );
  NAND2_X1 U7433 ( .A1(n7853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7854) );
  OR2_X1 U7434 ( .A1(n10001), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n10021) );
  OAI21_X1 U7435 ( .B1(n7871), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7868) );
  INV_X4 U7436 ( .A(n7955), .ZN(n7859) );
  AND4_X1 U7437 ( .A1(n7232), .A2(n6791), .A3(n7660), .A4(n8823), .ZN(n6790)
         );
  NAND2_X1 U7438 ( .A1(n8839), .A2(n8838), .ZN(n14675) );
  OR2_X1 U7439 ( .A1(n8057), .A2(n10669), .ZN(n8076) );
  OR2_X1 U7440 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10896), .ZN(n10897) );
  NOR2_X1 U7441 ( .A1(n7849), .A2(n6910), .ZN(n6909) );
  AND2_X1 U7442 ( .A1(n8820), .A2(n7474), .ZN(n7379) );
  AND3_X1 U7443 ( .A1(n8904), .A2(n6474), .A3(n8820), .ZN(n6789) );
  AND3_X2 U7444 ( .A1(n7867), .A2(n7841), .A3(n7866), .ZN(n7842) );
  XNOR2_X1 U7445 ( .A(n6830), .B(n9775), .ZN(n10943) );
  NAND4_X1 U7446 ( .A1(n14790), .A2(n7856), .A3(n7855), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7168) );
  NAND2_X1 U7447 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n8824), .ZN(n7486) );
  AND2_X1 U7448 ( .A1(n7080), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9135) );
  AND2_X1 U7449 ( .A1(n8819), .A2(n8882), .ZN(n8904) );
  AND2_X1 U7450 ( .A1(n7239), .A2(n8854), .ZN(n7231) );
  NAND4_X1 U7451 ( .A1(n7332), .A2(n7331), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7169) );
  NAND4_X1 U7452 ( .A1(n10223), .A2(n9689), .A3(n7105), .A4(n7104), .ZN(n9690)
         );
  AND3_X1 U7453 ( .A1(n9763), .A2(n9679), .A3(n9678), .ZN(n9683) );
  NAND2_X1 U7454 ( .A1(n9693), .A2(n9692), .ZN(n9694) );
  NOR2_X1 U7455 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8819) );
  NOR2_X1 U7456 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n9678) );
  NOR2_X1 U7457 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n9679) );
  INV_X1 U7458 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8885) );
  NOR2_X1 U7459 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8882) );
  NOR2_X1 U7460 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7234) );
  NOR2_X1 U7461 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7260) );
  NOR2_X1 U7462 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n9681) );
  NOR2_X1 U7463 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7259) );
  NOR2_X1 U7464 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n7261) );
  NOR2_X2 U7465 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n9686) );
  INV_X1 U7466 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9689) );
  NAND3_X1 U7467 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n8003) );
  INV_X1 U7468 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8516) );
  INV_X1 U7469 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7396) );
  INV_X4 U7470 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7471 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7856) );
  BUF_X1 U7472 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n15193) );
  XNOR2_X1 U7473 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n9132) );
  OAI21_X2 U7474 ( .B1(n7222), .B2(n14986), .A(n7219), .ZN(n14969) );
  NAND2_X1 U7475 ( .A1(n15003), .A2(n15011), .ZN(n7222) );
  NAND4_X2 U7476 ( .A1(n7400), .A2(n14146), .A3(n7172), .A4(n13941), .ZN(
        n13917) );
  NOR2_X4 U7477 ( .A1(n15030), .A2(n15151), .ZN(n15006) );
  NAND2_X1 U7478 ( .A1(n15181), .A2(n12468), .ZN(n6439) );
  NAND2_X1 U7479 ( .A1(n15181), .A2(n12468), .ZN(n6440) );
  AOI21_X2 U7480 ( .B1(n15021), .B2(n12413), .A(n12412), .ZN(n15003) );
  INV_X4 U7481 ( .A(n9604), .ZN(n9634) );
  NAND4_X2 U7482 ( .A1(n9242), .A2(n9241), .A3(n9240), .A4(n9239), .ZN(n11380)
         );
  INV_X1 U7483 ( .A(n12461), .ZN(n7073) );
  NAND2_X1 U7484 ( .A1(n8654), .A2(n8655), .ZN(n7646) );
  AND2_X1 U7485 ( .A1(n8793), .A2(n9049), .ZN(n9043) );
  NAND2_X1 U7486 ( .A1(n9725), .A2(n9728), .ZN(n9826) );
  NOR2_X1 U7487 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n9703) );
  NAND2_X1 U7488 ( .A1(n9686), .A2(n9680), .ZN(n7683) );
  NOR2_X1 U7489 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n9680) );
  OR2_X1 U7490 ( .A1(n14811), .A2(n9284), .ZN(n9607) );
  OR2_X1 U7491 ( .A1(n9636), .A2(n9635), .ZN(n9657) );
  AOI21_X1 U7492 ( .B1(n7753), .B2(n14863), .A(n6548), .ZN(n7752) );
  NOR2_X1 U7493 ( .A1(n14846), .A2(n7754), .ZN(n7753) );
  INV_X1 U7494 ( .A(n12457), .ZN(n7754) );
  INV_X1 U7495 ( .A(n14846), .ZN(n7632) );
  NAND2_X1 U7496 ( .A1(n7630), .A2(n7634), .ZN(n14847) );
  INV_X1 U7497 ( .A(n9716), .ZN(n9718) );
  OAI21_X1 U7498 ( .B1(n10369), .B2(n6927), .A(n6926), .ZN(n9716) );
  NAND2_X1 U7499 ( .A1(n11540), .A2(n12797), .ZN(n6926) );
  OR2_X1 U7500 ( .A1(n12404), .A2(n7879), .ZN(n7943) );
  INV_X1 U7501 ( .A(n7666), .ZN(n7665) );
  OAI21_X1 U7502 ( .B1(n13737), .B2(n7667), .A(n7669), .ZN(n7666) );
  NAND2_X1 U7503 ( .A1(n7681), .A2(n7680), .ZN(n9034) );
  AND2_X1 U7504 ( .A1(n7838), .A2(n9032), .ZN(n7680) );
  AND2_X1 U7505 ( .A1(n14527), .A2(n6590), .ZN(n6734) );
  OAI21_X1 U7506 ( .B1(n14525), .B2(n7468), .A(n7465), .ZN(n14527) );
  NAND2_X1 U7507 ( .A1(n8946), .A2(n8945), .ZN(n14550) );
  NOR2_X1 U7508 ( .A1(n14972), .A2(n7220), .ZN(n7219) );
  INV_X1 U7509 ( .A(n14466), .ZN(n7221) );
  NAND2_X2 U7510 ( .A1(n8843), .A2(n10436), .ZN(n8949) );
  OAI22_X1 U7511 ( .A1(n15279), .A2(n6450), .B1(P2_ADDR_REG_14__SCAN_IN), .B2(
        n15278), .ZN(n7601) );
  OAI211_X1 U7512 ( .C1(n14394), .C2(n7436), .A(n6951), .B(n14402), .ZN(n14407) );
  NAND2_X1 U7513 ( .A1(n8594), .A2(n8593), .ZN(n6929) );
  INV_X1 U7514 ( .A(n8595), .ZN(n6931) );
  NAND2_X1 U7515 ( .A1(n14421), .A2(n14420), .ZN(n6718) );
  AOI21_X1 U7516 ( .B1(n7479), .B2(n7478), .A(n7476), .ZN(n7475) );
  INV_X1 U7517 ( .A(n12818), .ZN(n7128) );
  NAND2_X1 U7518 ( .A1(n6953), .A2(n7440), .ZN(n7439) );
  OAI22_X1 U7519 ( .A1(n12282), .A2(n8650), .B1(n12295), .B2(n8726), .ZN(n8624) );
  NAND2_X1 U7520 ( .A1(n6553), .A2(n7138), .ZN(n7137) );
  NAND2_X1 U7521 ( .A1(n7138), .A2(n12917), .ZN(n7136) );
  NAND2_X1 U7522 ( .A1(n6903), .A2(n8652), .ZN(n6902) );
  INV_X1 U7523 ( .A(n7646), .ZN(n7644) );
  NAND2_X1 U7524 ( .A1(n8653), .A2(n7648), .ZN(n7647) );
  INV_X1 U7525 ( .A(n8655), .ZN(n7648) );
  INV_X1 U7526 ( .A(n8658), .ZN(n7645) );
  INV_X1 U7527 ( .A(n7353), .ZN(n7352) );
  OAI21_X1 U7528 ( .B1(n7355), .B2(n7354), .A(n8388), .ZN(n7353) );
  OR2_X1 U7529 ( .A1(n10195), .A2(n10194), .ZN(n10196) );
  OR2_X1 U7530 ( .A1(n12665), .A2(n12383), .ZN(n12865) );
  INV_X1 U7531 ( .A(n9862), .ZN(n6865) );
  INV_X1 U7532 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U7533 ( .A1(n6715), .A2(n14544), .ZN(n7457) );
  INV_X1 U7534 ( .A(n14543), .ZN(n6715) );
  NAND2_X1 U7535 ( .A1(n7635), .A2(n6481), .ZN(n7634) );
  INV_X1 U7536 ( .A(n14863), .ZN(n7635) );
  NOR2_X1 U7537 ( .A1(n8214), .A2(n8188), .ZN(n8189) );
  NAND2_X1 U7538 ( .A1(n8184), .A2(n10629), .ZN(n8251) );
  NAND2_X1 U7539 ( .A1(n8112), .A2(n10478), .ZN(n8140) );
  AND2_X1 U7540 ( .A1(n10280), .A2(n10279), .ZN(n10298) );
  XNOR2_X1 U7541 ( .A(n10259), .B(n15573), .ZN(n12809) );
  OR2_X1 U7542 ( .A1(n12556), .A2(n13176), .ZN(n12948) );
  AOI21_X1 U7543 ( .B1(n13210), .B2(n7205), .A(n7203), .ZN(n13172) );
  AND2_X1 U7544 ( .A1(n10346), .A2(n7207), .ZN(n7205) );
  NAND2_X1 U7545 ( .A1(n7204), .A2(n6545), .ZN(n7203) );
  NAND2_X1 U7546 ( .A1(n6850), .A2(n13193), .ZN(n12937) );
  NAND2_X1 U7547 ( .A1(n7715), .A2(n7713), .ZN(n7712) );
  INV_X1 U7548 ( .A(n12849), .ZN(n7713) );
  NAND2_X1 U7549 ( .A1(n9711), .A2(n9710), .ZN(n10204) );
  NAND2_X1 U7550 ( .A1(n9707), .A2(n12293), .ZN(n9711) );
  AOI21_X1 U7551 ( .B1(n7569), .B2(n7571), .A(n10035), .ZN(n7568) );
  INV_X1 U7552 ( .A(n10016), .ZN(n7569) );
  INV_X1 U7553 ( .A(n7571), .ZN(n7570) );
  INV_X1 U7554 ( .A(n7590), .ZN(n7589) );
  OAI21_X1 U7555 ( .B1(n9793), .B2(n7591), .A(n9835), .ZN(n7590) );
  INV_X1 U7556 ( .A(n8139), .ZN(n7562) );
  INV_X1 U7557 ( .A(n10528), .ZN(n6663) );
  NOR2_X1 U7558 ( .A1(n6494), .A2(n6938), .ZN(n13686) );
  AND2_X1 U7559 ( .A1(n15518), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U7560 ( .A1(n8434), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8459) );
  INV_X1 U7561 ( .A(n8436), .ZN(n8434) );
  OR2_X1 U7562 ( .A1(n13831), .A2(n13843), .ZN(n13790) );
  NAND2_X1 U7563 ( .A1(n9043), .A2(n9047), .ZN(n9048) );
  NAND2_X1 U7564 ( .A1(n6777), .A2(n6772), .ZN(n6771) );
  NOR2_X1 U7565 ( .A1(n6475), .A2(n6773), .ZN(n6772) );
  INV_X1 U7566 ( .A(n6775), .ZN(n6773) );
  NOR2_X1 U7567 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7525) );
  NOR2_X1 U7568 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7524) );
  AND3_X2 U7569 ( .A1(n6686), .A2(n7523), .A3(n7396), .ZN(n7910) );
  INV_X1 U7570 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U7571 ( .A1(n6556), .A2(n15070), .ZN(n7489) );
  OR2_X1 U7572 ( .A1(n15077), .A2(n14637), .ZN(n12523) );
  NAND2_X1 U7573 ( .A1(n15077), .A2(n14637), .ZN(n12526) );
  INV_X1 U7574 ( .A(n9596), .ZN(n9595) );
  NOR2_X1 U7575 ( .A1(n14886), .A2(n7748), .ZN(n7747) );
  INV_X1 U7576 ( .A(n14476), .ZN(n7748) );
  OR2_X1 U7577 ( .A1(n15128), .A2(n14944), .ZN(n14474) );
  NAND2_X1 U7578 ( .A1(n15128), .A2(n14944), .ZN(n14475) );
  AND2_X1 U7579 ( .A1(n12451), .A2(n14974), .ZN(n14598) );
  AND2_X1 U7580 ( .A1(n7225), .A2(n15219), .ZN(n7224) );
  AND2_X1 U7581 ( .A1(n11929), .A2(n11924), .ZN(n7613) );
  AND2_X1 U7582 ( .A1(n7619), .A2(n14590), .ZN(n7618) );
  NAND2_X1 U7583 ( .A1(n11925), .A2(n11924), .ZN(n7619) );
  XNOR2_X1 U7584 ( .A(n11381), .B(n15330), .ZN(n7611) );
  NOR2_X1 U7585 ( .A1(n7633), .A2(n14601), .ZN(n7629) );
  INV_X1 U7586 ( .A(n7634), .ZN(n7633) );
  NAND2_X1 U7587 ( .A1(n6834), .A2(n6833), .ZN(n8473) );
  NAND2_X1 U7588 ( .A1(n6835), .A2(n8452), .ZN(n6834) );
  NAND2_X1 U7589 ( .A1(n6831), .A2(n6467), .ZN(n6835) );
  NAND2_X1 U7590 ( .A1(n6831), .A2(n8445), .ZN(n8453) );
  NAND2_X1 U7591 ( .A1(n8296), .A2(n8295), .ZN(n8303) );
  NAND2_X1 U7592 ( .A1(n8230), .A2(n8229), .ZN(n6777) );
  NAND2_X1 U7593 ( .A1(n8163), .A2(n8211), .ZN(n8213) );
  NAND2_X1 U7594 ( .A1(n7594), .A2(n7593), .ZN(n9129) );
  AND2_X1 U7595 ( .A1(n7595), .A2(n7597), .ZN(n7594) );
  NAND2_X1 U7596 ( .A1(n7600), .A2(n6513), .ZN(n7593) );
  NAND2_X1 U7597 ( .A1(n9114), .A2(n6941), .ZN(n9116) );
  NAND2_X1 U7598 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(n6942), .ZN(n6941) );
  INV_X1 U7599 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6942) );
  NAND2_X1 U7600 ( .A1(n9165), .A2(n6945), .ZN(n9169) );
  NAND2_X1 U7601 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n6946), .ZN(n6945) );
  NAND2_X1 U7602 ( .A1(n12364), .A2(n6512), .ZN(n7428) );
  INV_X1 U7603 ( .A(n11863), .ZN(n7463) );
  NAND2_X1 U7604 ( .A1(n9897), .A2(n7463), .ZN(n7460) );
  AOI21_X1 U7605 ( .B1(n12695), .B2(n12694), .A(n7829), .ZN(n12643) );
  NAND2_X1 U7606 ( .A1(n6888), .A2(n12669), .ZN(n12668) );
  NAND2_X1 U7607 ( .A1(n6883), .A2(n6882), .ZN(n6888) );
  AND2_X1 U7608 ( .A1(n6884), .A2(n12479), .ZN(n6882) );
  OR2_X1 U7609 ( .A1(n12738), .A2(n13355), .ZN(n10033) );
  INV_X1 U7610 ( .A(n10051), .ZN(n7450) );
  NOR2_X1 U7611 ( .A1(n7453), .A2(n10049), .ZN(n7452) );
  NAND2_X1 U7612 ( .A1(n7433), .A2(n12652), .ZN(n7432) );
  NAND2_X1 U7613 ( .A1(n9973), .A2(n9974), .ZN(n7433) );
  AOI21_X1 U7614 ( .B1(n13181), .B2(n12093), .A(n10355), .ZN(n12551) );
  NAND2_X1 U7615 ( .A1(n6653), .A2(n11089), .ZN(n11125) );
  NAND2_X1 U7616 ( .A1(n10987), .A2(n10946), .ZN(n6653) );
  NAND2_X1 U7617 ( .A1(n11815), .A2(n11814), .ZN(n11888) );
  XNOR2_X1 U7618 ( .A(n13057), .B(n13066), .ZN(n13052) );
  AND2_X1 U7619 ( .A1(n10956), .A2(n10913), .ZN(n10953) );
  OAI21_X1 U7620 ( .B1(n13096), .B2(n13095), .A(n13094), .ZN(n13097) );
  NOR2_X1 U7621 ( .A1(n13097), .A2(n13098), .ZN(n13103) );
  OR2_X1 U7622 ( .A1(n13088), .A2(n7503), .ZN(n7500) );
  INV_X1 U7623 ( .A(n7206), .ZN(n6985) );
  XNOR2_X1 U7624 ( .A(n12843), .B(n12842), .ZN(n12773) );
  NAND2_X1 U7625 ( .A1(n12943), .A2(n12948), .ZN(n12784) );
  NAND2_X1 U7626 ( .A1(n13427), .A2(n12551), .ZN(n12939) );
  OR2_X1 U7627 ( .A1(n13236), .A2(n7806), .ZN(n7805) );
  AND2_X1 U7628 ( .A1(n12918), .A2(n13251), .ZN(n7806) );
  OR2_X1 U7629 ( .A1(n12918), .A2(n13227), .ZN(n13218) );
  AOI21_X1 U7630 ( .B1(n7707), .B2(n7704), .A(n6547), .ZN(n7703) );
  INV_X1 U7631 ( .A(n12890), .ZN(n7704) );
  XNOR2_X1 U7632 ( .A(n13391), .B(n13294), .ZN(n13271) );
  AND2_X1 U7633 ( .A1(n10263), .A2(n10330), .ZN(n13344) );
  INV_X1 U7634 ( .A(n15597), .ZN(n15580) );
  OR2_X1 U7635 ( .A1(n12946), .A2(n10356), .ZN(n15582) );
  AND2_X1 U7636 ( .A1(n13498), .A2(n10394), .ZN(n10909) );
  INV_X1 U7637 ( .A(n15638), .ZN(n15623) );
  INV_X1 U7638 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9733) );
  AND2_X1 U7639 ( .A1(n7690), .A2(n7689), .ZN(n7688) );
  OR2_X1 U7640 ( .A1(n10200), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n10222) );
  NAND2_X1 U7641 ( .A1(n10039), .A2(n6479), .ZN(n10072) );
  AND2_X1 U7642 ( .A1(n9921), .A2(n9902), .ZN(n9919) );
  NAND2_X1 U7643 ( .A1(n10409), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9814) );
  NAND2_X1 U7644 ( .A1(n9794), .A2(n9793), .ZN(n9815) );
  INV_X1 U7645 ( .A(n6879), .ZN(n6880) );
  NAND2_X1 U7646 ( .A1(n9740), .A2(n9739), .ZN(n9760) );
  OR2_X1 U7647 ( .A1(n8531), .A2(n9191), .ZN(n8540) );
  AND2_X1 U7648 ( .A1(n8269), .A2(n8268), .ZN(n13549) );
  CLKBUF_X1 U7649 ( .A(n7979), .Z(n6947) );
  OR2_X1 U7650 ( .A1(n11840), .A2(n11841), .ZN(n7389) );
  AND2_X1 U7651 ( .A1(n7389), .A2(n7388), .ZN(n12471) );
  NAND2_X1 U7652 ( .A1(n12392), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7388) );
  NAND2_X1 U7653 ( .A1(n12389), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6673) );
  NOR2_X1 U7654 ( .A1(n13694), .A2(n13695), .ZN(n13696) );
  OR2_X1 U7655 ( .A1(n13720), .A2(n13723), .ZN(n13718) );
  AND2_X1 U7656 ( .A1(n13779), .A2(n6692), .ZN(n13761) );
  NAND2_X1 U7657 ( .A1(n13760), .A2(n13968), .ZN(n7023) );
  AND2_X1 U7658 ( .A1(n13784), .A2(n13795), .ZN(n9038) );
  NAND2_X1 U7659 ( .A1(n7175), .A2(n6527), .ZN(n7662) );
  NOR2_X1 U7660 ( .A1(n13806), .A2(n7664), .ZN(n7663) );
  INV_X1 U7661 ( .A(n7785), .ZN(n7784) );
  NAND2_X1 U7662 ( .A1(n13856), .A2(n13839), .ZN(n7783) );
  OAI21_X1 U7663 ( .B1(n7787), .B2(n7786), .A(n13838), .ZN(n7785) );
  NAND2_X1 U7664 ( .A1(n13884), .A2(n9031), .ZN(n7681) );
  AND2_X1 U7665 ( .A1(n6765), .A2(n6515), .ZN(n7679) );
  OR2_X1 U7666 ( .A1(n6762), .A2(n13913), .ZN(n6765) );
  NAND2_X1 U7667 ( .A1(n6766), .A2(n13911), .ZN(n6762) );
  NAND2_X1 U7668 ( .A1(n13945), .A2(n9028), .ZN(n7678) );
  AND3_X1 U7669 ( .A1(n6764), .A2(n6766), .A3(n6763), .ZN(n9028) );
  INV_X1 U7670 ( .A(n13913), .ZN(n6764) );
  OR2_X1 U7671 ( .A1(n13911), .A2(n13910), .ZN(n6763) );
  XNOR2_X1 U7672 ( .A(n13920), .B(n13893), .ZN(n13913) );
  OR2_X1 U7673 ( .A1(n14084), .A2(n13659), .ZN(n8789) );
  NAND2_X1 U7674 ( .A1(n6659), .A2(n11614), .ZN(n13896) );
  XNOR2_X1 U7675 ( .A(n8560), .B(n9039), .ZN(n6659) );
  NAND2_X1 U7676 ( .A1(n14165), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7878) );
  INV_X1 U7677 ( .A(n14363), .ZN(n7367) );
  INV_X1 U7678 ( .A(n9594), .ZN(n7366) );
  AND2_X1 U7679 ( .A1(n9594), .A2(n9592), .ZN(n14261) );
  OR2_X1 U7680 ( .A1(n9539), .A2(n14206), .ZN(n9561) );
  NAND2_X1 U7681 ( .A1(n9521), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9539) );
  INV_X1 U7682 ( .A(n9523), .ZN(n9521) );
  AND2_X1 U7683 ( .A1(n9632), .A2(n9631), .ZN(n11263) );
  INV_X1 U7684 ( .A(n6434), .ZN(n9664) );
  XNOR2_X1 U7685 ( .A(n12343), .B(n12350), .ZN(n15304) );
  NOR2_X1 U7686 ( .A1(n12593), .A2(n15077), .ZN(n12596) );
  OR2_X1 U7687 ( .A1(n15082), .A2(n14365), .ZN(n12407) );
  AND2_X1 U7688 ( .A1(n7070), .A2(n12460), .ZN(n7069) );
  NAND2_X1 U7689 ( .A1(n7072), .A2(n7071), .ZN(n7070) );
  NAND2_X1 U7690 ( .A1(n12207), .A2(n8948), .ZN(n8936) );
  NAND2_X1 U7691 ( .A1(n15111), .A2(n14241), .ZN(n12422) );
  OR2_X1 U7692 ( .A1(n14889), .A2(n14901), .ZN(n12420) );
  XNOR2_X1 U7693 ( .A(n14889), .B(n14870), .ZN(n14886) );
  OR2_X1 U7694 ( .A1(n15131), .A2(n14957), .ZN(n14492) );
  AND2_X1 U7695 ( .A1(n12446), .A2(n12445), .ZN(n7739) );
  INV_X1 U7696 ( .A(n15011), .ZN(n12446) );
  OR2_X2 U7697 ( .A1(n9331), .A2(n10871), .ZN(n9353) );
  XNOR2_X1 U7698 ( .A(n14428), .B(n11949), .ZN(n14592) );
  NOR2_X1 U7699 ( .A1(n7650), .A2(n6543), .ZN(n7649) );
  NAND2_X1 U7700 ( .A1(n11482), .A2(n14584), .ZN(n7652) );
  INV_X1 U7701 ( .A(n14534), .ZN(n14624) );
  AND2_X1 U7702 ( .A1(n10723), .A2(n10722), .ZN(n15325) );
  NAND2_X1 U7703 ( .A1(n11302), .A2(n8948), .ZN(n8909) );
  OR2_X1 U7704 ( .A1(n10721), .A2(n8961), .ZN(n15363) );
  NAND2_X1 U7705 ( .A1(n8474), .A2(n7007), .ZN(n8683) );
  NAND2_X1 U7706 ( .A1(n7008), .A2(SI_27_), .ZN(n7007) );
  NAND2_X1 U7707 ( .A1(n8472), .A2(n8471), .ZN(n8474) );
  INV_X1 U7708 ( .A(n8473), .ZN(n7008) );
  NAND2_X1 U7709 ( .A1(n8827), .A2(n8953), .ZN(n7416) );
  OR2_X1 U7710 ( .A1(n8954), .A2(n7415), .ZN(n7414) );
  NAND2_X1 U7711 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n7415) );
  XNOR2_X1 U7712 ( .A(n9110), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n9128) );
  XNOR2_X1 U7713 ( .A(n9116), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U7714 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n6944), .ZN(n6943) );
  INV_X1 U7715 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6944) );
  INV_X1 U7716 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7332) );
  NOR2_X1 U7717 ( .A1(n9179), .A2(n9178), .ZN(n9183) );
  AND2_X1 U7718 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n9177), .ZN(n9178) );
  NAND2_X1 U7719 ( .A1(n6858), .A2(n13146), .ZN(n6857) );
  OAI21_X1 U7720 ( .B1(n7090), .B2(n13104), .A(n13110), .ZN(n13088) );
  AOI21_X1 U7721 ( .B1(n7542), .B2(n7539), .A(n6510), .ZN(n7538) );
  NOR2_X1 U7722 ( .A1(n11204), .A2(n7540), .ZN(n7539) );
  INV_X1 U7723 ( .A(n7993), .ZN(n7540) );
  NAND2_X1 U7724 ( .A1(n7542), .A2(n7993), .ZN(n7541) );
  INV_X1 U7725 ( .A(n13549), .ZN(n13657) );
  NAND2_X1 U7726 ( .A1(n7776), .A2(n7775), .ZN(n7774) );
  NAND2_X1 U7727 ( .A1(n13794), .A2(n13966), .ZN(n7775) );
  NAND2_X1 U7728 ( .A1(n14531), .A2(n14533), .ZN(n7417) );
  OAI21_X1 U7729 ( .B1(n14529), .B2(n14528), .A(n6734), .ZN(n6725) );
  NAND2_X1 U7730 ( .A1(n12588), .A2(n6517), .ZN(n6982) );
  XNOR2_X1 U7731 ( .A(n9155), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15659) );
  OAI21_X1 U7732 ( .B1(n7082), .B2(n6815), .A(n15275), .ZN(n6813) );
  NAND2_X1 U7733 ( .A1(n9172), .A2(n15507), .ZN(n7605) );
  NAND2_X1 U7734 ( .A1(n6917), .A2(n6916), .ZN(n7606) );
  INV_X1 U7735 ( .A(n15287), .ZN(n6916) );
  INV_X1 U7736 ( .A(n15286), .ZN(n6917) );
  XNOR2_X1 U7737 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n9177), .ZN(n15247) );
  AOI21_X1 U7738 ( .B1(n13670), .B2(n8707), .A(n8583), .ZN(n8591) );
  NAND2_X1 U7739 ( .A1(n7012), .A2(n7011), .ZN(n7010) );
  INV_X1 U7740 ( .A(n8590), .ZN(n7012) );
  INV_X1 U7741 ( .A(n8591), .ZN(n7011) );
  INV_X1 U7742 ( .A(n14410), .ZN(n6722) );
  NOR2_X1 U7743 ( .A1(n14412), .A2(n14410), .ZN(n6723) );
  NAND2_X1 U7744 ( .A1(n14409), .A2(n14408), .ZN(n6724) );
  NOR2_X1 U7745 ( .A1(n14414), .A2(n14417), .ZN(n7479) );
  INV_X1 U7746 ( .A(n12806), .ZN(n7149) );
  OAI21_X1 U7747 ( .B1(n14415), .B2(n7479), .A(n6954), .ZN(n14423) );
  AND2_X1 U7748 ( .A1(n7476), .A2(n7478), .ZN(n6954) );
  INV_X1 U7749 ( .A(n8600), .ZN(n7006) );
  OAI21_X1 U7750 ( .B1(n12814), .B2(n7128), .A(n7126), .ZN(n7125) );
  INV_X1 U7751 ( .A(n7127), .ZN(n7126) );
  NAND2_X1 U7752 ( .A1(n7658), .A2(n7657), .ZN(n7656) );
  OAI211_X1 U7753 ( .C1(n6721), .C2(n6720), .A(n14473), .B(n6719), .ZN(n14488)
         );
  INV_X1 U7754 ( .A(n14469), .ZN(n6720) );
  NAND2_X1 U7755 ( .A1(n6569), .A2(n14469), .ZN(n6719) );
  NAND2_X1 U7756 ( .A1(n7145), .A2(n7144), .ZN(n7143) );
  INV_X1 U7757 ( .A(n12864), .ZN(n7144) );
  NAND2_X1 U7758 ( .A1(n7146), .A2(n12865), .ZN(n7145) );
  NOR2_X1 U7759 ( .A1(n12867), .A2(n12868), .ZN(n7142) );
  NAND2_X1 U7760 ( .A1(n6904), .A2(n6538), .ZN(n8634) );
  NAND2_X1 U7761 ( .A1(n7627), .A2(n6499), .ZN(n7625) );
  INV_X1 U7762 ( .A(n7141), .ZN(n7138) );
  INV_X1 U7763 ( .A(n8647), .ZN(n7655) );
  AOI21_X1 U7764 ( .B1(n14026), .B2(n8707), .A(n8668), .ZN(n8731) );
  NAND2_X1 U7765 ( .A1(n7449), .A2(n14517), .ZN(n7448) );
  NOR2_X1 U7766 ( .A1(n8190), .A2(n7338), .ZN(n7337) );
  INV_X1 U7767 ( .A(n8161), .ZN(n7338) );
  NOR2_X1 U7768 ( .A1(n8212), .A2(SI_14_), .ZN(n8190) );
  INV_X1 U7769 ( .A(n12977), .ZN(n10316) );
  NOR2_X1 U7770 ( .A1(n12835), .A2(n12771), .ZN(n7801) );
  AOI21_X1 U7771 ( .B1(n7641), .B2(n7643), .A(n6564), .ZN(n7638) );
  NOR2_X1 U7772 ( .A1(n7641), .A2(n6482), .ZN(n7640) );
  AND2_X1 U7773 ( .A1(n8745), .A2(n8678), .ZN(n8752) );
  NAND2_X1 U7774 ( .A1(n7273), .A2(n7274), .ZN(n7272) );
  INV_X1 U7775 ( .A(n10618), .ZN(n7318) );
  AOI21_X1 U7776 ( .B1(n7352), .B2(n7354), .A(n7349), .ZN(n7348) );
  INV_X1 U7777 ( .A(n8395), .ZN(n7349) );
  AOI21_X1 U7778 ( .B1(n8301), .B2(n8300), .A(n8299), .ZN(n8302) );
  INV_X1 U7779 ( .A(n8335), .ZN(n8334) );
  OAI21_X1 U7780 ( .B1(n6443), .B2(n7186), .A(n7337), .ZN(n6768) );
  NAND2_X1 U7781 ( .A1(n8193), .A2(n8192), .ZN(n8250) );
  AND2_X1 U7782 ( .A1(n6471), .A2(n8140), .ZN(n6443) );
  NOR2_X1 U7783 ( .A1(n8120), .A2(n8118), .ZN(n8121) );
  INV_X1 U7784 ( .A(n8086), .ZN(n8087) );
  INV_X1 U7785 ( .A(n8030), .ZN(n8032) );
  NAND2_X1 U7786 ( .A1(n6980), .A2(n6738), .ZN(n6737) );
  OAI21_X1 U7787 ( .B1(n7955), .B2(n10441), .A(n6846), .ZN(n7996) );
  OAI21_X1 U7788 ( .B1(n7955), .B2(n10447), .A(n6950), .ZN(n7974) );
  NAND2_X1 U7789 ( .A1(n7955), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6950) );
  OAI21_X1 U7790 ( .B1(n12702), .B2(n7422), .A(n7421), .ZN(n10172) );
  NAND2_X1 U7791 ( .A1(n10193), .A2(n13264), .ZN(n7422) );
  NAND2_X1 U7792 ( .A1(n10155), .A2(n10193), .ZN(n7421) );
  NAND2_X1 U7793 ( .A1(n10191), .A2(n6887), .ZN(n6883) );
  NOR2_X1 U7794 ( .A1(n10196), .A2(n6520), .ZN(n6887) );
  NOR2_X1 U7795 ( .A1(n10134), .A2(n13252), .ZN(n10135) );
  NOR2_X1 U7796 ( .A1(n11041), .A2(n15593), .ZN(n9745) );
  NAND2_X1 U7797 ( .A1(n10987), .A2(n6522), .ZN(n7515) );
  OAI21_X1 U7798 ( .B1(n11126), .B2(n7519), .A(n7517), .ZN(n10948) );
  INV_X1 U7799 ( .A(n7518), .ZN(n7517) );
  OAI21_X1 U7800 ( .B1(n11125), .B2(n7519), .A(n10947), .ZN(n7518) );
  INV_X1 U7801 ( .A(n11215), .ZN(n7096) );
  AOI21_X1 U7802 ( .B1(n6822), .B2(n12245), .A(n12981), .ZN(n6818) );
  NOR2_X1 U7803 ( .A1(n13033), .A2(n13032), .ZN(n13034) );
  NAND2_X1 U7804 ( .A1(n13042), .A2(n13041), .ZN(n13064) );
  INV_X1 U7805 ( .A(n13109), .ZN(n7504) );
  NAND2_X1 U7806 ( .A1(n6881), .A2(n7154), .ZN(n10290) );
  INV_X1 U7807 ( .A(n10272), .ZN(n7154) );
  AND2_X1 U7808 ( .A1(n10232), .A2(n10231), .ZN(n10280) );
  AND2_X1 U7809 ( .A1(n10096), .A2(n7161), .ZN(n7160) );
  INV_X1 U7810 ( .A(n10098), .ZN(n10097) );
  AND2_X1 U7811 ( .A1(n10026), .A2(n7158), .ZN(n7157) );
  INV_X1 U7812 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n7158) );
  INV_X1 U7813 ( .A(n10028), .ZN(n10027) );
  NOR2_X1 U7814 ( .A1(n9949), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7155) );
  INV_X1 U7815 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7163) );
  INV_X1 U7816 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9847) );
  INV_X1 U7817 ( .A(n9882), .ZN(n9848) );
  NOR2_X1 U7818 ( .A1(n11780), .A2(n10318), .ZN(n7193) );
  OAI21_X1 U7819 ( .B1(n12819), .B2(n7698), .A(n12824), .ZN(n7697) );
  INV_X1 U7820 ( .A(n12821), .ZN(n7698) );
  AND3_X1 U7821 ( .A1(n10317), .A2(n12768), .A3(n11777), .ZN(n11780) );
  OR2_X1 U7822 ( .A1(n12819), .A2(n7839), .ZN(n10317) );
  NAND2_X1 U7823 ( .A1(n12827), .A2(n12826), .ZN(n12768) );
  AND2_X1 U7824 ( .A1(n11045), .A2(n7150), .ZN(n10998) );
  NAND2_X1 U7825 ( .A1(n9757), .A2(n15593), .ZN(n12807) );
  NAND2_X1 U7826 ( .A1(n10310), .A2(n10311), .ZN(n6871) );
  AND2_X1 U7827 ( .A1(n13451), .A2(n13264), .ZN(n12912) );
  NOR2_X1 U7828 ( .A1(n13262), .A2(n7792), .ZN(n7791) );
  INV_X1 U7829 ( .A(n10339), .ZN(n7792) );
  INV_X1 U7830 ( .A(n12911), .ZN(n7700) );
  AND2_X1 U7831 ( .A1(n12901), .A2(n13287), .ZN(n12890) );
  NAND2_X1 U7832 ( .A1(n13302), .A2(n13305), .ZN(n13286) );
  INV_X1 U7833 ( .A(n7726), .ZN(n7722) );
  AND2_X1 U7834 ( .A1(n13344), .A2(n13348), .ZN(n10329) );
  NAND2_X1 U7835 ( .A1(n7795), .A2(n12335), .ZN(n7794) );
  NAND2_X1 U7836 ( .A1(n7796), .A2(n10325), .ZN(n7795) );
  AND2_X1 U7837 ( .A1(n12865), .A2(n12866), .ZN(n12775) );
  INV_X1 U7838 ( .A(n9814), .ZN(n7591) );
  AOI21_X1 U7839 ( .B1(n13571), .B2(n8228), .A(n8227), .ZN(n13584) );
  INV_X1 U7840 ( .A(n13546), .ZN(n7544) );
  NAND2_X1 U7841 ( .A1(n8725), .A2(n8783), .ZN(n8768) );
  NAND2_X1 U7842 ( .A1(n6692), .A2(n13773), .ZN(n8785) );
  AND2_X1 U7843 ( .A1(n7177), .A2(n7178), .ZN(n7176) );
  XNOR2_X1 U7844 ( .A(n7410), .B(n13655), .ZN(n13838) );
  NOR2_X1 U7845 ( .A1(n8240), .A2(n8239), .ZN(n6693) );
  INV_X1 U7846 ( .A(n9067), .ZN(n6632) );
  NOR2_X1 U7847 ( .A1(n7676), .A2(n7673), .ZN(n7672) );
  INV_X1 U7848 ( .A(n9017), .ZN(n7673) );
  INV_X1 U7849 ( .A(n9022), .ZN(n7676) );
  INV_X1 U7850 ( .A(n9021), .ZN(n7675) );
  INV_X1 U7851 ( .A(n12110), .ZN(n9020) );
  INV_X1 U7852 ( .A(n8003), .ZN(n6689) );
  NAND2_X1 U7853 ( .A1(n12119), .A2(n8571), .ZN(n11327) );
  NAND2_X1 U7854 ( .A1(n7767), .A2(n9065), .ZN(n13929) );
  NAND2_X1 U7855 ( .A1(n13948), .A2(n9064), .ZN(n7767) );
  NOR2_X1 U7856 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n7257) );
  NOR2_X1 U7857 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7258) );
  AOI21_X1 U7858 ( .B1(n9626), .B2(n9625), .A(n9655), .ZN(n10381) );
  INV_X1 U7859 ( .A(n14330), .ZN(n9557) );
  INV_X1 U7860 ( .A(n7466), .ZN(n7465) );
  OAI21_X1 U7861 ( .B1(n7469), .B2(n7467), .A(n14526), .ZN(n7466) );
  INV_X1 U7862 ( .A(n14529), .ZN(n7467) );
  NAND2_X1 U7863 ( .A1(n7318), .A2(n7314), .ZN(n7313) );
  INV_X1 U7864 ( .A(n7316), .ZN(n7314) );
  AOI21_X1 U7865 ( .B1(n14706), .B2(n14707), .A(n7317), .ZN(n7316) );
  INV_X1 U7866 ( .A(n10619), .ZN(n7317) );
  INV_X1 U7867 ( .A(n11110), .ZN(n7292) );
  NAND2_X1 U7868 ( .A1(n12418), .A2(n12454), .ZN(n7065) );
  NAND2_X1 U7869 ( .A1(n6496), .A2(n7066), .ZN(n7063) );
  INV_X1 U7870 ( .A(n12454), .ZN(n7066) );
  NOR2_X1 U7871 ( .A1(n14921), .A2(n7246), .ZN(n7245) );
  INV_X1 U7872 ( .A(n14492), .ZN(n7246) );
  NOR2_X1 U7873 ( .A1(n7484), .A2(n15131), .ZN(n14924) );
  NAND2_X1 U7874 ( .A1(n9355), .A2(n9354), .ZN(n9368) );
  INV_X1 U7875 ( .A(n9353), .ZN(n9355) );
  NAND2_X1 U7876 ( .A1(n15058), .A2(n7493), .ZN(n7492) );
  INV_X1 U7877 ( .A(n11590), .ZN(n7241) );
  INV_X1 U7878 ( .A(n7742), .ZN(n7741) );
  OAI21_X1 U7879 ( .B1(n12449), .B2(n7743), .A(n12450), .ZN(n7742) );
  NAND2_X1 U7880 ( .A1(n6844), .A2(n6842), .ZN(n7347) );
  AND2_X1 U7881 ( .A1(n6843), .A2(n8716), .ZN(n6842) );
  NAND2_X1 U7882 ( .A1(n8683), .A2(n8681), .ZN(n6844) );
  NAND2_X1 U7883 ( .A1(n8682), .A2(n8681), .ZN(n6843) );
  AND2_X1 U7884 ( .A1(n7346), .A2(n8685), .ZN(n7345) );
  INV_X1 U7885 ( .A(n8700), .ZN(n7346) );
  INV_X1 U7886 ( .A(n7237), .ZN(n7232) );
  AND4_X1 U7887 ( .A1(n7229), .A2(n7228), .A3(n7227), .A4(n6641), .ZN(n7233)
         );
  NOR2_X1 U7888 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n7229) );
  NOR2_X1 U7889 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7228) );
  NOR2_X1 U7890 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7227) );
  INV_X1 U7891 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7056) );
  AND2_X1 U7892 ( .A1(n8822), .A2(n8821), .ZN(n6791) );
  INV_X1 U7893 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7660) );
  AND3_X1 U7894 ( .A1(n6791), .A2(n8823), .A3(n6474), .ZN(n7832) );
  NAND2_X1 U7895 ( .A1(n8303), .A2(n8302), .ZN(n8339) );
  INV_X1 U7896 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7236) );
  INV_X1 U7897 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7235) );
  NAND2_X1 U7898 ( .A1(n8275), .A2(SI_19_), .ZN(n8300) );
  NAND2_X1 U7899 ( .A1(n8257), .A2(n8256), .ZN(n8296) );
  AOI21_X1 U7900 ( .B1(n7334), .B2(n7336), .A(n6561), .ZN(n7333) );
  NAND2_X1 U7901 ( .A1(n8273), .A2(n8297), .ZN(n6736) );
  XNOR2_X1 U7902 ( .A(n8296), .B(SI_18_), .ZN(n8273) );
  NAND2_X1 U7903 ( .A1(n8889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8893) );
  OR2_X1 U7904 ( .A1(n8888), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U7905 ( .A1(n8036), .A2(SI_8_), .ZN(n8037) );
  XNOR2_X1 U7906 ( .A(n8070), .B(SI_9_), .ZN(n8069) );
  XNOR2_X1 U7907 ( .A(n7996), .B(SI_5_), .ZN(n7994) );
  NAND2_X1 U7908 ( .A1(n7954), .A2(n7953), .ZN(n7973) );
  NAND2_X1 U7909 ( .A1(n9100), .A2(n9099), .ZN(n9102) );
  NAND2_X1 U7910 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n9098), .ZN(n9099) );
  NAND2_X1 U7911 ( .A1(n10998), .A2(n12807), .ZN(n10258) );
  NAND2_X1 U7912 ( .A1(n11136), .A2(n7458), .ZN(n11404) );
  AND2_X1 U7913 ( .A1(n9812), .A2(n9789), .ZN(n7458) );
  INV_X1 U7914 ( .A(n7460), .ZN(n7462) );
  OR2_X1 U7915 ( .A1(n9826), .A2(n11050), .ZN(n9726) );
  OR2_X1 U7916 ( .A1(n9822), .A2(n9724), .ZN(n9727) );
  NAND2_X1 U7917 ( .A1(n12668), .A2(n12482), .ZN(n12728) );
  NAND2_X1 U7918 ( .A1(n7428), .A2(n7426), .ZN(n12618) );
  NOR2_X1 U7919 ( .A1(n7430), .A2(n7427), .ZN(n7426) );
  NOR4_X1 U7920 ( .A1(n12784), .A2(n12783), .A3(n10346), .A4(n13173), .ZN(
        n12787) );
  OR2_X1 U7921 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  AND4_X1 U7922 ( .A1(n9933), .A2(n9932), .A3(n9931), .A4(n9930), .ZN(n12369)
         );
  OAI21_X1 U7923 ( .B1(n13039), .B2(P3_REG2_REG_1__SCAN_IN), .A(n6956), .ZN(
        n10915) );
  NAND2_X1 U7924 ( .A1(n13039), .A2(n10968), .ZN(n6956) );
  OR2_X1 U7925 ( .A1(n10943), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7327) );
  NAND2_X1 U7926 ( .A1(n7088), .A2(n10983), .ZN(n10987) );
  NAND2_X1 U7927 ( .A1(n11001), .A2(n10984), .ZN(n7088) );
  INV_X1 U7928 ( .A(n11081), .ZN(n6755) );
  NAND2_X1 U7929 ( .A1(n11061), .A2(n11060), .ZN(n11066) );
  NAND2_X1 U7930 ( .A1(n11229), .A2(n7096), .ZN(n7095) );
  NAND2_X1 U7931 ( .A1(n11216), .A2(n7094), .ZN(n7093) );
  NOR2_X1 U7932 ( .A1(n11229), .A2(n7096), .ZN(n7094) );
  AOI21_X1 U7933 ( .B1(n11213), .B2(n11212), .A(n11211), .ZN(n11653) );
  NAND2_X1 U7934 ( .A1(n6816), .A2(n7320), .ZN(n11873) );
  OR2_X1 U7935 ( .A1(n7322), .A2(n6444), .ZN(n7320) );
  NAND2_X1 U7936 ( .A1(n11653), .A2(n7321), .ZN(n6816) );
  AND2_X1 U7937 ( .A1(n11806), .A2(n6462), .ZN(n7322) );
  NAND2_X1 U7938 ( .A1(n11888), .A2(n11885), .ZN(n12993) );
  NOR2_X1 U7939 ( .A1(n11809), .A2(n11884), .ZN(n11877) );
  NOR2_X1 U7940 ( .A1(n13010), .A2(n7098), .ZN(n12987) );
  NAND2_X1 U7941 ( .A1(n13023), .A2(n6747), .ZN(n13042) );
  NOR2_X1 U7942 ( .A1(n6749), .A2(n6748), .ZN(n6747) );
  INV_X1 U7943 ( .A(n13021), .ZN(n6748) );
  INV_X1 U7944 ( .A(n13022), .ZN(n6749) );
  AND2_X1 U7945 ( .A1(n7099), .A2(n13004), .ZN(n13010) );
  XNOR2_X1 U7946 ( .A(n13064), .B(n13058), .ZN(n13044) );
  NOR2_X1 U7947 ( .A1(n13044), .A2(n13043), .ZN(n13065) );
  OAI21_X1 U7948 ( .B1(n13051), .B2(n13050), .A(n13049), .ZN(n13057) );
  NAND2_X1 U7949 ( .A1(n13052), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n13059) );
  NAND2_X1 U7950 ( .A1(n13086), .A2(n13085), .ZN(n7090) );
  OR2_X1 U7951 ( .A1(n12483), .A2(n13212), .ZN(n12931) );
  AND2_X1 U7952 ( .A1(n12936), .A2(n12937), .ZN(n12934) );
  OAI21_X1 U7953 ( .B1(n13210), .B2(n13209), .A(n7210), .ZN(n13192) );
  NAND2_X1 U7954 ( .A1(n13218), .A2(n10344), .ZN(n13235) );
  OR2_X1 U7955 ( .A1(n10147), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n10163) );
  NAND2_X1 U7956 ( .A1(n10097), .A2(n10096), .ZN(n10113) );
  OR2_X1 U7957 ( .A1(n10077), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n10098) );
  AOI21_X1 U7958 ( .B1(n10329), .B2(n6572), .A(n7800), .ZN(n7798) );
  INV_X1 U7959 ( .A(n10330), .ZN(n7800) );
  OR2_X1 U7960 ( .A1(n10005), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n10028) );
  NAND2_X1 U7961 ( .A1(n7155), .A2(n10829), .ZN(n9989) );
  AOI21_X1 U7962 ( .B1(n6437), .B2(n7718), .A(n6563), .ZN(n7715) );
  NOR2_X1 U7963 ( .A1(n12773), .A2(n7717), .ZN(n7716) );
  INV_X1 U7964 ( .A(n6498), .ZN(n7718) );
  NAND2_X1 U7965 ( .A1(n11492), .A2(n12820), .ZN(n11730) );
  AND3_X1 U7966 ( .A1(n9821), .A2(n9820), .A3(n9819), .ZN(n11774) );
  AND4_X1 U7967 ( .A1(n9808), .A2(n9807), .A3(n9806), .A4(n9805), .ZN(n11784)
         );
  AND4_X1 U7968 ( .A1(n9784), .A2(n9783), .A3(n9782), .A4(n9781), .ZN(n15581)
         );
  AND3_X1 U7969 ( .A1(n6575), .A2(n12555), .A3(n12554), .ZN(n12559) );
  INV_X1 U7970 ( .A(n13166), .ZN(n7200) );
  AND2_X1 U7971 ( .A1(n10306), .A2(n10305), .ZN(n13193) );
  NAND2_X1 U7972 ( .A1(n12939), .A2(n7581), .ZN(n13173) );
  AND3_X1 U7973 ( .A1(n6871), .A2(n6870), .A3(n6508), .ZN(n12544) );
  NAND2_X1 U7974 ( .A1(n10296), .A2(n10295), .ZN(n6850) );
  NAND2_X1 U7975 ( .A1(n10270), .A2(n10269), .ZN(n13376) );
  NOR2_X1 U7976 ( .A1(n13234), .A2(n13235), .ZN(n13233) );
  AND2_X1 U7977 ( .A1(n7214), .A2(n7212), .ZN(n13236) );
  AND2_X1 U7978 ( .A1(n13235), .A2(n7213), .ZN(n7212) );
  NAND2_X1 U7979 ( .A1(n10161), .A2(n10160), .ZN(n12918) );
  OAI211_X1 U7980 ( .C1(n13277), .C2(n10338), .A(n13280), .B(n10337), .ZN(
        n10340) );
  NAND2_X1 U7981 ( .A1(n10340), .A2(n7791), .ZN(n13259) );
  INV_X1 U7982 ( .A(n7707), .ZN(n7705) );
  AND2_X1 U7983 ( .A1(n7700), .A2(n12909), .ZN(n13262) );
  AND2_X1 U7984 ( .A1(n13271), .A2(n12900), .ZN(n7707) );
  NAND2_X1 U7985 ( .A1(n6925), .A2(n12890), .ZN(n7708) );
  OR2_X1 U7986 ( .A1(n13470), .A2(n13316), .ZN(n13287) );
  INV_X1 U7987 ( .A(n12710), .ZN(n13307) );
  AOI21_X1 U7988 ( .B1(n13312), .B2(n12885), .A(n12889), .ZN(n13302) );
  NAND2_X1 U7989 ( .A1(n10025), .A2(n10024), .ZN(n13410) );
  NOR2_X1 U7990 ( .A1(n12874), .A2(n12869), .ZN(n7726) );
  NAND2_X1 U7991 ( .A1(n6571), .A2(n7729), .ZN(n7727) );
  NAND2_X1 U7992 ( .A1(n12870), .A2(n12377), .ZN(n7728) );
  AND3_X1 U7993 ( .A1(n10032), .A2(n10031), .A3(n10030), .ZN(n13355) );
  AND4_X1 U7994 ( .A1(n9994), .A2(n9993), .A3(n9992), .A4(n9991), .ZN(n13354)
         );
  AOI21_X1 U7995 ( .B1(n12150), .B2(n12851), .A(n12853), .ZN(n12241) );
  AND3_X1 U7996 ( .A1(n9800), .A2(n9799), .A3(n9798), .ZN(n15624) );
  NAND2_X1 U7997 ( .A1(n12801), .A2(n6928), .ZN(n15638) );
  INV_X1 U7998 ( .A(n10204), .ZN(n10545) );
  OAI22_X1 U7999 ( .A1(n10204), .A2(P3_D_REG_0__SCAN_IN), .B1(n9710), .B2(
        n9712), .ZN(n10369) );
  AND2_X1 U8000 ( .A1(n9720), .A2(n9733), .ZN(n7808) );
  OAI21_X1 U8001 ( .B1(n12581), .B2(n12580), .A(n12582), .ZN(n12753) );
  NAND2_X1 U8002 ( .A1(n7809), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U8003 ( .A1(n6878), .A2(n10275), .ZN(n10292) );
  NAND2_X1 U8004 ( .A1(n10274), .A2(n10273), .ZN(n6878) );
  NOR2_X1 U8005 ( .A1(n9690), .A2(n9694), .ZN(n7687) );
  NOR2_X1 U8006 ( .A1(n9691), .A2(n9690), .ZN(n9705) );
  NOR2_X1 U8007 ( .A1(n9695), .A2(n9694), .ZN(n9704) );
  NAND2_X1 U8008 ( .A1(n10179), .A2(n12212), .ZN(n7592) );
  OR2_X1 U8009 ( .A1(n10122), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n10124) );
  INV_X1 U8010 ( .A(n9691), .ZN(n7480) );
  INV_X1 U8011 ( .A(n10001), .ZN(n7481) );
  AOI21_X1 U8012 ( .B1(n10016), .B2(n10017), .A(n7572), .ZN(n7571) );
  INV_X1 U8013 ( .A(n10019), .ZN(n7572) );
  NAND2_X1 U8014 ( .A1(n6876), .A2(n9980), .ZN(n10018) );
  OAI21_X1 U8015 ( .B1(n9956), .B2(n6875), .A(n6873), .ZN(n6876) );
  INV_X1 U8016 ( .A(n6874), .ZN(n6873) );
  OAI21_X1 U8017 ( .B1(n9955), .B2(n6875), .A(n9978), .ZN(n6874) );
  NAND2_X1 U8018 ( .A1(n9997), .A2(n9981), .ZN(n9998) );
  OR2_X1 U8019 ( .A1(n10018), .A2(n10681), .ZN(n9981) );
  NAND2_X1 U8020 ( .A1(n6863), .A2(n6861), .ZN(n9940) );
  AOI21_X1 U8021 ( .B1(n6495), .B2(n6866), .A(n6862), .ZN(n6861) );
  INV_X1 U8022 ( .A(n9921), .ZN(n6862) );
  AND2_X1 U8023 ( .A1(n9941), .A2(n9922), .ZN(n9939) );
  AOI21_X1 U8024 ( .B1(n9899), .B2(n7586), .A(n7585), .ZN(n7584) );
  INV_X1 U8025 ( .A(n9901), .ZN(n7585) );
  INV_X1 U8026 ( .A(n9840), .ZN(n7586) );
  AND2_X1 U8027 ( .A1(n9840), .A2(n9839), .ZN(n9862) );
  OAI21_X1 U8028 ( .B1(n9876), .B2(n9875), .A(n9838), .ZN(n9863) );
  AND2_X1 U8029 ( .A1(n9814), .A2(n9792), .ZN(n9793) );
  NAND2_X1 U8030 ( .A1(n10738), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9790) );
  XNOR2_X1 U8031 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9772) );
  INV_X1 U8032 ( .A(n9759), .ZN(n7580) );
  INV_X1 U8033 ( .A(n9761), .ZN(n7575) );
  XNOR2_X1 U8034 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9740) );
  NAND2_X1 U8035 ( .A1(n9737), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9753) );
  INV_X1 U8036 ( .A(n11144), .ZN(n7542) );
  INV_X1 U8037 ( .A(n13773), .ZN(n13744) );
  NAND2_X1 U8038 ( .A1(n6654), .A2(n6519), .ZN(n13525) );
  INV_X1 U8039 ( .A(n13528), .ZN(n6939) );
  OAI21_X1 U8040 ( .B1(n13621), .B2(n7549), .A(n8272), .ZN(n7548) );
  NAND2_X1 U8041 ( .A1(n7552), .A2(n8249), .ZN(n7551) );
  INV_X1 U8042 ( .A(n13621), .ZN(n7552) );
  AND2_X1 U8043 ( .A1(n8373), .A2(n7534), .ZN(n7532) );
  NAND2_X1 U8044 ( .A1(n7553), .A2(n7554), .ZN(n10885) );
  NOR2_X1 U8045 ( .A1(n10887), .A2(n7555), .ZN(n7554) );
  INV_X1 U8046 ( .A(n7558), .ZN(n7555) );
  NAND2_X1 U8047 ( .A1(n6694), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U8048 ( .A1(n8062), .A2(n11751), .ZN(n7528) );
  INV_X1 U8049 ( .A(n11751), .ZN(n7529) );
  OR2_X1 U8050 ( .A1(n7943), .A2(n13989), .ZN(n7883) );
  NOR2_X1 U8051 ( .A1(n8810), .A2(n8809), .ZN(n8814) );
  AND4_X1 U8052 ( .A1(n8106), .A2(n8105), .A3(n8104), .A4(n8103), .ZN(n12195)
         );
  AND4_X1 U8053 ( .A1(n8045), .A2(n8044), .A3(n8043), .A4(n8042), .ZN(n11754)
         );
  OR2_X1 U8054 ( .A1(n7980), .A2(n12028), .ZN(n7945) );
  OAI21_X1 U8055 ( .B1(n6667), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6666), .ZN(
        n15449) );
  NAND2_X1 U8056 ( .A1(n6667), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6666) );
  OAI21_X1 U8057 ( .B1(n15470), .B2(n6663), .A(n6661), .ZN(n6665) );
  INV_X1 U8058 ( .A(n6662), .ZN(n6661) );
  OAI21_X1 U8059 ( .B1(n10526), .B2(n6663), .A(n6560), .ZN(n6662) );
  OR2_X1 U8060 ( .A1(n11165), .A2(n11166), .ZN(n7385) );
  AND2_X1 U8061 ( .A1(n7385), .A2(n7384), .ZN(n11467) );
  NAND2_X1 U8062 ( .A1(n11465), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7384) );
  OR2_X1 U8063 ( .A1(n11467), .A2(n11466), .ZN(n7383) );
  NAND2_X1 U8064 ( .A1(n6685), .A2(n6684), .ZN(n7387) );
  INV_X1 U8065 ( .A(n12470), .ZN(n6684) );
  AND2_X1 U8066 ( .A1(n7387), .A2(n7386), .ZN(n13682) );
  NAND2_X1 U8067 ( .A1(n12474), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7386) );
  NAND2_X1 U8068 ( .A1(n15500), .A2(n6620), .ZN(n7390) );
  NAND2_X1 U8069 ( .A1(n6448), .A2(n6673), .ZN(n6672) );
  NAND2_X1 U8070 ( .A1(n6683), .A2(n13699), .ZN(n13693) );
  AND3_X1 U8071 ( .A1(n13693), .A2(n7380), .A3(P2_REG1_REG_18__SCAN_IN), .ZN(
        n13694) );
  NAND2_X1 U8072 ( .A1(n6431), .A2(n7405), .ZN(n13727) );
  NAND2_X1 U8073 ( .A1(n13758), .A2(n13759), .ZN(n13738) );
  AND2_X1 U8074 ( .A1(n8437), .A2(n8459), .ZN(n13763) );
  INV_X1 U8075 ( .A(n9081), .ZN(n13759) );
  AOI21_X1 U8076 ( .B1(n7268), .B2(n7271), .A(n7265), .ZN(n7264) );
  INV_X1 U8077 ( .A(n13810), .ZN(n13775) );
  AND2_X1 U8078 ( .A1(n13806), .A2(n13790), .ZN(n7789) );
  NAND2_X1 U8079 ( .A1(n14137), .A2(n13860), .ZN(n7178) );
  OR2_X1 U8080 ( .A1(n13852), .A2(n13838), .ZN(n7179) );
  NAND2_X1 U8081 ( .A1(n7179), .A2(n7176), .ZN(n13824) );
  NAND2_X1 U8082 ( .A1(n13889), .A2(n9030), .ZN(n13884) );
  AOI21_X1 U8083 ( .B1(n7765), .B2(n7278), .A(n6542), .ZN(n7277) );
  INV_X1 U8084 ( .A(n9064), .ZN(n7278) );
  NAND2_X1 U8085 ( .A1(n12299), .A2(n13980), .ZN(n13973) );
  NOR2_X1 U8086 ( .A1(n13982), .A2(n7756), .ZN(n7755) );
  INV_X1 U8087 ( .A(n7759), .ZN(n7756) );
  AND4_X1 U8088 ( .A1(n8081), .A2(n8080), .A3(n8079), .A4(n8078), .ZN(n12168)
         );
  CLKBUF_X1 U8089 ( .A(n11974), .Z(n7031) );
  INV_X1 U8090 ( .A(n13669), .ZN(n12036) );
  AND2_X1 U8091 ( .A1(n7262), .A2(n9048), .ZN(n7833) );
  AND2_X1 U8092 ( .A1(n10491), .A2(n8542), .ZN(n13966) );
  INV_X1 U8093 ( .A(n13966), .ZN(n13930) );
  INV_X1 U8094 ( .A(n13968), .ZN(n13932) );
  AND2_X1 U8095 ( .A1(n9084), .A2(n9083), .ZN(n13951) );
  OR2_X1 U8096 ( .A1(n9088), .A2(n15536), .ZN(n7820) );
  NAND2_X1 U8097 ( .A1(n6492), .A2(n6760), .ZN(n6759) );
  INV_X1 U8098 ( .A(n9087), .ZN(n6760) );
  NAND2_X1 U8099 ( .A1(n8238), .A2(n8237), .ZN(n13920) );
  OAI211_X1 U8100 ( .C1(n6777), .C2(n6774), .A(n8718), .B(n6771), .ZN(n8238)
         );
  NAND2_X1 U8101 ( .A1(n6775), .A2(n8254), .ZN(n6774) );
  NOR2_X1 U8102 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7840) );
  INV_X1 U8103 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6908) );
  NAND2_X1 U8104 ( .A1(n6911), .A2(n7875), .ZN(n6910) );
  INV_X1 U8105 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U8106 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n7850) );
  INV_X1 U8107 ( .A(n7843), .ZN(n8196) );
  OR2_X1 U8108 ( .A1(n7969), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7998) );
  OR2_X1 U8109 ( .A1(n7937), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7958) );
  INV_X1 U8110 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9737) );
  NAND2_X1 U8111 ( .A1(n7370), .A2(n7368), .ZN(n6711) );
  NOR2_X1 U8112 ( .A1(n9556), .A2(n7369), .ZN(n7368) );
  INV_X1 U8113 ( .A(n7371), .ZN(n7369) );
  OR2_X1 U8114 ( .A1(n14199), .A2(n9559), .ZN(n9556) );
  AOI21_X1 U8115 ( .B1(n7365), .B2(n7367), .A(n7362), .ZN(n7361) );
  INV_X1 U8116 ( .A(n10381), .ZN(n7362) );
  XNOR2_X1 U8117 ( .A(n9247), .B(n6706), .ZN(n14231) );
  NAND2_X1 U8118 ( .A1(n6708), .A2(n6707), .ZN(n14232) );
  NAND2_X1 U8119 ( .A1(n10654), .A2(n10653), .ZN(n6708) );
  NOR2_X1 U8120 ( .A1(n11947), .A2(n7375), .ZN(n7374) );
  INV_X1 U8121 ( .A(n7376), .ZN(n7375) );
  NAND2_X1 U8122 ( .A1(n14212), .A2(n6531), .ZN(n14339) );
  INV_X1 U8123 ( .A(n11601), .ZN(n9300) );
  OAI21_X1 U8124 ( .B1(n10398), .B2(n11516), .A(n7377), .ZN(n9301) );
  INV_X1 U8125 ( .A(n7378), .ZN(n7377) );
  AND2_X1 U8126 ( .A1(n9609), .A2(n9608), .ZN(n7045) );
  NAND2_X1 U8127 ( .A1(n14259), .A2(n14260), .ZN(n9593) );
  AND2_X1 U8128 ( .A1(n11266), .A2(n9667), .ZN(n14577) );
  AOI21_X1 U8129 ( .B1(n12518), .B2(n9664), .A(n9663), .ZN(n14548) );
  OR2_X1 U8130 ( .A1(n14841), .A2(n6434), .ZN(n9568) );
  NAND2_X1 U8131 ( .A1(n9658), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9294) );
  NOR2_X1 U8132 ( .A1(n7294), .A2(n7293), .ZN(n14656) );
  NAND2_X1 U8133 ( .A1(n15193), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7293) );
  OAI21_X1 U8134 ( .B1(n14654), .B2(P1_REG1_REG_1__SCAN_IN), .A(n7041), .ZN(
        n14663) );
  NAND2_X1 U8135 ( .A1(n14654), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7041) );
  NAND2_X1 U8136 ( .A1(n6646), .A2(n7018), .ZN(n10686) );
  INV_X1 U8137 ( .A(n10605), .ZN(n7018) );
  INV_X1 U8138 ( .A(n10604), .ZN(n6646) );
  NAND2_X1 U8139 ( .A1(n10876), .A2(n10875), .ZN(n10877) );
  NAND2_X1 U8140 ( .A1(n10877), .A2(n10878), .ZN(n11104) );
  NAND2_X1 U8141 ( .A1(n11291), .A2(n11290), .ZN(n11292) );
  NAND2_X1 U8142 ( .A1(n7285), .A2(n7284), .ZN(n11436) );
  AND2_X1 U8143 ( .A1(n6463), .A2(n11283), .ZN(n7284) );
  NAND2_X1 U8144 ( .A1(n11292), .A2(n11293), .ZN(n11443) );
  OR2_X1 U8145 ( .A1(n11715), .A2(n11716), .ZN(n12349) );
  NAND2_X1 U8146 ( .A1(n12341), .A2(n6532), .ZN(n12343) );
  NOR2_X1 U8147 ( .A1(n15304), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n15303) );
  OAI21_X1 U8148 ( .B1(n14761), .B2(n14760), .A(n7279), .ZN(n14778) );
  NAND2_X1 U8149 ( .A1(n14765), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7279) );
  NOR2_X1 U8150 ( .A1(n7489), .A2(n12435), .ZN(n14796) );
  AND2_X1 U8151 ( .A1(n9637), .A2(n9657), .ZN(n12597) );
  NAND2_X1 U8152 ( .A1(n7250), .A2(n7252), .ZN(n7247) );
  NAND2_X1 U8153 ( .A1(n14825), .A2(n6794), .ZN(n12593) );
  NOR2_X1 U8154 ( .A1(n15082), .A2(n15087), .ZN(n6794) );
  NAND2_X1 U8155 ( .A1(n14811), .A2(n14639), .ZN(n12431) );
  NAND2_X1 U8156 ( .A1(n12429), .A2(n12430), .ZN(n7249) );
  XNOR2_X1 U8157 ( .A(n14811), .B(n14639), .ZN(n14814) );
  AND2_X1 U8158 ( .A1(n8938), .A2(n8937), .ZN(n14603) );
  AND2_X1 U8159 ( .A1(n9529), .A2(n9528), .ZN(n14241) );
  NAND2_X1 U8160 ( .A1(n7064), .A2(n12454), .ZN(n14908) );
  NAND2_X1 U8161 ( .A1(n14917), .A2(n14921), .ZN(n7064) );
  OR2_X1 U8162 ( .A1(n14908), .A2(n14909), .ZN(n14911) );
  NAND2_X1 U8163 ( .A1(n14918), .A2(n14475), .ZN(n14900) );
  NOR2_X1 U8164 ( .A1(n14899), .A2(n7654), .ZN(n7653) );
  INV_X1 U8165 ( .A(n14475), .ZN(n7654) );
  NAND2_X1 U8166 ( .A1(n14946), .A2(n7245), .ZN(n14918) );
  AND2_X1 U8167 ( .A1(n9478), .A2(n9477), .ZN(n14944) );
  INV_X1 U8168 ( .A(n9444), .ZN(n9446) );
  OR2_X1 U8169 ( .A1(n14598), .A2(n14597), .ZN(n14962) );
  AND4_X1 U8170 ( .A1(n9434), .A2(n9433), .A3(n9432), .A4(n9431), .ZN(n14975)
         );
  AND3_X1 U8171 ( .A1(n9450), .A2(n9449), .A3(n9448), .ZN(n14974) );
  OR2_X1 U8172 ( .A1(n15146), .A2(n14975), .ZN(n14471) );
  INV_X1 U8173 ( .A(n15223), .ZN(n14976) );
  NAND2_X1 U8174 ( .A1(n12448), .A2(n14986), .ZN(n14997) );
  INV_X1 U8175 ( .A(n14996), .ZN(n12448) );
  NAND2_X1 U8176 ( .A1(n7612), .A2(n7614), .ZN(n12409) );
  AOI21_X1 U8177 ( .B1(n11929), .B2(n7616), .A(n7615), .ZN(n7614) );
  AND2_X1 U8178 ( .A1(n11932), .A2(n11931), .ZN(n7615) );
  AOI21_X1 U8179 ( .B1(n14592), .B2(n7736), .A(n6539), .ZN(n7735) );
  INV_X1 U8180 ( .A(n11922), .ZN(n7736) );
  NOR2_X1 U8181 ( .A1(n7737), .A2(n14590), .ZN(n7734) );
  INV_X1 U8182 ( .A(n14592), .ZN(n7737) );
  NAND2_X1 U8183 ( .A1(n8868), .A2(n8867), .ZN(n14419) );
  NAND2_X1 U8184 ( .A1(n15324), .A2(n7611), .ZN(n6782) );
  XNOR2_X1 U8185 ( .A(n14652), .B(n11629), .ZN(n14584) );
  INV_X1 U8186 ( .A(n15052), .ZN(n15222) );
  NAND2_X1 U8187 ( .A1(n14176), .A2(n8948), .ZN(n8944) );
  NAND2_X1 U8188 ( .A1(n6786), .A2(n7631), .ZN(n14845) );
  NAND2_X1 U8189 ( .A1(n14869), .A2(n7629), .ZN(n6786) );
  NAND2_X1 U8190 ( .A1(n11613), .A2(n8948), .ZN(n6735) );
  INV_X1 U8191 ( .A(n15395), .ZN(n15404) );
  OAI21_X1 U8192 ( .B1(n8683), .B2(n8682), .A(n8681), .ZN(n8717) );
  AOI21_X1 U8193 ( .B1(n7345), .B2(n7343), .A(n7342), .ZN(n7341) );
  INV_X1 U8194 ( .A(n8687), .ZN(n7342) );
  INV_X1 U8195 ( .A(n8716), .ZN(n7343) );
  INV_X1 U8196 ( .A(n7345), .ZN(n7344) );
  XNOR2_X1 U8197 ( .A(n8826), .B(n8825), .ZN(n8969) );
  NAND2_X1 U8198 ( .A1(n8962), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8826) );
  XNOR2_X1 U8199 ( .A(n8453), .B(n8446), .ZN(n14183) );
  NOR2_X1 U8200 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6698) );
  NOR2_X1 U8201 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6697) );
  XNOR2_X1 U8202 ( .A(n8216), .B(n8215), .ZN(n11302) );
  OAI21_X1 U8203 ( .B1(n8213), .B2(n8212), .A(n8211), .ZN(n8216) );
  NAND2_X1 U8204 ( .A1(n8874), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U8205 ( .A1(n7955), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7927) );
  AND2_X1 U8206 ( .A1(n8831), .A2(n6641), .ZN(n8845) );
  NOR2_X1 U8207 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7296) );
  XNOR2_X1 U8208 ( .A(n9129), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n9143) );
  INV_X1 U8209 ( .A(n6809), .ZN(n9152) );
  NAND2_X1 U8210 ( .A1(n9107), .A2(n9108), .ZN(n9151) );
  OR2_X1 U8211 ( .A1(n9146), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U8212 ( .A1(n7081), .A2(n9117), .ZN(n9160) );
  NAND2_X1 U8213 ( .A1(n9158), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n7081) );
  INV_X1 U8214 ( .A(n15273), .ZN(n6815) );
  AOI22_X1 U8215 ( .A1(n9122), .A2(n9120), .B1(P3_ADDR_REG_13__SCAN_IN), .B2(
        n9121), .ZN(n9163) );
  AND4_X1 U8216 ( .A1(n9853), .A2(n9852), .A3(n9851), .A4(n9850), .ZN(n12843)
         );
  AND3_X1 U8217 ( .A1(n9779), .A2(n9778), .A3(n9777), .ZN(n11498) );
  OAI21_X1 U8218 ( .B1(n12727), .B2(n6890), .A(n6889), .ZN(n6891) );
  AOI21_X1 U8219 ( .B1(n12612), .B2(n12485), .A(n12489), .ZN(n6889) );
  INV_X1 U8220 ( .A(n12612), .ZN(n6890) );
  NAND2_X1 U8221 ( .A1(n9742), .A2(n7730), .ZN(n11047) );
  OAI21_X1 U8222 ( .B1(n7731), .B2(n7732), .A(n10911), .ZN(n7730) );
  NOR2_X1 U8223 ( .A1(n9755), .A2(n10414), .ZN(n7731) );
  AND2_X1 U8224 ( .A1(n10188), .A2(n10187), .ZN(n13238) );
  NAND2_X1 U8225 ( .A1(n7454), .A2(n10034), .ZN(n12680) );
  NAND2_X1 U8226 ( .A1(n12740), .A2(n10033), .ZN(n7454) );
  AOI21_X1 U8227 ( .B1(n13258), .B2(n12093), .A(n10133), .ZN(n13283) );
  AND2_X1 U8228 ( .A1(n10171), .A2(n10170), .ZN(n13227) );
  NAND2_X1 U8229 ( .A1(n7188), .A2(n7926), .ZN(n9765) );
  NAND2_X1 U8230 ( .A1(n15577), .A2(n10230), .ZN(n12720) );
  AND2_X1 U8231 ( .A1(n10240), .A2(n10239), .ZN(n13228) );
  OR3_X1 U8232 ( .A1(n12953), .A2(n10356), .A3(n10243), .ZN(n12733) );
  AND3_X1 U8233 ( .A1(n10048), .A2(n10047), .A3(n10046), .ZN(n13337) );
  OR3_X1 U8234 ( .A1(n12953), .A2(n10241), .A3(n10243), .ZN(n12743) );
  NAND2_X1 U8235 ( .A1(n10249), .A2(n10248), .ZN(n12747) );
  NAND2_X1 U8236 ( .A1(n6854), .A2(n7102), .ZN(n6853) );
  NAND2_X1 U8237 ( .A1(n7103), .A2(n15575), .ZN(n7102) );
  NAND2_X1 U8238 ( .A1(n6860), .A2(n6859), .ZN(n6854) );
  INV_X1 U8239 ( .A(n12800), .ZN(n6859) );
  INV_X1 U8240 ( .A(n13283), .ZN(n13252) );
  NAND2_X1 U8241 ( .A1(n10119), .A2(n10118), .ZN(n13294) );
  INV_X1 U8242 ( .A(n15581), .ZN(n12979) );
  NAND2_X1 U8243 ( .A1(n10964), .A2(n10963), .ZN(n11030) );
  NAND2_X1 U8244 ( .A1(n10991), .A2(n10932), .ZN(n11083) );
  NAND2_X1 U8245 ( .A1(n7516), .A2(n11124), .ZN(n11128) );
  NAND2_X1 U8246 ( .A1(n11126), .A2(n11125), .ZN(n7516) );
  NAND2_X1 U8247 ( .A1(n11069), .A2(n11070), .ZN(n11216) );
  NAND2_X1 U8248 ( .A1(n7101), .A2(n11071), .ZN(n11069) );
  NAND2_X1 U8249 ( .A1(n7089), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13111) );
  INV_X1 U8250 ( .A(n13088), .ZN(n7089) );
  NAND2_X1 U8251 ( .A1(n6829), .A2(n13122), .ZN(n6828) );
  XNOR2_X1 U8252 ( .A(n13117), .B(n13403), .ZN(n6829) );
  NOR2_X1 U8253 ( .A1(n13099), .A2(n6825), .ZN(n6824) );
  INV_X1 U8254 ( .A(n6826), .ZN(n6825) );
  AOI21_X1 U8255 ( .B1(n13100), .B2(n13116), .A(n6827), .ZN(n6826) );
  XNOR2_X1 U8256 ( .A(n13141), .B(n13142), .ZN(n7329) );
  INV_X1 U8257 ( .A(n6657), .ZN(n6656) );
  OAI211_X1 U8258 ( .C1(n13133), .C2(n7499), .A(n7495), .B(n13112), .ZN(n6657)
         );
  AND2_X1 U8259 ( .A1(n7501), .A2(n13127), .ZN(n7499) );
  OR2_X1 U8260 ( .A1(n13088), .A2(n7496), .ZN(n7495) );
  NAND2_X1 U8261 ( .A1(n6568), .A2(n7500), .ZN(n7494) );
  AND2_X1 U8262 ( .A1(n13133), .A2(n13127), .ZN(n7498) );
  NAND2_X1 U8263 ( .A1(n10360), .A2(n10359), .ZN(n13184) );
  NOR2_X1 U8264 ( .A1(n10358), .A2(n10357), .ZN(n10359) );
  NOR2_X1 U8265 ( .A1(n13212), .A2(n15582), .ZN(n10357) );
  OAI21_X1 U8266 ( .B1(n7036), .B2(n15601), .A(n7034), .ZN(n13371) );
  INV_X1 U8267 ( .A(n7035), .ZN(n7034) );
  XNOR2_X1 U8268 ( .A(n13199), .B(n13192), .ZN(n7036) );
  OAI22_X1 U8269 ( .A1(n13193), .A2(n15580), .B1(n15582), .B2(n13228), .ZN(
        n7035) );
  NAND2_X1 U8270 ( .A1(n10181), .A2(n10180), .ZN(n13223) );
  NAND2_X1 U8271 ( .A1(n10112), .A2(n10111), .ZN(n13391) );
  INV_X1 U8272 ( .A(n12559), .ZN(n7198) );
  INV_X1 U8273 ( .A(n13416), .ZN(n13382) );
  INV_X1 U8274 ( .A(n12939), .ZN(n12545) );
  INV_X1 U8275 ( .A(n6850), .ZN(n13187) );
  NAND2_X1 U8276 ( .A1(n10128), .A2(n10127), .ZN(n13457) );
  NAND2_X1 U8277 ( .A1(n11650), .A2(n12758), .ZN(n10128) );
  NAND2_X1 U8278 ( .A1(n10004), .A2(n10003), .ZN(n13487) );
  NAND2_X1 U8279 ( .A1(n9964), .A2(n9963), .ZN(n12665) );
  NAND2_X1 U8280 ( .A1(n9910), .A2(n9909), .ZN(n12069) );
  OR2_X1 U8281 ( .A1(n15643), .A2(n15638), .ZN(n13443) );
  OR2_X1 U8282 ( .A1(n9732), .A2(n13502), .ZN(n7682) );
  AND2_X1 U8283 ( .A1(n9734), .A2(n9720), .ZN(n9732) );
  XNOR2_X1 U8284 ( .A(n10201), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12957) );
  NAND2_X1 U8285 ( .A1(n6892), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U8286 ( .A1(n10039), .A2(n6537), .ZN(n6892) );
  NAND2_X1 U8287 ( .A1(n6650), .A2(n6455), .ZN(n9205) );
  NAND2_X1 U8288 ( .A1(n13565), .A2(n6505), .ZN(n6650) );
  NAND2_X1 U8289 ( .A1(n8348), .A2(n8347), .ZN(n13541) );
  AND2_X1 U8290 ( .A1(n8554), .A2(n6503), .ZN(n6649) );
  NAND2_X1 U8291 ( .A1(n14176), .A2(n8718), .ZN(n8479) );
  NAND2_X1 U8292 ( .A1(n9205), .A2(n9204), .ZN(n9203) );
  NAND2_X1 U8293 ( .A1(n7535), .A2(n7536), .ZN(n6648) );
  NAND2_X1 U8294 ( .A1(n11187), .A2(n7556), .ZN(n7553) );
  NOR2_X1 U8295 ( .A1(n11179), .A2(n7557), .ZN(n7556) );
  INV_X1 U8296 ( .A(n7919), .ZN(n7557) );
  NAND2_X1 U8297 ( .A1(n8152), .A2(n8151), .ZN(n14089) );
  AND2_X1 U8298 ( .A1(n8288), .A2(n8287), .ZN(n13859) );
  AND2_X1 U8299 ( .A1(n10631), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13631) );
  INV_X1 U8300 ( .A(n13610), .ZN(n13649) );
  INV_X1 U8301 ( .A(n13631), .ZN(n13645) );
  OR2_X1 U8302 ( .A1(n13749), .A2(n8424), .ZN(n8465) );
  OR2_X1 U8303 ( .A1(n13782), .A2(n8424), .ZN(n8429) );
  AOI21_X1 U8304 ( .B1(n6947), .B2(P2_REG1_REG_17__SCAN_IN), .A(n7768), .ZN(
        n8243) );
  AND4_X1 U8305 ( .A1(n8177), .A2(n8176), .A3(n8175), .A4(n8174), .ZN(n13659)
         );
  NAND2_X1 U8306 ( .A1(n8282), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7889) );
  INV_X1 U8307 ( .A(n6667), .ZN(n15453) );
  NAND2_X1 U8308 ( .A1(n15470), .A2(n10526), .ZN(n10527) );
  AOI21_X1 U8309 ( .B1(n13702), .B2(n15508), .A(n13705), .ZN(n6679) );
  NAND2_X1 U8310 ( .A1(n13704), .A2(n15471), .ZN(n6682) );
  NOR2_X1 U8311 ( .A1(n13703), .A2(n7028), .ZN(n7027) );
  NAND2_X1 U8312 ( .A1(n12570), .A2(n12569), .ZN(n13710) );
  XNOR2_X1 U8313 ( .A(n13711), .B(n14116), .ZN(n12570) );
  INV_X1 U8314 ( .A(n14007), .ZN(n14004) );
  XNOR2_X1 U8315 ( .A(n14007), .B(n6761), .ZN(n9201) );
  INV_X1 U8316 ( .A(n14008), .ZN(n6761) );
  NAND2_X1 U8317 ( .A1(n6759), .A2(n9086), .ZN(n9189) );
  AND2_X1 U8318 ( .A1(n8484), .A2(n8483), .ZN(n9190) );
  NAND2_X1 U8319 ( .A1(n7678), .A2(n7679), .ZN(n13891) );
  OR2_X1 U8320 ( .A1(n7948), .A2(n10468), .ZN(n7912) );
  NAND2_X1 U8321 ( .A1(n14041), .A2(n6977), .ZN(n14128) );
  INV_X1 U8322 ( .A(n6978), .ZN(n6977) );
  OAI21_X1 U8323 ( .B1(n14042), .B2(n15557), .A(n14040), .ZN(n6978) );
  NAND2_X1 U8324 ( .A1(n13710), .A2(n14000), .ZN(n14115) );
  NAND2_X1 U8325 ( .A1(n14180), .A2(n8718), .ZN(n8456) );
  NAND2_X1 U8326 ( .A1(n14024), .A2(n7182), .ZN(n14120) );
  AND2_X1 U8327 ( .A1(n14023), .A2(n14022), .ZN(n7182) );
  NAND2_X1 U8328 ( .A1(n14038), .A2(n6518), .ZN(n14127) );
  OR2_X1 U8329 ( .A1(n14039), .A2(n15557), .ZN(n7773) );
  NAND2_X1 U8330 ( .A1(n14128), .A2(n15561), .ZN(n6976) );
  NAND2_X1 U8331 ( .A1(n8902), .A2(n8901), .ZN(n15151) );
  NAND2_X1 U8332 ( .A1(n12134), .A2(n8948), .ZN(n8934) );
  NAND2_X1 U8333 ( .A1(n14214), .A2(n14213), .ZN(n14212) );
  AND2_X1 U8334 ( .A1(n9491), .A2(n9490), .ZN(n14923) );
  AND3_X1 U8335 ( .A1(n9466), .A2(n9465), .A3(n9464), .ZN(n14957) );
  NAND2_X1 U8336 ( .A1(n6705), .A2(n9443), .ZN(n14290) );
  NAND2_X1 U8337 ( .A1(n11708), .A2(n8948), .ZN(n8928) );
  AND3_X1 U8338 ( .A1(n9665), .A2(n14577), .A3(n11263), .ZN(n14368) );
  AND2_X1 U8339 ( .A1(n9633), .A2(n11263), .ZN(n14370) );
  INV_X1 U8340 ( .A(n14560), .ZN(n14627) );
  NAND2_X1 U8341 ( .A1(n6733), .A2(n14567), .ZN(n14632) );
  NAND2_X1 U8342 ( .A1(n14551), .A2(n6528), .ZN(n6733) );
  INV_X1 U8343 ( .A(n14365), .ZN(n14638) );
  NAND2_X1 U8344 ( .A1(n9584), .A2(n9583), .ZN(n14640) );
  NAND2_X1 U8345 ( .A1(n9546), .A2(n9545), .ZN(n14871) );
  NAND2_X1 U8346 ( .A1(n9514), .A2(n9513), .ZN(n14870) );
  INV_X1 U8347 ( .A(n14923), .ZN(n14643) );
  AND4_X1 U8348 ( .A1(n9227), .A2(n9226), .A3(n9225), .A4(n9224), .ZN(n11949)
         );
  OAI21_X1 U8349 ( .B1(n14786), .B2(n6633), .A(n6460), .ZN(n7280) );
  NOR2_X1 U8350 ( .A1(n14783), .A2(n14958), .ZN(n7282) );
  OR2_X1 U8351 ( .A1(n14784), .A2(n15305), .ZN(n7281) );
  NAND2_X1 U8352 ( .A1(n8951), .A2(n8950), .ZN(n14534) );
  INV_X1 U8353 ( .A(n15325), .ZN(n15024) );
  INV_X1 U8354 ( .A(n15090), .ZN(n7751) );
  AOI211_X1 U8355 ( .C1(n15087), .C2(n14807), .A(n15365), .B(n14806), .ZN(
        n15086) );
  OR2_X1 U8356 ( .A1(n8843), .A2(n14675), .ZN(n7052) );
  INV_X1 U8357 ( .A(n7051), .ZN(n7050) );
  OAI22_X1 U8358 ( .A1(n10467), .A2(n8949), .B1(n8859), .B2(n10468), .ZN(n7051) );
  NOR2_X1 U8359 ( .A1(n15072), .A2(n15071), .ZN(n6796) );
  NAND2_X1 U8360 ( .A1(n15067), .A2(n15395), .ZN(n7055) );
  OAI21_X1 U8361 ( .B1(n15659), .B2(n15658), .A(n6485), .ZN(n6812) );
  NAND2_X1 U8362 ( .A1(n15208), .A2(n6955), .ZN(n15213) );
  OAI21_X1 U8363 ( .B1(n15209), .B2(n15210), .A(P2_ADDR_REG_9__SCAN_IN), .ZN(
        n6955) );
  NAND2_X1 U8364 ( .A1(n6803), .A2(n15215), .ZN(n7609) );
  NAND2_X1 U8365 ( .A1(n15213), .A2(n15214), .ZN(n6803) );
  NAND2_X1 U8366 ( .A1(n6802), .A2(n6806), .ZN(n7610) );
  INV_X1 U8367 ( .A(n15213), .ZN(n6802) );
  XNOR2_X1 U8368 ( .A(n9160), .B(n9159), .ZN(n15267) );
  XNOR2_X1 U8369 ( .A(n9162), .B(n9161), .ZN(n15271) );
  NAND2_X1 U8370 ( .A1(n7082), .A2(n6815), .ZN(n6814) );
  OAI21_X1 U8371 ( .B1(n7601), .B2(n6552), .A(n7083), .ZN(n15286) );
  NAND2_X1 U8372 ( .A1(n9168), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U8373 ( .A1(n6801), .A2(n7602), .ZN(n9181) );
  NAND2_X1 U8374 ( .A1(n15247), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7602) );
  XNOR2_X1 U8375 ( .A(n9186), .B(n7332), .ZN(n9188) );
  XNOR2_X1 U8376 ( .A(n9181), .B(n9180), .ZN(n15195) );
  NOR2_X1 U8377 ( .A1(n7435), .A2(n7611), .ZN(n7434) );
  AOI21_X1 U8378 ( .B1(n8790), .B2(n8707), .A(n8566), .ZN(n8574) );
  OR2_X1 U8379 ( .A1(n8585), .A2(n8584), .ZN(n8586) );
  NAND2_X1 U8380 ( .A1(n14414), .A2(n14417), .ZN(n7478) );
  AOI22_X1 U8381 ( .A1(n13666), .A2(n8770), .B1(n15552), .B2(n8707), .ZN(n8600) );
  OAI21_X1 U8382 ( .B1(n12813), .B2(n7128), .A(n7131), .ZN(n7127) );
  OAI211_X1 U8383 ( .C1(n6928), .C2(n12802), .A(n12805), .B(n7148), .ZN(n12810) );
  AOI21_X1 U8384 ( .B1(n10998), .B2(n6928), .A(n7149), .ZN(n7148) );
  NAND2_X1 U8385 ( .A1(n6717), .A2(n6716), .ZN(n14431) );
  NAND2_X1 U8386 ( .A1(n14425), .A2(n14427), .ZN(n6716) );
  INV_X1 U8387 ( .A(n8604), .ZN(n6961) );
  NAND2_X1 U8388 ( .A1(n14431), .A2(n14432), .ZN(n14430) );
  INV_X1 U8389 ( .A(n14440), .ZN(n7444) );
  INV_X1 U8390 ( .A(n14441), .ZN(n7443) );
  NAND2_X1 U8391 ( .A1(n7129), .A2(n12825), .ZN(n7124) );
  NOR2_X1 U8392 ( .A1(n7442), .A2(n7441), .ZN(n7440) );
  NOR2_X1 U8393 ( .A1(n14440), .A2(n14441), .ZN(n7441) );
  NOR2_X1 U8394 ( .A1(n14448), .A2(n14447), .ZN(n7442) );
  AND2_X1 U8395 ( .A1(n8613), .A2(n8612), .ZN(n6912) );
  NAND2_X1 U8396 ( .A1(n7147), .A2(n12862), .ZN(n7146) );
  NAND2_X1 U8397 ( .A1(n12859), .A2(n6504), .ZN(n7147) );
  OR3_X1 U8398 ( .A1(n14921), .A2(n14498), .A3(n14497), .ZN(n14499) );
  NAND2_X1 U8399 ( .A1(n12884), .A2(n7121), .ZN(n7115) );
  INV_X1 U8400 ( .A(n12882), .ZN(n7121) );
  AOI21_X1 U8401 ( .B1(n12876), .B2(n7123), .A(n12880), .ZN(n7122) );
  NAND2_X1 U8402 ( .A1(n8631), .A2(n8630), .ZN(n7627) );
  OR2_X1 U8403 ( .A1(n8631), .A2(n8630), .ZN(n7626) );
  NAND2_X1 U8404 ( .A1(n7143), .A2(n7142), .ZN(n12873) );
  INV_X1 U8405 ( .A(n7109), .ZN(n7108) );
  OAI22_X1 U8406 ( .A1(n7122), .A2(n7111), .B1(n7116), .B2(n7110), .ZN(n7109)
         );
  INV_X1 U8407 ( .A(n7115), .ZN(n7111) );
  NAND2_X1 U8408 ( .A1(n7115), .A2(n7118), .ZN(n7110) );
  NAND2_X1 U8409 ( .A1(n7106), .A2(n7115), .ZN(n7114) );
  NAND2_X1 U8410 ( .A1(n7122), .A2(n7107), .ZN(n7106) );
  NAND2_X1 U8411 ( .A1(n7117), .A2(n7118), .ZN(n7107) );
  INV_X1 U8412 ( .A(n7120), .ZN(n7119) );
  AOI21_X1 U8413 ( .B1(n7122), .B2(n13334), .A(n7121), .ZN(n7120) );
  NAND2_X1 U8414 ( .A1(n12915), .A2(n12916), .ZN(n7141) );
  MUX2_X1 U8415 ( .A(n12914), .B(n12913), .S(n12946), .Z(n12915) );
  NAND2_X1 U8416 ( .A1(n14511), .A2(n14513), .ZN(n6731) );
  NAND2_X1 U8417 ( .A1(n14518), .A2(n7447), .ZN(n7446) );
  INV_X1 U8418 ( .A(n14517), .ZN(n7447) );
  INV_X1 U8419 ( .A(n13224), .ZN(n7140) );
  NAND2_X1 U8420 ( .A1(n6900), .A2(n8651), .ZN(n6899) );
  NAND2_X1 U8421 ( .A1(n6490), .A2(n6902), .ZN(n6901) );
  INV_X1 U8422 ( .A(n8652), .ZN(n6900) );
  AOI21_X1 U8423 ( .B1(n7642), .B2(n7644), .A(n8657), .ZN(n7641) );
  INV_X1 U8424 ( .A(n7647), .ZN(n7639) );
  INV_X1 U8425 ( .A(n8338), .ZN(n7354) );
  NOR2_X1 U8426 ( .A1(n6840), .A2(n6739), .ZN(n6738) );
  INV_X1 U8427 ( .A(n7997), .ZN(n6739) );
  OR2_X1 U8428 ( .A1(n7211), .A2(n10345), .ZN(n7208) );
  NOR2_X1 U8429 ( .A1(n12782), .A2(n13195), .ZN(n6881) );
  NAND2_X1 U8430 ( .A1(n7206), .A2(n10346), .ZN(n7204) );
  OR2_X1 U8431 ( .A1(n13228), .A2(n13376), .ZN(n12926) );
  NOR2_X1 U8432 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7685) );
  NOR2_X1 U8433 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7686) );
  NOR2_X1 U8434 ( .A1(n11969), .A2(n7779), .ZN(n7778) );
  INV_X1 U8435 ( .A(n9056), .ZN(n7779) );
  AND2_X1 U8436 ( .A1(n14581), .A2(n7611), .ZN(n14585) );
  AOI21_X1 U8437 ( .B1(n7335), .B2(n8189), .A(n6559), .ZN(n7334) );
  INV_X1 U8438 ( .A(n7337), .ZN(n7335) );
  INV_X1 U8439 ( .A(n8189), .ZN(n7336) );
  INV_X1 U8440 ( .A(n7185), .ZN(n7184) );
  OAI21_X1 U8441 ( .B1(n6443), .B2(n7186), .A(n8161), .ZN(n7185) );
  AND2_X1 U8442 ( .A1(n8037), .A2(n8034), .ZN(n6838) );
  OAI21_X1 U8443 ( .B1(n7859), .B2(P1_DATAO_REG_6__SCAN_IN), .A(n6779), .ZN(
        n8011) );
  NAND2_X1 U8444 ( .A1(n7859), .A2(n10439), .ZN(n6779) );
  INV_X1 U8445 ( .A(n7975), .ZN(n7167) );
  INV_X1 U8446 ( .A(n7994), .ZN(n6845) );
  AND2_X1 U8447 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n9141), .ZN(n7596) );
  NAND2_X1 U8448 ( .A1(n7598), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n7597) );
  INV_X1 U8449 ( .A(n9103), .ZN(n7598) );
  INV_X1 U8450 ( .A(n10155), .ZN(n7420) );
  NAND2_X1 U8451 ( .A1(n6928), .A2(n12952), .ZN(n6927) );
  INV_X1 U8452 ( .A(n11041), .ZN(n12487) );
  INV_X1 U8453 ( .A(n10034), .ZN(n7453) );
  NAND2_X1 U8454 ( .A1(n6886), .A2(n6885), .ZN(n6884) );
  INV_X1 U8455 ( .A(n10197), .ZN(n6885) );
  INV_X1 U8456 ( .A(n10196), .ZN(n6886) );
  NOR4_X1 U8457 ( .A1(n13235), .A2(n13249), .A3(n13292), .A4(n12779), .ZN(
        n12780) );
  NAND2_X1 U8458 ( .A1(n9763), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10942) );
  NAND2_X1 U8459 ( .A1(n10980), .A2(n10902), .ZN(n10903) );
  OR2_X1 U8460 ( .A1(n10948), .A2(n11056), .ZN(n10949) );
  NOR2_X1 U8461 ( .A1(n6444), .A2(n7325), .ZN(n7321) );
  NAND2_X1 U8462 ( .A1(n13090), .A2(n7319), .ZN(n13114) );
  OR2_X1 U8463 ( .A1(n13091), .A2(n13407), .ZN(n7319) );
  NAND2_X1 U8464 ( .A1(n7504), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7503) );
  INV_X1 U8465 ( .A(n7208), .ZN(n7207) );
  OAI21_X1 U8466 ( .B1(n7208), .B2(n12782), .A(n7209), .ZN(n7206) );
  NAND2_X1 U8467 ( .A1(n13212), .A2(n13433), .ZN(n7209) );
  NOR2_X1 U8468 ( .A1(n13193), .A2(n6849), .ZN(n6848) );
  INV_X1 U8469 ( .A(n10295), .ZN(n6849) );
  NOR2_X1 U8470 ( .A1(n10182), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U8471 ( .A1(n11506), .A2(n10320), .ZN(n11761) );
  NAND2_X1 U8472 ( .A1(n11761), .A2(n7717), .ZN(n11795) );
  INV_X1 U8473 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9823) );
  INV_X1 U8474 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9802) );
  NOR2_X1 U8475 ( .A1(n7215), .A2(n10342), .ZN(n7213) );
  NOR2_X1 U8476 ( .A1(n10341), .A2(n7216), .ZN(n7215) );
  INV_X1 U8477 ( .A(n10343), .ZN(n7216) );
  AND2_X1 U8478 ( .A1(n7791), .A2(n10343), .ZN(n7217) );
  OR2_X1 U8479 ( .A1(n13451), .A2(n13264), .ZN(n12914) );
  AND2_X1 U8480 ( .A1(n10265), .A2(n12893), .ZN(n12885) );
  INV_X1 U8481 ( .A(n13344), .ZN(n13350) );
  OR2_X1 U8482 ( .A1(n12381), .A2(n6572), .ZN(n13349) );
  NAND2_X1 U8483 ( .A1(n7717), .A2(n7803), .ZN(n7802) );
  INV_X1 U8484 ( .A(n10320), .ZN(n7803) );
  INV_X1 U8485 ( .A(n10319), .ZN(n7195) );
  NAND2_X1 U8486 ( .A1(n7193), .A2(n7801), .ZN(n7192) );
  OR2_X1 U8487 ( .A1(n12252), .A2(n12973), .ZN(n12860) );
  NOR2_X1 U8488 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7412) );
  NOR2_X1 U8489 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n7411) );
  INV_X1 U8490 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7105) );
  INV_X1 U8491 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7104) );
  INV_X1 U8492 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n10223) );
  OAI21_X1 U8493 ( .B1(P1_DATAO_REG_20__SCAN_IN), .B2(n11710), .A(n10140), 
        .ZN(n10137) );
  INV_X1 U8494 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9684) );
  INV_X1 U8495 ( .A(n9957), .ZN(n6875) );
  INV_X1 U8496 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9693) );
  INV_X1 U8497 ( .A(n9695), .ZN(n9682) );
  AOI21_X1 U8498 ( .B1(n7584), .B2(n9898), .A(n7583), .ZN(n7582) );
  NAND2_X1 U8499 ( .A1(n7584), .A2(n6865), .ZN(n6864) );
  INV_X1 U8500 ( .A(n9919), .ZN(n7583) );
  INV_X1 U8501 ( .A(n7584), .ZN(n6866) );
  OAI21_X1 U8502 ( .B1(n7579), .B2(n6879), .A(n9772), .ZN(n7578) );
  NAND2_X1 U8503 ( .A1(n10467), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6879) );
  INV_X1 U8504 ( .A(n13583), .ZN(n7550) );
  NOR2_X1 U8505 ( .A1(n6472), .A2(n13593), .ZN(n8420) );
  NOR2_X1 U8506 ( .A1(n8101), .A2(n6695), .ZN(n6694) );
  NOR2_X1 U8507 ( .A1(n8205), .A2(n12390), .ZN(n6996) );
  NOR2_X1 U8508 ( .A1(n8661), .A2(n8660), .ZN(n8680) );
  NAND2_X1 U8509 ( .A1(n6934), .A2(n6933), .ZN(n7016) );
  INV_X1 U8510 ( .A(n8659), .ZN(n6933) );
  NAND2_X1 U8511 ( .A1(n8661), .A2(n8660), .ZN(n6934) );
  AND2_X1 U8512 ( .A1(n8771), .A2(n8699), .ZN(n8783) );
  INV_X1 U8513 ( .A(n14016), .ZN(n7405) );
  INV_X1 U8514 ( .A(n7834), .ZN(n7667) );
  NAND2_X1 U8515 ( .A1(n13751), .A2(n13760), .ZN(n7669) );
  INV_X1 U8516 ( .A(n7835), .ZN(n7668) );
  AOI21_X1 U8517 ( .B1(n9078), .B2(n7270), .A(n7269), .ZN(n7268) );
  INV_X1 U8518 ( .A(n9079), .ZN(n7269) );
  INV_X1 U8519 ( .A(n9075), .ZN(n7270) );
  INV_X1 U8520 ( .A(n9078), .ZN(n7271) );
  INV_X1 U8521 ( .A(n9035), .ZN(n7664) );
  NAND2_X1 U8522 ( .A1(n7176), .A2(n13838), .ZN(n7174) );
  NOR2_X1 U8523 ( .A1(n13831), .A2(n7410), .ZN(n7409) );
  NOR2_X1 U8524 ( .A1(n8308), .A2(n8307), .ZN(n6995) );
  NAND2_X1 U8525 ( .A1(n13941), .A2(n13641), .ZN(n6766) );
  INV_X1 U8526 ( .A(n6693), .ZN(n8263) );
  NAND2_X1 U8527 ( .A1(n6996), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U8528 ( .A1(n7172), .A2(n13931), .ZN(n13910) );
  INV_X1 U8529 ( .A(n9060), .ZN(n7762) );
  AND2_X1 U8530 ( .A1(n12298), .A2(n12303), .ZN(n12299) );
  OR2_X1 U8531 ( .A1(n8076), .A2(n11755), .ZN(n8101) );
  NAND2_X1 U8532 ( .A1(n11980), .A2(n6507), .ZN(n11962) );
  AND2_X1 U8533 ( .A1(n12011), .A2(n12015), .ZN(n11980) );
  AND2_X1 U8534 ( .A1(n8536), .A2(n12562), .ZN(n10632) );
  AND2_X1 U8535 ( .A1(n9039), .A2(n11770), .ZN(n8536) );
  NAND2_X1 U8536 ( .A1(n6489), .A2(n6639), .ZN(n13719) );
  NAND2_X1 U8537 ( .A1(n13758), .A2(n7273), .ZN(n6639) );
  AND2_X1 U8538 ( .A1(n14008), .A2(n9085), .ZN(n9082) );
  INV_X1 U8539 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7875) );
  AND2_X1 U8540 ( .A1(n8495), .A2(n8494), .ZN(n8501) );
  INV_X1 U8541 ( .A(n8493), .ZN(n8495) );
  NAND2_X1 U8542 ( .A1(n7843), .A2(n6658), .ZN(n7871) );
  AND2_X1 U8543 ( .A1(n7867), .A2(n7866), .ZN(n6658) );
  NOR2_X1 U8544 ( .A1(n9368), .A2(n9367), .ZN(n9385) );
  NOR2_X1 U8545 ( .A1(n9400), .A2(n11725), .ZN(n9415) );
  NOR2_X1 U8546 ( .A1(n9471), .A2(n9470), .ZN(n7046) );
  OAI21_X1 U8547 ( .B1(n10396), .B2(n10397), .A(n9287), .ZN(n7378) );
  AND2_X1 U8548 ( .A1(n9587), .A2(n9586), .ZN(n9589) );
  OR2_X1 U8549 ( .A1(n14603), .A2(n9284), .ZN(n9587) );
  NAND2_X1 U8550 ( .A1(n7473), .A2(n14529), .ZN(n7468) );
  NAND2_X1 U8551 ( .A1(n7471), .A2(n7470), .ZN(n7469) );
  INV_X1 U8552 ( .A(n14523), .ZN(n7470) );
  INV_X1 U8553 ( .A(n14524), .ZN(n7471) );
  NAND2_X1 U8554 ( .A1(n6744), .A2(n14521), .ZN(n6743) );
  NAND2_X1 U8555 ( .A1(n7457), .A2(n14387), .ZN(n14540) );
  AND2_X1 U8556 ( .A1(n7318), .A2(n14706), .ZN(n7312) );
  AOI21_X1 U8557 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14765), .A(n14764), .ZN(
        n14774) );
  NAND2_X1 U8558 ( .A1(n7254), .A2(n7253), .ZN(n7252) );
  INV_X1 U8559 ( .A(n12430), .ZN(n7253) );
  AOI21_X1 U8560 ( .B1(n7254), .B2(n12428), .A(n7251), .ZN(n7250) );
  INV_X1 U8561 ( .A(n12587), .ZN(n7251) );
  INV_X1 U8562 ( .A(n7753), .ZN(n7071) );
  NOR2_X1 U8563 ( .A1(n12462), .A2(n7255), .ZN(n7254) );
  INV_X1 U8564 ( .A(n12431), .ZN(n7255) );
  NOR2_X1 U8565 ( .A1(n9430), .A2(n9416), .ZN(n9444) );
  NAND2_X1 U8566 ( .A1(n15146), .A2(n14975), .ZN(n14466) );
  INV_X1 U8567 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9367) );
  INV_X1 U8568 ( .A(n9385), .ZN(n9387) );
  INV_X1 U8569 ( .A(n7618), .ZN(n7616) );
  INV_X1 U8570 ( .A(n11928), .ZN(n11929) );
  AND2_X1 U8571 ( .A1(n6586), .A2(n8302), .ZN(n7355) );
  NAND2_X1 U8572 ( .A1(n8954), .A2(n8953), .ZN(n8985) );
  INV_X1 U8573 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7474) );
  INV_X1 U8574 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7238) );
  NAND2_X1 U8575 ( .A1(n6776), .A2(n8234), .ZN(n6775) );
  INV_X1 U8576 ( .A(n8250), .ZN(n6776) );
  NAND2_X1 U8577 ( .A1(n6769), .A2(n8189), .ZN(n8252) );
  INV_X1 U8578 ( .A(n6768), .ZN(n6767) );
  NAND2_X1 U8579 ( .A1(n8251), .A2(n8186), .ZN(n8214) );
  NAND2_X1 U8580 ( .A1(n7187), .A2(n6443), .ZN(n8145) );
  NAND2_X1 U8581 ( .A1(n8140), .A2(n8114), .ZN(n8120) );
  NAND2_X1 U8582 ( .A1(n8113), .A2(SI_12_), .ZN(n8114) );
  XNOR2_X1 U8583 ( .A(n8089), .B(SI_10_), .ZN(n8086) );
  XNOR2_X1 U8584 ( .A(n8033), .B(SI_7_), .ZN(n8030) );
  NOR2_X1 U8585 ( .A1(n8905), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6913) );
  INV_X1 U8586 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7331) );
  NAND2_X1 U8587 ( .A1(n9096), .A2(n7001), .ZN(n9131) );
  NAND2_X1 U8588 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7002), .ZN(n7001) );
  INV_X1 U8589 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7002) );
  XOR2_X1 U8590 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n11022), .Z(n9130) );
  OAI21_X1 U8591 ( .B1(n9129), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9105), .ZN(
        n9106) );
  XNOR2_X1 U8592 ( .A(n9106), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U8593 ( .A1(n9109), .A2(n7086), .ZN(n9110) );
  NAND2_X1 U8594 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n7087), .ZN(n7086) );
  NAND2_X1 U8595 ( .A1(n9151), .A2(n9150), .ZN(n9109) );
  INV_X1 U8596 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7087) );
  AND2_X1 U8597 ( .A1(n7608), .A2(n6805), .ZN(n6804) );
  NAND2_X1 U8598 ( .A1(n6806), .A2(n15215), .ZN(n6805) );
  OR2_X1 U8599 ( .A1(n15267), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7608) );
  OAI21_X1 U8600 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n11817), .A(n9118), .ZN(
        n9125) );
  OAI21_X1 U8601 ( .B1(n9175), .B2(n9174), .A(n9173), .ZN(n9176) );
  NOR2_X1 U8602 ( .A1(n7733), .A2(n10413), .ZN(n7732) );
  NAND2_X1 U8603 ( .A1(n6883), .A2(n6884), .ZN(n12671) );
  NAND2_X1 U8604 ( .A1(n12642), .A2(n10136), .ZN(n10191) );
  INV_X1 U8605 ( .A(n12761), .ZN(n7188) );
  AND4_X1 U8606 ( .A1(n9886), .A2(n9885), .A3(n9884), .A4(n9883), .ZN(n11785)
         );
  OAI21_X1 U8607 ( .B1(n10978), .B2(n11434), .A(n10897), .ZN(n10967) );
  AND2_X1 U8608 ( .A1(n6752), .A2(n6751), .ZN(n11426) );
  NAND2_X1 U8609 ( .A1(n13134), .A2(n11428), .ZN(n6752) );
  NAND2_X1 U8610 ( .A1(n13039), .A2(n10918), .ZN(n6751) );
  INV_X1 U8611 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n11022) );
  NAND2_X1 U8612 ( .A1(n10928), .A2(n11011), .ZN(n11013) );
  NAND2_X1 U8613 ( .A1(n11013), .A2(n10929), .ZN(n10993) );
  NAND2_X1 U8614 ( .A1(n11019), .A2(n10944), .ZN(n7514) );
  NAND2_X1 U8615 ( .A1(n10981), .A2(n10982), .ZN(n10980) );
  AND2_X1 U8616 ( .A1(n11125), .A2(n7515), .ZN(n11085) );
  NAND2_X1 U8617 ( .A1(n10993), .A2(n10992), .ZN(n10991) );
  NAND2_X1 U8618 ( .A1(n6570), .A2(n11125), .ZN(n11126) );
  NAND2_X1 U8619 ( .A1(n10949), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7101) );
  NAND2_X1 U8620 ( .A1(n7100), .A2(n11071), .ZN(n11073) );
  INV_X1 U8621 ( .A(n7101), .ZN(n7100) );
  AOI21_X1 U8622 ( .B1(n11216), .B2(n11215), .A(n11654), .ZN(n11667) );
  NAND2_X1 U8623 ( .A1(n11233), .A2(n11234), .ZN(n11665) );
  NAND2_X1 U8624 ( .A1(n6746), .A2(n11662), .ZN(n11813) );
  NAND2_X1 U8625 ( .A1(n11665), .A2(n11664), .ZN(n6746) );
  NAND2_X1 U8626 ( .A1(n11813), .A2(n11812), .ZN(n11815) );
  NOR2_X1 U8627 ( .A1(n9959), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U8628 ( .A1(n9683), .A2(n9682), .ZN(n9959) );
  NAND2_X1 U8629 ( .A1(n11874), .A2(n11875), .ZN(n6822) );
  NAND2_X1 U8630 ( .A1(n12993), .A2(n12990), .ZN(n13023) );
  NAND2_X1 U8631 ( .A1(n6817), .A2(n6821), .ZN(n13005) );
  NAND2_X1 U8632 ( .A1(n12988), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6821) );
  OAI21_X1 U8633 ( .B1(n6819), .B2(n11876), .A(n6818), .ZN(n6817) );
  INV_X1 U8634 ( .A(n6822), .ZN(n6819) );
  NAND2_X1 U8635 ( .A1(n7522), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7521) );
  NAND2_X1 U8636 ( .A1(n6652), .A2(n13058), .ZN(n7520) );
  NAND2_X1 U8637 ( .A1(n6651), .A2(n13075), .ZN(n13086) );
  NAND2_X1 U8638 ( .A1(n7521), .A2(n7520), .ZN(n6651) );
  INV_X1 U8639 ( .A(n7520), .ZN(n13077) );
  AOI21_X1 U8640 ( .B1(n13067), .B2(n13066), .A(n13065), .ZN(n13096) );
  NAND2_X1 U8641 ( .A1(n13092), .A2(n13093), .ZN(n6827) );
  NOR2_X1 U8642 ( .A1(n13103), .A2(n6621), .ZN(n13132) );
  NAND2_X1 U8643 ( .A1(n7497), .A2(n13135), .ZN(n7496) );
  INV_X1 U8644 ( .A(n7503), .ZN(n7497) );
  INV_X1 U8645 ( .A(n13110), .ZN(n7502) );
  INV_X1 U8646 ( .A(n12784), .ZN(n12548) );
  AOI21_X1 U8647 ( .B1(n13427), .B2(n12960), .A(n15601), .ZN(n6991) );
  NAND2_X1 U8648 ( .A1(n12542), .A2(n12541), .ZN(n12556) );
  NAND2_X1 U8649 ( .A1(n10298), .A2(n10297), .ZN(n10351) );
  OR2_X1 U8650 ( .A1(n10351), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12092) );
  NOR2_X1 U8651 ( .A1(n12551), .A2(n15580), .ZN(n10358) );
  OR2_X1 U8652 ( .A1(n12782), .A2(n10272), .ZN(n13194) );
  NAND2_X1 U8653 ( .A1(n13376), .A2(n13228), .ZN(n13196) );
  NAND2_X1 U8654 ( .A1(n13438), .A2(n13238), .ZN(n7804) );
  OR2_X1 U8655 ( .A1(n10163), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n10182) );
  NAND2_X1 U8656 ( .A1(n10097), .A2(n7160), .ZN(n10129) );
  INV_X1 U8657 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7159) );
  OR2_X1 U8658 ( .A1(n13304), .A2(n13278), .ZN(n13291) );
  NAND2_X1 U8659 ( .A1(n10027), .A2(n6468), .ZN(n10077) );
  INV_X1 U8660 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7156) );
  NAND2_X1 U8661 ( .A1(n10027), .A2(n7157), .ZN(n10062) );
  NAND2_X1 U8662 ( .A1(n10027), .A2(n10026), .ZN(n10044) );
  NAND2_X1 U8663 ( .A1(n9988), .A2(n9987), .ZN(n10005) );
  INV_X1 U8664 ( .A(n9989), .ZN(n9988) );
  INV_X1 U8665 ( .A(n7155), .ZN(n9966) );
  AND2_X1 U8666 ( .A1(n6493), .A2(n9911), .ZN(n7162) );
  OR2_X1 U8667 ( .A1(n9928), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U8668 ( .A1(n9848), .A2(n6493), .ZN(n9912) );
  NAND4_X1 U8669 ( .A1(n9802), .A2(n11499), .A3(n7164), .A4(n9823), .ZN(n9882)
         );
  INV_X1 U8670 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7164) );
  NAND2_X1 U8671 ( .A1(n9848), .A2(n9847), .ZN(n9856) );
  NAND2_X1 U8672 ( .A1(n7191), .A2(n6612), .ZN(n11508) );
  INV_X1 U8673 ( .A(n7193), .ZN(n7191) );
  NAND2_X1 U8674 ( .A1(n11508), .A2(n11507), .ZN(n11506) );
  AOI21_X1 U8675 ( .B1(n7696), .B2(n7698), .A(n7694), .ZN(n7693) );
  INV_X1 U8676 ( .A(n12827), .ZN(n7694) );
  INV_X1 U8677 ( .A(n12819), .ZN(n11733) );
  NAND2_X1 U8678 ( .A1(n11499), .A2(n9802), .ZN(n9824) );
  NAND2_X1 U8679 ( .A1(n7218), .A2(n10315), .ZN(n11495) );
  NAND2_X1 U8680 ( .A1(n15578), .A2(n15579), .ZN(n7218) );
  INV_X1 U8681 ( .A(n10259), .ZN(n11494) );
  INV_X1 U8682 ( .A(n12809), .ZN(n15578) );
  INV_X1 U8683 ( .A(n10998), .ZN(n15598) );
  INV_X1 U8684 ( .A(n11047), .ZN(n15593) );
  NAND2_X1 U8685 ( .A1(n7581), .A2(n12543), .ZN(n6867) );
  NOR2_X1 U8686 ( .A1(n7705), .A2(n12910), .ZN(n7701) );
  OAI21_X1 U8687 ( .B1(n7703), .B2(n12910), .A(n7700), .ZN(n7699) );
  NOR2_X1 U8688 ( .A1(n13277), .A2(n13305), .ZN(n13304) );
  AND2_X1 U8689 ( .A1(n13287), .A2(n12894), .ZN(n13305) );
  INV_X1 U8690 ( .A(n12885), .ZN(n13314) );
  NAND2_X1 U8691 ( .A1(n10043), .A2(n10042), .ZN(n13406) );
  NAND2_X1 U8692 ( .A1(n7724), .A2(n12881), .ZN(n7719) );
  NOR2_X1 U8693 ( .A1(n7722), .A2(n10264), .ZN(n7721) );
  NAND2_X1 U8694 ( .A1(n13349), .A2(n10329), .ZN(n13353) );
  AND4_X1 U8695 ( .A1(n9971), .A2(n9970), .A3(n9969), .A4(n9968), .ZN(n12383)
         );
  INV_X1 U8696 ( .A(n7797), .ZN(n7796) );
  OAI21_X1 U8697 ( .B1(n10325), .B2(n7830), .A(n10326), .ZN(n7797) );
  AND2_X1 U8698 ( .A1(n12860), .A2(n12863), .ZN(n12858) );
  INV_X1 U8699 ( .A(n7716), .ZN(n7710) );
  INV_X1 U8700 ( .A(n7712), .ZN(n7711) );
  NAND2_X1 U8701 ( .A1(n12540), .A2(n12539), .ZN(n12581) );
  NAND2_X1 U8702 ( .A1(n7592), .A2(n12209), .ZN(n6877) );
  OAI21_X1 U8703 ( .B1(n10156), .B2(n10157), .A(n10159), .ZN(n10174) );
  INV_X1 U8704 ( .A(n9713), .ZN(n9687) );
  INV_X1 U8705 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n6893) );
  INV_X1 U8706 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n10798) );
  INV_X1 U8707 ( .A(n10037), .ZN(n7565) );
  OR2_X1 U8708 ( .A1(n9923), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9944) );
  INV_X1 U8709 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9907) );
  XNOR2_X1 U8710 ( .A(n9844), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11225) );
  AOI21_X1 U8711 ( .B1(n7589), .B2(n7591), .A(n6558), .ZN(n7588) );
  OR2_X1 U8712 ( .A1(n9796), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U8713 ( .A1(n9763), .A2(n9775), .ZN(n9796) );
  NOR2_X1 U8714 ( .A1(n9763), .A2(n13502), .ZN(n6830) );
  AND2_X1 U8715 ( .A1(n8467), .A2(n8466), .ZN(n8535) );
  AOI21_X1 U8716 ( .B1(n6441), .B2(n12193), .A(n6458), .ZN(n7561) );
  NAND2_X1 U8717 ( .A1(n12192), .A2(n6441), .ZN(n6654) );
  OR2_X1 U8718 ( .A1(n8375), .A2(n13615), .ZN(n8377) );
  NAND2_X1 U8719 ( .A1(n11695), .A2(n8068), .ZN(n7530) );
  INV_X1 U8720 ( .A(n11342), .ZN(n7537) );
  INV_X1 U8721 ( .A(n13673), .ZN(n10642) );
  INV_X1 U8722 ( .A(n6694), .ZN(n8128) );
  NAND2_X1 U8723 ( .A1(n8420), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8436) );
  AOI21_X1 U8724 ( .B1(n13556), .B2(n8370), .A(n8365), .ZN(n13535) );
  OR2_X1 U8725 ( .A1(n13536), .A2(n13539), .ZN(n8357) );
  NOR2_X1 U8726 ( .A1(n7551), .A2(n6606), .ZN(n7545) );
  OAI21_X1 U8727 ( .B1(n7547), .B2(n6606), .A(n7544), .ZN(n7543) );
  OR2_X1 U8728 ( .A1(n8153), .A2(n11849), .ZN(n8171) );
  OR2_X1 U8729 ( .A1(n12120), .A2(n10632), .ZN(n7897) );
  NAND2_X1 U8730 ( .A1(n13583), .A2(n6993), .ZN(n13582) );
  NOR2_X1 U8731 ( .A1(n13629), .A2(n8432), .ZN(n7559) );
  NAND2_X1 U8732 ( .A1(n8169), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8205) );
  INV_X1 U8733 ( .A(n8171), .ZN(n8169) );
  INV_X1 U8734 ( .A(n6996), .ZN(n8207) );
  AND4_X1 U8735 ( .A1(n8025), .A2(n8024), .A3(n8023), .A4(n8022), .ZN(n11475)
         );
  INV_X1 U8736 ( .A(n15483), .ZN(n6664) );
  NAND2_X1 U8737 ( .A1(n10666), .A2(n10667), .ZN(n11164) );
  OR2_X1 U8738 ( .A1(n10661), .A2(n10662), .ZN(n11170) );
  OR2_X1 U8739 ( .A1(n11172), .A2(n11173), .ZN(n11460) );
  AND2_X1 U8740 ( .A1(n7383), .A2(n7382), .ZN(n11574) );
  NAND2_X1 U8741 ( .A1(n11573), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7382) );
  NAND2_X1 U8742 ( .A1(n11574), .A2(n11575), .ZN(n11839) );
  NAND2_X1 U8743 ( .A1(n13684), .A2(n13685), .ZN(n7391) );
  OR2_X1 U8744 ( .A1(n15519), .A2(n11614), .ZN(n7028) );
  AND2_X1 U8745 ( .A1(n8480), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13729) );
  NAND2_X1 U8746 ( .A1(n8457), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8482) );
  INV_X1 U8747 ( .A(n8459), .ZN(n8457) );
  NAND2_X1 U8748 ( .A1(n13761), .A2(n14121), .ZN(n13747) );
  NAND2_X1 U8749 ( .A1(n7263), .A2(n7268), .ZN(n13771) );
  OR2_X1 U8750 ( .A1(n13841), .A2(n7271), .ZN(n7263) );
  NAND2_X1 U8751 ( .A1(n9079), .A2(n8787), .ZN(n13802) );
  NAND2_X1 U8752 ( .A1(n7267), .A2(n9078), .ZN(n13792) );
  NAND2_X1 U8753 ( .A1(n13841), .A2(n9075), .ZN(n7267) );
  NAND2_X1 U8754 ( .A1(n13795), .A2(n13968), .ZN(n7776) );
  NAND2_X1 U8755 ( .A1(n6447), .A2(n13865), .ZN(n13814) );
  NAND2_X1 U8756 ( .A1(n6523), .A2(n13826), .ZN(n13825) );
  AND2_X1 U8757 ( .A1(n13865), .A2(n14137), .ZN(n13849) );
  AND2_X1 U8758 ( .A1(n13865), .A2(n7409), .ZN(n13829) );
  NAND2_X1 U8759 ( .A1(n6995), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U8760 ( .A1(n7788), .A2(n7787), .ZN(n13858) );
  NAND2_X1 U8761 ( .A1(n6693), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8308) );
  INV_X1 U8762 ( .A(n6995), .ZN(n8319) );
  NAND2_X1 U8763 ( .A1(n9068), .A2(n6631), .ZN(n6630) );
  NOR2_X1 U8764 ( .A1(n9070), .A2(n6632), .ZN(n6631) );
  NAND2_X1 U8765 ( .A1(n7678), .A2(n6478), .ZN(n13889) );
  INV_X1 U8766 ( .A(n13892), .ZN(n9029) );
  INV_X1 U8767 ( .A(n7013), .ZN(n13899) );
  AND2_X1 U8768 ( .A1(n7399), .A2(n7172), .ZN(n13939) );
  NOR2_X1 U8769 ( .A1(n7398), .A2(n14074), .ZN(n7399) );
  AND2_X1 U8770 ( .A1(n13945), .A2(n13910), .ZN(n13927) );
  NAND2_X1 U8771 ( .A1(n7401), .A2(n7172), .ZN(n13953) );
  NAND2_X1 U8772 ( .A1(n7757), .A2(n6516), .ZN(n6643) );
  INV_X1 U8773 ( .A(n9061), .ZN(n7763) );
  AND2_X1 U8774 ( .A1(n7760), .A2(n7764), .ZN(n7759) );
  OR2_X1 U8775 ( .A1(n14089), .A2(n13530), .ZN(n7764) );
  OR2_X1 U8776 ( .A1(n9062), .A2(n7761), .ZN(n7760) );
  NAND2_X1 U8777 ( .A1(n7762), .A2(n9061), .ZN(n7761) );
  NOR2_X2 U8778 ( .A1(n12281), .A2(n14154), .ZN(n12298) );
  AOI21_X1 U8779 ( .B1(n7675), .B2(n9022), .A(n6541), .ZN(n7674) );
  AND4_X1 U8780 ( .A1(n8133), .A2(n8132), .A3(n8131), .A4(n8130), .ZN(n12295)
         );
  NAND2_X1 U8781 ( .A1(n9055), .A2(n7781), .ZN(n7780) );
  CLKBUF_X1 U8782 ( .A(n11962), .Z(n12170) );
  AND2_X1 U8783 ( .A1(n12012), .A2(n11984), .ZN(n11981) );
  NOR2_X1 U8784 ( .A1(n8020), .A2(n6690), .ZN(n6688) );
  CLKBUF_X1 U8785 ( .A(n11980), .Z(n12012) );
  NOR2_X2 U8786 ( .A1(n12041), .A2(n15552), .ZN(n12011) );
  OR2_X1 U8787 ( .A1(n13974), .A2(n11614), .ZN(n9091) );
  AND2_X1 U8788 ( .A1(n15533), .A2(n9090), .ZN(n9192) );
  INV_X1 U8789 ( .A(n11356), .ZN(n11350) );
  AND2_X2 U8790 ( .A1(n8567), .A2(n11353), .ZN(n12123) );
  NAND2_X1 U8791 ( .A1(n13824), .A2(n9035), .ZN(n13817) );
  NAND2_X1 U8792 ( .A1(n8419), .A2(n8418), .ZN(n13784) );
  NAND2_X1 U8793 ( .A1(n7767), .A2(n7765), .ZN(n13935) );
  INV_X2 U8794 ( .A(n12126), .ZN(n15537) );
  OR2_X1 U8795 ( .A1(n8503), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n8506) );
  OR2_X1 U8796 ( .A1(n8095), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8097) );
  OR2_X1 U8797 ( .A1(n8097), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n8147) );
  OR2_X1 U8798 ( .A1(n8196), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U8799 ( .A1(n9385), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9400) );
  INV_X1 U8800 ( .A(n9415), .ZN(n9428) );
  NAND2_X1 U8801 ( .A1(n14320), .A2(n6446), .ZN(n14189) );
  AND2_X1 U8802 ( .A1(n14297), .A2(n9555), .ZN(n14203) );
  AND2_X1 U8803 ( .A1(n9624), .A2(n9623), .ZN(n9655) );
  OR2_X1 U8804 ( .A1(n9329), .A2(n11952), .ZN(n9331) );
  NAND2_X1 U8805 ( .A1(n9326), .A2(n9327), .ZN(n7376) );
  AOI21_X1 U8806 ( .B1(n7372), .B2(n9500), .A(n6557), .ZN(n7371) );
  NAND2_X1 U8807 ( .A1(n9415), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9430) );
  INV_X1 U8808 ( .A(n6703), .ZN(n6702) );
  OAI21_X1 U8809 ( .B1(n6446), .B2(n6704), .A(n6484), .ZN(n6703) );
  OR2_X1 U8810 ( .A1(n14276), .A2(n14274), .ZN(n9439) );
  INV_X1 U8811 ( .A(n9412), .ZN(n6704) );
  NAND2_X1 U8812 ( .A1(n6712), .A2(n14298), .ZN(n14259) );
  NAND2_X1 U8813 ( .A1(n9256), .A2(n9255), .ZN(n10653) );
  NAND2_X1 U8814 ( .A1(n7046), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9507) );
  INV_X1 U8815 ( .A(n7046), .ZN(n9484) );
  NAND2_X1 U8816 ( .A1(n9505), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9523) );
  INV_X1 U8817 ( .A(n9507), .ZN(n9505) );
  OR2_X1 U8818 ( .A1(n9557), .A2(n14329), .ZN(n14200) );
  AND2_X1 U8819 ( .A1(n14202), .A2(n9538), .ZN(n14330) );
  NAND2_X1 U8820 ( .A1(n14231), .A2(n14232), .ZN(n14230) );
  NAND2_X1 U8821 ( .A1(n9459), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9471) );
  INV_X1 U8822 ( .A(n9461), .ZN(n9459) );
  NAND2_X1 U8823 ( .A1(n14189), .A2(n9412), .ZN(n14275) );
  AND2_X1 U8824 ( .A1(n9596), .A2(n9579), .ZN(n14268) );
  OAI22_X1 U8825 ( .A1(n10615), .A2(n12508), .B1(n6434), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n6781) );
  INV_X1 U8826 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U8827 ( .A1(n14663), .A2(n14662), .ZN(n14661) );
  INV_X1 U8828 ( .A(n14716), .ZN(n7310) );
  AOI21_X1 U8829 ( .B1(n7308), .B2(n7307), .A(n7306), .ZN(n7305) );
  INV_X1 U8830 ( .A(n14715), .ZN(n7306) );
  INV_X1 U8831 ( .A(n7312), .ZN(n7307) );
  NAND2_X1 U8832 ( .A1(n7311), .A2(n7313), .ZN(n14717) );
  NAND2_X1 U8833 ( .A1(n14708), .A2(n7312), .ZN(n7311) );
  AND2_X1 U8834 ( .A1(n10686), .A2(n10685), .ZN(n14722) );
  OAI21_X1 U8835 ( .B1(n7305), .B2(n7302), .A(n7301), .ZN(n7300) );
  INV_X1 U8836 ( .A(n10706), .ZN(n7302) );
  INV_X1 U8837 ( .A(n10705), .ZN(n7301) );
  NAND2_X1 U8838 ( .A1(n6635), .A2(n6634), .ZN(n10876) );
  INV_X1 U8839 ( .A(n10692), .ZN(n6634) );
  INV_X1 U8840 ( .A(n10691), .ZN(n6635) );
  INV_X1 U8841 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10871) );
  NAND2_X1 U8842 ( .A1(n6637), .A2(n6636), .ZN(n11291) );
  INV_X1 U8843 ( .A(n11108), .ZN(n6636) );
  INV_X1 U8844 ( .A(n11107), .ZN(n6637) );
  NAND2_X1 U8845 ( .A1(n7289), .A2(n14729), .ZN(n14733) );
  OR2_X1 U8846 ( .A1(n14731), .A2(n14730), .ZN(n7289) );
  NAND2_X1 U8847 ( .A1(n7288), .A2(n7292), .ZN(n7287) );
  INV_X1 U8848 ( .A(n7290), .ZN(n7288) );
  AOI21_X1 U8849 ( .B1(n14729), .B2(n14730), .A(n7291), .ZN(n7290) );
  INV_X1 U8850 ( .A(n11111), .ZN(n7291) );
  AND2_X1 U8851 ( .A1(n7292), .A2(n14729), .ZN(n7286) );
  NAND2_X1 U8852 ( .A1(n12349), .A2(n12348), .ZN(n12351) );
  XNOR2_X1 U8853 ( .A(n14782), .B(n9475), .ZN(n14784) );
  NOR2_X1 U8854 ( .A1(n7489), .A2(n14800), .ZN(n7488) );
  NAND2_X1 U8855 ( .A1(n12523), .A2(n12526), .ZN(n14605) );
  INV_X1 U8856 ( .A(n14864), .ZN(n7068) );
  XNOR2_X1 U8857 ( .A(n9636), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n12437) );
  OAI21_X1 U8858 ( .B1(n14847), .B2(n12430), .A(n12429), .ZN(n7256) );
  NAND2_X1 U8859 ( .A1(n14864), .A2(n7753), .ZN(n7074) );
  OR2_X1 U8860 ( .A1(n6788), .A2(n7629), .ZN(n6787) );
  INV_X1 U8861 ( .A(n7631), .ZN(n6788) );
  XNOR2_X1 U8862 ( .A(n14603), .B(n14640), .ZN(n14830) );
  INV_X1 U8863 ( .A(n7485), .ZN(n7814) );
  AND2_X1 U8864 ( .A1(n9561), .A2(n9540), .ZN(n14857) );
  AND2_X1 U8865 ( .A1(n7063), .A2(n7746), .ZN(n7062) );
  AOI21_X1 U8866 ( .B1(n14909), .B2(n7747), .A(n6459), .ZN(n7746) );
  INV_X1 U8867 ( .A(n7653), .ZN(n6785) );
  NAND2_X1 U8868 ( .A1(n6784), .A2(n7653), .ZN(n6783) );
  CLKBUF_X1 U8869 ( .A(n14905), .Z(n14926) );
  NOR2_X1 U8870 ( .A1(n7483), .A2(n15137), .ZN(n6800) );
  NAND2_X1 U8871 ( .A1(n9444), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9461) );
  INV_X1 U8872 ( .A(n7483), .ZN(n7482) );
  NAND2_X1 U8873 ( .A1(n15006), .A2(n14995), .ZN(n14989) );
  NOR2_X1 U8874 ( .A1(n12411), .A2(n15019), .ZN(n12412) );
  NAND2_X1 U8875 ( .A1(n7223), .A2(n12408), .ZN(n15220) );
  OR2_X1 U8876 ( .A1(n12409), .A2(n14593), .ZN(n7223) );
  NOR2_X1 U8877 ( .A1(n7492), .A2(n15230), .ZN(n7490) );
  OAI21_X1 U8878 ( .B1(n7735), .B2(n7078), .A(n11923), .ZN(n7076) );
  NAND2_X1 U8879 ( .A1(n7620), .A2(n7618), .ZN(n12215) );
  NAND2_X1 U8880 ( .A1(n11926), .A2(n11924), .ZN(n7620) );
  NOR2_X1 U8881 ( .A1(n12222), .A2(n14428), .ZN(n15051) );
  NAND2_X1 U8882 ( .A1(n9222), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9314) );
  INV_X1 U8883 ( .A(n9312), .ZN(n9222) );
  NAND2_X1 U8884 ( .A1(n7044), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9329) );
  INV_X1 U8885 ( .A(n9314), .ZN(n7044) );
  NAND2_X1 U8886 ( .A1(n11628), .A2(n11679), .ZN(n7057) );
  NAND2_X1 U8887 ( .A1(n11632), .A2(n11679), .ZN(n7058) );
  OR2_X1 U8888 ( .A1(n14650), .A2(n11635), .ZN(n7242) );
  NOR2_X1 U8889 ( .A1(n11636), .A2(n7241), .ZN(n7240) );
  AND2_X1 U8890 ( .A1(n8851), .A2(n6795), .ZN(n11645) );
  INV_X2 U8891 ( .A(n8949), .ZN(n8925) );
  NAND2_X1 U8892 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9289) );
  NAND2_X1 U8893 ( .A1(n9221), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9312) );
  INV_X1 U8894 ( .A(n9289), .ZN(n9221) );
  NAND2_X1 U8895 ( .A1(n8851), .A2(n11622), .ZN(n11587) );
  INV_X1 U8896 ( .A(n14550), .ZN(n15070) );
  NAND2_X1 U8897 ( .A1(n14180), .A2(n8948), .ZN(n8942) );
  OR2_X1 U8898 ( .A1(n14826), .A2(n14825), .ZN(n15094) );
  CLKBUF_X1 U8899 ( .A(n14961), .Z(n14963) );
  INV_X1 U8900 ( .A(n14438), .ZN(n15259) );
  OR2_X1 U8901 ( .A1(n11926), .A2(n11925), .ZN(n7617) );
  INV_X1 U8902 ( .A(n15363), .ZN(n15400) );
  AND2_X1 U8903 ( .A1(n6948), .A2(n8702), .ZN(n12403) );
  NAND2_X1 U8904 ( .A1(n7347), .A2(n7345), .ZN(n8702) );
  NAND2_X1 U8905 ( .A1(n7347), .A2(n8685), .ZN(n8701) );
  XNOR2_X1 U8906 ( .A(n8717), .B(n8716), .ZN(n14172) );
  AND2_X1 U8907 ( .A1(n7660), .A2(n8824), .ZN(n7659) );
  XNOR2_X1 U8908 ( .A(n8975), .B(P1_IR_REG_25__SCAN_IN), .ZN(n8984) );
  XNOR2_X1 U8909 ( .A(n8977), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8983) );
  XNOR2_X1 U8910 ( .A(n8396), .B(n8410), .ZN(n12207) );
  NAND2_X1 U8911 ( .A1(n7351), .A2(n8338), .ZN(n8389) );
  NAND2_X1 U8912 ( .A1(n8303), .A2(n7355), .ZN(n7351) );
  XNOR2_X1 U8913 ( .A(n8330), .B(n8329), .ZN(n11769) );
  NAND2_X1 U8914 ( .A1(n8328), .A2(n8327), .ZN(n8330) );
  XNOR2_X1 U8915 ( .A(n8278), .B(n8277), .ZN(n11613) );
  NAND2_X1 U8916 ( .A1(n6736), .A2(n8274), .ZN(n8278) );
  OAI211_X1 U8917 ( .C1(n6777), .C2(n8254), .A(n6775), .B(n6770), .ZN(n11365)
         );
  NAND2_X1 U8918 ( .A1(n6777), .A2(n6475), .ZN(n6770) );
  XNOR2_X1 U8919 ( .A(n6918), .B(n8069), .ZN(n10469) );
  XNOR2_X1 U8920 ( .A(n8047), .B(n8046), .ZN(n10448) );
  NAND2_X1 U8921 ( .A1(n6913), .A2(n8854), .ZN(n8863) );
  NAND2_X1 U8922 ( .A1(n7165), .A2(n7975), .ZN(n7995) );
  NAND2_X1 U8923 ( .A1(n7973), .A2(n7972), .ZN(n7165) );
  INV_X1 U8924 ( .A(n6913), .ZN(n8853) );
  AOI21_X1 U8925 ( .B1(n7931), .B2(n7932), .A(n7930), .ZN(n7936) );
  INV_X1 U8926 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9141) );
  XNOR2_X1 U8927 ( .A(n9102), .B(n9101), .ZN(n9140) );
  INV_X1 U8928 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9101) );
  NOR2_X1 U8929 ( .A1(n9144), .A2(n9145), .ZN(n9148) );
  NAND2_X1 U8930 ( .A1(n9154), .A2(n9153), .ZN(n9155) );
  OAI21_X1 U8931 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n9113), .A(n9112), .ZN(
        n9126) );
  NAND2_X1 U8932 ( .A1(n6808), .A2(n7607), .ZN(n9162) );
  NAND2_X1 U8933 ( .A1(n15267), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7607) );
  OAI21_X1 U8934 ( .B1(n15213), .B2(n6807), .A(n6804), .ZN(n6808) );
  NOR2_X1 U8935 ( .A1(n6806), .A2(n15215), .ZN(n6807) );
  INV_X1 U8936 ( .A(n15247), .ZN(n7604) );
  NAND2_X1 U8937 ( .A1(n12610), .A2(n12612), .ZN(n12611) );
  NAND2_X1 U8938 ( .A1(n12727), .A2(n12486), .ZN(n12610) );
  NOR2_X1 U8939 ( .A1(n7425), .A2(n7424), .ZN(n12619) );
  NAND2_X1 U8940 ( .A1(n7431), .A2(n6449), .ZN(n7424) );
  INV_X1 U8941 ( .A(n7428), .ZN(n7425) );
  OAI211_X1 U8942 ( .C1(n11559), .C2(n7460), .A(n9936), .B(n7459), .ZN(n11906)
         );
  INV_X1 U8943 ( .A(n9889), .ZN(n7461) );
  NAND3_X1 U8944 ( .A1(n7455), .A2(n9746), .A3(n6477), .ZN(n11043) );
  NAND2_X1 U8945 ( .A1(n11404), .A2(n9813), .ZN(n11560) );
  AND2_X1 U8946 ( .A1(n10083), .A2(n10082), .ZN(n13316) );
  INV_X1 U8947 ( .A(n7451), .ZN(n6896) );
  AOI21_X1 U8948 ( .B1(n10012), .B2(n7451), .A(n6566), .ZN(n6895) );
  AND2_X1 U8949 ( .A1(n10033), .A2(n10051), .ZN(n7451) );
  NAND2_X1 U8950 ( .A1(n9897), .A2(n7464), .ZN(n11864) );
  AND3_X2 U8951 ( .A1(n9731), .A2(n9730), .A3(n9729), .ZN(n15583) );
  INV_X1 U8952 ( .A(n7429), .ZN(n12326) );
  AOI21_X1 U8953 ( .B1(n12364), .B2(n9973), .A(n7432), .ZN(n7429) );
  INV_X1 U8954 ( .A(n12733), .ZN(n12741) );
  INV_X1 U8955 ( .A(n12749), .ZN(n12730) );
  NAND2_X1 U8956 ( .A1(n12618), .A2(n10013), .ZN(n12740) );
  AND2_X1 U8957 ( .A1(n12272), .A2(n12103), .ZN(n13153) );
  INV_X1 U8958 ( .A(n13193), .ZN(n12961) );
  INV_X1 U8959 ( .A(n13228), .ZN(n12963) );
  NAND2_X1 U8960 ( .A1(n10104), .A2(n10103), .ZN(n12710) );
  INV_X1 U8961 ( .A(n13316), .ZN(n12967) );
  INV_X1 U8962 ( .A(n12369), .ZN(n12974) );
  INV_X1 U8963 ( .A(n11785), .ZN(n12976) );
  INV_X1 U8964 ( .A(n11784), .ZN(n12978) );
  OAI22_X1 U8965 ( .A1(n13125), .A2(n6750), .B1(n11428), .B2(n13151), .ZN(
        n11430) );
  INV_X1 U8966 ( .A(n11426), .ZN(n6750) );
  AND2_X1 U8967 ( .A1(n11031), .A2(n10917), .ZN(n10964) );
  NOR2_X1 U8968 ( .A1(n11426), .A2(n11429), .ZN(n10963) );
  NAND2_X1 U8969 ( .A1(n7512), .A2(n7513), .ZN(n11001) );
  NAND2_X1 U8970 ( .A1(n10924), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7510) );
  AND2_X1 U8971 ( .A1(n7513), .A2(n10984), .ZN(n11002) );
  AOI21_X1 U8972 ( .B1(n11120), .B2(n6755), .A(n6555), .ZN(n6754) );
  INV_X1 U8973 ( .A(n11120), .ZN(n6756) );
  AND3_X1 U8974 ( .A1(n7093), .A2(n7095), .A3(n7091), .ZN(n11217) );
  XNOR2_X1 U8975 ( .A(n11653), .B(n11654), .ZN(n11655) );
  NAND2_X1 U8976 ( .A1(n11653), .A2(n7324), .ZN(n7323) );
  INV_X1 U8977 ( .A(n7506), .ZN(n7508) );
  AND2_X1 U8978 ( .A1(n6820), .A2(n6822), .ZN(n12982) );
  NAND2_X1 U8979 ( .A1(n11876), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n6820) );
  XNOR2_X1 U8980 ( .A(n13005), .B(n13018), .ZN(n12983) );
  AOI21_X1 U8981 ( .B1(n13013), .B2(n13012), .A(n13011), .ZN(n13033) );
  NOR2_X1 U8982 ( .A1(n7521), .A2(n13077), .ZN(n13076) );
  NAND2_X1 U8983 ( .A1(n13059), .A2(n13060), .ZN(n13062) );
  NAND2_X1 U8984 ( .A1(n7500), .A2(n7501), .ZN(n13128) );
  XNOR2_X1 U8985 ( .A(n13132), .B(n13131), .ZN(n13106) );
  NOR2_X1 U8986 ( .A1(n13106), .A2(n13107), .ZN(n13130) );
  NAND2_X1 U8987 ( .A1(n12763), .A2(n12762), .ZN(n13158) );
  NAND2_X1 U8988 ( .A1(n10095), .A2(n10094), .ZN(n13299) );
  NAND2_X1 U8989 ( .A1(n10061), .A2(n10060), .ZN(n13400) );
  NAND2_X1 U8990 ( .A1(n7799), .A2(n7798), .ZN(n13333) );
  NAND2_X1 U8991 ( .A1(n9927), .A2(n9926), .ZN(n12852) );
  NAND2_X1 U8992 ( .A1(n7714), .A2(n7715), .ZN(n11793) );
  NAND2_X1 U8993 ( .A1(n7014), .A2(n7716), .ZN(n7714) );
  AOI21_X1 U8994 ( .B1(n7014), .B2(n12835), .A(n7718), .ZN(n12070) );
  NAND2_X1 U8995 ( .A1(n7695), .A2(n12821), .ZN(n11772) );
  NAND2_X1 U8996 ( .A1(n11730), .A2(n12819), .ZN(n7695) );
  INV_X1 U8997 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11499) );
  OR2_X1 U8998 ( .A1(n11776), .A2(n15638), .ZN(n13340) );
  INV_X1 U8999 ( .A(n15577), .ZN(n15604) );
  NOR2_X1 U9000 ( .A1(n12544), .A2(n12543), .ZN(n13171) );
  AND2_X1 U9001 ( .A1(n13376), .A2(n15623), .ZN(n6937) );
  INV_X1 U9002 ( .A(n7805), .ZN(n13225) );
  AOI21_X1 U9003 ( .B1(n13224), .B2(n13221), .A(n13220), .ZN(n13439) );
  NAND2_X1 U9004 ( .A1(n13259), .A2(n10341), .ZN(n13250) );
  NAND2_X1 U9005 ( .A1(n10340), .A2(n10339), .ZN(n13261) );
  OAI21_X1 U9006 ( .B1(n6925), .B2(n7705), .A(n7703), .ZN(n13257) );
  NAND2_X1 U9007 ( .A1(n7708), .A2(n7707), .ZN(n13270) );
  NOR2_X1 U9008 ( .A1(n7706), .A2(n12888), .ZN(n13272) );
  INV_X1 U9009 ( .A(n7708), .ZN(n7706) );
  NAND2_X1 U9010 ( .A1(n10076), .A2(n10075), .ZN(n13470) );
  NAND2_X1 U9011 ( .A1(n7725), .A2(n7727), .ZN(n13332) );
  NAND2_X1 U9012 ( .A1(n12378), .A2(n7726), .ZN(n7725) );
  OAI21_X1 U9013 ( .B1(n12378), .B2(n12870), .A(n12377), .ZN(n13345) );
  NAND2_X1 U9014 ( .A1(n9986), .A2(n9985), .ZN(n13492) );
  INV_X1 U9015 ( .A(n13443), .ZN(n13493) );
  AND2_X1 U9016 ( .A1(n10207), .A2(n10206), .ZN(n13497) );
  AND2_X1 U9017 ( .A1(n10910), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13498) );
  AND2_X1 U9018 ( .A1(n7808), .A2(n7152), .ZN(n7807) );
  MUX2_X1 U9019 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9696), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9700) );
  NAND2_X1 U9020 ( .A1(n10267), .A2(n7592), .ZN(n10266) );
  XNOR2_X1 U9021 ( .A(n10126), .B(n10125), .ZN(n11650) );
  NAND2_X1 U9022 ( .A1(n7567), .A2(n7571), .ZN(n10036) );
  NAND2_X1 U9023 ( .A1(n10018), .A2(n10016), .ZN(n7567) );
  OAI21_X1 U9024 ( .B1(n9998), .B2(n10679), .A(n9997), .ZN(n10000) );
  NAND2_X1 U9025 ( .A1(n6872), .A2(n9957), .ZN(n9979) );
  NAND2_X1 U9026 ( .A1(n9956), .A2(n9955), .ZN(n6872) );
  OAI21_X1 U9027 ( .B1(n9865), .B2(n9898), .A(n7584), .ZN(n9920) );
  NAND2_X1 U9028 ( .A1(n9865), .A2(n9840), .ZN(n9900) );
  NAND2_X1 U9029 ( .A1(n9815), .A2(n9814), .ZN(n9836) );
  OAI21_X1 U9030 ( .B1(n9760), .B2(n7575), .A(n7574), .ZN(n9773) );
  AOI21_X1 U9031 ( .B1(n9761), .B2(n7580), .A(n7579), .ZN(n7574) );
  NAND2_X1 U9032 ( .A1(n9761), .A2(n9762), .ZN(n9771) );
  NAND2_X1 U9033 ( .A1(n9760), .A2(n9759), .ZN(n9762) );
  CLKBUF_X1 U9034 ( .A(n10943), .Z(n7009) );
  INV_X1 U9035 ( .A(n9740), .ZN(n9738) );
  NAND2_X1 U9036 ( .A1(n6654), .A2(n7561), .ZN(n13527) );
  NAND2_X1 U9037 ( .A1(n8167), .A2(n8166), .ZN(n14084) );
  NAND2_X1 U9038 ( .A1(n7530), .A2(n6608), .ZN(n11750) );
  OAI21_X1 U9039 ( .B1(n6993), .B2(n7551), .A(n7547), .ZN(n13548) );
  XNOR2_X1 U9040 ( .A(n12015), .B(n8490), .ZN(n11694) );
  INV_X1 U9041 ( .A(n12015), .ZN(n14111) );
  NOR2_X1 U9042 ( .A1(n8358), .A2(n8359), .ZN(n13558) );
  NAND2_X1 U9043 ( .A1(n13558), .A2(n13557), .ZN(n13556) );
  AND2_X1 U9044 ( .A1(n13643), .A2(n13968), .ZN(n13568) );
  INV_X1 U9045 ( .A(n11353), .ZN(n10637) );
  NAND2_X1 U9046 ( .A1(n12190), .A2(n8139), .ZN(n12310) );
  AND3_X1 U9047 ( .A1(n7533), .A2(n8374), .A3(n8373), .ZN(n13613) );
  NAND2_X1 U9048 ( .A1(n11472), .A2(n6608), .ZN(n6647) );
  OAI21_X1 U9049 ( .B1(n8067), .B2(n7528), .A(n8085), .ZN(n7527) );
  NAND2_X1 U9050 ( .A1(n13582), .A2(n8249), .ZN(n13622) );
  NAND2_X1 U9051 ( .A1(n13563), .A2(n8433), .ZN(n13628) );
  NAND2_X1 U9052 ( .A1(n14183), .A2(n8718), .ZN(n8448) );
  NAND2_X1 U9053 ( .A1(n11302), .A2(n8718), .ZN(n7173) );
  INV_X1 U9054 ( .A(n8772), .ZN(n7356) );
  OR2_X1 U9055 ( .A1(n8775), .A2(n8792), .ZN(n8813) );
  NOR2_X1 U9056 ( .A1(n8814), .A2(n8811), .ZN(n8812) );
  NAND2_X1 U9057 ( .A1(n8489), .A2(n8488), .ZN(n13742) );
  NAND2_X1 U9058 ( .A1(n6691), .A2(n8442), .ZN(n13773) );
  NAND2_X1 U9059 ( .A1(n13763), .A2(n8282), .ZN(n6691) );
  NAND2_X1 U9060 ( .A1(n8405), .A2(n8404), .ZN(n13810) );
  OR2_X1 U9061 ( .A1(n13798), .A2(n8424), .ZN(n8405) );
  NAND2_X1 U9062 ( .A1(n8356), .A2(n8355), .ZN(n13794) );
  INV_X1 U9063 ( .A(n11475), .ZN(n13666) );
  AND2_X1 U9064 ( .A1(n8006), .A2(n6965), .ZN(n6964) );
  AND3_X1 U9065 ( .A1(n7986), .A2(n7984), .A3(n7985), .ZN(n6979) );
  NAND2_X1 U9066 ( .A1(n7920), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7987) );
  OR2_X1 U9067 ( .A1(n7019), .A2(n7020), .ZN(n7947) );
  NAND2_X1 U9068 ( .A1(n8002), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7923) );
  INV_X1 U9069 ( .A(n12120), .ZN(n13672) );
  NAND2_X1 U9070 ( .A1(n11164), .A2(n6674), .ZN(n11165) );
  NAND2_X1 U9071 ( .A1(n6676), .A2(n6675), .ZN(n6674) );
  INV_X1 U9072 ( .A(n7385), .ZN(n11464) );
  OR2_X1 U9073 ( .A1(n11462), .A2(n11463), .ZN(n11570) );
  INV_X1 U9074 ( .A(n7383), .ZN(n11572) );
  NAND2_X1 U9075 ( .A1(n11839), .A2(n7042), .ZN(n11840) );
  OR2_X1 U9076 ( .A1(n11842), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7042) );
  INV_X1 U9077 ( .A(n7389), .ZN(n12388) );
  INV_X1 U9078 ( .A(n7387), .ZN(n12469) );
  XNOR2_X1 U9079 ( .A(n13682), .B(n13685), .ZN(n12389) );
  INV_X1 U9080 ( .A(n6673), .ZN(n13683) );
  NOR2_X1 U9081 ( .A1(n13683), .A2(n7392), .ZN(n15501) );
  INV_X1 U9082 ( .A(n7391), .ZN(n7392) );
  NOR2_X1 U9083 ( .A1(n15514), .A2(n6671), .ZN(n6670) );
  INV_X1 U9084 ( .A(n7390), .ZN(n6671) );
  NAND2_X1 U9085 ( .A1(n6672), .A2(n7390), .ZN(n15515) );
  OR2_X1 U9086 ( .A1(n10515), .A2(P2_U3088), .ZN(n15522) );
  NAND2_X1 U9087 ( .A1(n13693), .A2(n7380), .ZN(n13687) );
  NAND2_X1 U9088 ( .A1(n7023), .A2(n7022), .ZN(n7021) );
  OAI21_X1 U9089 ( .B1(n13759), .B2(n13758), .A(n13738), .ZN(n7024) );
  NAND2_X1 U9090 ( .A1(n13795), .A2(n13966), .ZN(n7022) );
  NAND2_X1 U9091 ( .A1(n7179), .A2(n7178), .ZN(n13822) );
  NAND2_X1 U9092 ( .A1(n7681), .A2(n9032), .ZN(n13872) );
  NAND2_X1 U9093 ( .A1(n9068), .A2(n9067), .ZN(n13888) );
  OAI21_X1 U9094 ( .B1(n13948), .B2(n7766), .A(n7277), .ZN(n13914) );
  INV_X1 U9095 ( .A(n14084), .ZN(n13980) );
  NAND2_X1 U9096 ( .A1(n7758), .A2(n9061), .ZN(n12294) );
  NAND2_X1 U9097 ( .A1(n12277), .A2(n9060), .ZN(n7758) );
  NAND2_X1 U9098 ( .A1(n7677), .A2(n9021), .ZN(n12160) );
  NAND2_X1 U9099 ( .A1(n7031), .A2(n9017), .ZN(n7677) );
  NAND2_X1 U9100 ( .A1(n13987), .A2(n9196), .ZN(n13979) );
  INV_X1 U9101 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6972) );
  AND2_X1 U9102 ( .A1(n14001), .A2(n14000), .ZN(n14117) );
  AND2_X1 U9103 ( .A1(n14018), .A2(n14017), .ZN(n14019) );
  OAI211_X1 U9104 ( .C1(n9201), .C2(n15557), .A(n6759), .B(n6757), .ZN(n9217)
         );
  NOR2_X1 U9105 ( .A1(n6533), .A2(n6758), .ZN(n6757) );
  INV_X1 U9106 ( .A(n9086), .ZN(n6758) );
  INV_X1 U9107 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6975) );
  INV_X1 U9108 ( .A(n12282), .ZN(n14154) );
  NAND2_X1 U9109 ( .A1(n6907), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7877) );
  NOR2_X1 U9110 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7847) );
  CLKBUF_X1 U9111 ( .A(n7886), .Z(n12562) );
  INV_X1 U9112 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10579) );
  OR2_X1 U9113 ( .A1(n8048), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8049) );
  INV_X1 U9114 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10412) );
  AND2_X1 U9115 ( .A1(n7970), .A2(n7998), .ZN(n15466) );
  INV_X1 U9116 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10409) );
  AOI21_X1 U9117 ( .B1(n7937), .B2(n6506), .A(n6669), .ZN(n6668) );
  NOR2_X1 U9118 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n6669) );
  NAND2_X1 U9119 ( .A1(n14166), .A2(n7396), .ZN(n7395) );
  NAND2_X1 U9120 ( .A1(n6470), .A2(n7394), .ZN(n7393) );
  NOR2_X1 U9121 ( .A1(n14166), .A2(n7396), .ZN(n7394) );
  INV_X1 U9122 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10416) );
  INV_X1 U9123 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10415) );
  NAND2_X1 U9124 ( .A1(n7862), .A2(n6470), .ZN(n15427) );
  NAND2_X1 U9126 ( .A1(n11541), .A2(n9325), .ZN(n11742) );
  AOI22_X1 U9127 ( .A1(n7361), .A2(n7364), .B1(n7363), .B2(n7367), .ZN(n7359)
         );
  NAND2_X1 U9128 ( .A1(n14320), .A2(n9398), .ZN(n14191) );
  NAND2_X1 U9129 ( .A1(n12257), .A2(n7003), .ZN(n14214) );
  NAND2_X1 U9130 ( .A1(n7005), .A2(n7004), .ZN(n7003) );
  INV_X1 U9131 ( .A(n9340), .ZN(n7004) );
  INV_X1 U9132 ( .A(n9339), .ZN(n7005) );
  INV_X1 U9133 ( .A(n11949), .ZN(n15048) );
  NAND2_X1 U9134 ( .A1(n7357), .A2(n7361), .ZN(n10380) );
  INV_X1 U9135 ( .A(n7373), .ZN(n11945) );
  NAND2_X1 U9136 ( .A1(n11740), .A2(n7376), .ZN(n11946) );
  NAND2_X1 U9137 ( .A1(n7370), .A2(n7371), .ZN(n14240) );
  NAND2_X1 U9138 ( .A1(n14339), .A2(n9366), .ZN(n14251) );
  AND2_X1 U9139 ( .A1(n7373), .A2(n6461), .ZN(n12259) );
  NAND2_X1 U9140 ( .A1(n14252), .A2(n9383), .ZN(n14322) );
  NAND2_X1 U9141 ( .A1(n14212), .A2(n7836), .ZN(n14341) );
  NAND2_X1 U9142 ( .A1(n9309), .A2(n9308), .ZN(n11543) );
  INV_X1 U9143 ( .A(n9307), .ZN(n9308) );
  OAI21_X1 U9144 ( .B1(n9306), .B2(n11603), .A(n9305), .ZN(n9307) );
  NAND2_X1 U9145 ( .A1(n11543), .A2(n11542), .ZN(n11541) );
  NAND2_X1 U9146 ( .A1(n9643), .A2(n9642), .ZN(n14637) );
  OR2_X1 U9147 ( .A1(n14808), .A2(n6433), .ZN(n9603) );
  INV_X1 U9148 ( .A(n14241), .ZN(n14642) );
  OR2_X1 U9149 ( .A1(n9420), .A2(n9419), .ZN(n14987) );
  INV_X1 U9150 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10487) );
  AND4_X1 U9151 ( .A1(n9361), .A2(n9360), .A3(n9359), .A4(n9358), .ZN(n15053)
         );
  AND4_X1 U9152 ( .A1(n9345), .A2(n9344), .A3(n9343), .A4(n9342), .ZN(n14439)
         );
  INV_X1 U9153 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10480) );
  OR2_X1 U9154 ( .A1(n12508), .A2(n14676), .ZN(n9260) );
  OR2_X1 U9155 ( .A1(n12508), .A2(n14655), .ZN(n9242) );
  OR2_X1 U9156 ( .A1(n12508), .A2(n11450), .ZN(n9251) );
  NAND2_X1 U9157 ( .A1(n7315), .A2(n14706), .ZN(n14710) );
  OR2_X1 U9158 ( .A1(n14708), .A2(n14707), .ZN(n7315) );
  NAND2_X1 U9159 ( .A1(n7298), .A2(n7305), .ZN(n14719) );
  OR2_X1 U9160 ( .A1(n14708), .A2(n7309), .ZN(n7298) );
  AND2_X1 U9161 ( .A1(n7303), .A2(n7299), .ZN(n10717) );
  OR2_X1 U9162 ( .A1(n14708), .A2(n7304), .ZN(n7303) );
  INV_X1 U9163 ( .A(n7300), .ZN(n7299) );
  NAND2_X1 U9164 ( .A1(n7308), .A2(n10706), .ZN(n7304) );
  AND2_X1 U9165 ( .A1(n11104), .A2(n11103), .ZN(n14738) );
  AND2_X1 U9166 ( .A1(n11443), .A2(n11442), .ZN(n11445) );
  NAND2_X1 U9167 ( .A1(n11445), .A2(n11444), .ZN(n11713) );
  NOR2_X1 U9168 ( .A1(n11438), .A2(n11437), .ZN(n11724) );
  NOR2_X1 U9169 ( .A1(n15303), .A2(n12344), .ZN(n14745) );
  NAND2_X1 U9170 ( .A1(n14751), .A2(n14750), .ZN(n14753) );
  XNOR2_X1 U9171 ( .A(n14778), .B(n14773), .ZN(n14763) );
  NAND2_X1 U9172 ( .A1(n14763), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14781) );
  INV_X1 U9173 ( .A(n15305), .ZN(n14785) );
  AOI21_X1 U9174 ( .B1(n12505), .B2(n14550), .A(n6797), .ZN(n15072) );
  OR2_X1 U9175 ( .A1(n14796), .A2(n15365), .ZN(n6797) );
  NAND2_X1 U9176 ( .A1(n12590), .A2(n15024), .ZN(n12592) );
  INV_X1 U9177 ( .A(n14603), .ZN(n14829) );
  NAND2_X1 U9178 ( .A1(n14868), .A2(n12422), .ZN(n14852) );
  NAND2_X1 U9179 ( .A1(n14911), .A2(n14476), .ZN(n14884) );
  NAND2_X1 U9180 ( .A1(n14918), .A2(n7653), .ZN(n14904) );
  NAND2_X1 U9181 ( .A1(n14946), .A2(n14492), .ZN(n14920) );
  NAND2_X1 U9182 ( .A1(n7623), .A2(n12416), .ZN(n14943) );
  NAND2_X1 U9183 ( .A1(n7624), .A2(n14471), .ZN(n14971) );
  NAND2_X1 U9184 ( .A1(n14997), .A2(n12449), .ZN(n14968) );
  NAND2_X1 U9185 ( .A1(n7740), .A2(n12445), .ZN(n15012) );
  INV_X1 U9186 ( .A(n15399), .ZN(n15058) );
  NAND2_X1 U9187 ( .A1(n7734), .A2(n12179), .ZN(n7079) );
  NAND2_X1 U9188 ( .A1(n12179), .A2(n12183), .ZN(n7738) );
  NAND2_X1 U9189 ( .A1(n7651), .A2(n11590), .ZN(n11637) );
  OAI21_X1 U9190 ( .B1(n14624), .B2(n15363), .A(n15064), .ZN(n8971) );
  AND4_X1 U9191 ( .A1(n15101), .A2(n15100), .A3(n15099), .A4(n15098), .ZN(
        n15102) );
  AND2_X1 U9192 ( .A1(n6452), .A2(n7745), .ZN(n7744) );
  INV_X1 U9193 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7745) );
  XNOR2_X1 U9194 ( .A(n8690), .B(n8689), .ZN(n14164) );
  OAI21_X1 U9195 ( .B1(n8717), .B2(n7344), .A(n7341), .ZN(n8690) );
  CLKBUF_X1 U9196 ( .A(n8969), .Z(n14671) );
  XNOR2_X1 U9197 ( .A(n8932), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15191) );
  OR2_X1 U9198 ( .A1(n8931), .A2(n9755), .ZN(n8932) );
  INV_X1 U9199 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11710) );
  NAND2_X1 U9200 ( .A1(n8958), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8957) );
  INV_X1 U9201 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11528) );
  INV_X1 U9202 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10681) );
  INV_X1 U9203 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10581) );
  INV_X1 U9204 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10451) );
  INV_X1 U9205 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10445) );
  INV_X1 U9206 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10439) );
  INV_X1 U9207 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10443) );
  OAI21_X1 U9208 ( .B1(n7955), .B2(n10467), .A(n7927), .ZN(n7904) );
  NAND2_X1 U9209 ( .A1(n6642), .A2(n6640), .ZN(n8839) );
  NAND2_X1 U9210 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6641), .ZN(n6640) );
  OAI21_X1 U9211 ( .B1(n7955), .B2(n10452), .A(n6793), .ZN(n6792) );
  INV_X1 U9212 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7297) );
  NOR2_X1 U9213 ( .A1(n8831), .A2(n7296), .ZN(n7295) );
  INV_X1 U9214 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9133) );
  AOI21_X1 U9215 ( .B1(n15201), .B2(n15198), .A(n15199), .ZN(n15661) );
  OAI21_X1 U9216 ( .B1(n6812), .B2(n6811), .A(n6810), .ZN(n15209) );
  NAND2_X1 U9217 ( .A1(n15206), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6810) );
  NOR2_X1 U9218 ( .A1(n15206), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6811) );
  XNOR2_X1 U9219 ( .A(n6891), .B(n12497), .ZN(n12502) );
  NAND2_X1 U9220 ( .A1(n11136), .A2(n9789), .ZN(n11407) );
  NAND2_X1 U9221 ( .A1(n6853), .A2(n10908), .ZN(n6852) );
  NAND2_X1 U9222 ( .A1(n10936), .A2(n11081), .ZN(n11119) );
  AND2_X1 U9223 ( .A1(n6828), .A2(n6824), .ZN(n13101) );
  AOI21_X1 U9224 ( .B1(n7494), .B2(n6656), .A(n13148), .ZN(n6655) );
  NAND2_X1 U9225 ( .A1(n7329), .A2(n13122), .ZN(n7328) );
  NAND2_X1 U9226 ( .A1(n7202), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7201) );
  NOR2_X1 U9227 ( .A1(n6609), .A2(n6988), .ZN(n6987) );
  NOR2_X1 U9228 ( .A1(n15652), .A2(n10379), .ZN(n6988) );
  INV_X1 U9229 ( .A(n7040), .ZN(n7039) );
  OAI22_X1 U9230 ( .A1(n13433), .A2(n13382), .B1(n15652), .B2(n13374), .ZN(
        n7040) );
  NOR2_X1 U9231 ( .A1(n6610), .A2(n6990), .ZN(n6989) );
  NOR2_X1 U9232 ( .A1(n15645), .A2(n10830), .ZN(n6990) );
  INV_X1 U9233 ( .A(n7038), .ZN(n7037) );
  OAI22_X1 U9234 ( .A1(n13433), .A2(n13443), .B1(n15645), .B2(n13432), .ZN(
        n7038) );
  OAI21_X1 U9235 ( .B1(n11203), .B2(n7541), .A(n7538), .ZN(n11343) );
  NAND2_X1 U9236 ( .A1(n11187), .A2(n7919), .ZN(n11180) );
  NAND2_X1 U9237 ( .A1(n9203), .A2(n6649), .ZN(n8558) );
  NAND2_X1 U9238 ( .A1(n7553), .A2(n7558), .ZN(n10888) );
  NAND2_X1 U9239 ( .A1(n11202), .A2(n7993), .ZN(n11145) );
  AND2_X1 U9240 ( .A1(n10527), .A2(n10528), .ZN(n10663) );
  NAND2_X1 U9241 ( .A1(n6681), .A2(n6678), .ZN(n6677) );
  NAND2_X1 U9242 ( .A1(n6680), .A2(n6679), .ZN(n6678) );
  INV_X1 U9243 ( .A(n9202), .ZN(n6973) );
  AOI22_X1 U9244 ( .A1(n13751), .A2(n14096), .B1(P2_REG1_REG_27__SCAN_IN), 
        .B2(n15567), .ZN(n7180) );
  INV_X1 U9245 ( .A(n6969), .ZN(P2_U3522) );
  AOI21_X1 U9246 ( .B1(n14128), .B2(n14101), .A(n6970), .ZN(n6969) );
  NAND2_X1 U9247 ( .A1(n6605), .A2(n6971), .ZN(n6970) );
  OR2_X1 U9248 ( .A1(n14101), .A2(n6972), .ZN(n6971) );
  AOI21_X1 U9249 ( .B1(n12577), .B2(n14153), .A(n7403), .ZN(n7402) );
  AOI22_X1 U9250 ( .A1(n13751), .A2(n14153), .B1(P2_REG0_REG_27__SCAN_IN), 
        .B2(n15559), .ZN(n7032) );
  NAND2_X1 U9251 ( .A1(n14127), .A2(n15561), .ZN(n7772) );
  INV_X1 U9252 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n7771) );
  OR2_X1 U9253 ( .A1(n15561), .A2(n6975), .ZN(n6974) );
  NAND2_X1 U9254 ( .A1(n15087), .A2(n14357), .ZN(n6920) );
  OAI21_X1 U9255 ( .B1(n14629), .B2(n14628), .A(n14627), .ZN(n14630) );
  INV_X1 U9256 ( .A(n6923), .ZN(n6922) );
  OAI211_X1 U9257 ( .C1(n15089), .C2(n15340), .A(n7750), .B(n7749), .ZN(
        P1_U3267) );
  AOI21_X1 U9258 ( .B1(n15086), .B2(n15235), .A(n14816), .ZN(n7749) );
  NAND2_X1 U9259 ( .A1(n7751), .A2(n14865), .ZN(n7750) );
  INV_X1 U9260 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7053) );
  NAND2_X1 U9261 ( .A1(n15205), .A2(n15206), .ZN(n15204) );
  INV_X1 U9262 ( .A(n6812), .ZN(n15205) );
  INV_X1 U9263 ( .A(n7610), .ZN(n15212) );
  NOR2_X1 U9264 ( .A1(n15268), .A2(n15267), .ZN(n15266) );
  AND2_X1 U9265 ( .A1(n7610), .A2(n7609), .ZN(n15268) );
  INV_X1 U9266 ( .A(n7082), .ZN(n15274) );
  INV_X1 U9267 ( .A(n6814), .ZN(n15272) );
  NOR2_X1 U9268 ( .A1(n15279), .A2(n15278), .ZN(n15277) );
  NOR2_X1 U9269 ( .A1(n7601), .A2(n7085), .ZN(n15282) );
  AND2_X1 U9270 ( .A1(n7601), .A2(n7085), .ZN(n15283) );
  INV_X1 U9271 ( .A(n7606), .ZN(n15285) );
  NOR2_X1 U9272 ( .A1(n15248), .A2(n15247), .ZN(n15246) );
  AND2_X1 U9273 ( .A1(n7606), .A2(n7605), .ZN(n15248) );
  OAI21_X1 U9274 ( .B1(n15195), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6486), .ZN(
        n6940) );
  CLKBUF_X3 U9276 ( .A(n8579), .Z(n8707) );
  INV_X2 U9277 ( .A(n8579), .ZN(n8650) );
  NOR2_X1 U9278 ( .A1(n12309), .A2(n7562), .ZN(n6441) );
  NAND2_X1 U9279 ( .A1(n8721), .A2(n8720), .ZN(n14016) );
  INV_X1 U9280 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14166) );
  INV_X1 U9281 ( .A(n14467), .ZN(n14446) );
  INV_X2 U9282 ( .A(n14541), .ZN(n14530) );
  INV_X1 U9283 ( .A(n11370), .ZN(n15343) );
  NOR2_X1 U9284 ( .A1(n6880), .A2(n7579), .ZN(n9761) );
  NAND2_X1 U9285 ( .A1(n9863), .A2(n9862), .ZN(n9865) );
  AND2_X1 U9286 ( .A1(n11808), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U9287 ( .A1(n6529), .A2(n6711), .ZN(n6445) );
  INV_X1 U9288 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10738) );
  AND2_X1 U9289 ( .A1(n9409), .A2(n9398), .ZN(n6446) );
  AND2_X1 U9290 ( .A1(n14129), .A2(n7409), .ZN(n6447) );
  INV_X1 U9291 ( .A(n13860), .ZN(n13655) );
  AND2_X1 U9292 ( .A1(n8325), .A2(n8324), .ZN(n13860) );
  AND2_X1 U9293 ( .A1(n7391), .A2(n6620), .ZN(n6448) );
  AOI21_X1 U9294 ( .B1(n7366), .B2(n14363), .A(n9610), .ZN(n7365) );
  INV_X1 U9295 ( .A(n7365), .ZN(n7364) );
  INV_X1 U9296 ( .A(n13334), .ZN(n7123) );
  XNOR2_X1 U9297 ( .A(n13751), .B(n13760), .ZN(n13737) );
  INV_X1 U9298 ( .A(n13737), .ZN(n6696) );
  NAND2_X1 U9299 ( .A1(n9995), .A2(n12971), .ZN(n6449) );
  INV_X1 U9300 ( .A(n7766), .ZN(n7765) );
  AND2_X1 U9301 ( .A1(n15278), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6450) );
  INV_X1 U9302 ( .A(n12483), .ZN(n13433) );
  INV_X1 U9303 ( .A(n7581), .ZN(n12941) );
  OR2_X1 U9304 ( .A1(n13427), .A2(n12551), .ZN(n7581) );
  INV_X1 U9305 ( .A(n14137), .ZN(n7410) );
  AND3_X1 U9306 ( .A1(n8903), .A2(n7379), .A3(n6549), .ZN(n6451) );
  AND2_X1 U9307 ( .A1(n8824), .A2(n8825), .ZN(n6452) );
  AND3_X1 U9308 ( .A1(n8820), .A2(n10744), .A3(n7474), .ZN(n6453) );
  AND2_X1 U9309 ( .A1(n7979), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6454) );
  INV_X1 U9310 ( .A(n7643), .ZN(n7642) );
  OAI21_X1 U9311 ( .B1(n7647), .B2(n7644), .A(n8658), .ZN(n7643) );
  OR2_X1 U9312 ( .A1(n7559), .A2(n7822), .ZN(n6455) );
  AND2_X1 U9313 ( .A1(n6447), .A2(n7408), .ZN(n6456) );
  AND2_X1 U9314 ( .A1(n6976), .A2(n6974), .ZN(n6457) );
  NOR2_X1 U9315 ( .A1(n8160), .A2(n8159), .ZN(n6458) );
  NOR2_X1 U9316 ( .A1(n14889), .A2(n14870), .ZN(n6459) );
  AND2_X1 U9317 ( .A1(n7281), .A2(n7282), .ZN(n6460) );
  NAND2_X1 U9318 ( .A1(n9338), .A2(n9337), .ZN(n6461) );
  OR2_X1 U9319 ( .A1(n11229), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n6462) );
  AND2_X1 U9320 ( .A1(n7287), .A2(n6544), .ZN(n6463) );
  NAND2_X1 U9321 ( .A1(n8704), .A2(n8703), .ZN(n13999) );
  INV_X1 U9322 ( .A(n13999), .ZN(n7406) );
  AND2_X1 U9323 ( .A1(n7505), .A2(n6614), .ZN(n6464) );
  OR2_X1 U9324 ( .A1(n14649), .A2(n14413), .ZN(n6465) );
  INV_X1 U9325 ( .A(n15569), .ZN(n15567) );
  XNOR2_X1 U9326 ( .A(n8959), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U9327 ( .A1(n11937), .A2(n15259), .ZN(n11938) );
  OR2_X1 U9328 ( .A1(n15645), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n6466) );
  AND2_X1 U9329 ( .A1(n8445), .A2(SI_26_), .ZN(n6467) );
  AND2_X1 U9330 ( .A1(n7157), .A2(n7156), .ZN(n6468) );
  AND2_X1 U9331 ( .A1(n8940), .A2(n8939), .ZN(n14811) );
  AND2_X1 U9332 ( .A1(n7530), .A2(n8066), .ZN(n6469) );
  INV_X1 U9333 ( .A(n14639), .ZN(n14522) );
  INV_X1 U9334 ( .A(n7943), .ZN(n8002) );
  AND2_X2 U9335 ( .A1(n13718), .A2(n8784), .ZN(n14008) );
  NAND2_X1 U9336 ( .A1(n10146), .A2(n10145), .ZN(n13451) );
  NAND2_X1 U9337 ( .A1(n6686), .A2(n7523), .ZN(n6470) );
  OR2_X1 U9338 ( .A1(n8120), .A2(n8119), .ZN(n6471) );
  OR2_X1 U9339 ( .A1(n8377), .A2(n8349), .ZN(n6472) );
  AND2_X1 U9340 ( .A1(n8899), .A2(n8896), .ZN(n11711) );
  NAND2_X1 U9341 ( .A1(n8881), .A2(n8880), .ZN(n15399) );
  INV_X1 U9342 ( .A(n15214), .ZN(n6806) );
  AND2_X1 U9343 ( .A1(n15307), .A2(n6638), .ZN(n6473) );
  AND2_X1 U9344 ( .A1(n13525), .A2(n8183), .ZN(n13571) );
  AND3_X1 U9345 ( .A1(n7056), .A2(n8973), .A3(n8953), .ZN(n6474) );
  OR2_X1 U9346 ( .A1(n14864), .A2(n14863), .ZN(n14862) );
  AND2_X1 U9347 ( .A1(n10416), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7579) );
  AND2_X1 U9348 ( .A1(n8254), .A2(n8250), .ZN(n6475) );
  OR2_X1 U9349 ( .A1(n14838), .A2(n14266), .ZN(n6476) );
  AND2_X1 U9350 ( .A1(n9758), .A2(n15594), .ZN(n6477) );
  NAND2_X1 U9351 ( .A1(n6710), .A2(n8984), .ZN(n10393) );
  AND2_X1 U9352 ( .A1(n9029), .A2(n7679), .ZN(n6478) );
  NAND2_X1 U9353 ( .A1(n10278), .A2(n10277), .ZN(n12483) );
  INV_X1 U9354 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8827) );
  INV_X1 U9355 ( .A(n8611), .ZN(n7657) );
  INV_X1 U9356 ( .A(n9043), .ZN(n11309) );
  INV_X1 U9357 ( .A(n12835), .ZN(n7717) );
  INV_X1 U9358 ( .A(n12884), .ZN(n7118) );
  AND2_X1 U9359 ( .A1(n10798), .A2(n10058), .ZN(n6479) );
  OR2_X1 U9360 ( .A1(n13541), .A2(n13794), .ZN(n6480) );
  NAND2_X1 U9361 ( .A1(n15104), .A2(n12423), .ZN(n6481) );
  AND2_X1 U9362 ( .A1(n7646), .A2(n7645), .ZN(n6482) );
  AND2_X1 U9363 ( .A1(n7778), .A2(n6628), .ZN(n6483) );
  AND2_X1 U9364 ( .A1(n9440), .A2(n9439), .ZN(n6484) );
  OR2_X1 U9365 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9155), .ZN(n6485) );
  OR2_X1 U9366 ( .A1(n9181), .A2(n9180), .ZN(n6486) );
  OR2_X1 U9367 ( .A1(n9162), .A2(n9161), .ZN(n6487) );
  AND3_X1 U9368 ( .A1(n7946), .A2(n7944), .A3(n7945), .ZN(n6488) );
  AND2_X1 U9369 ( .A1(n9082), .A2(n7272), .ZN(n6489) );
  NOR2_X1 U9370 ( .A1(n7655), .A2(n8648), .ZN(n6490) );
  NAND2_X2 U9371 ( .A1(n7790), .A2(n13507), .ZN(n9822) );
  AND2_X1 U9372 ( .A1(n13223), .A2(n12964), .ZN(n6491) );
  INV_X1 U9373 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6641) );
  INV_X1 U9374 ( .A(n13871), .ZN(n7787) );
  AND2_X1 U9375 ( .A1(n13719), .A2(n13971), .ZN(n6492) );
  AND2_X1 U9376 ( .A1(n9847), .A2(n7163), .ZN(n6493) );
  AND2_X1 U9377 ( .A1(n6672), .A2(n6670), .ZN(n6494) );
  NAND2_X1 U9378 ( .A1(n8919), .A2(n8918), .ZN(n15137) );
  INV_X1 U9379 ( .A(n15131), .ZN(n14941) );
  NAND2_X1 U9380 ( .A1(n7313), .A2(n7310), .ZN(n7309) );
  INV_X1 U9381 ( .A(n10934), .ZN(n11089) );
  AND2_X1 U9382 ( .A1(n7582), .A2(n6864), .ZN(n6495) );
  AND2_X1 U9383 ( .A1(n7747), .A2(n7065), .ZN(n6496) );
  INV_X1 U9384 ( .A(n6837), .ZN(n8010) );
  XNOR2_X1 U9385 ( .A(n8011), .B(n6778), .ZN(n6837) );
  INV_X1 U9386 ( .A(n14972), .ZN(n7743) );
  INV_X1 U9387 ( .A(n11423), .ZN(n7150) );
  INV_X1 U9388 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U9389 ( .A1(n8898), .A2(n8897), .ZN(n15036) );
  AND4_X1 U9390 ( .A1(n9763), .A2(n9703), .A3(n9679), .A4(n9678), .ZN(n6497)
         );
  AND3_X1 U9391 ( .A1(n8204), .A2(n8203), .A3(n8202), .ZN(n13641) );
  INV_X1 U9392 ( .A(n10924), .ZN(n11018) );
  XNOR2_X1 U9393 ( .A(n9776), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10924) );
  OR2_X1 U9394 ( .A1(n12837), .A2(n12838), .ZN(n6498) );
  AND2_X1 U9395 ( .A1(n8627), .A2(n8628), .ZN(n6499) );
  NAND2_X1 U9396 ( .A1(n15006), .A2(n7482), .ZN(n7811) );
  AOI21_X1 U9397 ( .B1(n12403), .B2(n8948), .A(n8947), .ZN(n15066) );
  INV_X1 U9398 ( .A(n13134), .ZN(n13039) );
  BUF_X1 U9399 ( .A(n13517), .Z(n7029) );
  INV_X1 U9400 ( .A(n8651), .ZN(n6903) );
  AND2_X1 U9401 ( .A1(n13132), .A2(n13131), .ZN(n6500) );
  NAND2_X1 U9402 ( .A1(n8914), .A2(n8913), .ZN(n15142) );
  NAND2_X1 U9403 ( .A1(n7502), .A2(n7504), .ZN(n7501) );
  AND2_X1 U9404 ( .A1(n7524), .A2(n7525), .ZN(n8014) );
  AND2_X1 U9405 ( .A1(n12258), .A2(n6461), .ZN(n6501) );
  AND2_X1 U9406 ( .A1(n6665), .A2(n6664), .ZN(n6502) );
  AND2_X1 U9407 ( .A1(n8553), .A2(n13610), .ZN(n6503) );
  AND3_X1 U9408 ( .A1(n12857), .A2(n12856), .A3(n12858), .ZN(n6504) );
  AND2_X1 U9409 ( .A1(n7560), .A2(n13564), .ZN(n6505) );
  AND2_X1 U9410 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6506) );
  NAND2_X1 U9411 ( .A1(n12495), .A2(n12494), .ZN(n13427) );
  AND2_X1 U9412 ( .A1(n12110), .A2(n11984), .ZN(n6507) );
  AND2_X1 U9413 ( .A1(n12934), .A2(n12931), .ZN(n6508) );
  INV_X1 U9414 ( .A(n13882), .ZN(n14059) );
  AND2_X1 U9415 ( .A1(n8281), .A2(n8280), .ZN(n13882) );
  NOR2_X1 U9416 ( .A1(n13410), .A2(n12969), .ZN(n6509) );
  NAND2_X1 U9417 ( .A1(n7661), .A2(n7832), .ZN(n8978) );
  AND2_X1 U9418 ( .A1(n8009), .A2(n8008), .ZN(n6510) );
  NOR2_X1 U9419 ( .A1(n6440), .A2(n9266), .ZN(n6511) );
  INV_X1 U9420 ( .A(n14161), .ZN(n12171) );
  AND2_X1 U9421 ( .A1(n8100), .A2(n8099), .ZN(n14161) );
  AND2_X1 U9422 ( .A1(n9973), .A2(n9996), .ZN(n6512) );
  INV_X1 U9423 ( .A(n13760), .ZN(n13635) );
  NAND2_X1 U9424 ( .A1(n8465), .A2(n8464), .ZN(n13760) );
  AND2_X1 U9425 ( .A1(n9103), .A2(n7599), .ZN(n6513) );
  NOR2_X1 U9426 ( .A1(n15501), .A2(n15500), .ZN(n6514) );
  NAND2_X1 U9427 ( .A1(n13920), .A2(n13893), .ZN(n6515) );
  INV_X1 U9428 ( .A(n12046), .ZN(n15543) );
  AND2_X1 U9429 ( .A1(n8001), .A2(n8000), .ZN(n12046) );
  NOR2_X1 U9430 ( .A1(n9062), .A2(n7763), .ZN(n6516) );
  OR2_X1 U9431 ( .A1(n12504), .A2(n14637), .ZN(n6517) );
  INV_X1 U9432 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8844) );
  AND2_X1 U9433 ( .A1(n7773), .A2(n14037), .ZN(n6518) );
  AND2_X1 U9434 ( .A1(n6939), .A2(n7561), .ZN(n6519) );
  NOR2_X1 U9435 ( .A1(n10192), .A2(n13264), .ZN(n6520) );
  INV_X1 U9436 ( .A(n14422), .ZN(n7476) );
  NAND2_X1 U9437 ( .A1(n14474), .A2(n14475), .ZN(n14921) );
  OR2_X1 U9438 ( .A1(n13737), .A2(n7668), .ZN(n6521) );
  AND2_X1 U9439 ( .A1(n10946), .A2(n10934), .ZN(n6522) );
  INV_X1 U9440 ( .A(n7030), .ZN(n14906) );
  NOR2_X1 U9441 ( .A1(n14905), .A2(n15122), .ZN(n7030) );
  AND2_X1 U9442 ( .A1(n13841), .A2(n13789), .ZN(n6523) );
  AND2_X1 U9443 ( .A1(n13563), .A2(n7559), .ZN(n6524) );
  INV_X1 U9444 ( .A(n13839), .ZN(n7786) );
  INV_X1 U9445 ( .A(n9168), .ZN(n7085) );
  AND2_X1 U9446 ( .A1(n8413), .A2(n6832), .ZN(n6525) );
  NAND3_X1 U9447 ( .A1(n12929), .A2(n12928), .A3(n12927), .ZN(n6526) );
  AND2_X1 U9448 ( .A1(n7663), .A2(n7174), .ZN(n6527) );
  AND2_X1 U9449 ( .A1(n14562), .A2(n14563), .ZN(n6528) );
  OR2_X1 U9450 ( .A1(n9559), .A2(n9558), .ZN(n6529) );
  AND2_X1 U9451 ( .A1(n12417), .A2(n12416), .ZN(n6530) );
  AND2_X1 U9452 ( .A1(n9363), .A2(n7836), .ZN(n6531) );
  AND2_X1 U9453 ( .A1(n12422), .A2(n12421), .ZN(n14880) );
  INV_X1 U9454 ( .A(n7637), .ZN(n7636) );
  NAND2_X1 U9455 ( .A1(n6481), .A2(n12422), .ZN(n7637) );
  OR2_X1 U9456 ( .A1(n12342), .A2(n11717), .ZN(n6532) );
  NAND2_X1 U9457 ( .A1(n9089), .A2(n7820), .ZN(n6533) );
  AND2_X1 U9458 ( .A1(n6480), .A2(n13802), .ZN(n6534) );
  INV_X1 U9459 ( .A(n12462), .ZN(n14607) );
  NAND2_X1 U9460 ( .A1(n12407), .A2(n12587), .ZN(n12462) );
  AND2_X1 U9461 ( .A1(n7506), .A2(n7097), .ZN(n6535) );
  INV_X1 U9462 ( .A(n11622), .ZN(n14404) );
  AND2_X1 U9463 ( .A1(n7069), .A2(n12462), .ZN(n6536) );
  AND2_X1 U9464 ( .A1(n6479), .A2(n6893), .ZN(n6537) );
  INV_X1 U9465 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9692) );
  INV_X1 U9466 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8824) );
  AND2_X1 U9467 ( .A1(n7626), .A2(n7625), .ZN(n6538) );
  AND2_X1 U9468 ( .A1(n12832), .A2(n12833), .ZN(n12771) );
  INV_X1 U9469 ( .A(n12874), .ZN(n7729) );
  NOR2_X1 U9470 ( .A1(n14428), .A2(n15048), .ZN(n6539) );
  NOR2_X1 U9471 ( .A1(n13980), .A2(n13659), .ZN(n6540) );
  NOR2_X1 U9472 ( .A1(n14161), .A2(n12195), .ZN(n6541) );
  INV_X1 U9473 ( .A(n12782), .ZN(n13209) );
  NAND2_X1 U9474 ( .A1(n12926), .A2(n13196), .ZN(n12782) );
  AND2_X1 U9475 ( .A1(n13941), .A2(n13658), .ZN(n6542) );
  AND2_X1 U9476 ( .A1(n7752), .A2(n7073), .ZN(n7072) );
  NOR2_X1 U9477 ( .A1(n14651), .A2(n11622), .ZN(n6543) );
  INV_X1 U9478 ( .A(n7325), .ZN(n7324) );
  NOR2_X1 U9479 ( .A1(n11654), .A2(n12064), .ZN(n7325) );
  NAND2_X1 U9480 ( .A1(n11289), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6544) );
  INV_X1 U9481 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10708) );
  OR2_X1 U9482 ( .A1(n8628), .A2(n8627), .ZN(n7628) );
  NAND2_X1 U9483 ( .A1(n13187), .A2(n13193), .ZN(n6545) );
  INV_X1 U9484 ( .A(n13739), .ZN(n7274) );
  NAND2_X1 U9485 ( .A1(n8448), .A2(n8447), .ZN(n14026) );
  INV_X1 U9486 ( .A(n14026), .ZN(n6692) );
  AND2_X1 U9487 ( .A1(n7256), .A2(n12431), .ZN(n6546) );
  NOR2_X1 U9488 ( .A1(n13391), .A2(n13265), .ZN(n6547) );
  NOR2_X1 U9489 ( .A1(n14838), .A2(n14641), .ZN(n6548) );
  AND4_X1 U9490 ( .A1(n8956), .A2(n8955), .A3(n10744), .A4(n8952), .ZN(n6549)
         );
  INV_X1 U9491 ( .A(n7822), .ZN(n7560) );
  OR2_X1 U9492 ( .A1(n8869), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6550) );
  AND2_X1 U9493 ( .A1(n7166), .A2(n6845), .ZN(n6551) );
  INV_X1 U9494 ( .A(n12577), .ZN(n14116) );
  NAND2_X1 U9495 ( .A1(n8693), .A2(n8692), .ZN(n12577) );
  AND2_X1 U9496 ( .A1(n7085), .A2(n7084), .ZN(n6552) );
  AND2_X1 U9497 ( .A1(n13262), .A2(n12906), .ZN(n6553) );
  AND2_X1 U9498 ( .A1(n7067), .A2(n7069), .ZN(n6554) );
  INV_X1 U9499 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10441) );
  NOR2_X1 U9500 ( .A1(n9609), .A2(n9608), .ZN(n9610) );
  INV_X1 U9501 ( .A(n13212), .ZN(n12962) );
  AND2_X1 U9502 ( .A1(n10288), .A2(n10287), .ZN(n13212) );
  AND2_X1 U9503 ( .A1(n10939), .A2(n10938), .ZN(n6555) );
  NOR2_X1 U9504 ( .A1(n15077), .A2(n15082), .ZN(n6556) );
  AND2_X1 U9505 ( .A1(n9080), .A2(n8786), .ZN(n13772) );
  INV_X1 U9506 ( .A(n13772), .ZN(n7265) );
  INV_X1 U9507 ( .A(n6869), .ZN(n12796) );
  AND2_X1 U9508 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  AND2_X1 U9509 ( .A1(n9504), .A2(n9503), .ZN(n6557) );
  AND2_X1 U9510 ( .A1(n10412), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U9511 ( .A1(n8251), .A2(n8250), .ZN(n6559) );
  NAND2_X1 U9512 ( .A1(n10664), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6560) );
  OR2_X1 U9513 ( .A1(n8255), .A2(n8254), .ZN(n6561) );
  INV_X1 U9514 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10418) );
  NAND2_X1 U9515 ( .A1(n14986), .A2(n14972), .ZN(n6562) );
  AND2_X1 U9516 ( .A1(n12843), .A2(n12842), .ZN(n6563) );
  AND2_X1 U9517 ( .A1(n6482), .A2(n7639), .ZN(n6564) );
  XOR2_X1 U9518 ( .A(n9188), .B(n9187), .Z(n6565) );
  NOR2_X1 U9519 ( .A1(n7452), .A2(n7450), .ZN(n6566) );
  AND2_X1 U9520 ( .A1(n12069), .A2(n12975), .ZN(n6567) );
  AND2_X1 U9521 ( .A1(n7501), .A2(n7498), .ZN(n6568) );
  NAND3_X1 U9522 ( .A1(n7438), .A2(n14465), .A3(n7437), .ZN(n6569) );
  AND2_X1 U9523 ( .A1(n7515), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U9524 ( .A1(n15082), .A2(n14365), .ZN(n12587) );
  INV_X1 U9525 ( .A(n14425), .ZN(n7456) );
  NAND2_X1 U9526 ( .A1(n7728), .A2(n13350), .ZN(n6571) );
  INV_X1 U9527 ( .A(n14511), .ZN(n7413) );
  INV_X1 U9528 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10467) );
  INV_X1 U9529 ( .A(n7724), .ZN(n7723) );
  NAND2_X1 U9530 ( .A1(n7727), .A2(n7123), .ZN(n7724) );
  INV_X1 U9531 ( .A(n7309), .ZN(n7308) );
  INV_X1 U9532 ( .A(n7117), .ZN(n7116) );
  NAND2_X1 U9533 ( .A1(n13334), .A2(n12884), .ZN(n7117) );
  INV_X1 U9534 ( .A(n7473), .ZN(n7472) );
  NAND2_X1 U9535 ( .A1(n14524), .A2(n14523), .ZN(n7473) );
  INV_X1 U9536 ( .A(n14518), .ZN(n7449) );
  NAND2_X1 U9537 ( .A1(n14862), .A2(n12457), .ZN(n14836) );
  AND2_X1 U9538 ( .A1(n13492), .A2(n12971), .ZN(n6572) );
  AND2_X1 U9539 ( .A1(n8370), .A2(n8365), .ZN(n6573) );
  OR2_X1 U9540 ( .A1(n9148), .A2(n9147), .ZN(n6574) );
  NAND2_X1 U9541 ( .A1(n14825), .A2(n14811), .ZN(n12435) );
  AND2_X1 U9542 ( .A1(n7831), .A2(n7200), .ZN(n6575) );
  NOR2_X1 U9543 ( .A1(n7019), .A2(n8005), .ZN(n6576) );
  INV_X1 U9544 ( .A(n15046), .ZN(n7078) );
  AND2_X1 U9545 ( .A1(n8121), .A2(n8144), .ZN(n6577) );
  NOR2_X1 U9546 ( .A1(n8018), .A2(n7887), .ZN(n6578) );
  AND2_X1 U9547 ( .A1(n12784), .A2(n6991), .ZN(n6579) );
  AND2_X1 U9548 ( .A1(n13920), .A2(n13933), .ZN(n6580) );
  AND2_X1 U9549 ( .A1(n14458), .A2(n14449), .ZN(n6581) );
  AND2_X1 U9550 ( .A1(n8161), .A2(n8143), .ZN(n8144) );
  INV_X1 U9551 ( .A(n8144), .ZN(n7186) );
  AND2_X1 U9552 ( .A1(n11242), .A2(n11240), .ZN(n6582) );
  AND2_X1 U9553 ( .A1(n10944), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6583) );
  AND2_X1 U9554 ( .A1(n13395), .A2(n13307), .ZN(n12888) );
  AND2_X1 U9555 ( .A1(n7214), .A2(n7213), .ZN(n6584) );
  AND2_X1 U9556 ( .A1(n13790), .A2(n9072), .ZN(n13826) );
  INV_X1 U9557 ( .A(n13826), .ZN(n7177) );
  AND2_X1 U9558 ( .A1(n13005), .A2(n13004), .ZN(n6585) );
  AND2_X1 U9559 ( .A1(n7837), .A2(n7818), .ZN(n6586) );
  AND2_X1 U9560 ( .A1(n7187), .A2(n6471), .ZN(n6587) );
  INV_X1 U9561 ( .A(n7211), .ZN(n7210) );
  NOR2_X1 U9562 ( .A1(n13228), .A2(n13215), .ZN(n7211) );
  AND2_X1 U9563 ( .A1(n9379), .A2(n9366), .ZN(n6588) );
  AND2_X1 U9564 ( .A1(n7662), .A2(n6480), .ZN(n6589) );
  NAND2_X1 U9565 ( .A1(n14532), .A2(n7418), .ZN(n6590) );
  OR2_X1 U9566 ( .A1(n7658), .A2(n7657), .ZN(n6591) );
  AND2_X1 U9567 ( .A1(n6901), .A2(n6899), .ZN(n6592) );
  AND2_X1 U9568 ( .A1(n9693), .A2(n9692), .ZN(n6593) );
  AND2_X1 U9569 ( .A1(n7802), .A2(n10322), .ZN(n6594) );
  AND2_X1 U9570 ( .A1(n7095), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6595) );
  NOR2_X1 U9571 ( .A1(n8647), .A2(n8649), .ZN(n6596) );
  INV_X1 U9572 ( .A(n7130), .ZN(n7129) );
  INV_X1 U9573 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8955) );
  INV_X1 U9574 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6686) );
  AND2_X1 U9575 ( .A1(n7627), .A2(n7628), .ZN(n6597) );
  OR2_X1 U9576 ( .A1(n7444), .A2(n7443), .ZN(n6598) );
  NAND2_X1 U9577 ( .A1(n14426), .A2(n7456), .ZN(n6599) );
  NAND2_X1 U9578 ( .A1(n14512), .A2(n7413), .ZN(n6600) );
  NAND2_X1 U9579 ( .A1(n7254), .A2(n7249), .ZN(n6601) );
  AND2_X2 U9580 ( .A1(n9194), .A2(n13956), .ZN(n13909) );
  NOR2_X1 U9581 ( .A1(n13146), .A2(n10218), .ZN(n6602) );
  NAND2_X1 U9582 ( .A1(n11740), .A2(n7374), .ZN(n7373) );
  NAND2_X1 U9583 ( .A1(n11560), .A2(n11561), .ZN(n11559) );
  AND4_X1 U9584 ( .A1(n7233), .A2(n7232), .A3(n8904), .A4(n8820), .ZN(n7661)
         );
  INV_X1 U9585 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6675) );
  NOR2_X1 U9586 ( .A1(n12222), .A2(n7492), .ZN(n11937) );
  NAND2_X1 U9587 ( .A1(n7197), .A2(n10323), .ZN(n11797) );
  INV_X1 U9588 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n7511) );
  NAND3_X1 U9589 ( .A1(n6442), .A2(n7379), .A3(n8903), .ZN(n6603) );
  OR2_X1 U9590 ( .A1(n8003), .A2(n6994), .ZN(n6604) );
  NAND2_X1 U9591 ( .A1(n11906), .A2(n9938), .ZN(n12364) );
  INV_X2 U9592 ( .A(n15643), .ZN(n15645) );
  INV_X1 U9593 ( .A(n11879), .ZN(n7097) );
  NAND2_X1 U9594 ( .A1(n7464), .A2(n7462), .ZN(n11862) );
  INV_X1 U9595 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7239) );
  INV_X1 U9596 ( .A(SI_6_), .ZN(n6778) );
  NAND2_X1 U9597 ( .A1(n6799), .A2(n7242), .ZN(n11681) );
  OAI21_X1 U9598 ( .B1(n12618), .B2(n6896), .A(n6895), .ZN(n12687) );
  NAND2_X1 U9599 ( .A1(n9053), .A2(n9052), .ZN(n12006) );
  NAND2_X1 U9600 ( .A1(n7222), .A2(n14442), .ZN(n14985) );
  NAND2_X1 U9601 ( .A1(n7617), .A2(n11924), .ZN(n12182) );
  NAND2_X1 U9602 ( .A1(n7079), .A2(n7735), .ZN(n15039) );
  NAND2_X1 U9603 ( .A1(n7738), .A2(n11922), .ZN(n12213) );
  NAND2_X1 U9604 ( .A1(n7652), .A2(n11483), .ZN(n11589) );
  OR2_X1 U9605 ( .A1(n12766), .A2(n12912), .ZN(n13249) );
  INV_X1 U9606 ( .A(n14036), .ZN(n7408) );
  INV_X1 U9607 ( .A(n7398), .ZN(n7401) );
  OR2_X1 U9608 ( .A1(n14129), .A2(n14104), .ZN(n6605) );
  AND2_X1 U9609 ( .A1(n8290), .A2(n8289), .ZN(n6606) );
  OR2_X1 U9610 ( .A1(n14129), .A2(n14160), .ZN(n6607) );
  OR2_X1 U9611 ( .A1(n11495), .A2(n12767), .ZN(n11779) );
  INV_X1 U9612 ( .A(n13264), .ZN(n12966) );
  AND2_X1 U9613 ( .A1(n10153), .A2(n10152), .ZN(n13264) );
  NAND2_X1 U9614 ( .A1(n6648), .A2(n8029), .ZN(n11472) );
  NOR2_X1 U9615 ( .A1(n8067), .A2(n7529), .ZN(n6608) );
  NOR2_X1 U9616 ( .A1(n13187), .A2(n13382), .ZN(n6609) );
  NOR2_X1 U9617 ( .A1(n13187), .A2(n13443), .ZN(n6610) );
  AND2_X1 U9618 ( .A1(n7780), .A2(n9056), .ZN(n6611) );
  INV_X1 U9619 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6994) );
  INV_X1 U9620 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6690) );
  INV_X1 U9621 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6695) );
  OR2_X1 U9622 ( .A1(n11779), .A2(n10319), .ZN(n6612) );
  OR2_X1 U9623 ( .A1(n12192), .A2(n12193), .ZN(n12190) );
  INV_X1 U9624 ( .A(n13751), .ZN(n14121) );
  AND2_X1 U9625 ( .A1(n7725), .A2(n7723), .ZN(n6613) );
  OR2_X1 U9626 ( .A1(n12980), .A2(n12338), .ZN(n6614) );
  NAND2_X1 U9627 ( .A1(n10039), .A2(n10798), .ZN(n6615) );
  AND2_X1 U9628 ( .A1(n6643), .A2(n7759), .ZN(n6616) );
  NOR3_X1 U9629 ( .A1(n13406), .A2(n13337), .A3(n12946), .ZN(n6617) );
  INV_X1 U9630 ( .A(n7431), .ZN(n7430) );
  NAND2_X1 U9631 ( .A1(n7432), .A2(n9996), .ZN(n7431) );
  AND2_X1 U9632 ( .A1(n14369), .A2(n6920), .ZN(n6618) );
  AND2_X1 U9633 ( .A1(n7160), .A2(n7159), .ZN(n6619) );
  INV_X1 U9634 ( .A(n15310), .ZN(n6633) );
  NAND2_X1 U9635 ( .A1(n15504), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6620) );
  AND3_X1 U9636 ( .A1(n8851), .A2(n6795), .A3(n15364), .ZN(n11644) );
  INV_X1 U9637 ( .A(n14428), .ZN(n7493) );
  AND2_X1 U9638 ( .A1(n13105), .A2(n13104), .ZN(n6621) );
  XNOR2_X1 U9639 ( .A(n9152), .B(n9149), .ZN(n15202) );
  NAND2_X1 U9640 ( .A1(n6782), .A2(n11383), .ZN(n11482) );
  OR2_X1 U9641 ( .A1(n15408), .A2(n7053), .ZN(n6622) );
  NAND2_X1 U9642 ( .A1(n11203), .A2(n11204), .ZN(n11202) );
  NAND2_X1 U9643 ( .A1(n14230), .A2(n6709), .ZN(n11152) );
  AND2_X1 U9644 ( .A1(n7455), .A2(n9746), .ZN(n6623) );
  AND2_X1 U9645 ( .A1(n7285), .A2(n6463), .ZN(n6624) );
  AND2_X1 U9646 ( .A1(n7285), .A2(n7287), .ZN(n6625) );
  INV_X1 U9647 ( .A(n15652), .ZN(n7202) );
  AND3_X2 U9648 ( .A1(n10377), .A2(n11416), .A3(n10376), .ZN(n15652) );
  AND2_X1 U9649 ( .A1(n7323), .A2(n6462), .ZN(n6626) );
  INV_X1 U9650 ( .A(n11168), .ZN(n6676) );
  INV_X1 U9651 ( .A(n13705), .ZN(n11614) );
  XNOR2_X1 U9652 ( .A(n9688), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12797) );
  INV_X1 U9653 ( .A(n11124), .ZN(n7519) );
  INV_X1 U9654 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n7161) );
  INV_X1 U9655 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7152) );
  NAND2_X1 U9656 ( .A1(n13146), .A2(n11540), .ZN(n12800) );
  INV_X1 U9657 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U9658 ( .A1(n7514), .A2(n11018), .ZN(n10984) );
  NAND2_X1 U9659 ( .A1(n7958), .A2(n6668), .ZN(n6667) );
  AND2_X1 U9660 ( .A1(n10908), .A2(n12952), .ZN(n6627) );
  INV_X1 U9661 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7084) );
  INV_X1 U9662 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7020) );
  INV_X1 U9663 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7622) );
  INV_X1 U9664 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7599) );
  INV_X1 U9665 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7621) );
  INV_X1 U9666 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7769) );
  AOI211_X1 U9667 ( .C1(n15081), .C2(n15235), .A(n12465), .B(n12464), .ZN(
        n12466) );
  AND2_X1 U9668 ( .A1(n10393), .A2(n10464), .ZN(n11266) );
  XNOR2_X1 U9669 ( .A(n13114), .B(n13104), .ZN(n13117) );
  NAND2_X1 U9670 ( .A1(n7090), .A2(n13104), .ZN(n13110) );
  AOI21_X1 U9671 ( .B1(n13746), .B2(n13971), .A(n13745), .ZN(n14023) );
  AOI21_X1 U9672 ( .B1(n7777), .B2(n13971), .A(n7774), .ZN(n14038) );
  AOI21_X1 U9673 ( .B1(n13813), .B2(n13971), .A(n13812), .ZN(n14041) );
  AOI21_X1 U9674 ( .B1(n7024), .B2(n13971), .A(n7021), .ZN(n14028) );
  OAI21_X4 U9675 ( .B1(n15550), .B2(n11823), .A(n13987), .ZN(n13983) );
  OAI21_X2 U9676 ( .B1(n12006), .B2(n6629), .A(n6483), .ZN(n11958) );
  NAND2_X1 U9677 ( .A1(n12004), .A2(n7781), .ZN(n6628) );
  INV_X1 U9678 ( .A(n7781), .ZN(n6629) );
  NAND2_X1 U9679 ( .A1(n12006), .A2(n12007), .ZN(n9055) );
  NAND2_X1 U9680 ( .A1(n6630), .A2(n9069), .ZN(n13875) );
  OAI22_X2 U9681 ( .A1(n13875), .A2(n9071), .B1(n13859), .B2(n14059), .ZN(
        n13856) );
  XNOR2_X1 U9682 ( .A(n14777), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14786) );
  NOR2_X2 U9683 ( .A1(n7873), .A2(n7849), .ZN(n8508) );
  AND3_X4 U9684 ( .A1(n8014), .A2(n7840), .A3(n7910), .ZN(n7843) );
  AND2_X1 U9685 ( .A1(n7257), .A2(n7258), .ZN(n7866) );
  AND3_X2 U9686 ( .A1(n7260), .A2(n7259), .A3(n7261), .ZN(n7867) );
  NAND2_X1 U9687 ( .A1(n12351), .A2(n15314), .ZN(n6638) );
  OAI21_X2 U9688 ( .B1(n6949), .B2(n9014), .A(n9013), .ZN(n11989) );
  NAND2_X2 U9689 ( .A1(n11322), .A2(n9008), .ZN(n6949) );
  NAND2_X1 U9690 ( .A1(n7266), .A2(n7264), .ZN(n13770) );
  OAI21_X1 U9691 ( .B1(n8831), .B2(n8827), .A(P1_IR_REG_2__SCAN_IN), .ZN(n6642) );
  NOR2_X2 U9692 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8831) );
  OAI22_X2 U9693 ( .A1(n13769), .A2(n9038), .B1(n13795), .B2(n13784), .ZN(
        n13757) );
  INV_X2 U9694 ( .A(n7967), .ZN(n8691) );
  NAND2_X2 U9695 ( .A1(n14181), .A2(n8541), .ZN(n10492) );
  XNOR2_X2 U9696 ( .A(n7854), .B(n7875), .ZN(n8541) );
  NAND2_X1 U9697 ( .A1(n11348), .A2(n11356), .ZN(n11352) );
  XNOR2_X2 U9698 ( .A(n6645), .B(n12120), .ZN(n11356) );
  AND3_X2 U9699 ( .A1(n7885), .A2(n7882), .A3(n6644), .ZN(n12120) );
  AND2_X1 U9700 ( .A1(n7884), .A2(n7883), .ZN(n6644) );
  INV_X2 U9701 ( .A(n8567), .ZN(n6645) );
  AND3_X4 U9702 ( .A1(n7864), .A2(n7865), .A3(n7863), .ZN(n8567) );
  NAND2_X1 U9703 ( .A1(n14703), .A2(n10602), .ZN(n10604) );
  NAND3_X1 U9704 ( .A1(n7262), .A2(n9049), .A3(n9048), .ZN(n12049) );
  NAND3_X1 U9705 ( .A1(n9043), .A2(n9042), .A3(n11246), .ZN(n7262) );
  NAND2_X1 U9706 ( .A1(n6647), .A2(n7526), .ZN(n11898) );
  INV_X1 U9707 ( .A(n13034), .ZN(n6652) );
  NAND2_X1 U9708 ( .A1(n13034), .A2(n13066), .ZN(n7522) );
  NAND3_X1 U9709 ( .A1(n7328), .A2(n7017), .A3(n6655), .ZN(P3_U3201) );
  NAND2_X1 U9710 ( .A1(n10885), .A2(n7966), .ZN(n11203) );
  NAND2_X1 U9711 ( .A1(n11188), .A2(n11189), .ZN(n11187) );
  NAND2_X1 U9712 ( .A1(n6660), .A2(n7505), .ZN(n12986) );
  NAND2_X1 U9713 ( .A1(n6464), .A2(n6660), .ZN(n7099) );
  NAND2_X1 U9714 ( .A1(n6535), .A2(n7507), .ZN(n6660) );
  NOR2_X4 U9715 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9763) );
  INV_X1 U9716 ( .A(n6665), .ZN(n15484) );
  NAND2_X1 U9717 ( .A1(n6677), .A2(n13707), .ZN(P2_U3233) );
  NAND2_X1 U9718 ( .A1(n13697), .A2(n15471), .ZN(n6680) );
  NAND2_X1 U9719 ( .A1(n6682), .A2(n7027), .ZN(n6681) );
  INV_X1 U9720 ( .A(n13686), .ZN(n6683) );
  INV_X1 U9721 ( .A(n12471), .ZN(n6685) );
  MUX2_X1 U9722 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n6687), .S(n15564), .Z(
        P2_U3528) );
  MUX2_X1 U9723 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n6687), .S(n15561), .Z(
        P2_U3496) );
  OAI211_X1 U9724 ( .C1(n14015), .C2(n14014), .A(n14020), .B(n14019), .ZN(
        n6687) );
  NAND3_X1 U9725 ( .A1(n6689), .A2(P2_REG3_REG_7__SCAN_IN), .A3(
        P2_REG3_REG_6__SCAN_IN), .ZN(n8055) );
  NAND3_X1 U9726 ( .A1(n6689), .A2(n6688), .A3(P2_REG3_REG_6__SCAN_IN), .ZN(
        n8057) );
  AOI21_X2 U9727 ( .B1(n13739), .B2(n9081), .A(n6696), .ZN(n7273) );
  OAI21_X2 U9728 ( .B1(n11543), .B2(n6701), .A(n6699), .ZN(n11740) );
  OR2_X1 U9729 ( .A1(n11542), .A2(n6701), .ZN(n6700) );
  INV_X1 U9730 ( .A(n9325), .ZN(n6701) );
  INV_X1 U9731 ( .A(n9246), .ZN(n6706) );
  NAND3_X1 U9732 ( .A1(n9256), .A2(n9255), .A3(n10720), .ZN(n6707) );
  AND2_X1 U9733 ( .A1(n9252), .A2(n9253), .ZN(n10654) );
  NAND2_X1 U9734 ( .A1(n9247), .A2(n9246), .ZN(n6709) );
  NAND2_X2 U9735 ( .A1(n10393), .A2(n6714), .ZN(n9284) );
  NAND3_X1 U9736 ( .A1(n6529), .A2(n6711), .A3(n14297), .ZN(n6712) );
  NAND3_X1 U9737 ( .A1(n6442), .A2(n6453), .A3(n8903), .ZN(n8923) );
  NAND4_X1 U9738 ( .A1(n6442), .A2(n6453), .A3(n8903), .A4(n8955), .ZN(n8958)
         );
  NAND2_X2 U9739 ( .A1(n7457), .A2(n6713), .ZN(n14467) );
  AOI21_X1 U9740 ( .B1(n14543), .B2(n14384), .A(n6714), .ZN(n6713) );
  INV_X1 U9741 ( .A(n14387), .ZN(n6714) );
  NAND3_X1 U9742 ( .A1(n6718), .A2(n14423), .A3(n6599), .ZN(n6717) );
  NAND2_X1 U9743 ( .A1(n7439), .A2(n6581), .ZN(n6721) );
  OAI22_X1 U9744 ( .A1(n6724), .A2(n6723), .B1(n14411), .B2(n6722), .ZN(n14415) );
  NOR2_X2 U9745 ( .A1(n7230), .A2(n7237), .ZN(n8903) );
  NAND3_X1 U9746 ( .A1(n6728), .A2(n7446), .A3(n6726), .ZN(n7445) );
  NAND2_X1 U9747 ( .A1(n6727), .A2(n14516), .ZN(n6726) );
  INV_X1 U9748 ( .A(n6730), .ZN(n6727) );
  NAND2_X1 U9749 ( .A1(n6729), .A2(n14514), .ZN(n6728) );
  NAND2_X1 U9750 ( .A1(n6730), .A2(n14515), .ZN(n6729) );
  NAND2_X1 U9751 ( .A1(n6732), .A2(n6731), .ZN(n6730) );
  NAND3_X1 U9752 ( .A1(n14510), .A2(n14509), .A3(n6600), .ZN(n6732) );
  NAND2_X1 U9753 ( .A1(n6980), .A2(n7997), .ZN(n6740) );
  NAND3_X1 U9754 ( .A1(n8032), .A2(n6836), .A3(n6737), .ZN(n7171) );
  NAND2_X1 U9755 ( .A1(n6740), .A2(n8010), .ZN(n6839) );
  XNOR2_X1 U9756 ( .A(n6740), .B(n6837), .ZN(n10417) );
  NAND2_X1 U9757 ( .A1(n6743), .A2(n6741), .ZN(n14525) );
  NAND2_X1 U9758 ( .A1(n6742), .A2(n14519), .ZN(n6741) );
  NAND2_X1 U9759 ( .A1(n6745), .A2(n14520), .ZN(n6742) );
  INV_X1 U9760 ( .A(n6745), .ZN(n6744) );
  NAND2_X1 U9761 ( .A1(n7445), .A2(n7448), .ZN(n6745) );
  XNOR2_X2 U9762 ( .A(n6753), .B(P3_IR_REG_27__SCAN_IN), .ZN(n13134) );
  AND3_X2 U9763 ( .A1(n7688), .A2(n7691), .A3(n6497), .ZN(n9734) );
  OAI21_X1 U9764 ( .B1(n7187), .B2(n7186), .A(n6767), .ZN(n6769) );
  INV_X2 U9765 ( .A(n7859), .ZN(n9755) );
  NOR2_X1 U9766 ( .A1(n6511), .A2(n6781), .ZN(n6780) );
  INV_X1 U9767 ( .A(n7245), .ZN(n6784) );
  OAI211_X2 U9768 ( .C1(n14946), .C2(n6785), .A(n6783), .B(n12419), .ZN(n14887) );
  NAND2_X2 U9769 ( .A1(n7623), .A2(n6530), .ZN(n14946) );
  OAI211_X1 U9770 ( .C1(n14869), .C2(n6788), .A(n6476), .B(n6787), .ZN(n14817)
         );
  AND2_X2 U9771 ( .A1(n14885), .A2(n12420), .ZN(n14869) );
  NAND2_X1 U9772 ( .A1(n8828), .A2(n6452), .ZN(n7244) );
  INV_X1 U9773 ( .A(n7661), .ZN(n8916) );
  XNOR2_X1 U9774 ( .A(n7860), .B(n6792), .ZN(n10453) );
  NAND2_X1 U9775 ( .A1(n7955), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6793) );
  NOR2_X1 U9776 ( .A1(n15355), .A2(n14404), .ZN(n6795) );
  INV_X1 U9777 ( .A(n11376), .ZN(n8851) );
  NAND2_X1 U9778 ( .A1(n11681), .A2(n14589), .ZN(n6798) );
  NAND2_X1 U9779 ( .A1(n7651), .A2(n7240), .ZN(n6799) );
  NAND2_X1 U9780 ( .A1(n14924), .A2(n14931), .ZN(n14905) );
  NAND2_X1 U9781 ( .A1(n6800), .A2(n15006), .ZN(n7484) );
  NOR2_X2 U9782 ( .A1(n14855), .A2(n15104), .ZN(n7485) );
  AND2_X2 U9783 ( .A1(n7030), .A2(n14895), .ZN(n14892) );
  NAND3_X1 U9784 ( .A1(n7605), .A2(n7603), .A3(n7606), .ZN(n6801) );
  XNOR2_X1 U9785 ( .A(n9148), .B(n9147), .ZN(n15655) );
  OAI21_X1 U9786 ( .B1(n15655), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6574), .ZN(
        n6809) );
  NAND2_X1 U9787 ( .A1(n11059), .A2(n11058), .ZN(n11213) );
  NAND2_X1 U9788 ( .A1(n6823), .A2(n10900), .ZN(n10981) );
  NAND2_X1 U9789 ( .A1(n11004), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U9790 ( .A1(n8414), .A2(n8413), .ZN(n8444) );
  INV_X1 U9791 ( .A(n8443), .ZN(n6832) );
  NAND2_X1 U9792 ( .A1(n8453), .A2(n13521), .ZN(n6833) );
  NAND2_X1 U9793 ( .A1(n6837), .A2(n8013), .ZN(n6836) );
  NAND2_X1 U9794 ( .A1(n7171), .A2(n6838), .ZN(n6981) );
  NAND2_X1 U9795 ( .A1(n6839), .A2(n8013), .ZN(n8031) );
  INV_X1 U9796 ( .A(n8013), .ZN(n6840) );
  NAND2_X1 U9797 ( .A1(n6841), .A2(n7333), .ZN(n8257) );
  NAND2_X1 U9798 ( .A1(n8162), .A2(n7334), .ZN(n6841) );
  NAND2_X1 U9799 ( .A1(n7955), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U9800 ( .A1(n8773), .A2(n6847), .ZN(n6897) );
  NAND4_X1 U9801 ( .A1(n8768), .A2(n6968), .A3(n8759), .A4(n8758), .ZN(n6847)
         );
  NAND2_X1 U9802 ( .A1(n10296), .A2(n6848), .ZN(n12936) );
  XNOR2_X1 U9803 ( .A(n6850), .B(n12487), .ZN(n12488) );
  INV_X1 U9804 ( .A(n6999), .ZN(n6858) );
  NAND3_X1 U9805 ( .A1(n6852), .A2(n6851), .A3(n12958), .ZN(P3_U3296) );
  NAND4_X1 U9806 ( .A1(n6857), .A2(n6627), .A3(n6856), .A4(n6855), .ZN(n6851)
         );
  NAND3_X1 U9807 ( .A1(n6997), .A2(n12799), .A3(n6999), .ZN(n6855) );
  OR2_X1 U9808 ( .A1(n6997), .A2(n12799), .ZN(n6856) );
  INV_X1 U9809 ( .A(n7103), .ZN(n6860) );
  NAND2_X1 U9810 ( .A1(n9863), .A2(n6495), .ZN(n6863) );
  NAND4_X1 U9811 ( .A1(n6871), .A2(n6508), .A3(n7581), .A4(n6870), .ZN(n6868)
         );
  OR2_X1 U9812 ( .A1(n10309), .A2(n10308), .ZN(n6870) );
  NAND2_X1 U9813 ( .A1(n9786), .A2(n11094), .ZN(n11136) );
  XNOR2_X2 U9814 ( .A(n6894), .B(n9717), .ZN(n13146) );
  NAND3_X1 U9815 ( .A1(n9682), .A2(n9683), .A3(n6593), .ZN(n10001) );
  NAND2_X1 U9816 ( .A1(n6898), .A2(n6592), .ZN(n8656) );
  NAND3_X1 U9817 ( .A1(n7025), .A2(n7026), .A3(n6902), .ZN(n6898) );
  OAI211_X1 U9818 ( .C1(n8625), .C2(n8626), .A(n6905), .B(n6597), .ZN(n6904)
         );
  NAND2_X1 U9819 ( .A1(n6906), .A2(n8624), .ZN(n6905) );
  NAND2_X1 U9820 ( .A1(n8625), .A2(n8626), .ZN(n6906) );
  NOR2_X1 U9821 ( .A1(n7849), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n7874) );
  NAND3_X1 U9822 ( .A1(n6909), .A2(n7842), .A3(n7843), .ZN(n14165) );
  NAND4_X1 U9823 ( .A1(n6909), .A2(n7842), .A3(n7843), .A4(n6908), .ZN(n6907)
         );
  OAI22_X1 U9824 ( .A1(n8614), .A2(n6912), .B1(n8613), .B2(n8612), .ZN(n8618)
         );
  NAND2_X1 U9825 ( .A1(n8618), .A2(n8619), .ZN(n8617) );
  NAND3_X1 U9826 ( .A1(n8609), .A2(n7813), .A3(n6591), .ZN(n6963) );
  AOI22_X1 U9827 ( .A1(n8642), .A2(n8641), .B1(n8640), .B2(n8639), .ZN(n8646)
         );
  NAND2_X1 U9828 ( .A1(n11357), .A2(n12116), .ZN(n9041) );
  NAND2_X1 U9829 ( .A1(n9040), .A2(n11350), .ZN(n11357) );
  NAND2_X2 U9830 ( .A1(n14174), .A2(n12404), .ZN(n7019) );
  INV_X1 U9831 ( .A(n9046), .ZN(n9047) );
  NAND2_X1 U9832 ( .A1(n12166), .A2(n9059), .ZN(n12277) );
  NAND2_X1 U9833 ( .A1(n14969), .A2(n12414), .ZN(n14954) );
  NOR2_X1 U9834 ( .A1(n14817), .A2(n14830), .ZN(n14819) );
  NAND2_X2 U9835 ( .A1(n8876), .A2(n8875), .ZN(n14428) );
  NAND2_X1 U9836 ( .A1(n7171), .A2(n8034), .ZN(n8047) );
  NAND2_X1 U9837 ( .A1(n7224), .A2(n7226), .ZN(n15021) );
  NAND2_X1 U9838 ( .A1(n7339), .A2(n8037), .ZN(n6918) );
  NAND3_X1 U9839 ( .A1(n6914), .A2(n12795), .A3(n12794), .ZN(n12798) );
  NAND2_X1 U9840 ( .A1(n6869), .A2(n6959), .ZN(n6914) );
  NOR2_X1 U9841 ( .A1(n7580), .A2(n7579), .ZN(n7573) );
  INV_X1 U9842 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7855) );
  NAND2_X1 U9843 ( .A1(n7955), .A2(SI_0_), .ZN(n7891) );
  NAND2_X1 U9844 ( .A1(n14593), .A2(n12408), .ZN(n7225) );
  OR2_X1 U9845 ( .A1(n12538), .A2(n12537), .ZN(n12540) );
  NOR2_X1 U9846 ( .A1(n12793), .A2(n12788), .ZN(n6959) );
  OAI21_X1 U9847 ( .B1(n12786), .B2(n13153), .A(n12765), .ZN(n12793) );
  NAND2_X1 U9848 ( .A1(n10177), .A2(n10176), .ZN(n10179) );
  NAND2_X1 U9849 ( .A1(n9791), .A2(n9790), .ZN(n9794) );
  NAND2_X1 U9850 ( .A1(n14120), .A2(n14101), .ZN(n7181) );
  NAND2_X1 U9851 ( .A1(n14120), .A2(n15561), .ZN(n7033) );
  NAND2_X1 U9852 ( .A1(n12003), .A2(n9016), .ZN(n11974) );
  NAND2_X1 U9853 ( .A1(n11323), .A2(n11328), .ZN(n11322) );
  OAI21_X2 U9854 ( .B1(n12275), .B2(n9025), .A(n9024), .ZN(n12305) );
  NAND2_X1 U9855 ( .A1(n11243), .A2(n9007), .ZN(n11323) );
  NAND2_X1 U9856 ( .A1(n7577), .A2(n7576), .ZN(n9791) );
  NAND2_X1 U9857 ( .A1(n9942), .A2(n9941), .ZN(n9956) );
  NOR2_X1 U9858 ( .A1(n13158), .A2(n12764), .ZN(n12789) );
  NAND2_X1 U9859 ( .A1(n7587), .A2(n7588), .ZN(n9876) );
  NAND2_X1 U9860 ( .A1(n10139), .A2(n10138), .ZN(n6915) );
  NAND2_X1 U9861 ( .A1(n10110), .A2(n10109), .ZN(n10139) );
  XNOR2_X1 U9862 ( .A(n6940), .B(n6565), .ZN(SUB_1596_U4) );
  OAI22_X1 U9863 ( .A1(n12687), .A2(n12688), .B1(n13326), .B2(n10067), .ZN(
        n12709) );
  NAND2_X1 U9864 ( .A1(n12620), .A2(n6449), .ZN(n7427) );
  OAI22_X2 U9865 ( .A1(n14290), .A2(n9458), .B1(n9457), .B2(n9456), .ZN(n14352) );
  NAND2_X1 U9866 ( .A1(n6921), .A2(n6618), .ZN(P1_U3240) );
  NAND2_X1 U9867 ( .A1(n14364), .A2(n14370), .ZN(n6921) );
  NOR2_X1 U9868 ( .A1(n14766), .A2(n14767), .ZN(n14776) );
  XNOR2_X1 U9869 ( .A(n14774), .B(n14773), .ZN(n14766) );
  NAND2_X1 U9870 ( .A1(n14789), .A2(n6922), .ZN(P1_U3262) );
  OAI21_X1 U9871 ( .B1(n15319), .B2(n14790), .A(n14788), .ZN(n6923) );
  NAND2_X1 U9872 ( .A1(n12005), .A2(n12004), .ZN(n12003) );
  NAND2_X1 U9873 ( .A1(n12559), .A2(n15645), .ZN(n6992) );
  NAND2_X1 U9874 ( .A1(n6992), .A2(n6466), .ZN(n12560) );
  XNOR2_X1 U9875 ( .A(n8840), .B(n8844), .ZN(n10616) );
  NAND2_X1 U9876 ( .A1(n7692), .A2(n7693), .ZN(n11505) );
  INV_X1 U9877 ( .A(n7697), .ZN(n7696) );
  NAND2_X1 U9878 ( .A1(n13062), .A2(n13061), .ZN(n13090) );
  NOR2_X1 U9879 ( .A1(n13003), .A2(n6585), .ZN(n13051) );
  NAND2_X1 U9880 ( .A1(n11023), .A2(n10898), .ZN(n10899) );
  INV_X1 U9881 ( .A(n8605), .ZN(n6962) );
  NAND2_X1 U9882 ( .A1(n6930), .A2(n6929), .ZN(n8598) );
  NAND2_X1 U9883 ( .A1(n6932), .A2(n6931), .ZN(n6930) );
  NAND2_X1 U9884 ( .A1(n7049), .A2(n8587), .ZN(n6932) );
  NOR2_X1 U9885 ( .A1(n6578), .A2(n7888), .ZN(n7890) );
  NAND2_X1 U9886 ( .A1(n13378), .A2(n6935), .ZN(P3_U3484) );
  NAND2_X1 U9887 ( .A1(n6936), .A2(n12246), .ZN(n6935) );
  INV_X1 U9888 ( .A(n13437), .ZN(n6936) );
  NOR2_X1 U9889 ( .A1(n13375), .A2(n6937), .ZN(n13434) );
  INV_X1 U9890 ( .A(n7190), .ZN(n7189) );
  NAND2_X1 U9891 ( .A1(n11251), .A2(n12126), .ZN(n11248) );
  NAND2_X1 U9892 ( .A1(n7550), .A2(n8249), .ZN(n7549) );
  INV_X1 U9893 ( .A(n7548), .ZN(n7547) );
  NAND2_X1 U9894 ( .A1(n7812), .A2(n13946), .ZN(n13945) );
  AOI21_X1 U9895 ( .B1(n7546), .B2(n7545), .A(n7543), .ZN(n13602) );
  NAND2_X1 U9896 ( .A1(n8111), .A2(n11896), .ZN(n12192) );
  AOI21_X1 U9897 ( .B1(n7538), .B2(n7541), .A(n7537), .ZN(n7536) );
  NAND2_X1 U9898 ( .A1(n9066), .A2(n9065), .ZN(n7766) );
  NAND2_X1 U9899 ( .A1(n9131), .A2(n9130), .ZN(n9100) );
  NAND2_X1 U9900 ( .A1(n7604), .A2(n15523), .ZN(n7603) );
  NAND2_X1 U9901 ( .A1(n9157), .A2(n9156), .ZN(n9112) );
  OAI22_X2 U9902 ( .A1(n9169), .A2(n9170), .B1(P1_ADDR_REG_15__SCAN_IN), .B2(
        n13038), .ZN(n9174) );
  NAND2_X2 U9903 ( .A1(n12456), .A2(n12455), .ZN(n14864) );
  NAND2_X1 U9904 ( .A1(n8047), .A2(n8035), .ZN(n7339) );
  INV_X1 U9905 ( .A(n7076), .ZN(n7075) );
  OAI21_X1 U9906 ( .B1(n14961), .B2(n14598), .A(n14596), .ZN(n14934) );
  INV_X1 U9907 ( .A(n7879), .ZN(n14174) );
  OAI22_X1 U9908 ( .A1(n8603), .A2(n8602), .B1(n8601), .B2(n7006), .ZN(n8605)
         );
  NAND2_X1 U9909 ( .A1(n8623), .A2(n8622), .ZN(n8625) );
  NAND2_X1 U9910 ( .A1(n9058), .A2(n12161), .ZN(n12166) );
  NAND2_X1 U9911 ( .A1(n8701), .A2(n8700), .ZN(n6948) );
  NAND2_X1 U9912 ( .A1(n6962), .A2(n6961), .ZN(n7813) );
  OAI21_X1 U9913 ( .B1(n9195), .B2(n13909), .A(n6973), .ZN(P2_U3237) );
  NAND2_X1 U9914 ( .A1(n14995), .A2(n14470), .ZN(n7483) );
  NAND2_X1 U9915 ( .A1(n7183), .A2(n7184), .ZN(n8191) );
  NAND2_X1 U9916 ( .A1(n7971), .A2(n7975), .ZN(n7166) );
  OR2_X1 U9917 ( .A1(n7141), .A2(n12908), .ZN(n7135) );
  NAND2_X1 U9918 ( .A1(n7151), .A2(n6526), .ZN(n12945) );
  NAND2_X1 U9919 ( .A1(n6960), .A2(n12951), .ZN(n7000) );
  NAND2_X1 U9920 ( .A1(n7000), .A2(n12950), .ZN(n7103) );
  NAND2_X1 U9921 ( .A1(n7133), .A2(n7137), .ZN(n7132) );
  OAI211_X1 U9922 ( .C1(n12907), .C2(n7134), .A(n7132), .B(n7140), .ZN(n7139)
         );
  NAND2_X1 U9923 ( .A1(n7434), .A2(n14397), .ZN(n6951) );
  INV_X1 U9924 ( .A(n14584), .ZN(n7435) );
  NAND3_X1 U9925 ( .A1(n14436), .A2(n14435), .A3(n6598), .ZN(n6953) );
  NAND2_X1 U9926 ( .A1(n7563), .A2(n10070), .ZN(n10088) );
  OAI21_X1 U9927 ( .B1(n14525), .B2(n7472), .A(n7469), .ZN(n14528) );
  NAND2_X1 U9928 ( .A1(n6998), .A2(n6928), .ZN(n6997) );
  NAND3_X1 U9929 ( .A1(n12949), .A2(n12948), .A3(n12947), .ZN(n6960) );
  NAND2_X1 U9930 ( .A1(n11352), .A2(n6582), .ZN(n9006) );
  NAND2_X1 U9931 ( .A1(n15664), .A2(n15665), .ZN(n9136) );
  NAND2_X1 U9932 ( .A1(n13150), .A2(n13149), .ZN(n7017) );
  NAND4_X1 U9933 ( .A1(n9770), .A2(n9769), .A3(n9768), .A4(n9767), .ZN(n10259)
         );
  OAI21_X2 U9934 ( .B1(n13247), .B2(n12912), .A(n12914), .ZN(n10311) );
  NAND2_X4 U9935 ( .A1(n13513), .A2(n13517), .ZN(n10911) );
  XNOR2_X2 U9936 ( .A(n7682), .B(n9733), .ZN(n13513) );
  AND2_X1 U9937 ( .A1(n10093), .A2(n11225), .ZN(n6958) );
  OAI21_X1 U9938 ( .B1(n13321), .B2(n13324), .A(n12882), .ZN(n13312) );
  AOI21_X1 U9939 ( .B1(n7711), .B2(n7710), .A(n6567), .ZN(n7709) );
  XNOR2_X2 U9940 ( .A(n7153), .B(P3_IR_REG_29__SCAN_IN), .ZN(n9728) );
  NAND2_X1 U9941 ( .A1(n11493), .A2(n12767), .ZN(n11492) );
  AOI21_X2 U9942 ( .B1(n12332), .B2(n12775), .A(n10262), .ZN(n12378) );
  NAND2_X1 U9943 ( .A1(n11504), .A2(n12832), .ZN(n11760) );
  OR2_X1 U9944 ( .A1(n8508), .A2(n7850), .ZN(n7851) );
  OR2_X2 U9945 ( .A1(n7948), .A2(n10453), .ZN(n7865) );
  NAND2_X1 U9946 ( .A1(n11247), .A2(n11248), .ZN(n11246) );
  NAND2_X1 U9947 ( .A1(n7566), .A2(n7564), .ZN(n10054) );
  OR2_X1 U9948 ( .A1(n7980), .A2(n10649), .ZN(n7884) );
  NAND2_X1 U9949 ( .A1(n12049), .A2(n12048), .ZN(n12047) );
  NAND2_X1 U9950 ( .A1(n6963), .A2(n7656), .ZN(n8614) );
  XNOR2_X2 U9951 ( .A(n7877), .B(n7876), .ZN(n12404) );
  OAI22_X1 U9952 ( .A1(n7943), .A2(n7622), .B1(n7019), .B2(n7621), .ZN(n7888)
         );
  NAND2_X1 U9953 ( .A1(n11991), .A2(n9015), .ZN(n12005) );
  NAND2_X1 U9954 ( .A1(n7033), .A2(n7032), .ZN(P2_U3494) );
  NAND2_X1 U9955 ( .A1(n11989), .A2(n11988), .ZN(n11991) );
  OR3_X2 U9956 ( .A1(n13719), .A2(n13951), .A3(n14011), .ZN(n7828) );
  AOI21_X1 U9957 ( .B1(n7277), .B2(n7766), .A(n6580), .ZN(n7276) );
  NOR2_X1 U9958 ( .A1(n6576), .A2(n6454), .ZN(n6965) );
  NAND2_X1 U9959 ( .A1(n6967), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U9960 ( .A1(n7015), .A2(n7016), .ZN(n6968) );
  NOR2_X1 U9961 ( .A1(n8680), .A2(n8679), .ZN(n7015) );
  NAND2_X1 U9962 ( .A1(n13825), .A2(n13790), .ZN(n13807) );
  NAND2_X1 U9963 ( .A1(n6457), .A2(n6607), .ZN(P2_U3490) );
  NAND2_X1 U9964 ( .A1(n9005), .A2(n9006), .ZN(n11243) );
  NAND2_X1 U9965 ( .A1(n7857), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7330) );
  NAND2_X1 U9966 ( .A1(n6981), .A2(n7340), .ZN(n7170) );
  NAND2_X1 U9967 ( .A1(n14868), .A2(n7636), .ZN(n7630) );
  NAND2_X1 U9968 ( .A1(n14887), .A2(n14886), .ZN(n14885) );
  NAND2_X1 U9969 ( .A1(n7671), .A2(n7674), .ZN(n12275) );
  NAND2_X1 U9970 ( .A1(n6983), .A2(n7186), .ZN(n8146) );
  INV_X1 U9971 ( .A(n8145), .ZN(n6983) );
  NAND2_X1 U9972 ( .A1(n7217), .A2(n10340), .ZN(n7214) );
  XNOR2_X1 U9973 ( .A(n6984), .B(n10346), .ZN(n10350) );
  NAND2_X1 U9974 ( .A1(n6986), .A2(n6985), .ZN(n6984) );
  NAND2_X1 U9975 ( .A1(n13210), .A2(n7207), .ZN(n6986) );
  OAI21_X1 U9976 ( .B1(n10378), .B2(n7202), .A(n6987), .ZN(P3_U3486) );
  OAI21_X1 U9977 ( .B1(n10378), .B2(n15643), .A(n6989), .ZN(P3_U3454) );
  INV_X1 U9978 ( .A(n7527), .ZN(n7526) );
  NAND4_X1 U9979 ( .A1(n12787), .A2(n12950), .A3(n12947), .A4(n12951), .ZN(
        n6998) );
  NAND2_X1 U9980 ( .A1(n12798), .A2(n12797), .ZN(n6999) );
  OAI21_X1 U9981 ( .B1(n12753), .B2(n12752), .A(n12751), .ZN(n12755) );
  NAND2_X1 U9982 ( .A1(n8974), .A2(n8973), .ZN(n8976) );
  NAND2_X1 U9983 ( .A1(n7234), .A2(n7231), .ZN(n7230) );
  NAND2_X1 U9984 ( .A1(n11152), .A2(n11154), .ZN(n11153) );
  OR2_X1 U9985 ( .A1(n10967), .A2(n10968), .ZN(n10965) );
  NAND2_X1 U9986 ( .A1(n11025), .A2(n11024), .ZN(n11023) );
  OAI21_X1 U9987 ( .B1(n8828), .B2(n8827), .A(P1_IR_REG_27__SCAN_IN), .ZN(
        n7487) );
  NAND2_X1 U9988 ( .A1(n14362), .A2(n14363), .ZN(n14361) );
  XNOR2_X1 U9989 ( .A(n8412), .B(n12089), .ZN(n8411) );
  OAI22_X1 U9990 ( .A1(n12636), .A2(n12635), .B1(n13307), .B2(n10106), .ZN(
        n12695) );
  INV_X1 U9991 ( .A(n8610), .ZN(n7658) );
  AOI22_X1 U9992 ( .A1(n13955), .A2(n8707), .B1(n8650), .B2(n13969), .ZN(n8633) );
  NAND2_X1 U9993 ( .A1(n12987), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n13013) );
  NOR2_X1 U9994 ( .A1(n7099), .A2(n13004), .ZN(n7098) );
  NAND2_X1 U9995 ( .A1(n7092), .A2(n11229), .ZN(n7091) );
  AOI21_X1 U9996 ( .B1(n11670), .B2(n11668), .A(n11669), .ZN(n11807) );
  NAND2_X1 U9997 ( .A1(n10178), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n10267) );
  NAND2_X1 U9998 ( .A1(n12945), .A2(n12942), .ZN(n12944) );
  OAI21_X1 U9999 ( .B1(n8634), .B2(n8633), .A(n8632), .ZN(n8636) );
  AND2_X1 U10000 ( .A1(n8586), .A2(n7010), .ZN(n8587) );
  NAND2_X1 U10001 ( .A1(n12047), .A2(n9050), .ZN(n11993) );
  NAND2_X1 U10002 ( .A1(n6436), .A2(n11318), .ZN(n12043) );
  NOR2_X2 U10003 ( .A1(n13796), .A2(n13784), .ZN(n13779) );
  NAND2_X2 U10004 ( .A1(n13865), .A2(n6456), .ZN(n13796) );
  NAND2_X2 U10005 ( .A1(n7013), .A2(n13882), .ZN(n13878) );
  NOR2_X2 U10006 ( .A1(n13917), .A2(n14064), .ZN(n7013) );
  NAND2_X1 U10007 ( .A1(n12240), .A2(n12860), .ZN(n12332) );
  AOI21_X1 U10008 ( .B1(n7702), .B2(n7701), .A(n7699), .ZN(n13247) );
  NAND2_X1 U10009 ( .A1(n7720), .A2(n7719), .ZN(n13321) );
  NAND2_X1 U10010 ( .A1(n15572), .A2(n12809), .ZN(n10260) );
  NAND2_X1 U10011 ( .A1(n7350), .A2(n7348), .ZN(n8412) );
  OR2_X1 U10012 ( .A1(n14568), .A2(n14571), .ZN(n14562) );
  AND2_X1 U10013 ( .A1(n14566), .A2(n14565), .ZN(n14567) );
  OAI211_X1 U10014 ( .C1(n8780), .C2(n8775), .A(n8782), .B(n12105), .ZN(n7048)
         );
  AND2_X2 U10015 ( .A1(n8560), .A2(n13705), .ZN(n11823) );
  AND2_X2 U10016 ( .A1(n7886), .A2(n8776), .ZN(n8560) );
  INV_X1 U10017 ( .A(n8358), .ZN(n13600) );
  NAND3_X1 U10018 ( .A1(n8386), .A2(n8384), .A3(n7531), .ZN(n13592) );
  NAND2_X1 U10019 ( .A1(n14787), .A2(n14958), .ZN(n7283) );
  NAND2_X2 U10020 ( .A1(n9593), .A2(n14261), .ZN(n14263) );
  AOI21_X1 U10022 ( .B1(n8646), .B2(n8645), .A(n6596), .ZN(n7025) );
  NAND2_X1 U10023 ( .A1(n7275), .A2(n7276), .ZN(n9068) );
  OAI21_X1 U10024 ( .B1(n8646), .B2(n8645), .A(n8644), .ZN(n7026) );
  NAND2_X1 U10025 ( .A1(n8562), .A2(n13673), .ZN(n8563) );
  NAND2_X1 U10026 ( .A1(n8813), .A2(n8812), .ZN(n7047) );
  AOI22_X1 U10027 ( .A1(n8650), .A2(n8571), .B1(n13671), .B2(n8726), .ZN(n8584) );
  NAND2_X2 U10028 ( .A1(n11823), .A2(n9039), .ZN(n8579) );
  OR2_X1 U10029 ( .A1(n7967), .A2(n10738), .ZN(n7939) );
  XNOR2_X2 U10030 ( .A(n12056), .B(n13671), .ZN(n11249) );
  AOI22_X2 U10031 ( .A1(n9896), .A2(n9895), .B1(n9894), .B2(n11855), .ZN(n9897) );
  NOR2_X1 U10032 ( .A1(n15653), .A2(n15654), .ZN(n9144) );
  AOI21_X1 U10033 ( .B1(n7568), .B2(n7570), .A(n7565), .ZN(n7564) );
  INV_X1 U10034 ( .A(n15232), .ZN(n7043) );
  INV_X1 U10035 ( .A(n12222), .ZN(n7491) );
  OR2_X1 U10036 ( .A1(n8949), .A2(n10452), .ZN(n8834) );
  OR4_X2 U10037 ( .A1(n13199), .A2(n12782), .A3(n13224), .A4(n12781), .ZN(
        n12783) );
  INV_X1 U10038 ( .A(n7578), .ZN(n7577) );
  NAND2_X1 U10039 ( .A1(n7487), .A2(n7486), .ZN(n8829) );
  NOR2_X1 U10040 ( .A1(n13130), .A2(n6500), .ZN(n13137) );
  AOI21_X1 U10041 ( .B1(n7670), .B2(n7835), .A(n7834), .ZN(n13736) );
  OAI21_X1 U10042 ( .B1(n13431), .B2(n15643), .A(n7037), .ZN(P3_U3453) );
  OAI21_X1 U10043 ( .B1(n13431), .B2(n7202), .A(n7039), .ZN(P3_U3485) );
  NAND2_X1 U10044 ( .A1(n7283), .A2(n7280), .ZN(n14789) );
  INV_X1 U10045 ( .A(n13697), .ZN(n13704) );
  XNOR2_X1 U10046 ( .A(n13696), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13697) );
  INV_X1 U10047 ( .A(n7361), .ZN(n7360) );
  NAND2_X1 U10048 ( .A1(n9560), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U10049 ( .A1(n15156), .A2(n15408), .ZN(n7054) );
  NAND3_X1 U10050 ( .A1(n7048), .A2(n7047), .A3(n7810), .ZN(P2_U3328) );
  OAI21_X1 U10051 ( .B1(n8577), .B2(n8578), .A(n8576), .ZN(n7049) );
  NAND2_X1 U10052 ( .A1(n10056), .A2(n10055), .ZN(n10069) );
  NAND2_X2 U10053 ( .A1(n8969), .A2(n15291), .ZN(n8843) );
  NAND2_X1 U10054 ( .A1(n7054), .A2(n6622), .ZN(P1_U3525) );
  NAND2_X1 U10055 ( .A1(n12533), .A2(n12532), .ZN(n15067) );
  INV_X1 U10056 ( .A(n11633), .ZN(n7059) );
  NAND2_X1 U10057 ( .A1(n7060), .A2(n11634), .ZN(n11680) );
  NAND2_X1 U10058 ( .A1(n11633), .A2(n11632), .ZN(n7060) );
  NAND2_X1 U10059 ( .A1(n14917), .A2(n6496), .ZN(n7061) );
  NAND2_X1 U10060 ( .A1(n7061), .A2(n7062), .ZN(n14879) );
  NAND2_X1 U10061 ( .A1(n7077), .A2(n7075), .ZN(n12440) );
  NAND3_X1 U10062 ( .A1(n12179), .A2(n7734), .A3(n15046), .ZN(n7077) );
  OAI21_X2 U10063 ( .B1(n14996), .B2(n6562), .A(n7741), .ZN(n14961) );
  INV_X1 U10064 ( .A(n7611), .ZN(n15323) );
  NAND2_X1 U10065 ( .A1(n9132), .A2(n9135), .ZN(n9096) );
  INV_X1 U10066 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7080) );
  OAI21_X2 U10067 ( .B1(n15271), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6487), .ZN(
        n7082) );
  NAND2_X1 U10068 ( .A1(n15286), .A2(n15287), .ZN(n9172) );
  INV_X1 U10069 ( .A(n11216), .ZN(n7092) );
  NAND3_X1 U10070 ( .A1(n7093), .A2(n6595), .A3(n7091), .ZN(n11670) );
  INV_X1 U10071 ( .A(n11877), .ZN(n11878) );
  NAND2_X1 U10072 ( .A1(n11877), .A2(n7097), .ZN(n7505) );
  AND2_X1 U10073 ( .A1(n10949), .A2(n11071), .ZN(n10950) );
  NAND2_X1 U10074 ( .A1(n10948), .A2(n11056), .ZN(n11071) );
  NAND2_X1 U10075 ( .A1(n12877), .A2(n7108), .ZN(n7113) );
  NAND2_X1 U10076 ( .A1(n7113), .A2(n7112), .ZN(n12886) );
  AOI21_X1 U10077 ( .B1(n7119), .B2(n7114), .A(n6617), .ZN(n7112) );
  OAI211_X1 U10078 ( .C1(n7130), .C2(n7125), .A(n12831), .B(n7124), .ZN(n12836) );
  NAND2_X1 U10079 ( .A1(n12823), .A2(n12824), .ZN(n7130) );
  INV_X1 U10080 ( .A(n12817), .ZN(n7131) );
  INV_X1 U10081 ( .A(n7134), .ZN(n7133) );
  NAND3_X1 U10082 ( .A1(n7136), .A2(n7135), .A3(n12919), .ZN(n7134) );
  INV_X1 U10083 ( .A(n7139), .ZN(n12925) );
  NOR2_X1 U10084 ( .A1(n13173), .A2(n12935), .ZN(n7151) );
  NAND2_X1 U10085 ( .A1(n9725), .A2(n13507), .ZN(n9723) );
  NAND2_X1 U10086 ( .A1(n10097), .A2(n6619), .ZN(n10147) );
  NAND2_X1 U10087 ( .A1(n9848), .A2(n7162), .ZN(n9928) );
  NAND3_X1 U10088 ( .A1(n9823), .A2(n11499), .A3(n9802), .ZN(n9880) );
  INV_X1 U10089 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14790) );
  AND2_X4 U10090 ( .A1(n7168), .A2(n7169), .ZN(n7955) );
  NAND2_X1 U10091 ( .A1(n13852), .A2(n7176), .ZN(n7175) );
  NAND2_X1 U10092 ( .A1(n7181), .A2(n7180), .ZN(P2_U3526) );
  NAND2_X1 U10093 ( .A1(n8122), .A2(n6577), .ZN(n7183) );
  OAI21_X1 U10094 ( .B1(n7798), .B2(n6509), .A(n10331), .ZN(n7190) );
  NAND2_X1 U10095 ( .A1(n13323), .A2(n13324), .ZN(n10333) );
  INV_X1 U10096 ( .A(n11779), .ZN(n7196) );
  NAND3_X1 U10097 ( .A1(n7194), .A2(n7192), .A3(n6594), .ZN(n7197) );
  NAND3_X1 U10098 ( .A1(n7196), .A2(n7801), .A3(n7195), .ZN(n7194) );
  NAND2_X1 U10099 ( .A1(n7198), .A2(n15652), .ZN(n7199) );
  NAND3_X1 U10100 ( .A1(n12558), .A2(n7201), .A3(n7199), .ZN(P3_U3488) );
  NAND3_X1 U10101 ( .A1(n12555), .A2(n12554), .A3(n7831), .ZN(n13167) );
  OAI21_X1 U10102 ( .B1(n14442), .B2(n7221), .A(n14471), .ZN(n7220) );
  AND2_X1 U10103 ( .A1(n14471), .A2(n14466), .ZN(n14999) );
  NAND2_X1 U10104 ( .A1(n14985), .A2(n14999), .ZN(n7624) );
  NAND2_X1 U10105 ( .A1(n12409), .A2(n12408), .ZN(n7226) );
  NAND3_X1 U10106 ( .A1(n8885), .A2(n7238), .A3(n8864), .ZN(n7237) );
  XNOR2_X2 U10107 ( .A(n7243), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U10108 ( .A1(n14847), .A2(n7250), .ZN(n7248) );
  AOI21_X1 U10109 ( .B1(n14847), .B2(n12429), .A(n6601), .ZN(n12503) );
  NAND2_X1 U10110 ( .A1(n13841), .A2(n7268), .ZN(n7266) );
  NAND2_X1 U10111 ( .A1(n13948), .A2(n7277), .ZN(n7275) );
  NAND2_X1 U10112 ( .A1(n14731), .A2(n7286), .ZN(n7285) );
  MUX2_X1 U10113 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n14655), .S(n14654), .Z(
        n7294) );
  XNOR2_X1 U10114 ( .A(n11873), .B(n11875), .ZN(n11876) );
  NAND2_X1 U10115 ( .A1(n10943), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7326) );
  NAND2_X1 U10116 ( .A1(n7327), .A2(n7326), .ZN(n11025) );
  NAND2_X1 U10117 ( .A1(n7892), .A2(n7330), .ZN(n14187) );
  NAND2_X1 U10118 ( .A1(n8303), .A2(n7352), .ZN(n7350) );
  NAND2_X1 U10119 ( .A1(n14263), .A2(n7365), .ZN(n7357) );
  NAND2_X1 U10120 ( .A1(n14263), .A2(n7363), .ZN(n7358) );
  NAND2_X1 U10121 ( .A1(n14263), .A2(n9594), .ZN(n14362) );
  OAI211_X1 U10122 ( .C1(n14263), .C2(n7360), .A(n7359), .B(n7358), .ZN(n10382) );
  NAND2_X1 U10123 ( .A1(n14352), .A2(n7372), .ZN(n7370) );
  AND2_X1 U10124 ( .A1(n9499), .A2(n14311), .ZN(n7372) );
  AND2_X1 U10125 ( .A1(n10397), .A2(n10396), .ZN(n11516) );
  NAND2_X2 U10126 ( .A1(n10393), .A2(n14387), .ZN(n9604) );
  NAND2_X1 U10127 ( .A1(n14339), .A2(n6588), .ZN(n14252) );
  NAND2_X1 U10128 ( .A1(n13686), .A2(n7381), .ZN(n7380) );
  INV_X1 U10129 ( .A(n13699), .ZN(n7381) );
  NAND3_X1 U10130 ( .A1(n7937), .A2(n7395), .A3(n7393), .ZN(n10598) );
  NAND3_X1 U10131 ( .A1(n7843), .A2(n7842), .A3(n7874), .ZN(n7853) );
  CLKBUF_X1 U10132 ( .A(n13973), .Z(n7398) );
  INV_X1 U10133 ( .A(n13973), .ZN(n7400) );
  NAND2_X1 U10134 ( .A1(n7404), .A2(n7402), .ZN(P2_U3498) );
  NOR2_X1 U10135 ( .A1(n15561), .A2(n8695), .ZN(n7403) );
  NAND2_X1 U10136 ( .A1(n14115), .A2(n15561), .ZN(n7404) );
  NAND3_X1 U10137 ( .A1(n6431), .A2(n7405), .A3(n7406), .ZN(n13711) );
  NAND4_X1 U10138 ( .A1(n7412), .A2(n7411), .A3(n9842), .A4(n9907), .ZN(n9695)
         );
  NAND3_X1 U10139 ( .A1(n8985), .A2(n7416), .A3(n7414), .ZN(n14575) );
  INV_X1 U10140 ( .A(n14531), .ZN(n7418) );
  NOR2_X2 U10141 ( .A1(n12701), .A2(n7419), .ZN(n7423) );
  NOR2_X2 U10142 ( .A1(n12702), .A2(n12966), .ZN(n12701) );
  NOR2_X2 U10143 ( .A1(n10172), .A2(n7423), .ZN(n12628) );
  NAND2_X1 U10144 ( .A1(n14397), .A2(n14584), .ZN(n7436) );
  OAI21_X1 U10145 ( .B1(n14407), .B2(n14406), .A(n14405), .ZN(n14409) );
  NAND2_X1 U10146 ( .A1(n14455), .A2(n14456), .ZN(n7437) );
  NAND2_X1 U10147 ( .A1(n14458), .A2(n14457), .ZN(n7438) );
  NAND2_X1 U10148 ( .A1(n9743), .A2(n9744), .ZN(n7455) );
  NAND2_X1 U10149 ( .A1(n11043), .A2(n7455), .ZN(n11095) );
  NAND2_X1 U10150 ( .A1(n14382), .A2(n14383), .ZN(n14543) );
  NAND3_X1 U10151 ( .A1(n7461), .A2(n9897), .A3(n7463), .ZN(n7459) );
  NAND2_X1 U10152 ( .A1(n11559), .A2(n9889), .ZN(n7464) );
  NAND2_X1 U10153 ( .A1(n7477), .A2(n7475), .ZN(n14421) );
  NAND2_X1 U10154 ( .A1(n14415), .A2(n7478), .ZN(n7477) );
  NAND2_X1 U10155 ( .A1(n7481), .A2(n7480), .ZN(n9713) );
  INV_X1 U10156 ( .A(n7484), .ZN(n14935) );
  NAND2_X1 U10157 ( .A1(n14806), .A2(n7488), .ZN(n14795) );
  NAND3_X1 U10158 ( .A1(n7491), .A2(n15259), .A3(n7490), .ZN(n15232) );
  NAND2_X1 U10159 ( .A1(n11809), .A2(n11884), .ZN(n7506) );
  NAND2_X1 U10160 ( .A1(n7507), .A2(n7506), .ZN(n11880) );
  NOR2_X1 U10161 ( .A1(n7508), .A2(n11877), .ZN(n11810) );
  NOR2_X1 U10162 ( .A1(n11877), .A2(n12251), .ZN(n7507) );
  NAND2_X1 U10163 ( .A1(n7509), .A2(n7510), .ZN(n7512) );
  NAND2_X1 U10164 ( .A1(n6583), .A2(n11019), .ZN(n7509) );
  NAND3_X1 U10165 ( .A1(n11019), .A2(n10944), .A3(n10924), .ZN(n7513) );
  NAND2_X1 U10166 ( .A1(n7520), .A2(n7522), .ZN(n13035) );
  INV_X1 U10167 ( .A(n11472), .ZN(n11695) );
  NAND3_X1 U10168 ( .A1(n7533), .A2(n8374), .A3(n7532), .ZN(n7531) );
  NAND2_X1 U10169 ( .A1(n8358), .A2(n6573), .ZN(n7533) );
  AND2_X1 U10170 ( .A1(n13613), .A2(n13612), .ZN(n13609) );
  INV_X1 U10171 ( .A(n8385), .ZN(n7534) );
  NAND2_X1 U10172 ( .A1(n11203), .A2(n7538), .ZN(n7535) );
  INV_X1 U10173 ( .A(n13584), .ZN(n7546) );
  OR2_X1 U10174 ( .A1(n7942), .A2(n7941), .ZN(n7558) );
  NAND2_X1 U10175 ( .A1(n13565), .A2(n13564), .ZN(n13563) );
  NAND2_X1 U10176 ( .A1(n10088), .A2(n10087), .ZN(n10090) );
  NAND2_X1 U10177 ( .A1(n10069), .A2(n10068), .ZN(n7563) );
  NAND2_X1 U10178 ( .A1(n10018), .A2(n7568), .ZN(n7566) );
  NAND2_X1 U10179 ( .A1(n9760), .A2(n7573), .ZN(n7576) );
  NAND2_X1 U10180 ( .A1(n9794), .A2(n7589), .ZN(n7587) );
  NAND2_X1 U10181 ( .A1(n9140), .A2(n7596), .ZN(n7595) );
  NAND2_X1 U10182 ( .A1(n9140), .A2(n9141), .ZN(n7600) );
  NAND2_X1 U10183 ( .A1(n7600), .A2(n9103), .ZN(n9104) );
  NAND2_X2 U10184 ( .A1(n8829), .A2(n8962), .ZN(n15291) );
  NAND2_X1 U10185 ( .A1(n11926), .A2(n7613), .ZN(n7612) );
  AOI21_X2 U10186 ( .B1(n7634), .B2(n7637), .A(n7632), .ZN(n7631) );
  NAND2_X1 U10187 ( .A1(n7652), .A2(n7649), .ZN(n7651) );
  INV_X1 U10188 ( .A(n11483), .ZN(n7650) );
  NAND3_X1 U10189 ( .A1(n7661), .A2(n7659), .A3(n7832), .ZN(n8962) );
  INV_X1 U10190 ( .A(n13757), .ZN(n7670) );
  OAI21_X2 U10191 ( .B1(n13757), .B2(n6521), .A(n7665), .ZN(n14007) );
  NAND2_X1 U10192 ( .A1(n11974), .A2(n7672), .ZN(n7671) );
  NAND4_X1 U10193 ( .A1(n9686), .A2(n10798), .A3(n9684), .A4(n9685), .ZN(n9691) );
  NOR2_X2 U10194 ( .A1(n7684), .A2(n7683), .ZN(n7691) );
  NAND4_X1 U10195 ( .A1(n7686), .A2(n7685), .A3(n9685), .A4(n9681), .ZN(n7684)
         );
  NOR2_X1 U10196 ( .A1(n9694), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7689) );
  INV_X1 U10197 ( .A(n9690), .ZN(n7690) );
  NAND3_X1 U10198 ( .A1(n6497), .A2(n7691), .A3(n7687), .ZN(n9719) );
  INV_X1 U10199 ( .A(n9683), .ZN(n9872) );
  NAND2_X1 U10200 ( .A1(n11730), .A2(n7696), .ZN(n7692) );
  INV_X1 U10201 ( .A(n13286), .ZN(n7702) );
  NAND2_X1 U10202 ( .A1(n12378), .A2(n7721), .ZN(n7720) );
  NAND2_X1 U10203 ( .A1(n10911), .A2(n7733), .ZN(n9877) );
  NAND2_X1 U10204 ( .A1(n7740), .A2(n7739), .ZN(n15014) );
  NAND2_X1 U10205 ( .A1(n15018), .A2(n15022), .ZN(n7740) );
  NAND2_X1 U10206 ( .A1(n8828), .A2(n7744), .ZN(n15172) );
  XNOR2_X2 U10207 ( .A(n14815), .B(n14814), .ZN(n15090) );
  INV_X1 U10208 ( .A(n12277), .ZN(n7757) );
  NAND2_X1 U10209 ( .A1(n7920), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U10210 ( .A1(n7920), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U10211 ( .A1(n7920), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8156) );
  NAND2_X1 U10212 ( .A1(n7920), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U10213 ( .A1(n7920), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10214 ( .A1(n7920), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U10215 ( .A1(n7920), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10216 ( .A1(n6967), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10217 ( .A1(n7920), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U10218 ( .A1(n6967), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8547) );
  NOR2_X1 U10219 ( .A1(n7019), .A2(n7769), .ZN(n7768) );
  NAND2_X1 U10220 ( .A1(n7772), .A2(n7770), .ZN(P2_U3491) );
  OR2_X1 U10221 ( .A1(n15561), .A2(n7771), .ZN(n7770) );
  NAND2_X1 U10222 ( .A1(n13793), .A2(n13792), .ZN(n7777) );
  NAND2_X1 U10223 ( .A1(n9055), .A2(n9054), .ZN(n11975) );
  NOR2_X1 U10224 ( .A1(n9057), .A2(n7782), .ZN(n7781) );
  INV_X1 U10225 ( .A(n9054), .ZN(n7782) );
  NAND2_X1 U10226 ( .A1(n11958), .A2(n12162), .ZN(n9058) );
  INV_X1 U10227 ( .A(n13856), .ZN(n7788) );
  NAND2_X2 U10228 ( .A1(n7783), .A2(n7784), .ZN(n13841) );
  NAND2_X1 U10229 ( .A1(n13825), .A2(n7789), .ZN(n13809) );
  INV_X2 U10230 ( .A(n9828), .ZN(n9854) );
  NAND2_X2 U10231 ( .A1(n9728), .A2(n7790), .ZN(n9828) );
  NAND3_X1 U10232 ( .A1(n7790), .A2(P3_REG1_REG_1__SCAN_IN), .A3(n9728), .ZN(
        n9729) );
  OAI21_X1 U10233 ( .B1(n11797), .B2(n10325), .A(n7796), .ZN(n12334) );
  INV_X1 U10234 ( .A(n7793), .ZN(n10328) );
  AOI21_X1 U10235 ( .B1(n11797), .B2(n7796), .A(n7794), .ZN(n7793) );
  NAND2_X1 U10236 ( .A1(n12381), .A2(n10329), .ZN(n7799) );
  NAND2_X1 U10237 ( .A1(n9734), .A2(n7808), .ZN(n9722) );
  NAND2_X1 U10238 ( .A1(n9734), .A2(n7807), .ZN(n7809) );
  CLKBUF_X1 U10239 ( .A(n12299), .Z(n13972) );
  NAND2_X1 U10240 ( .A1(n12575), .A2(n12574), .ZN(n12576) );
  NAND2_X1 U10241 ( .A1(n14115), .A2(n15564), .ZN(n12575) );
  OR2_X1 U10242 ( .A1(n13170), .A2(n13495), .ZN(n12561) );
  CLKBUF_X1 U10243 ( .A(n14924), .Z(n14937) );
  NAND2_X1 U10244 ( .A1(n15063), .A2(n15408), .ZN(n9003) );
  INV_X1 U10245 ( .A(n6431), .ZN(n13726) );
  NAND2_X1 U10246 ( .A1(n14794), .A2(n8972), .ZN(n15063) );
  OR2_X1 U10247 ( .A1(n14652), .A2(n11629), .ZN(n11627) );
  INV_X1 U10248 ( .A(n12605), .ZN(n12604) );
  CLKBUF_X1 U10249 ( .A(n11958), .Z(n12164) );
  INV_X4 U10250 ( .A(n10301), .ZN(n12269) );
  AND3_X1 U10251 ( .A1(n15091), .A2(n15395), .A3(n15092), .ZN(n15096) );
  NAND2_X1 U10252 ( .A1(n12602), .A2(n12601), .ZN(n12605) );
  OAI21_X1 U10253 ( .B1(n12462), .B2(n6554), .A(n12602), .ZN(n12463) );
  OR2_X1 U10254 ( .A1(n11380), .A2(n15343), .ZN(n14391) );
  NAND2_X1 U10255 ( .A1(n13178), .A2(n6579), .ZN(n12554) );
  NAND2_X1 U10256 ( .A1(n13172), .A2(n13173), .ZN(n13178) );
  NAND2_X1 U10257 ( .A1(n9217), .A2(n14101), .ZN(n9095) );
  NAND2_X1 U10258 ( .A1(n12807), .A2(n12806), .ZN(n11040) );
  AOI21_X1 U10259 ( .B1(n9190), .B2(n13990), .A(n9189), .ZN(n9195) );
  NAND2_X1 U10260 ( .A1(n7873), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7869) );
  OR2_X1 U10261 ( .A1(n7019), .A2(n7881), .ZN(n7882) );
  OAI21_X2 U10262 ( .B1(n14934), .B2(n12453), .A(n12452), .ZN(n14917) );
  OR2_X1 U10263 ( .A1(n9214), .A2(n9213), .ZN(n15559) );
  AND2_X1 U10264 ( .A1(n8818), .A2(n8817), .ZN(n7810) );
  INV_X1 U10265 ( .A(n13806), .ZN(n9036) );
  NAND2_X1 U10266 ( .A1(n13592), .A2(n13591), .ZN(n13590) );
  NOR2_X1 U10267 ( .A1(n14937), .A2(n14936), .ZN(n7815) );
  AND2_X1 U10268 ( .A1(n10085), .A2(n12967), .ZN(n7816) );
  INV_X1 U10269 ( .A(n15601), .ZN(n10349) );
  NOR2_X1 U10270 ( .A1(n14240), .A2(n14239), .ZN(n7817) );
  OR2_X1 U10271 ( .A1(n8336), .A2(SI_21_), .ZN(n7818) );
  OR2_X1 U10272 ( .A1(n8774), .A2(n11614), .ZN(n7819) );
  NAND2_X1 U10273 ( .A1(n11375), .A2(n14399), .ZN(n11376) );
  AND3_X1 U10274 ( .A1(n9654), .A2(n9653), .A3(n14370), .ZN(n7821) );
  AND2_X1 U10275 ( .A1(n8451), .A2(n8450), .ZN(n7822) );
  AND2_X1 U10276 ( .A1(n10190), .A2(n10195), .ZN(n7823) );
  AND2_X1 U10277 ( .A1(n12548), .A2(n10349), .ZN(n7824) );
  NAND2_X2 U10278 ( .A1(n12506), .A2(n15055), .ZN(n15049) );
  INV_X1 U10279 ( .A(n14242), .ZN(n14291) );
  AND2_X1 U10280 ( .A1(n9830), .A2(n9829), .ZN(n7825) );
  INV_X1 U10281 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n9097) );
  INV_X1 U10282 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9149) );
  XNOR2_X1 U10283 ( .A(n11380), .B(n15343), .ZN(n11259) );
  INV_X1 U10284 ( .A(n9066), .ZN(n13928) );
  OR4_X1 U10285 ( .A1(n14011), .A2(n13951), .A3(n13723), .A4(n13720), .ZN(
        n7826) );
  NAND4_X1 U10286 ( .A1(n13719), .A2(n13718), .A3(n13971), .A4(n14011), .ZN(
        n7827) );
  AND2_X1 U10287 ( .A1(n10121), .A2(n13294), .ZN(n7829) );
  AND2_X1 U10288 ( .A1(n12151), .A2(n12235), .ZN(n7830) );
  NOR2_X1 U10289 ( .A1(n12553), .A2(n12552), .ZN(n7831) );
  INV_X1 U10290 ( .A(n12934), .ZN(n10346) );
  INV_X1 U10291 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13502) );
  INV_X1 U10292 ( .A(n12105), .ZN(n8781) );
  AND2_X1 U10293 ( .A1(n14026), .A2(n13773), .ZN(n7834) );
  OR2_X1 U10294 ( .A1(n14026), .A2(n13773), .ZN(n7835) );
  OR2_X1 U10295 ( .A1(n9350), .A2(n9349), .ZN(n7836) );
  OR2_X1 U10296 ( .A1(n8334), .A2(SI_20_), .ZN(n7837) );
  OR2_X1 U10297 ( .A1(n14140), .A2(n13656), .ZN(n7838) );
  NAND2_X1 U10298 ( .A1(n12979), .A2(n11498), .ZN(n7839) );
  AND2_X1 U10299 ( .A1(n8650), .A2(n11353), .ZN(n8562) );
  AOI22_X1 U10300 ( .A1(n13669), .A2(n8650), .B1(n12038), .B2(n8726), .ZN(
        n8594) );
  OAI21_X1 U10301 ( .B1(n8594), .B2(n8593), .A(n8592), .ZN(n8595) );
  INV_X1 U10302 ( .A(n8606), .ZN(n8607) );
  INV_X1 U10303 ( .A(n8615), .ZN(n8616) );
  OAI22_X1 U10304 ( .A1(n13941), .A2(n8650), .B1(n13641), .B2(n8707), .ZN(
        n8641) );
  AOI22_X1 U10305 ( .A1(n13920), .A2(n8707), .B1(n8770), .B2(n13893), .ZN(
        n8645) );
  OAI22_X1 U10306 ( .A1(n13901), .A2(n8726), .B1(n13549), .B2(n8770), .ZN(
        n8648) );
  OAI22_X1 U10307 ( .A1(n13901), .A2(n8770), .B1(n13549), .B2(n8707), .ZN(
        n8647) );
  INV_X1 U10308 ( .A(n10324), .ZN(n10325) );
  OR3_X1 U10309 ( .A1(n8757), .A2(n8756), .A3(n8755), .ZN(n8758) );
  INV_X1 U10310 ( .A(n14203), .ZN(n9559) );
  NAND2_X1 U10311 ( .A1(n14603), .A2(n14640), .ZN(n12424) );
  NAND2_X1 U10312 ( .A1(n9072), .A2(n13789), .ZN(n9073) );
  NAND2_X1 U10313 ( .A1(n9303), .A2(n11519), .ZN(n9287) );
  NOR2_X1 U10314 ( .A1(n8187), .A2(n10675), .ZN(n8188) );
  AND2_X1 U10315 ( .A1(n12678), .A2(n13337), .ZN(n10049) );
  INV_X1 U10316 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U10317 ( .A1(n15583), .A2(n11047), .ZN(n12806) );
  INV_X1 U10318 ( .A(n10137), .ZN(n10138) );
  NOR2_X1 U10319 ( .A1(n9074), .A2(n9073), .ZN(n9075) );
  AOI22_X1 U10320 ( .A1(n11380), .A2(n9648), .B1(n11370), .B2(n9644), .ZN(
        n9246) );
  INV_X1 U10321 ( .A(n9561), .ZN(n9560) );
  AND2_X1 U10322 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_REG3_REG_11__SCAN_IN), 
        .ZN(n9354) );
  NAND2_X1 U10323 ( .A1(n9658), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9248) );
  NAND2_X1 U10324 ( .A1(n8231), .A2(n10682), .ZN(n8256) );
  NAND2_X1 U10325 ( .A1(n8141), .A2(n10626), .ZN(n8161) );
  INV_X1 U10326 ( .A(n8046), .ZN(n8035) );
  NOR2_X1 U10327 ( .A1(n12480), .A2(n12963), .ZN(n12481) );
  INV_X1 U10328 ( .A(n11406), .ZN(n9812) );
  OR2_X1 U10329 ( .A1(n13091), .A2(n13084), .ZN(n13085) );
  INV_X1 U10330 ( .A(n13523), .ZN(n9710) );
  OR2_X1 U10331 ( .A1(n10637), .A2(n7940), .ZN(n7894) );
  NAND2_X1 U10332 ( .A1(n10642), .A2(n10637), .ZN(n11355) );
  INV_X1 U10333 ( .A(n14192), .ZN(n9409) );
  OR2_X1 U10334 ( .A1(n14277), .A2(n14278), .ZN(n9441) );
  OR2_X1 U10335 ( .A1(n14239), .A2(n9557), .ZN(n14199) );
  INV_X1 U10336 ( .A(n12527), .ZN(n12528) );
  NAND2_X1 U10337 ( .A1(n8411), .A2(n8410), .ZN(n8414) );
  NAND2_X1 U10338 ( .A1(n9159), .A2(n9160), .ZN(n9118) );
  OR2_X1 U10339 ( .A1(n9822), .A2(n9801), .ZN(n9808) );
  NAND2_X1 U10340 ( .A1(n12547), .A2(n7824), .ZN(n12555) );
  AND2_X1 U10341 ( .A1(n12930), .A2(n10356), .ZN(n15597) );
  INV_X1 U10342 ( .A(n12768), .ZN(n12824) );
  AND2_X1 U10343 ( .A1(n10348), .A2(n10347), .ZN(n15601) );
  INV_X1 U10344 ( .A(n12957), .ZN(n12801) );
  INV_X1 U10345 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11755) );
  OR2_X1 U10346 ( .A1(n13616), .A2(n13930), .ZN(n13623) );
  INV_X1 U10347 ( .A(n13568), .ZN(n13634) );
  INV_X1 U10348 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10669) );
  AND2_X1 U10349 ( .A1(n11915), .A2(n8776), .ZN(n10491) );
  MUX2_X1 U10350 ( .A(n6686), .B(n14187), .S(n10492), .Z(n11353) );
  OR2_X1 U10351 ( .A1(n14013), .A2(n14012), .ZN(n14014) );
  INV_X1 U10352 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n11952) );
  INV_X1 U10353 ( .A(n14250), .ZN(n9379) );
  AND2_X1 U10354 ( .A1(n9442), .A2(n9441), .ZN(n9443) );
  AND2_X1 U10355 ( .A1(n14260), .A2(n9577), .ZN(n14298) );
  OR2_X1 U10356 ( .A1(n14564), .A2(n14563), .ZN(n14565) );
  INV_X1 U10357 ( .A(n9657), .ZN(n12518) );
  INV_X1 U10358 ( .A(n12508), .ZN(n9659) );
  NAND2_X1 U10359 ( .A1(n9638), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9241) );
  INV_X1 U10360 ( .A(n14987), .ZN(n14956) );
  NAND2_X1 U10361 ( .A1(n11266), .A2(n11265), .ZN(n15055) );
  NAND2_X1 U10362 ( .A1(n8344), .A2(n8343), .ZN(n8346) );
  NAND2_X1 U10363 ( .A1(n6550), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8873) );
  INV_X1 U10364 ( .A(n12743), .ZN(n12735) );
  INV_X1 U10365 ( .A(n11540), .ZN(n12952) );
  INV_X1 U10366 ( .A(n13151), .ZN(n13112) );
  INV_X1 U10367 ( .A(n13340), .ZN(n13347) );
  OR2_X1 U10368 ( .A1(n10229), .A2(n15603), .ZN(n15577) );
  AND3_X1 U10369 ( .A1(n10909), .A2(n10371), .A3(n10370), .ZN(n11416) );
  AND2_X1 U10370 ( .A1(n15652), .A2(n15623), .ZN(n13416) );
  INV_X1 U10371 ( .A(n12775), .ZN(n12335) );
  AND3_X1 U10372 ( .A1(n13499), .A2(n13497), .A3(n10370), .ZN(n10365) );
  AND2_X1 U10373 ( .A1(n9957), .A2(n9943), .ZN(n9955) );
  INV_X1 U10374 ( .A(n11984), .ZN(n14106) );
  AND2_X1 U10375 ( .A1(n8383), .A2(n8382), .ZN(n13843) );
  INV_X1 U10376 ( .A(n15421), .ZN(n15508) );
  AOI21_X1 U10377 ( .B1(n9199), .B2(n13995), .A(n9198), .ZN(n9200) );
  NAND2_X1 U10378 ( .A1(n15533), .A2(n8538), .ZN(n13956) );
  INV_X1 U10379 ( .A(n13951), .ZN(n13971) );
  INV_X1 U10380 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9093) );
  INV_X1 U10381 ( .A(n15536), .ZN(n15553) );
  AND2_X1 U10382 ( .A1(n8511), .A2(n8515), .ZN(n15524) );
  AND2_X1 U10383 ( .A1(n10496), .A2(n10490), .ZN(n8543) );
  OAI21_X1 U10384 ( .B1(n12439), .B2(n14380), .A(n10387), .ZN(n10388) );
  NAND2_X1 U10385 ( .A1(n9674), .A2(n9673), .ZN(n9675) );
  INV_X1 U10386 ( .A(n14353), .ZN(n14242) );
  AOI22_X1 U10387 ( .A1(n15223), .A2(n14638), .B1(n14636), .B2(n15222), .ZN(
        n12591) );
  AND2_X1 U10388 ( .A1(n10458), .A2(n10608), .ZN(n15223) );
  INV_X1 U10389 ( .A(n8971), .ZN(n8972) );
  NAND2_X1 U10390 ( .A1(n9001), .A2(n10463), .ZN(n11262) );
  OR4_X1 U10391 ( .A1(n15393), .A2(n15392), .A3(n15391), .A4(n15390), .ZN(
        n15394) );
  INV_X1 U10392 ( .A(n11262), .ZN(n9665) );
  NAND2_X1 U10393 ( .A1(n8981), .A2(n8980), .ZN(n10460) );
  INV_X1 U10394 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n11425) );
  AND2_X1 U10395 ( .A1(n10956), .A2(n10955), .ZN(n15570) );
  INV_X1 U10396 ( .A(n12747), .ZN(n12662) );
  INV_X1 U10397 ( .A(n12720), .ZN(n12744) );
  AND2_X1 U10398 ( .A1(n12272), .A2(n12097), .ZN(n13176) );
  INV_X1 U10399 ( .A(n13227), .ZN(n13251) );
  INV_X1 U10400 ( .A(n13354), .ZN(n12971) );
  AND2_X1 U10401 ( .A1(n11503), .A2(n11773), .ZN(n13363) );
  OR2_X1 U10402 ( .A1(n15610), .A2(n15571), .ZN(n11773) );
  OR2_X1 U10403 ( .A1(n13170), .A2(n13418), .ZN(n12558) );
  NAND2_X1 U10404 ( .A1(n13372), .A2(n15652), .ZN(n13418) );
  INV_X1 U10405 ( .A(n13158), .ZN(n13424) );
  NAND2_X1 U10406 ( .A1(n9948), .A2(n9947), .ZN(n12252) );
  NAND2_X1 U10407 ( .A1(n15645), .A2(n13372), .ZN(n13495) );
  AOI21_X2 U10408 ( .B1(n10366), .B2(n10365), .A(n10364), .ZN(n15643) );
  INV_X1 U10409 ( .A(n9210), .ZN(n9211) );
  INV_X1 U10410 ( .A(n13647), .ZN(n13620) );
  INV_X1 U10411 ( .A(n13641), .ZN(n13658) );
  INV_X1 U10412 ( .A(n11754), .ZN(n13664) );
  OAI21_X1 U10413 ( .B1(n9201), .B2(n13983), .A(n9200), .ZN(n9202) );
  OR2_X1 U10414 ( .A1(n14101), .A2(n9093), .ZN(n9094) );
  INV_X1 U10415 ( .A(n15567), .ZN(n14101) );
  INV_X1 U10416 ( .A(n15567), .ZN(n15564) );
  INV_X1 U10417 ( .A(n13920), .ZN(n14146) );
  INV_X1 U10418 ( .A(n15526), .ZN(n15527) );
  AND2_X1 U10419 ( .A1(n8543), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15533) );
  INV_X1 U10420 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10679) );
  INV_X1 U10421 ( .A(n10388), .ZN(n10389) );
  OR2_X1 U10422 ( .A1(n14603), .A2(n15363), .ZN(n15093) );
  INV_X1 U10423 ( .A(n15111), .ZN(n14878) );
  INV_X1 U10424 ( .A(n14370), .ZN(n14359) );
  OR2_X1 U10425 ( .A1(n14308), .A2(n15363), .ZN(n14380) );
  AND2_X1 U10426 ( .A1(n15231), .A2(n11529), .ZN(n14952) );
  INV_X1 U10427 ( .A(n14865), .ZN(n15062) );
  OR2_X1 U10428 ( .A1(n10718), .A2(n11262), .ZN(n15418) );
  OR2_X1 U10429 ( .A1(n10718), .A2(n9665), .ZN(n15406) );
  AND2_X1 U10430 ( .A1(n10457), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10464) );
  INV_X1 U10431 ( .A(n9219), .ZN(n14544) );
  INV_X1 U10432 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11303) );
  INV_X1 U10433 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10489) );
  XNOR2_X1 U10434 ( .A(n9134), .B(n9133), .ZN(n15664) );
  NAND2_X1 U10435 ( .A1(n10255), .A2(n10254), .ZN(P3_U3169) );
  INV_X1 U10436 ( .A(n14653), .ZN(P1_U4016) );
  NAND2_X1 U10437 ( .A1(n9003), .A2(n9002), .ZN(P1_U3527) );
  NOR2_X1 U10438 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n7841) );
  NOR2_X1 U10439 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n7846) );
  NOR2_X1 U10440 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n7845) );
  INV_X1 U10441 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7844) );
  NAND4_X1 U10442 ( .A1(n7846), .A2(n7845), .A3(n7844), .A4(n8516), .ZN(n7849)
         );
  INV_X1 U10443 ( .A(n7853), .ZN(n7848) );
  NOR2_X1 U10444 ( .A1(n7848), .A2(n7847), .ZN(n7852) );
  INV_X1 U10445 ( .A(n7891), .ZN(n7857) );
  AND2_X1 U10446 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U10447 ( .A1(n7859), .A2(n7858), .ZN(n8837) );
  INV_X1 U10448 ( .A(SI_1_), .ZN(n10413) );
  XNOR2_X1 U10449 ( .A(n7934), .B(n10413), .ZN(n7860) );
  INV_X1 U10450 ( .A(n10492), .ZN(n7956) );
  NAND2_X1 U10451 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n7861) );
  MUX2_X1 U10452 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7861), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7862) );
  INV_X1 U10453 ( .A(n15427), .ZN(n10508) );
  NAND2_X1 U10454 ( .A1(n7956), .A2(n10508), .ZN(n7863) );
  INV_X1 U10455 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n10742) );
  XNOR2_X1 U10456 ( .A(n7868), .B(n10742), .ZN(n7886) );
  OR2_X2 U10457 ( .A1(n7873), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n8493) );
  INV_X1 U10458 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10459 ( .A1(n7871), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7872) );
  INV_X1 U10460 ( .A(n8560), .ZN(n8779) );
  XNOR2_X1 U10461 ( .A(n8567), .B(n7940), .ZN(n7895) );
  INV_X1 U10462 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7876) );
  XNOR2_X2 U10463 ( .A(n7878), .B(P2_IR_REG_29__SCAN_IN), .ZN(n7879) );
  NAND2_X1 U10464 ( .A1(n7979), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7885) );
  INV_X1 U10465 ( .A(n12404), .ZN(n7880) );
  INV_X1 U10466 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10649) );
  INV_X1 U10467 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n13989) );
  INV_X1 U10468 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7881) );
  INV_X1 U10469 ( .A(n8776), .ZN(n11770) );
  XNOR2_X1 U10470 ( .A(n7895), .B(n7897), .ZN(n10645) );
  INV_X1 U10471 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U10472 ( .A1(n13673), .A2(n13974), .ZN(n7893) );
  NAND2_X1 U10473 ( .A1(n7891), .A2(n9737), .ZN(n7892) );
  NAND2_X1 U10474 ( .A1(n7893), .A2(n10637), .ZN(n10633) );
  NAND2_X1 U10475 ( .A1(n10633), .A2(n7894), .ZN(n10644) );
  NAND2_X1 U10476 ( .A1(n10645), .A2(n10644), .ZN(n10643) );
  INV_X1 U10477 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U10478 ( .A1(n7897), .A2(n7896), .ZN(n7898) );
  NAND2_X1 U10479 ( .A1(n10643), .A2(n7898), .ZN(n11188) );
  NAND2_X1 U10480 ( .A1(n7979), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7903) );
  INV_X1 U10481 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n12121) );
  OR2_X1 U10482 ( .A1(n7980), .A2(n12121), .ZN(n7902) );
  INV_X1 U10483 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7899) );
  OR2_X1 U10484 ( .A1(n7943), .A2(n7899), .ZN(n7901) );
  INV_X1 U10485 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7900) );
  NOR2_X1 U10486 ( .A1(n11251), .A2(n10632), .ZN(n7914) );
  OR2_X1 U10487 ( .A1(n7967), .A2(n10416), .ZN(n7913) );
  INV_X1 U10488 ( .A(SI_2_), .ZN(n7926) );
  XNOR2_X1 U10489 ( .A(n7904), .B(n7926), .ZN(n7909) );
  INV_X1 U10490 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U10491 ( .A1(n7955), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7905) );
  OAI211_X1 U10492 ( .C1(n7955), .C2(n10452), .A(n7905), .B(n10413), .ZN(n7933) );
  NAND2_X1 U10493 ( .A1(n7934), .A2(n7933), .ZN(n7907) );
  NAND2_X1 U10494 ( .A1(n7955), .A2(n10415), .ZN(n7906) );
  OAI211_X1 U10495 ( .C1(n7955), .C2(P2_DATAO_REG_1__SCAN_IN), .A(n7906), .B(
        SI_1_), .ZN(n7925) );
  NAND2_X1 U10496 ( .A1(n7907), .A2(n7925), .ZN(n7908) );
  XNOR2_X1 U10497 ( .A(n7909), .B(n7908), .ZN(n10468) );
  INV_X1 U10498 ( .A(n7910), .ZN(n7937) );
  INV_X1 U10499 ( .A(n10598), .ZN(n10510) );
  NAND2_X1 U10500 ( .A1(n7956), .A2(n10510), .ZN(n7911) );
  XNOR2_X1 U10501 ( .A(n15537), .B(n7940), .ZN(n7915) );
  NAND2_X1 U10502 ( .A1(n7914), .A2(n7915), .ZN(n7918) );
  INV_X1 U10503 ( .A(n7914), .ZN(n7917) );
  INV_X1 U10504 ( .A(n7915), .ZN(n7916) );
  NAND2_X1 U10505 ( .A1(n7917), .A2(n7916), .ZN(n7919) );
  AND2_X1 U10506 ( .A1(n7918), .A2(n7919), .ZN(n11189) );
  NAND2_X1 U10507 ( .A1(n7979), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7924) );
  OR2_X1 U10508 ( .A1(n7980), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10509 ( .A1(n13671), .A2(n13974), .ZN(n7941) );
  MUX2_X1 U10510 ( .A(n10443), .B(n10738), .S(n7955), .Z(n7951) );
  XNOR2_X1 U10511 ( .A(n7951), .B(SI_3_), .ZN(n7949) );
  INV_X1 U10512 ( .A(n7925), .ZN(n7931) );
  OAI211_X1 U10513 ( .C1(n7955), .C2(n10467), .A(n7927), .B(n7926), .ZN(n7932)
         );
  NAND2_X1 U10514 ( .A1(n7955), .A2(n10416), .ZN(n7928) );
  OAI211_X1 U10515 ( .C1(P2_DATAO_REG_2__SCAN_IN), .C2(n7955), .A(n7928), .B(
        SI_2_), .ZN(n7929) );
  INV_X1 U10516 ( .A(n7929), .ZN(n7930) );
  NAND3_X1 U10517 ( .A1(n7934), .A2(n7933), .A3(n7932), .ZN(n7935) );
  NAND2_X1 U10518 ( .A1(n7936), .A2(n7935), .ZN(n7950) );
  XNOR2_X1 U10519 ( .A(n7950), .B(n7949), .ZN(n10442) );
  NAND2_X1 U10520 ( .A1(n7956), .A2(n15453), .ZN(n7938) );
  OAI211_X2 U10521 ( .C1(n7948), .C2(n10442), .A(n7939), .B(n7938), .ZN(n8571)
         );
  XNOR2_X1 U10522 ( .A(n8571), .B(n7940), .ZN(n7942) );
  XNOR2_X1 U10523 ( .A(n7941), .B(n7942), .ZN(n11179) );
  NAND2_X1 U10524 ( .A1(n7979), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7946) );
  XNOR2_X1 U10525 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n12028) );
  INV_X1 U10526 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n12027) );
  OR2_X1 U10527 ( .A1(n7943), .A2(n12027), .ZN(n7944) );
  NAND2_X1 U10528 ( .A1(n13670), .A2(n13974), .ZN(n7965) );
  INV_X1 U10529 ( .A(n7948), .ZN(n7976) );
  NAND2_X1 U10530 ( .A1(n7950), .A2(n7949), .ZN(n7954) );
  INV_X1 U10531 ( .A(n7951), .ZN(n7952) );
  NAND2_X1 U10532 ( .A1(n7952), .A2(SI_3_), .ZN(n7953) );
  XNOR2_X1 U10533 ( .A(n7974), .B(SI_4_), .ZN(n7971) );
  XNOR2_X1 U10534 ( .A(n7973), .B(n7971), .ZN(n10408) );
  NAND2_X1 U10535 ( .A1(n7976), .A2(n10408), .ZN(n7963) );
  NAND2_X1 U10536 ( .A1(n7958), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7957) );
  MUX2_X1 U10537 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7957), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7961) );
  INV_X1 U10538 ( .A(n7958), .ZN(n7960) );
  INV_X1 U10539 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U10540 ( .A1(n7960), .A2(n7959), .ZN(n7969) );
  NAND2_X1 U10541 ( .A1(n7961), .A2(n7969), .ZN(n10507) );
  INV_X1 U10542 ( .A(n10507), .ZN(n10532) );
  NAND2_X1 U10543 ( .A1(n7956), .A2(n10532), .ZN(n7962) );
  OAI211_X1 U10544 ( .C1(n8719), .C2(n10409), .A(n7963), .B(n7962), .ZN(n8582)
         );
  XNOR2_X1 U10545 ( .A(n6432), .B(n7940), .ZN(n7964) );
  NAND2_X1 U10546 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  OAI21_X1 U10547 ( .B1(n7965), .B2(n7964), .A(n7966), .ZN(n10887) );
  NAND2_X1 U10548 ( .A1(n7969), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7968) );
  MUX2_X1 U10549 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7968), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n7970) );
  AOI22_X1 U10550 ( .A1(n8691), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7956), .B2(
        n15466), .ZN(n7978) );
  INV_X1 U10551 ( .A(n7971), .ZN(n7972) );
  NAND2_X1 U10552 ( .A1(n7974), .A2(SI_4_), .ZN(n7975) );
  XNOR2_X1 U10553 ( .A(n7995), .B(n7994), .ZN(n10410) );
  NAND2_X1 U10554 ( .A1(n10410), .A2(n7976), .ZN(n7977) );
  XNOR2_X1 U10555 ( .A(n12038), .B(n7940), .ZN(n7988) );
  NAND2_X1 U10556 ( .A1(n7979), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10557 ( .A1(n8002), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7985) );
  INV_X1 U10558 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U10559 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7981) );
  NAND2_X1 U10560 ( .A1(n7982), .A2(n7981), .ZN(n7983) );
  NAND2_X1 U10561 ( .A1(n8003), .A2(n7983), .ZN(n12020) );
  OR2_X1 U10562 ( .A1(n8424), .A2(n12020), .ZN(n7984) );
  NAND2_X1 U10563 ( .A1(n13669), .A2(n13974), .ZN(n7989) );
  NAND2_X1 U10564 ( .A1(n7988), .A2(n7989), .ZN(n7993) );
  INV_X1 U10565 ( .A(n7988), .ZN(n7991) );
  INV_X1 U10566 ( .A(n7989), .ZN(n7990) );
  NAND2_X1 U10567 ( .A1(n7991), .A2(n7990), .ZN(n7992) );
  AND2_X1 U10568 ( .A1(n7993), .A2(n7992), .ZN(n11204) );
  NAND2_X1 U10569 ( .A1(n7996), .A2(SI_5_), .ZN(n7997) );
  NAND2_X1 U10570 ( .A1(n10417), .A2(n7976), .ZN(n8001) );
  NAND2_X1 U10571 ( .A1(n7998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7999) );
  XNOR2_X1 U10572 ( .A(n7999), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U10573 ( .A1(n8691), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8279), .B2(
        n10538), .ZN(n8000) );
  XNOR2_X1 U10574 ( .A(n12046), .B(n7940), .ZN(n8009) );
  INV_X1 U10575 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10537) );
  OR2_X1 U10576 ( .A1(n8708), .A2(n10537), .ZN(n8007) );
  NAND2_X1 U10577 ( .A1(n8003), .A2(n6994), .ZN(n8004) );
  NAND2_X1 U10578 ( .A1(n6604), .A2(n8004), .ZN(n11146) );
  OR2_X1 U10579 ( .A1(n8424), .A2(n11146), .ZN(n8006) );
  INV_X1 U10580 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8005) );
  NOR2_X1 U10581 ( .A1(n11312), .A2(n12569), .ZN(n8008) );
  XNOR2_X1 U10582 ( .A(n8008), .B(n8009), .ZN(n11144) );
  INV_X1 U10583 ( .A(n8011), .ZN(n8012) );
  NAND2_X1 U10584 ( .A1(n8012), .A2(SI_6_), .ZN(n8013) );
  MUX2_X1 U10585 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9755), .Z(n8033) );
  XNOR2_X1 U10586 ( .A(n8031), .B(n8030), .ZN(n10432) );
  NAND2_X1 U10587 ( .A1(n7910), .A2(n8014), .ZN(n8048) );
  NAND2_X1 U10588 ( .A1(n8048), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8015) );
  XNOR2_X1 U10589 ( .A(n8015), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U10590 ( .A1(n8691), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8279), .B2(
        n10664), .ZN(n8016) );
  INV_X1 U10591 ( .A(n8016), .ZN(n8017) );
  INV_X2 U10592 ( .A(n7940), .ZN(n8490) );
  XNOR2_X1 U10593 ( .A(n11999), .B(n8490), .ZN(n8026) );
  NAND2_X1 U10594 ( .A1(n7920), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8025) );
  INV_X1 U10595 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8019) );
  OR2_X1 U10596 ( .A1(n8018), .A2(n8019), .ZN(n8024) );
  INV_X1 U10597 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U10598 ( .A1(n6604), .A2(n8020), .ZN(n8021) );
  NAND2_X1 U10599 ( .A1(n8055), .A2(n8021), .ZN(n11998) );
  OR2_X1 U10600 ( .A1(n8424), .A2(n11998), .ZN(n8023) );
  INV_X1 U10601 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11997) );
  OR2_X1 U10602 ( .A1(n8708), .A2(n11997), .ZN(n8022) );
  NOR2_X1 U10603 ( .A1(n11475), .A2(n12569), .ZN(n8027) );
  XNOR2_X1 U10604 ( .A(n8026), .B(n8027), .ZN(n11342) );
  INV_X1 U10605 ( .A(n8026), .ZN(n8028) );
  NAND2_X1 U10606 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  NAND2_X1 U10607 ( .A1(n8033), .A2(SI_7_), .ZN(n8034) );
  MUX2_X1 U10608 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10436), .Z(n8036) );
  MUX2_X1 U10609 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10436), .Z(n8070) );
  NAND2_X1 U10610 ( .A1(n10469), .A2(n8718), .ZN(n8040) );
  NAND2_X1 U10611 ( .A1(n8196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8038) );
  XNOR2_X1 U10612 ( .A(n8038), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11168) );
  AOI22_X1 U10613 ( .A1(n8691), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8279), .B2(
        n11168), .ZN(n8039) );
  XNOR2_X1 U10614 ( .A(n11984), .B(n8490), .ZN(n11699) );
  NAND2_X1 U10615 ( .A1(n7920), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8045) );
  OR2_X1 U10616 ( .A1(n8018), .A2(n6675), .ZN(n8044) );
  NAND2_X1 U10617 ( .A1(n8057), .A2(n10669), .ZN(n8041) );
  NAND2_X1 U10618 ( .A1(n8076), .A2(n8041), .ZN(n11983) );
  OR2_X1 U10619 ( .A1(n8424), .A2(n11983), .ZN(n8043) );
  INV_X1 U10620 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11979) );
  OR2_X1 U10621 ( .A1(n8708), .A2(n11979), .ZN(n8042) );
  OR2_X1 U10622 ( .A1(n11754), .A2(n12569), .ZN(n11698) );
  NAND2_X1 U10623 ( .A1(n10448), .A2(n8718), .ZN(n8053) );
  NAND2_X1 U10624 ( .A1(n8049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8050) );
  MUX2_X1 U10625 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8050), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8051) );
  NAND2_X1 U10626 ( .A1(n8051), .A2(n8196), .ZN(n15489) );
  INV_X1 U10627 ( .A(n15489), .ZN(n10665) );
  AOI22_X1 U10628 ( .A1(n8691), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8279), .B2(
        n10665), .ZN(n8052) );
  INV_X1 U10629 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8054) );
  OR2_X1 U10630 ( .A1(n8018), .A2(n8054), .ZN(n8060) );
  NAND2_X1 U10631 ( .A1(n8055), .A2(n6690), .ZN(n8056) );
  NAND2_X1 U10632 ( .A1(n8057), .A2(n8056), .ZN(n12014) );
  OR2_X1 U10633 ( .A1(n8424), .A2(n12014), .ZN(n8059) );
  INV_X1 U10634 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n12010) );
  OR2_X1 U10635 ( .A1(n8708), .A2(n12010), .ZN(n8058) );
  OR2_X1 U10636 ( .A1(n11702), .A2(n12569), .ZN(n11693) );
  OAI22_X1 U10637 ( .A1(n11699), .A2(n11698), .B1(n11694), .B2(n11693), .ZN(
        n8062) );
  INV_X1 U10638 ( .A(n8062), .ZN(n8068) );
  INV_X1 U10639 ( .A(n11694), .ZN(n11697) );
  INV_X1 U10640 ( .A(n11693), .ZN(n11473) );
  INV_X1 U10641 ( .A(n11698), .ZN(n8063) );
  OAI21_X1 U10642 ( .B1(n11697), .B2(n11473), .A(n8063), .ZN(n8065) );
  AND3_X1 U10643 ( .A1(n11694), .A2(n11693), .A3(n11698), .ZN(n8064) );
  AOI21_X1 U10644 ( .B1(n11699), .B2(n8065), .A(n8064), .ZN(n8066) );
  INV_X1 U10645 ( .A(n8066), .ZN(n8067) );
  NAND2_X1 U10646 ( .A1(n8070), .A2(SI_9_), .ZN(n8071) );
  MUX2_X1 U10647 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10436), .Z(n8089) );
  XNOR2_X1 U10648 ( .A(n8088), .B(n8086), .ZN(n10472) );
  NAND2_X1 U10649 ( .A1(n10472), .A2(n8718), .ZN(n8074) );
  NAND2_X1 U10650 ( .A1(n8095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8072) );
  XNOR2_X1 U10651 ( .A(n8072), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U10652 ( .A1(n8691), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8279), 
        .B2(n11465), .ZN(n8073) );
  XNOR2_X1 U10653 ( .A(n12110), .B(n8490), .ZN(n8082) );
  INV_X1 U10654 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8075) );
  OR2_X1 U10655 ( .A1(n8018), .A2(n8075), .ZN(n8080) );
  NAND2_X1 U10656 ( .A1(n8076), .A2(n11755), .ZN(n8077) );
  NAND2_X1 U10657 ( .A1(n8101), .A2(n8077), .ZN(n11752) );
  OR2_X1 U10658 ( .A1(n8424), .A2(n11752), .ZN(n8079) );
  INV_X1 U10659 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11167) );
  OR2_X1 U10660 ( .A1(n8708), .A2(n11167), .ZN(n8078) );
  NOR2_X1 U10661 ( .A1(n12168), .A2(n12569), .ZN(n8083) );
  XNOR2_X1 U10662 ( .A(n8082), .B(n8083), .ZN(n11751) );
  INV_X1 U10663 ( .A(n8082), .ZN(n8084) );
  NAND2_X1 U10664 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  NAND2_X1 U10665 ( .A1(n8089), .A2(SI_10_), .ZN(n8117) );
  NAND2_X1 U10666 ( .A1(n8122), .A2(n8117), .ZN(n8093) );
  MUX2_X1 U10667 ( .A(n10489), .B(n10487), .S(n10436), .Z(n8090) );
  INV_X1 U10668 ( .A(SI_11_), .ZN(n10454) );
  NAND2_X1 U10669 ( .A1(n8090), .A2(n10454), .ZN(n8119) );
  INV_X1 U10670 ( .A(n8090), .ZN(n8091) );
  NAND2_X1 U10671 ( .A1(n8091), .A2(SI_11_), .ZN(n8116) );
  NAND2_X1 U10672 ( .A1(n8119), .A2(n8116), .ZN(n8092) );
  NAND2_X1 U10673 ( .A1(n8093), .A2(n8092), .ZN(n8094) );
  NAND2_X1 U10674 ( .A1(n8115), .A2(n8094), .ZN(n10486) );
  NAND2_X1 U10675 ( .A1(n10486), .A2(n8718), .ZN(n8100) );
  NAND2_X1 U10676 ( .A1(n8097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8096) );
  MUX2_X1 U10677 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8096), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n8098) );
  NAND2_X1 U10678 ( .A1(n8098), .A2(n8147), .ZN(n11568) );
  INV_X1 U10679 ( .A(n11568), .ZN(n11573) );
  AOI22_X1 U10680 ( .A1(n8691), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11573), 
        .B2(n8279), .ZN(n8099) );
  XNOR2_X1 U10681 ( .A(n14161), .B(n8490), .ZN(n8107) );
  NAND2_X1 U10682 ( .A1(n6947), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8106) );
  INV_X1 U10683 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14158) );
  OR2_X1 U10684 ( .A1(n7019), .A2(n14158), .ZN(n8105) );
  NAND2_X1 U10685 ( .A1(n8101), .A2(n6695), .ZN(n8102) );
  NAND2_X1 U10686 ( .A1(n8128), .A2(n8102), .ZN(n12172) );
  OR2_X1 U10687 ( .A1(n8424), .A2(n12172), .ZN(n8104) );
  INV_X1 U10688 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n12173) );
  OR2_X1 U10689 ( .A1(n8708), .A2(n12173), .ZN(n8103) );
  OR2_X1 U10690 ( .A1(n12195), .A2(n12569), .ZN(n8108) );
  NAND2_X1 U10691 ( .A1(n8107), .A2(n8108), .ZN(n11897) );
  NAND2_X1 U10692 ( .A1(n11898), .A2(n11897), .ZN(n8111) );
  INV_X1 U10693 ( .A(n8107), .ZN(n8110) );
  INV_X1 U10694 ( .A(n8108), .ZN(n8109) );
  NAND2_X1 U10695 ( .A1(n8110), .A2(n8109), .ZN(n11896) );
  MUX2_X1 U10696 ( .A(n10581), .B(n10579), .S(n10436), .Z(n8112) );
  INV_X1 U10697 ( .A(SI_12_), .ZN(n10478) );
  INV_X1 U10698 ( .A(n8112), .ZN(n8113) );
  NAND3_X1 U10699 ( .A1(n8115), .A2(n8120), .A3(n8119), .ZN(n8123) );
  NAND2_X1 U10700 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  NAND2_X1 U10701 ( .A1(n8123), .A2(n6587), .ZN(n10578) );
  NAND2_X1 U10702 ( .A1(n10578), .A2(n8718), .ZN(n8126) );
  NAND2_X1 U10703 ( .A1(n8147), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8124) );
  XNOR2_X1 U10704 ( .A(n8124), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U10705 ( .A1(n8691), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11842), 
        .B2(n8279), .ZN(n8125) );
  XNOR2_X1 U10706 ( .A(n12282), .B(n8490), .ZN(n8134) );
  NAND2_X1 U10707 ( .A1(n7920), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8133) );
  INV_X1 U10708 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11571) );
  OR2_X1 U10709 ( .A1(n8018), .A2(n11571), .ZN(n8132) );
  INV_X1 U10710 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U10711 ( .A1(n8128), .A2(n8127), .ZN(n8129) );
  NAND2_X1 U10712 ( .A1(n8153), .A2(n8129), .ZN(n12283) );
  OR2_X1 U10713 ( .A1(n8424), .A2(n12283), .ZN(n8131) );
  INV_X1 U10714 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12284) );
  OR2_X1 U10715 ( .A1(n8708), .A2(n12284), .ZN(n8130) );
  OR2_X1 U10716 ( .A1(n12295), .A2(n12569), .ZN(n8135) );
  NAND2_X1 U10717 ( .A1(n8134), .A2(n8135), .ZN(n8139) );
  INV_X1 U10718 ( .A(n8134), .ZN(n8137) );
  INV_X1 U10719 ( .A(n8135), .ZN(n8136) );
  NAND2_X1 U10720 ( .A1(n8137), .A2(n8136), .ZN(n8138) );
  NAND2_X1 U10721 ( .A1(n8139), .A2(n8138), .ZN(n12193) );
  MUX2_X1 U10722 ( .A(n10681), .B(n10679), .S(n9755), .Z(n8141) );
  INV_X1 U10723 ( .A(SI_13_), .ZN(n10626) );
  INV_X1 U10724 ( .A(n8141), .ZN(n8142) );
  NAND2_X1 U10725 ( .A1(n8142), .A2(SI_13_), .ZN(n8143) );
  NAND2_X1 U10726 ( .A1(n8162), .A2(n8146), .ZN(n10678) );
  NAND2_X1 U10727 ( .A1(n10678), .A2(n8718), .ZN(n8152) );
  INV_X1 U10728 ( .A(n8147), .ZN(n8149) );
  INV_X1 U10729 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U10730 ( .A1(n8149), .A2(n8148), .ZN(n8164) );
  NAND2_X1 U10731 ( .A1(n8164), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8150) );
  XNOR2_X1 U10732 ( .A(n8150), .B(P2_IR_REG_13__SCAN_IN), .ZN(n12392) );
  AOI22_X1 U10733 ( .A1(n12392), .A2(n8279), .B1(n8691), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n8151) );
  XNOR2_X1 U10734 ( .A(n14089), .B(n7940), .ZN(n8160) );
  NAND2_X1 U10735 ( .A1(n6947), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U10736 ( .A1(n8002), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8157) );
  INV_X1 U10737 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U10738 ( .A1(n8153), .A2(n11849), .ZN(n8154) );
  NAND2_X1 U10739 ( .A1(n8171), .A2(n8154), .ZN(n12314) );
  OR2_X1 U10740 ( .A1(n8424), .A2(n12314), .ZN(n8155) );
  NAND4_X1 U10741 ( .A1(n8158), .A2(n8157), .A3(n8156), .A4(n8155), .ZN(n13967) );
  NAND2_X1 U10742 ( .A1(n13967), .A2(n13974), .ZN(n8159) );
  XNOR2_X1 U10743 ( .A(n8160), .B(n8159), .ZN(n12309) );
  INV_X1 U10744 ( .A(SI_14_), .ZN(n10675) );
  NAND2_X1 U10745 ( .A1(n8191), .A2(n10675), .ZN(n8211) );
  OR2_X1 U10746 ( .A1(n8191), .A2(n10675), .ZN(n8163) );
  MUX2_X1 U10747 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10436), .Z(n8212) );
  XNOR2_X1 U10748 ( .A(n8213), .B(n8212), .ZN(n11198) );
  NAND2_X1 U10749 ( .A1(n11198), .A2(n8718), .ZN(n8167) );
  OAI21_X1 U10750 ( .B1(n8164), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8165) );
  XNOR2_X1 U10751 ( .A(n8165), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U10752 ( .A1(n12474), .A2(n8279), .B1(n8691), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n8166) );
  XNOR2_X1 U10753 ( .A(n13980), .B(n8490), .ZN(n8178) );
  NAND2_X1 U10754 ( .A1(n6947), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8177) );
  INV_X1 U10755 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8168) );
  OR2_X1 U10756 ( .A1(n8708), .A2(n8168), .ZN(n8176) );
  INV_X1 U10757 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U10758 ( .A1(n8171), .A2(n8170), .ZN(n8172) );
  NAND2_X1 U10759 ( .A1(n8205), .A2(n8172), .ZN(n13976) );
  OR2_X1 U10760 ( .A1(n8424), .A2(n13976), .ZN(n8175) );
  INV_X1 U10761 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8173) );
  OR2_X1 U10762 ( .A1(n7019), .A2(n8173), .ZN(n8174) );
  OR2_X1 U10763 ( .A1(n13659), .A2(n12569), .ZN(n8179) );
  NAND2_X1 U10764 ( .A1(n8178), .A2(n8179), .ZN(n8183) );
  INV_X1 U10765 ( .A(n8178), .ZN(n8181) );
  INV_X1 U10766 ( .A(n8179), .ZN(n8180) );
  NAND2_X1 U10767 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  NAND2_X1 U10768 ( .A1(n8183), .A2(n8182), .ZN(n13528) );
  INV_X1 U10769 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11305) );
  MUX2_X1 U10770 ( .A(n11303), .B(n11305), .S(n10436), .Z(n8184) );
  INV_X1 U10771 ( .A(SI_15_), .ZN(n10629) );
  INV_X1 U10772 ( .A(n8184), .ZN(n8185) );
  NAND2_X1 U10773 ( .A1(n8185), .A2(SI_15_), .ZN(n8186) );
  INV_X1 U10774 ( .A(n8212), .ZN(n8187) );
  INV_X1 U10775 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11298) );
  INV_X1 U10776 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11301) );
  MUX2_X1 U10777 ( .A(n11298), .B(n11301), .S(n10436), .Z(n8193) );
  INV_X1 U10778 ( .A(SI_16_), .ZN(n8192) );
  INV_X1 U10779 ( .A(n8193), .ZN(n8194) );
  NAND2_X1 U10780 ( .A1(n8194), .A2(SI_16_), .ZN(n8253) );
  AND2_X1 U10781 ( .A1(n8250), .A2(n8253), .ZN(n8229) );
  NAND2_X1 U10782 ( .A1(n11297), .A2(n8718), .ZN(n8199) );
  INV_X1 U10783 ( .A(n7867), .ZN(n8195) );
  OR2_X1 U10784 ( .A1(n8196), .A2(n8195), .ZN(n8217) );
  OR2_X1 U10785 ( .A1(n8217), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U10786 ( .A1(n8235), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8197) );
  XNOR2_X1 U10787 ( .A(n8197), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U10788 ( .A1(n8691), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8279), 
        .B2(n15504), .ZN(n8198) );
  XNOR2_X1 U10789 ( .A(n13941), .B(n8490), .ZN(n8222) );
  INV_X1 U10790 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n12390) );
  INV_X1 U10791 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10792 ( .A1(n8207), .A2(n8200), .ZN(n8201) );
  NAND2_X1 U10793 ( .A1(n8240), .A2(n8201), .ZN(n13937) );
  OR2_X1 U10794 ( .A1(n13937), .A2(n8424), .ZN(n8204) );
  AOI22_X1 U10795 ( .A1(n7920), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n6947), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U10796 ( .A1(n8002), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U10797 ( .A1(n13658), .A2(n13974), .ZN(n8223) );
  NAND2_X1 U10798 ( .A1(n8222), .A2(n8223), .ZN(n13575) );
  NAND2_X1 U10799 ( .A1(n8205), .A2(n12390), .ZN(n8206) );
  NAND2_X1 U10800 ( .A1(n8207), .A2(n8206), .ZN(n13957) );
  INV_X1 U10801 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n13958) );
  OAI22_X1 U10802 ( .A1(n13957), .A2(n8424), .B1(n8708), .B2(n13958), .ZN(
        n8210) );
  INV_X1 U10803 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14149) );
  NAND2_X1 U10804 ( .A1(n6947), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8208) );
  OAI21_X1 U10805 ( .B1(n14149), .B2(n7019), .A(n8208), .ZN(n8209) );
  OR2_X1 U10806 ( .A1(n8210), .A2(n8209), .ZN(n13969) );
  AND2_X1 U10807 ( .A1(n13969), .A2(n13974), .ZN(n13639) );
  NAND2_X1 U10808 ( .A1(n13575), .A2(n13639), .ZN(n8226) );
  INV_X1 U10809 ( .A(n8214), .ZN(n8215) );
  NAND2_X1 U10810 ( .A1(n8217), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8218) );
  MUX2_X1 U10811 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8218), .S(
        P2_IR_REG_15__SCAN_IN), .Z(n8219) );
  AND2_X1 U10812 ( .A1(n8219), .A2(n8235), .ZN(n13685) );
  AOI22_X1 U10813 ( .A1(n8691), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8279), 
        .B2(n13685), .ZN(n8220) );
  XNOR2_X1 U10814 ( .A(n13955), .B(n7940), .ZN(n13572) );
  INV_X1 U10815 ( .A(n13572), .ZN(n13573) );
  NAND2_X1 U10816 ( .A1(n13575), .A2(n13573), .ZN(n8221) );
  NAND2_X1 U10817 ( .A1(n8226), .A2(n8221), .ZN(n8228) );
  INV_X1 U10818 ( .A(n8222), .ZN(n8225) );
  INV_X1 U10819 ( .A(n8223), .ZN(n8224) );
  NAND2_X1 U10820 ( .A1(n8225), .A2(n8224), .ZN(n13574) );
  OAI21_X1 U10821 ( .B1(n8226), .B2(n13572), .A(n13574), .ZN(n8227) );
  INV_X1 U10822 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11366) );
  INV_X1 U10823 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11369) );
  MUX2_X1 U10824 ( .A(n11366), .B(n11369), .S(n9755), .Z(n8231) );
  INV_X1 U10825 ( .A(SI_17_), .ZN(n10682) );
  INV_X1 U10826 ( .A(n8231), .ZN(n8232) );
  NAND2_X1 U10827 ( .A1(n8232), .A2(SI_17_), .ZN(n8233) );
  NAND2_X1 U10828 ( .A1(n8256), .A2(n8233), .ZN(n8254) );
  INV_X1 U10829 ( .A(n8254), .ZN(n8234) );
  OR2_X1 U10830 ( .A1(n8235), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U10831 ( .A1(n8258), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8236) );
  XNOR2_X1 U10832 ( .A(n8236), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15518) );
  AOI22_X1 U10833 ( .A1(n8691), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n15518), 
        .B2(n8279), .ZN(n8237) );
  XNOR2_X1 U10834 ( .A(n13920), .B(n7940), .ZN(n8244) );
  INV_X1 U10835 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U10836 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  NAND2_X1 U10837 ( .A1(n8263), .A2(n8241), .ZN(n13586) );
  NAND2_X1 U10838 ( .A1(n8002), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8242) );
  OAI211_X1 U10839 ( .C1(n13586), .C2(n8424), .A(n8243), .B(n8242), .ZN(n13893) );
  NAND2_X1 U10840 ( .A1(n13893), .A2(n13974), .ZN(n8245) );
  NAND2_X1 U10841 ( .A1(n8244), .A2(n8245), .ZN(n8249) );
  INV_X1 U10842 ( .A(n8244), .ZN(n8247) );
  INV_X1 U10843 ( .A(n8245), .ZN(n8246) );
  NAND2_X1 U10844 ( .A1(n8247), .A2(n8246), .ZN(n8248) );
  AND2_X1 U10845 ( .A1(n8249), .A2(n8248), .ZN(n13583) );
  INV_X1 U10846 ( .A(n8253), .ZN(n8255) );
  INV_X1 U10847 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11526) );
  MUX2_X1 U10848 ( .A(n11528), .B(n11526), .S(n10436), .Z(n8293) );
  XNOR2_X1 U10849 ( .A(n8273), .B(n8293), .ZN(n11525) );
  NAND2_X1 U10850 ( .A1(n11525), .A2(n8718), .ZN(n8261) );
  OAI21_X1 U10851 ( .B1(n8258), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8259) );
  XNOR2_X1 U10852 ( .A(n8259), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U10853 ( .A1(n13699), .A2(n8279), .B1(n8691), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8260) );
  XNOR2_X1 U10854 ( .A(n13901), .B(n7940), .ZN(n8271) );
  INV_X1 U10855 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U10856 ( .A1(n8263), .A2(n8262), .ZN(n8264) );
  NAND2_X1 U10857 ( .A1(n8308), .A2(n8264), .ZN(n13902) );
  OR2_X1 U10858 ( .A1(n13902), .A2(n8424), .ZN(n8269) );
  INV_X1 U10859 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13903) );
  NAND2_X1 U10860 ( .A1(n6947), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8265) );
  OAI211_X1 U10861 ( .C1(n13903), .C2(n8708), .A(n8266), .B(n8265), .ZN(n8267)
         );
  INV_X1 U10862 ( .A(n8267), .ZN(n8268) );
  NOR2_X1 U10863 ( .A1(n13549), .A2(n12569), .ZN(n8270) );
  XNOR2_X1 U10864 ( .A(n8271), .B(n8270), .ZN(n13621) );
  NAND2_X1 U10865 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  INV_X1 U10866 ( .A(n8293), .ZN(n8297) );
  INV_X1 U10867 ( .A(SI_18_), .ZN(n11052) );
  OR2_X1 U10868 ( .A1(n8296), .A2(n11052), .ZN(n8274) );
  MUX2_X1 U10869 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10436), .Z(n8275) );
  INV_X1 U10870 ( .A(n8275), .ZN(n8276) );
  INV_X1 U10871 ( .A(SI_19_), .ZN(n12567) );
  NAND2_X1 U10872 ( .A1(n8276), .A2(n12567), .ZN(n8298) );
  NAND2_X1 U10873 ( .A1(n8300), .A2(n8298), .ZN(n8277) );
  NAND2_X1 U10874 ( .A1(n11613), .A2(n8718), .ZN(n8281) );
  AOI22_X1 U10875 ( .A1(n8691), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13705), 
        .B2(n8279), .ZN(n8280) );
  XNOR2_X1 U10876 ( .A(n13882), .B(n7940), .ZN(n8292) );
  INV_X1 U10877 ( .A(n8292), .ZN(n8290) );
  XNOR2_X1 U10878 ( .A(n8308), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n13880) );
  NAND2_X1 U10879 ( .A1(n13880), .A2(n8282), .ZN(n8288) );
  INV_X1 U10880 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8285) );
  NAND2_X1 U10881 ( .A1(n7920), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U10882 ( .A1(n6947), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8283) );
  OAI211_X1 U10883 ( .C1(n8285), .C2(n8708), .A(n8284), .B(n8283), .ZN(n8286)
         );
  INV_X1 U10884 ( .A(n8286), .ZN(n8287) );
  NOR2_X1 U10885 ( .A1(n13859), .A2(n12569), .ZN(n8291) );
  INV_X1 U10886 ( .A(n8291), .ZN(n8289) );
  AND2_X1 U10887 ( .A1(n8292), .A2(n8291), .ZN(n13546) );
  OAI21_X1 U10888 ( .B1(n8293), .B2(n11052), .A(n8300), .ZN(n8294) );
  INV_X1 U10889 ( .A(n8294), .ZN(n8295) );
  NOR2_X1 U10890 ( .A1(n8297), .A2(SI_18_), .ZN(n8301) );
  INV_X1 U10891 ( .A(n8298), .ZN(n8299) );
  XNOR2_X1 U10892 ( .A(n8339), .B(SI_20_), .ZN(n8326) );
  INV_X1 U10893 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12564) );
  MUX2_X1 U10894 ( .A(n11710), .B(n12564), .S(n10436), .Z(n8335) );
  XNOR2_X1 U10895 ( .A(n8326), .B(n8335), .ZN(n11708) );
  NAND2_X1 U10896 ( .A1(n11708), .A2(n8718), .ZN(n8305) );
  OR2_X1 U10897 ( .A1(n8719), .A2(n12564), .ZN(n8304) );
  XNOR2_X1 U10898 ( .A(n14140), .B(n8490), .ZN(n8315) );
  INV_X1 U10899 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n13550) );
  INV_X1 U10900 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8306) );
  OAI21_X1 U10901 ( .B1(n8308), .B2(n13550), .A(n8306), .ZN(n8309) );
  NAND2_X1 U10902 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n8307) );
  NAND2_X1 U10903 ( .A1(n8309), .A2(n8319), .ZN(n13863) );
  OR2_X1 U10904 ( .A1(n13863), .A2(n8424), .ZN(n8314) );
  INV_X1 U10905 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13864) );
  NAND2_X1 U10906 ( .A1(n7920), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8311) );
  NAND2_X1 U10907 ( .A1(n6947), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8310) );
  OAI211_X1 U10908 ( .C1(n13864), .C2(n8708), .A(n8311), .B(n8310), .ZN(n8312)
         );
  INV_X1 U10909 ( .A(n8312), .ZN(n8313) );
  NAND2_X1 U10910 ( .A1(n8314), .A2(n8313), .ZN(n13656) );
  NAND2_X1 U10911 ( .A1(n13656), .A2(n13974), .ZN(n8316) );
  XNOR2_X1 U10912 ( .A(n8315), .B(n8316), .ZN(n13601) );
  INV_X1 U10913 ( .A(n8315), .ZN(n8317) );
  AND2_X1 U10914 ( .A1(n8317), .A2(n8316), .ZN(n8359) );
  INV_X1 U10915 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10916 ( .A1(n8319), .A2(n8318), .ZN(n8320) );
  NAND2_X1 U10917 ( .A1(n8375), .A2(n8320), .ZN(n13846) );
  OR2_X1 U10918 ( .A1(n13846), .A2(n8424), .ZN(n8325) );
  INV_X1 U10919 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13847) );
  NAND2_X1 U10920 ( .A1(n6947), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8322) );
  OAI211_X1 U10921 ( .C1(n13847), .C2(n8708), .A(n8322), .B(n8321), .ZN(n8323)
         );
  INV_X1 U10922 ( .A(n8323), .ZN(n8324) );
  NAND2_X1 U10923 ( .A1(n13655), .A2(n13974), .ZN(n8333) );
  NAND2_X1 U10924 ( .A1(n8326), .A2(n8334), .ZN(n8328) );
  INV_X1 U10925 ( .A(SI_20_), .ZN(n11539) );
  OR2_X1 U10926 ( .A1(n8339), .A2(n11539), .ZN(n8327) );
  MUX2_X1 U10927 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9755), .Z(n8336) );
  XNOR2_X1 U10928 ( .A(n8336), .B(SI_21_), .ZN(n8329) );
  NAND2_X1 U10929 ( .A1(n11769), .A2(n8718), .ZN(n8332) );
  INV_X1 U10930 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11771) );
  OR2_X1 U10931 ( .A1(n8719), .A2(n11771), .ZN(n8331) );
  XNOR2_X1 U10932 ( .A(n14137), .B(n8490), .ZN(n8364) );
  XOR2_X1 U10933 ( .A(n8333), .B(n8364), .Z(n13557) );
  INV_X1 U10934 ( .A(n8364), .ZN(n8360) );
  INV_X1 U10935 ( .A(n8333), .ZN(n8368) );
  NAND2_X1 U10936 ( .A1(n8360), .A2(n8368), .ZN(n8370) );
  NOR2_X1 U10937 ( .A1(n8335), .A2(n11539), .ZN(n8337) );
  AOI22_X1 U10938 ( .A1(n8337), .A2(n7818), .B1(n8336), .B2(SI_21_), .ZN(n8338) );
  MUX2_X1 U10939 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10436), .Z(n8392) );
  XNOR2_X1 U10940 ( .A(n8931), .B(n8392), .ZN(n11916) );
  NAND2_X1 U10941 ( .A1(n11916), .A2(n8718), .ZN(n8341) );
  NAND2_X1 U10942 ( .A1(n8691), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8340) );
  XNOR2_X1 U10943 ( .A(n14133), .B(n8490), .ZN(n8365) );
  INV_X1 U10944 ( .A(n8931), .ZN(n8342) );
  NAND2_X1 U10945 ( .A1(n8342), .A2(n8392), .ZN(n8344) );
  NAND2_X1 U10946 ( .A1(n8389), .A2(SI_22_), .ZN(n8343) );
  INV_X1 U10947 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12136) );
  INV_X1 U10948 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10175) );
  MUX2_X1 U10949 ( .A(n12136), .B(n10175), .S(n10436), .Z(n8387) );
  INV_X1 U10950 ( .A(n8387), .ZN(n8393) );
  XNOR2_X1 U10951 ( .A(n8393), .B(SI_23_), .ZN(n8345) );
  XNOR2_X2 U10952 ( .A(n8346), .B(n8345), .ZN(n12134) );
  NAND2_X1 U10953 ( .A1(n12134), .A2(n8718), .ZN(n8348) );
  NAND2_X1 U10954 ( .A1(n8691), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8347) );
  XNOR2_X1 U10955 ( .A(n13541), .B(n8490), .ZN(n13536) );
  INV_X1 U10956 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13615) );
  INV_X1 U10957 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8349) );
  NAND2_X1 U10958 ( .A1(n8377), .A2(n8349), .ZN(n8350) );
  AND2_X1 U10959 ( .A1(n6472), .A2(n8350), .ZN(n13815) );
  NAND2_X1 U10960 ( .A1(n13815), .A2(n8282), .ZN(n8356) );
  INV_X1 U10961 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10962 ( .A1(n6947), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10963 ( .A1(n7920), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8351) );
  OAI211_X1 U10964 ( .C1(n8353), .C2(n8708), .A(n8352), .B(n8351), .ZN(n8354)
         );
  INV_X1 U10965 ( .A(n8354), .ZN(n8355) );
  AND2_X1 U10966 ( .A1(n13794), .A2(n13974), .ZN(n13539) );
  NAND2_X1 U10967 ( .A1(n13535), .A2(n8357), .ZN(n8386) );
  INV_X1 U10968 ( .A(n8359), .ZN(n8367) );
  INV_X1 U10969 ( .A(n8365), .ZN(n8369) );
  OAI211_X1 U10970 ( .C1(n8360), .C2(n8368), .A(n8367), .B(n8369), .ZN(n8361)
         );
  INV_X1 U10971 ( .A(n8361), .ZN(n8362) );
  NAND2_X1 U10972 ( .A1(n13600), .A2(n8362), .ZN(n8374) );
  NAND2_X1 U10973 ( .A1(n8367), .A2(n8368), .ZN(n8363) );
  NAND2_X1 U10974 ( .A1(n8364), .A2(n8363), .ZN(n8366) );
  OAI211_X1 U10975 ( .C1(n8368), .C2(n8367), .A(n8366), .B(n8365), .ZN(n8372)
         );
  NAND2_X1 U10976 ( .A1(n8370), .A2(n8369), .ZN(n8371) );
  NAND2_X1 U10977 ( .A1(n8372), .A2(n8371), .ZN(n8373) );
  NAND2_X1 U10978 ( .A1(n8375), .A2(n13615), .ZN(n8376) );
  NAND2_X1 U10979 ( .A1(n8377), .A2(n8376), .ZN(n13614) );
  OR2_X1 U10980 ( .A1(n13614), .A2(n8424), .ZN(n8383) );
  INV_X1 U10981 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U10982 ( .A1(n6947), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8379) );
  OAI211_X1 U10983 ( .C1(n8708), .C2(n8380), .A(n8379), .B(n8378), .ZN(n8381)
         );
  INV_X1 U10984 ( .A(n8381), .ZN(n8382) );
  NOR2_X1 U10985 ( .A1(n13843), .A2(n12569), .ZN(n13612) );
  OAI21_X1 U10986 ( .B1(n13536), .B2(n13794), .A(n13612), .ZN(n8385) );
  NAND2_X1 U10987 ( .A1(n13536), .A2(n13539), .ZN(n8384) );
  INV_X1 U10988 ( .A(SI_22_), .ZN(n10144) );
  INV_X1 U10989 ( .A(n8392), .ZN(n8390) );
  INV_X1 U10990 ( .A(SI_23_), .ZN(n11618) );
  AOI22_X1 U10991 ( .A1(n10144), .A2(n8390), .B1(n8387), .B2(n11618), .ZN(
        n8388) );
  OAI21_X1 U10992 ( .B1(n8390), .B2(n10144), .A(n11618), .ZN(n8394) );
  AND2_X1 U10993 ( .A1(SI_22_), .A2(SI_23_), .ZN(n8391) );
  AOI22_X1 U10994 ( .A1(n8394), .A2(n8393), .B1(n8392), .B2(n8391), .ZN(n8395)
         );
  INV_X1 U10995 ( .A(SI_24_), .ZN(n12089) );
  INV_X1 U10996 ( .A(n8411), .ZN(n8396) );
  MUX2_X1 U10997 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10436), .Z(n8410) );
  NAND2_X1 U10998 ( .A1(n12207), .A2(n8718), .ZN(n8398) );
  INV_X1 U10999 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12212) );
  OR2_X1 U11000 ( .A1(n8719), .A2(n12212), .ZN(n8397) );
  XNOR2_X1 U11001 ( .A(n14036), .B(n7940), .ZN(n8407) );
  INV_X1 U11002 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13593) );
  INV_X1 U11003 ( .A(n8420), .ZN(n8422) );
  NAND2_X1 U11004 ( .A1(n6472), .A2(n13593), .ZN(n8399) );
  NAND2_X1 U11005 ( .A1(n8422), .A2(n8399), .ZN(n13798) );
  INV_X1 U11006 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U11007 ( .A1(n6947), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8400) );
  OAI211_X1 U11008 ( .C1(n8402), .C2(n8708), .A(n8401), .B(n8400), .ZN(n8403)
         );
  INV_X1 U11009 ( .A(n8403), .ZN(n8404) );
  NAND2_X1 U11010 ( .A1(n13810), .A2(n13974), .ZN(n8406) );
  NOR2_X1 U11011 ( .A1(n8407), .A2(n8406), .ZN(n8408) );
  AOI21_X1 U11012 ( .B1(n8407), .B2(n8406), .A(n8408), .ZN(n13591) );
  INV_X1 U11013 ( .A(n8408), .ZN(n8409) );
  NAND2_X1 U11014 ( .A1(n8412), .A2(SI_24_), .ZN(n8413) );
  INV_X1 U11015 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12320) );
  INV_X1 U11016 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12323) );
  MUX2_X1 U11017 ( .A(n12320), .B(n12323), .S(n10436), .Z(n8415) );
  INV_X1 U11018 ( .A(SI_25_), .ZN(n12292) );
  NAND2_X1 U11019 ( .A1(n8415), .A2(n12292), .ZN(n8445) );
  INV_X1 U11020 ( .A(n8415), .ZN(n8416) );
  NAND2_X1 U11021 ( .A1(n8416), .A2(SI_25_), .ZN(n8417) );
  NAND2_X1 U11022 ( .A1(n8445), .A2(n8417), .ZN(n8443) );
  XNOR2_X1 U11023 ( .A(n8444), .B(n8443), .ZN(n12318) );
  NAND2_X1 U11024 ( .A1(n12318), .A2(n8718), .ZN(n8419) );
  OR2_X1 U11025 ( .A1(n8719), .A2(n12323), .ZN(n8418) );
  XNOR2_X1 U11026 ( .A(n13784), .B(n7940), .ZN(n8431) );
  INV_X1 U11027 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8421) );
  NAND2_X1 U11028 ( .A1(n8422), .A2(n8421), .ZN(n8423) );
  NAND2_X1 U11029 ( .A1(n8436), .A2(n8423), .ZN(n13782) );
  INV_X1 U11030 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13781) );
  NAND2_X1 U11031 ( .A1(n6947), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8426) );
  OAI211_X1 U11032 ( .C1(n8708), .C2(n13781), .A(n8426), .B(n8425), .ZN(n8427)
         );
  INV_X1 U11033 ( .A(n8427), .ZN(n8428) );
  NAND2_X1 U11034 ( .A1(n13795), .A2(n13974), .ZN(n8430) );
  NOR2_X1 U11035 ( .A1(n8431), .A2(n8430), .ZN(n8432) );
  AOI21_X1 U11036 ( .B1(n8431), .B2(n8430), .A(n8432), .ZN(n13564) );
  INV_X1 U11037 ( .A(n8432), .ZN(n8433) );
  INV_X1 U11038 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U11039 ( .A1(n8436), .A2(n8435), .ZN(n8437) );
  INV_X1 U11040 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U11041 ( .A1(n7920), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U11042 ( .A1(n6947), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8438) );
  OAI211_X1 U11043 ( .C1(n8440), .C2(n8708), .A(n8439), .B(n8438), .ZN(n8441)
         );
  INV_X1 U11044 ( .A(n8441), .ZN(n8442) );
  NAND2_X1 U11045 ( .A1(n13773), .A2(n13974), .ZN(n8450) );
  INV_X1 U11046 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15186) );
  INV_X1 U11047 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14185) );
  MUX2_X1 U11048 ( .A(n15186), .B(n14185), .S(n10436), .Z(n8452) );
  XNOR2_X1 U11049 ( .A(n8452), .B(SI_26_), .ZN(n8446) );
  OR2_X1 U11050 ( .A1(n8719), .A2(n14185), .ZN(n8447) );
  XNOR2_X1 U11051 ( .A(n14026), .B(n8490), .ZN(n8449) );
  XOR2_X1 U11052 ( .A(n8450), .B(n8449), .Z(n13629) );
  INV_X1 U11053 ( .A(n8449), .ZN(n8451) );
  INV_X1 U11054 ( .A(SI_26_), .ZN(n13521) );
  INV_X1 U11055 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15184) );
  INV_X1 U11056 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14182) );
  MUX2_X1 U11057 ( .A(n15184), .B(n14182), .S(n10436), .Z(n8470) );
  XNOR2_X1 U11058 ( .A(n8470), .B(SI_27_), .ZN(n8454) );
  OR2_X1 U11059 ( .A1(n8719), .A2(n14182), .ZN(n8455) );
  XNOR2_X1 U11060 ( .A(n13751), .B(n8490), .ZN(n8467) );
  INV_X1 U11061 ( .A(n8467), .ZN(n8469) );
  INV_X1 U11062 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U11063 ( .A1(n8459), .A2(n8458), .ZN(n8460) );
  NAND2_X1 U11064 ( .A1(n8482), .A2(n8460), .ZN(n13749) );
  INV_X1 U11065 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13748) );
  NAND2_X1 U11066 ( .A1(n6947), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U11067 ( .A1(n6967), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8461) );
  OAI211_X1 U11068 ( .C1(n8708), .C2(n13748), .A(n8462), .B(n8461), .ZN(n8463)
         );
  INV_X1 U11069 ( .A(n8463), .ZN(n8464) );
  AND2_X1 U11070 ( .A1(n13760), .A2(n13974), .ZN(n8466) );
  INV_X1 U11071 ( .A(n8466), .ZN(n8468) );
  AOI21_X1 U11072 ( .B1(n8469), .B2(n8468), .A(n8535), .ZN(n9204) );
  INV_X1 U11073 ( .A(SI_27_), .ZN(n13515) );
  NAND2_X1 U11074 ( .A1(n8473), .A2(n13515), .ZN(n8472) );
  INV_X1 U11075 ( .A(n8470), .ZN(n8471) );
  INV_X1 U11076 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12609) );
  INV_X1 U11077 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14179) );
  MUX2_X1 U11078 ( .A(n12609), .B(n14179), .S(n10436), .Z(n8475) );
  INV_X1 U11079 ( .A(SI_28_), .ZN(n13512) );
  NAND2_X1 U11080 ( .A1(n8475), .A2(n13512), .ZN(n8681) );
  INV_X1 U11081 ( .A(n8475), .ZN(n8476) );
  NAND2_X1 U11082 ( .A1(n8476), .A2(SI_28_), .ZN(n8477) );
  NAND2_X1 U11083 ( .A1(n8681), .A2(n8477), .ZN(n8682) );
  OR2_X1 U11084 ( .A1(n8719), .A2(n14179), .ZN(n8478) );
  INV_X1 U11085 ( .A(n8482), .ZN(n8480) );
  INV_X1 U11086 ( .A(n13729), .ZN(n8484) );
  INV_X1 U11087 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U11088 ( .A1(n8482), .A2(n8481), .ZN(n8483) );
  NAND2_X1 U11089 ( .A1(n9190), .A2(n8282), .ZN(n8489) );
  NAND2_X1 U11090 ( .A1(n8002), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8485) );
  OAI211_X1 U11091 ( .C1(n9093), .C2(n8018), .A(n8486), .B(n8485), .ZN(n8487)
         );
  INV_X1 U11092 ( .A(n8487), .ZN(n8488) );
  NAND2_X1 U11093 ( .A1(n13742), .A2(n13974), .ZN(n8491) );
  XNOR2_X1 U11094 ( .A(n8491), .B(n8490), .ZN(n8492) );
  XNOR2_X1 U11095 ( .A(n13720), .B(n8492), .ZN(n8554) );
  INV_X1 U11096 ( .A(n8554), .ZN(n8534) );
  INV_X1 U11097 ( .A(n8501), .ZN(n8496) );
  NAND2_X1 U11098 ( .A1(n8496), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U11099 ( .A1(n8517), .A2(n8516), .ZN(n8497) );
  NAND2_X1 U11100 ( .A1(n8497), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8499) );
  INV_X1 U11101 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8498) );
  XNOR2_X1 U11102 ( .A(n8499), .B(n8498), .ZN(n12210) );
  XNOR2_X1 U11103 ( .A(n12210), .B(P2_B_REG_SCAN_IN), .ZN(n8505) );
  NOR2_X1 U11104 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8500) );
  NAND2_X1 U11105 ( .A1(n8501), .A2(n8500), .ZN(n8503) );
  NAND2_X1 U11106 ( .A1(n8503), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8502) );
  MUX2_X1 U11107 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8502), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8504) );
  NAND2_X1 U11108 ( .A1(n8504), .A2(n8506), .ZN(n12321) );
  NAND2_X1 U11109 ( .A1(n8505), .A2(n12321), .ZN(n8511) );
  NAND2_X1 U11110 ( .A1(n8506), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8507) );
  MUX2_X1 U11111 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8507), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8510) );
  INV_X1 U11112 ( .A(n8508), .ZN(n8509) );
  NAND2_X1 U11113 ( .A1(n8510), .A2(n8509), .ZN(n14186) );
  INV_X1 U11114 ( .A(n14186), .ZN(n8515) );
  INV_X1 U11115 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15528) );
  NAND2_X1 U11116 ( .A1(n15524), .A2(n15528), .ZN(n8513) );
  NAND2_X1 U11117 ( .A1(n14186), .A2(n12210), .ZN(n8512) );
  NAND2_X1 U11118 ( .A1(n8513), .A2(n8512), .ZN(n15529) );
  INV_X1 U11119 ( .A(n15529), .ZN(n9213) );
  NOR2_X1 U11120 ( .A1(n12321), .A2(n12210), .ZN(n8514) );
  NAND2_X1 U11121 ( .A1(n8515), .A2(n8514), .ZN(n10496) );
  XNOR2_X1 U11122 ( .A(n8517), .B(n8516), .ZN(n10490) );
  NAND2_X1 U11123 ( .A1(n9213), .A2(n15533), .ZN(n8531) );
  INV_X1 U11124 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15531) );
  NAND2_X1 U11125 ( .A1(n15524), .A2(n15531), .ZN(n8519) );
  NAND2_X1 U11126 ( .A1(n14186), .A2(n12321), .ZN(n8518) );
  NAND2_X1 U11127 ( .A1(n8519), .A2(n8518), .ZN(n15532) );
  INV_X1 U11128 ( .A(n15532), .ZN(n8530) );
  NOR4_X1 U11129 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8523) );
  NOR4_X1 U11130 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8522) );
  NOR4_X1 U11131 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8521) );
  NOR4_X1 U11132 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8520) );
  NAND4_X1 U11133 ( .A1(n8523), .A2(n8522), .A3(n8521), .A4(n8520), .ZN(n8529)
         );
  NOR2_X1 U11134 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n8527) );
  NOR4_X1 U11135 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n8526) );
  NOR4_X1 U11136 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8525) );
  NOR4_X1 U11137 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8524) );
  NAND4_X1 U11138 ( .A1(n8527), .A2(n8526), .A3(n8525), .A4(n8524), .ZN(n8528)
         );
  OAI21_X1 U11139 ( .B1(n8529), .B2(n8528), .A(n15524), .ZN(n9092) );
  NAND2_X1 U11140 ( .A1(n8530), .A2(n9092), .ZN(n9191) );
  NAND2_X1 U11141 ( .A1(n12562), .A2(n11614), .ZN(n8777) );
  INV_X1 U11142 ( .A(n8777), .ZN(n8815) );
  INV_X1 U11143 ( .A(n8536), .ZN(n10584) );
  OR2_X1 U11144 ( .A1(n8815), .A2(n10584), .ZN(n15536) );
  INV_X1 U11145 ( .A(n9039), .ZN(n11915) );
  INV_X1 U11146 ( .A(n10491), .ZN(n8532) );
  NAND2_X1 U11147 ( .A1(n15536), .A2(n8532), .ZN(n8533) );
  NOR2_X2 U11148 ( .A1(n8540), .A2(n8533), .ZN(n13610) );
  NAND2_X1 U11149 ( .A1(n8534), .A2(n13610), .ZN(n8559) );
  INV_X1 U11150 ( .A(n8535), .ZN(n8553) );
  INV_X1 U11151 ( .A(n8540), .ZN(n8537) );
  INV_X1 U11152 ( .A(n12562), .ZN(n8792) );
  AND2_X1 U11153 ( .A1(n8536), .A2(n8792), .ZN(n9196) );
  NAND2_X1 U11154 ( .A1(n8537), .A2(n9196), .ZN(n8539) );
  INV_X1 U11155 ( .A(n9091), .ZN(n8538) );
  NAND2_X1 U11156 ( .A1(n8539), .A2(n13956), .ZN(n13647) );
  INV_X1 U11157 ( .A(n13643), .ZN(n13616) );
  INV_X1 U11158 ( .A(n8541), .ZN(n8542) );
  OAI21_X1 U11159 ( .B1(n9191), .B2(n15529), .A(n9091), .ZN(n8545) );
  NAND2_X1 U11160 ( .A1(n10491), .A2(n8777), .ZN(n9090) );
  AND2_X1 U11161 ( .A1(n8543), .A2(n9090), .ZN(n8544) );
  NAND2_X1 U11162 ( .A1(n8545), .A2(n8544), .ZN(n10631) );
  AOI22_X1 U11163 ( .A1(n9190), .A2(n13631), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n8552) );
  NAND2_X1 U11164 ( .A1(n13729), .A2(n8282), .ZN(n8550) );
  INV_X1 U11165 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10825) );
  NAND2_X1 U11166 ( .A1(n8002), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8546) );
  OAI211_X1 U11167 ( .C1(n8018), .C2(n10825), .A(n8547), .B(n8546), .ZN(n8548)
         );
  INV_X1 U11168 ( .A(n8548), .ZN(n8549) );
  NAND2_X1 U11169 ( .A1(n8550), .A2(n8549), .ZN(n13653) );
  AND2_X1 U11170 ( .A1(n8541), .A2(n10491), .ZN(n13968) );
  NAND2_X1 U11171 ( .A1(n13653), .A2(n13568), .ZN(n8551) );
  OAI211_X1 U11172 ( .C1(n13635), .C2(n13623), .A(n8552), .B(n8551), .ZN(n8556) );
  NOR3_X1 U11173 ( .A1(n8554), .A2(n8553), .A3(n13649), .ZN(n8555) );
  AOI211_X1 U11174 ( .C1(n13720), .C2(n13647), .A(n8556), .B(n8555), .ZN(n8557) );
  OAI211_X1 U11175 ( .C1(n9203), .C2(n8559), .A(n8558), .B(n8557), .ZN(
        P2_U3192) );
  AOI21_X1 U11176 ( .B1(n13705), .B2(n9039), .A(n8779), .ZN(n8561) );
  AOI21_X1 U11177 ( .B1(n10637), .B2(n8726), .A(n8561), .ZN(n8565) );
  NAND2_X1 U11178 ( .A1(n10637), .A2(n8561), .ZN(n8564) );
  OAI211_X1 U11179 ( .C1(n13673), .C2(n8565), .A(n8564), .B(n8563), .ZN(n8569)
         );
  OAI22_X1 U11180 ( .A1(n12120), .A2(n8707), .B1(n8567), .B2(n8650), .ZN(n8570) );
  OAI22_X1 U11181 ( .A1(n11251), .A2(n8707), .B1(n15537), .B2(n8650), .ZN(
        n8575) );
  AND2_X1 U11182 ( .A1(n12126), .A2(n8650), .ZN(n8566) );
  OAI22_X1 U11183 ( .A1(n8569), .A2(n8570), .B1(n8575), .B2(n8574), .ZN(n8578)
         );
  AOI22_X1 U11184 ( .A1(n13672), .A2(n8726), .B1(n8650), .B2(n6645), .ZN(n8568) );
  AOI21_X1 U11185 ( .B1(n8570), .B2(n8569), .A(n8568), .ZN(n8577) );
  NAND2_X1 U11186 ( .A1(n13671), .A2(n8650), .ZN(n8573) );
  NAND2_X1 U11187 ( .A1(n8571), .A2(n8707), .ZN(n8572) );
  NAND2_X1 U11188 ( .A1(n8573), .A2(n8572), .ZN(n8585) );
  AOI22_X1 U11189 ( .A1(n8575), .A2(n8574), .B1(n8584), .B2(n8585), .ZN(n8576)
         );
  NAND2_X1 U11190 ( .A1(n13670), .A2(n8650), .ZN(n8581) );
  NAND2_X1 U11191 ( .A1(n6432), .A2(n8579), .ZN(n8580) );
  NAND2_X1 U11192 ( .A1(n8581), .A2(n8580), .ZN(n8590) );
  AND2_X1 U11193 ( .A1(n6432), .A2(n8650), .ZN(n8583) );
  NAND2_X1 U11194 ( .A1(n13669), .A2(n8726), .ZN(n8589) );
  NAND2_X1 U11195 ( .A1(n12038), .A2(n8650), .ZN(n8588) );
  NAND2_X1 U11196 ( .A1(n8589), .A2(n8588), .ZN(n8593) );
  NAND2_X1 U11197 ( .A1(n8591), .A2(n8590), .ZN(n8592) );
  OAI22_X1 U11198 ( .A1(n12046), .A2(n8707), .B1(n11312), .B2(n8770), .ZN(
        n8597) );
  OAI22_X1 U11199 ( .A1(n11999), .A2(n8707), .B1(n11475), .B2(n8650), .ZN(
        n8599) );
  OAI22_X1 U11200 ( .A1(n8598), .A2(n8597), .B1(n8600), .B2(n8599), .ZN(n8603)
         );
  AOI22_X1 U11201 ( .A1(n15543), .A2(n8707), .B1(n13668), .B2(n8770), .ZN(
        n8596) );
  AOI21_X1 U11202 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(n8602) );
  INV_X1 U11203 ( .A(n8599), .ZN(n8601) );
  OAI22_X1 U11204 ( .A1(n12015), .A2(n8726), .B1(n11702), .B2(n8770), .ZN(
        n8604) );
  NAND2_X1 U11205 ( .A1(n8605), .A2(n8604), .ZN(n8608) );
  INV_X1 U11206 ( .A(n11702), .ZN(n13665) );
  AOI22_X1 U11207 ( .A1(n14111), .A2(n8707), .B1(n8770), .B2(n13665), .ZN(
        n8606) );
  NAND2_X1 U11208 ( .A1(n8608), .A2(n8607), .ZN(n8609) );
  OAI22_X1 U11209 ( .A1(n11984), .A2(n8650), .B1(n11754), .B2(n8726), .ZN(
        n8611) );
  AOI22_X1 U11210 ( .A1(n14106), .A2(n8770), .B1(n13664), .B2(n8726), .ZN(
        n8610) );
  OAI22_X1 U11211 ( .A1(n12110), .A2(n8707), .B1(n12168), .B2(n8650), .ZN(
        n8613) );
  INV_X1 U11212 ( .A(n12168), .ZN(n13663) );
  AOI22_X1 U11213 ( .A1(n9020), .A2(n8707), .B1(n8770), .B2(n13663), .ZN(n8612) );
  OAI22_X1 U11214 ( .A1(n14161), .A2(n8770), .B1(n12195), .B2(n8707), .ZN(
        n8619) );
  INV_X1 U11215 ( .A(n12195), .ZN(n13662) );
  AOI22_X1 U11216 ( .A1(n12171), .A2(n8770), .B1(n13662), .B2(n8707), .ZN(
        n8615) );
  NAND2_X1 U11217 ( .A1(n8617), .A2(n8616), .ZN(n8623) );
  INV_X1 U11218 ( .A(n8618), .ZN(n8621) );
  INV_X1 U11219 ( .A(n8619), .ZN(n8620) );
  NAND2_X1 U11220 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  OAI22_X1 U11221 ( .A1(n12282), .A2(n8707), .B1(n12295), .B2(n8770), .ZN(
        n8626) );
  AOI22_X1 U11222 ( .A1(n14089), .A2(n8707), .B1(n8770), .B2(n13967), .ZN(
        n8628) );
  INV_X1 U11223 ( .A(n14089), .ZN(n12303) );
  INV_X1 U11224 ( .A(n13967), .ZN(n13530) );
  OAI22_X1 U11225 ( .A1(n12303), .A2(n8707), .B1(n13530), .B2(n8770), .ZN(
        n8627) );
  OAI22_X1 U11226 ( .A1(n13980), .A2(n8726), .B1(n13659), .B2(n8770), .ZN(
        n8629) );
  OAI22_X1 U11227 ( .A1(n13980), .A2(n8770), .B1(n13659), .B2(n8707), .ZN(
        n8631) );
  INV_X1 U11228 ( .A(n8629), .ZN(n8630) );
  INV_X1 U11229 ( .A(n13969), .ZN(n13931) );
  OAI22_X1 U11230 ( .A1(n7172), .A2(n8707), .B1(n13931), .B2(n8770), .ZN(n8632) );
  NAND2_X1 U11231 ( .A1(n8634), .A2(n8633), .ZN(n8635) );
  NAND2_X1 U11232 ( .A1(n8636), .A2(n8635), .ZN(n8637) );
  OAI22_X1 U11233 ( .A1(n13941), .A2(n8707), .B1(n13641), .B2(n8650), .ZN(
        n8638) );
  NAND2_X1 U11234 ( .A1(n8637), .A2(n8638), .ZN(n8642) );
  INV_X1 U11235 ( .A(n8637), .ZN(n8640) );
  INV_X1 U11236 ( .A(n8638), .ZN(n8639) );
  AOI22_X1 U11237 ( .A1(n13920), .A2(n8770), .B1(n13893), .B2(n8707), .ZN(
        n8643) );
  INV_X1 U11238 ( .A(n8643), .ZN(n8644) );
  INV_X1 U11239 ( .A(n8648), .ZN(n8649) );
  OAI22_X1 U11240 ( .A1(n13882), .A2(n8650), .B1(n13859), .B2(n8707), .ZN(
        n8651) );
  OAI22_X1 U11241 ( .A1(n13882), .A2(n8726), .B1(n13859), .B2(n8770), .ZN(
        n8652) );
  AOI22_X1 U11242 ( .A1(n14140), .A2(n8770), .B1(n13656), .B2(n8707), .ZN(
        n8655) );
  AOI22_X1 U11243 ( .A1(n14140), .A2(n8707), .B1(n8770), .B2(n13656), .ZN(
        n8653) );
  INV_X1 U11244 ( .A(n8653), .ZN(n8654) );
  OAI22_X1 U11245 ( .A1(n14137), .A2(n8770), .B1(n13860), .B2(n8707), .ZN(
        n8658) );
  AOI22_X1 U11246 ( .A1(n7410), .A2(n8770), .B1(n13655), .B2(n8726), .ZN(n8657) );
  OAI22_X1 U11247 ( .A1(n14133), .A2(n8707), .B1(n13843), .B2(n8770), .ZN(
        n8660) );
  INV_X1 U11248 ( .A(n13843), .ZN(n13654) );
  AOI22_X1 U11249 ( .A1(n13831), .A2(n8707), .B1(n8770), .B2(n13654), .ZN(
        n8659) );
  AND2_X1 U11250 ( .A1(n13794), .A2(n8770), .ZN(n8662) );
  AOI21_X1 U11251 ( .B1(n13541), .B2(n8707), .A(n8662), .ZN(n8754) );
  NAND2_X1 U11252 ( .A1(n13541), .A2(n8770), .ZN(n8664) );
  NAND2_X1 U11253 ( .A1(n13794), .A2(n8726), .ZN(n8663) );
  NAND2_X1 U11254 ( .A1(n8664), .A2(n8663), .ZN(n8753) );
  AND2_X1 U11255 ( .A1(n13760), .A2(n8707), .ZN(n8665) );
  AOI21_X1 U11256 ( .B1(n13751), .B2(n8770), .A(n8665), .ZN(n8730) );
  NAND2_X1 U11257 ( .A1(n13751), .A2(n8707), .ZN(n8667) );
  NAND2_X1 U11258 ( .A1(n13760), .A2(n8770), .ZN(n8666) );
  NAND2_X1 U11259 ( .A1(n8667), .A2(n8666), .ZN(n8740) );
  AND2_X1 U11260 ( .A1(n13773), .A2(n8770), .ZN(n8668) );
  NAND2_X1 U11261 ( .A1(n14026), .A2(n8770), .ZN(n8670) );
  NAND2_X1 U11262 ( .A1(n13773), .A2(n8707), .ZN(n8669) );
  NAND2_X1 U11263 ( .A1(n8670), .A2(n8669), .ZN(n8734) );
  AND2_X1 U11264 ( .A1(n13795), .A2(n8770), .ZN(n8671) );
  AOI21_X1 U11265 ( .B1(n13784), .B2(n8726), .A(n8671), .ZN(n8733) );
  NAND2_X1 U11266 ( .A1(n13784), .A2(n8770), .ZN(n8673) );
  NAND2_X1 U11267 ( .A1(n13795), .A2(n8707), .ZN(n8672) );
  NAND2_X1 U11268 ( .A1(n8673), .A2(n8672), .ZN(n8732) );
  OAI22_X1 U11269 ( .A1(n8731), .A2(n8734), .B1(n8733), .B2(n8732), .ZN(n8674)
         );
  AOI21_X1 U11270 ( .B1(n8730), .B2(n8740), .A(n8674), .ZN(n8745) );
  AND2_X1 U11271 ( .A1(n13810), .A2(n8726), .ZN(n8675) );
  AOI21_X1 U11272 ( .B1(n14036), .B2(n8770), .A(n8675), .ZN(n8747) );
  NAND2_X1 U11273 ( .A1(n14036), .A2(n8707), .ZN(n8677) );
  NAND2_X1 U11274 ( .A1(n13810), .A2(n8770), .ZN(n8676) );
  NAND2_X1 U11275 ( .A1(n8677), .A2(n8676), .ZN(n8746) );
  NAND2_X1 U11276 ( .A1(n8747), .A2(n8746), .ZN(n8678) );
  OAI21_X1 U11277 ( .B1(n8754), .B2(n8753), .A(n8752), .ZN(n8679) );
  INV_X1 U11278 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15182) );
  INV_X1 U11279 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14173) );
  MUX2_X1 U11280 ( .A(n15182), .B(n14173), .S(n10436), .Z(n8684) );
  XNOR2_X1 U11281 ( .A(n8684), .B(SI_29_), .ZN(n8716) );
  INV_X1 U11282 ( .A(SI_29_), .ZN(n13509) );
  NAND2_X1 U11283 ( .A1(n8684), .A2(n13509), .ZN(n8685) );
  MUX2_X1 U11284 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10436), .Z(n8686) );
  NAND2_X1 U11285 ( .A1(n8686), .A2(SI_30_), .ZN(n8687) );
  OAI21_X1 U11286 ( .B1(SI_30_), .B2(n8686), .A(n8687), .ZN(n8700) );
  MUX2_X1 U11287 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10436), .Z(n8688) );
  XNOR2_X1 U11288 ( .A(n8688), .B(SI_31_), .ZN(n8689) );
  NAND2_X1 U11289 ( .A1(n14164), .A2(n8718), .ZN(n8693) );
  NAND2_X1 U11290 ( .A1(n8691), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8692) );
  INV_X1 U11291 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8694) );
  OR2_X1 U11292 ( .A1(n8018), .A2(n8694), .ZN(n8698) );
  INV_X1 U11293 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n10827) );
  OR2_X1 U11294 ( .A1(n8708), .A2(n10827), .ZN(n8697) );
  INV_X1 U11295 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8695) );
  OR2_X1 U11296 ( .A1(n7019), .A2(n8695), .ZN(n8696) );
  AND3_X1 U11297 ( .A1(n8698), .A2(n8697), .A3(n8696), .ZN(n8705) );
  NAND2_X1 U11298 ( .A1(n12577), .A2(n8705), .ZN(n8771) );
  OR2_X1 U11299 ( .A1(n12577), .A2(n8705), .ZN(n8699) );
  NAND2_X1 U11300 ( .A1(n12403), .A2(n8718), .ZN(n8704) );
  INV_X1 U11301 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12583) );
  OR2_X1 U11302 ( .A1(n8719), .A2(n12583), .ZN(n8703) );
  INV_X1 U11303 ( .A(n8705), .ZN(n13651) );
  NAND2_X1 U11304 ( .A1(n11915), .A2(n13705), .ZN(n9084) );
  OAI211_X1 U11305 ( .C1(n9084), .C2(n8792), .A(n8776), .B(n8777), .ZN(n8706)
         );
  AOI21_X1 U11306 ( .B1(n13651), .B2(n8707), .A(n8706), .ZN(n8712) );
  INV_X1 U11307 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14002) );
  OR2_X1 U11308 ( .A1(n8018), .A2(n14002), .ZN(n8711) );
  INV_X1 U11309 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13713) );
  OR2_X1 U11310 ( .A1(n8708), .A2(n13713), .ZN(n8710) );
  INV_X1 U11311 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14118) );
  OR2_X1 U11312 ( .A1(n7019), .A2(n14118), .ZN(n8709) );
  AND3_X1 U11313 ( .A1(n8711), .A2(n8710), .A3(n8709), .ZN(n13722) );
  NOR2_X1 U11314 ( .A1(n8712), .A2(n13722), .ZN(n8713) );
  AOI21_X1 U11315 ( .B1(n13999), .B2(n8770), .A(n8713), .ZN(n8766) );
  NAND2_X1 U11316 ( .A1(n13999), .A2(n8579), .ZN(n8715) );
  INV_X1 U11317 ( .A(n13722), .ZN(n13652) );
  NAND2_X1 U11318 ( .A1(n13652), .A2(n8770), .ZN(n8714) );
  NAND2_X1 U11319 ( .A1(n8715), .A2(n8714), .ZN(n8765) );
  NAND2_X1 U11320 ( .A1(n14172), .A2(n8718), .ZN(n8721) );
  OR2_X1 U11321 ( .A1(n8719), .A2(n14173), .ZN(n8720) );
  AND2_X1 U11322 ( .A1(n13653), .A2(n8707), .ZN(n8722) );
  AOI21_X1 U11323 ( .B1(n14016), .B2(n8770), .A(n8722), .ZN(n8763) );
  NAND2_X1 U11324 ( .A1(n14016), .A2(n8707), .ZN(n8724) );
  NAND2_X1 U11325 ( .A1(n13653), .A2(n8770), .ZN(n8723) );
  NAND2_X1 U11326 ( .A1(n8724), .A2(n8723), .ZN(n8762) );
  OAI22_X1 U11327 ( .A1(n8766), .A2(n8765), .B1(n8763), .B2(n8762), .ZN(n8725)
         );
  AND2_X1 U11328 ( .A1(n13742), .A2(n8726), .ZN(n8727) );
  AOI21_X1 U11329 ( .B1(n13720), .B2(n8770), .A(n8727), .ZN(n8761) );
  NAND2_X1 U11330 ( .A1(n13720), .A2(n8707), .ZN(n8729) );
  NAND2_X1 U11331 ( .A1(n13742), .A2(n8770), .ZN(n8728) );
  NAND2_X1 U11332 ( .A1(n8729), .A2(n8728), .ZN(n8760) );
  INV_X1 U11333 ( .A(n8730), .ZN(n8742) );
  INV_X1 U11334 ( .A(n8731), .ZN(n8737) );
  NAND2_X1 U11335 ( .A1(n8733), .A2(n8732), .ZN(n8736) );
  NAND2_X1 U11336 ( .A1(n8737), .A2(n8736), .ZN(n8735) );
  NAND2_X1 U11337 ( .A1(n8735), .A2(n8734), .ZN(n8739) );
  OR2_X1 U11338 ( .A1(n8737), .A2(n8736), .ZN(n8738) );
  NAND2_X1 U11339 ( .A1(n8739), .A2(n8738), .ZN(n8741) );
  OR2_X1 U11340 ( .A1(n8742), .A2(n8741), .ZN(n8744) );
  INV_X1 U11341 ( .A(n8740), .ZN(n8743) );
  AOI22_X1 U11342 ( .A1(n8744), .A2(n8743), .B1(n8742), .B2(n8741), .ZN(n8750)
         );
  INV_X1 U11343 ( .A(n8745), .ZN(n8748) );
  OR3_X1 U11344 ( .A1(n8748), .A2(n8747), .A3(n8746), .ZN(n8749) );
  OAI211_X1 U11345 ( .C1(n8761), .C2(n8760), .A(n8750), .B(n8749), .ZN(n8751)
         );
  INV_X1 U11346 ( .A(n8751), .ZN(n8759) );
  INV_X1 U11347 ( .A(n8752), .ZN(n8757) );
  INV_X1 U11348 ( .A(n8753), .ZN(n8756) );
  INV_X1 U11349 ( .A(n8754), .ZN(n8755) );
  AOI22_X1 U11350 ( .A1(n8763), .A2(n8762), .B1(n8761), .B2(n8760), .ZN(n8764)
         );
  NAND2_X1 U11351 ( .A1(n8783), .A2(n8764), .ZN(n8767) );
  AOI22_X1 U11352 ( .A1(n8768), .A2(n8767), .B1(n8766), .B2(n8765), .ZN(n8773)
         );
  NAND2_X1 U11353 ( .A1(n13651), .A2(n8770), .ZN(n8769) );
  OAI22_X1 U11354 ( .A1(n8771), .A2(n8770), .B1(n8769), .B2(n12577), .ZN(n8772) );
  MUX2_X1 U11355 ( .A(n9039), .B(n11770), .S(n8792), .Z(n8774) );
  NAND2_X1 U11356 ( .A1(n8775), .A2(n7819), .ZN(n8782) );
  NAND2_X1 U11357 ( .A1(n8776), .A2(n11614), .ZN(n8778) );
  OAI211_X1 U11358 ( .C1(n8779), .C2(n11915), .A(n8778), .B(n8777), .ZN(n8780)
         );
  INV_X1 U11359 ( .A(n10490), .ZN(n10495) );
  AND2_X1 U11360 ( .A1(n10495), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12105) );
  INV_X1 U11361 ( .A(n8783), .ZN(n8810) );
  XNOR2_X1 U11362 ( .A(n13999), .B(n13652), .ZN(n8808) );
  NAND2_X1 U11363 ( .A1(n13720), .A2(n13723), .ZN(n8784) );
  NAND2_X1 U11364 ( .A1(n14026), .A2(n13744), .ZN(n13739) );
  NAND2_X1 U11365 ( .A1(n13739), .A2(n8785), .ZN(n9081) );
  INV_X1 U11366 ( .A(n13795), .ZN(n13594) );
  NAND2_X1 U11367 ( .A1(n13784), .A2(n13594), .ZN(n9080) );
  OR2_X1 U11368 ( .A1(n13784), .A2(n13594), .ZN(n8786) );
  NAND2_X1 U11369 ( .A1(n14036), .A2(n13775), .ZN(n9079) );
  OR2_X1 U11370 ( .A1(n14036), .A2(n13775), .ZN(n8787) );
  NAND2_X1 U11371 ( .A1(n13831), .A2(n13843), .ZN(n9072) );
  INV_X1 U11372 ( .A(n13656), .ZN(n13842) );
  NAND2_X1 U11373 ( .A1(n14140), .A2(n13842), .ZN(n13839) );
  OR2_X1 U11374 ( .A1(n14140), .A2(n13842), .ZN(n8788) );
  NAND2_X1 U11375 ( .A1(n13839), .A2(n8788), .ZN(n13871) );
  NAND2_X1 U11376 ( .A1(n14084), .A2(n13659), .ZN(n9063) );
  NAND2_X1 U11377 ( .A1(n9063), .A2(n8789), .ZN(n13982) );
  INV_X1 U11378 ( .A(n12295), .ZN(n13661) );
  OR2_X1 U11379 ( .A1(n14154), .A2(n13661), .ZN(n9024) );
  NAND2_X1 U11380 ( .A1(n14154), .A2(n13661), .ZN(n9023) );
  NAND2_X1 U11381 ( .A1(n9024), .A2(n9023), .ZN(n12276) );
  INV_X1 U11382 ( .A(n11251), .ZN(n8790) );
  NAND2_X1 U11383 ( .A1(n13673), .A2(n11353), .ZN(n10634) );
  AND2_X1 U11384 ( .A1(n11355), .A2(n10634), .ZN(n10582) );
  NAND4_X1 U11385 ( .A1(n11241), .A2(n10582), .A3(n8792), .A4(n11350), .ZN(
        n8794) );
  NAND2_X1 U11386 ( .A1(n12036), .A2(n12038), .ZN(n9049) );
  NAND2_X1 U11387 ( .A1(n13669), .A2(n11318), .ZN(n8793) );
  NOR3_X1 U11388 ( .A1(n8794), .A2(n11249), .A3(n11309), .ZN(n8795) );
  XNOR2_X1 U11389 ( .A(n15552), .B(n13666), .ZN(n11992) );
  XNOR2_X1 U11390 ( .A(n13670), .B(n6432), .ZN(n11307) );
  XNOR2_X1 U11391 ( .A(n15543), .B(n13668), .ZN(n12048) );
  NAND4_X1 U11392 ( .A1(n8795), .A2(n11992), .A3(n11307), .A4(n12048), .ZN(
        n8796) );
  XNOR2_X1 U11393 ( .A(n14111), .B(n11702), .ZN(n12004) );
  NOR2_X1 U11394 ( .A1(n8796), .A2(n12004), .ZN(n8797) );
  XNOR2_X1 U11395 ( .A(n12171), .B(n13662), .ZN(n12161) );
  XNOR2_X1 U11396 ( .A(n14106), .B(n13664), .ZN(n11976) );
  NAND4_X1 U11397 ( .A1(n12276), .A2(n8797), .A3(n12161), .A4(n11976), .ZN(
        n8798) );
  XNOR2_X1 U11398 ( .A(n14089), .B(n13530), .ZN(n12304) );
  XNOR2_X1 U11399 ( .A(n9020), .B(n12168), .ZN(n11969) );
  OR3_X1 U11400 ( .A1(n8798), .A2(n12304), .A3(n11969), .ZN(n8799) );
  NOR2_X1 U11401 ( .A1(n13982), .A2(n8799), .ZN(n8800) );
  XNOR2_X1 U11402 ( .A(n13955), .B(n13969), .ZN(n13947) );
  XNOR2_X1 U11403 ( .A(n14074), .B(n13658), .ZN(n9066) );
  NAND4_X1 U11404 ( .A1(n13913), .A2(n8800), .A3(n13947), .A4(n9066), .ZN(
        n8801) );
  NOR2_X1 U11405 ( .A1(n13871), .A2(n8801), .ZN(n8802) );
  INV_X1 U11406 ( .A(n13859), .ZN(n13894) );
  XNOR2_X1 U11407 ( .A(n14059), .B(n13894), .ZN(n13883) );
  XNOR2_X1 U11408 ( .A(n14064), .B(n13657), .ZN(n13892) );
  NAND4_X1 U11409 ( .A1(n13826), .A2(n8802), .A3(n13883), .A4(n13892), .ZN(
        n8803) );
  NOR2_X1 U11410 ( .A1(n13802), .A2(n8803), .ZN(n8804) );
  XNOR2_X1 U11411 ( .A(n13541), .B(n13794), .ZN(n13806) );
  NAND4_X1 U11412 ( .A1(n13772), .A2(n8804), .A3(n13806), .A4(n13838), .ZN(
        n8805) );
  NOR2_X1 U11413 ( .A1(n9081), .A2(n8805), .ZN(n8806) );
  AND2_X1 U11414 ( .A1(n13737), .A2(n8806), .ZN(n8807) );
  NAND4_X1 U11415 ( .A1(n8808), .A2(n14008), .A3(n8807), .A4(n14011), .ZN(
        n8809) );
  NAND3_X1 U11416 ( .A1(n12105), .A2(n13705), .A3(n11770), .ZN(n8811) );
  NAND4_X1 U11417 ( .A1(n8814), .A2(n12105), .A3(n11614), .A4(n11770), .ZN(
        n8818) );
  INV_X1 U11418 ( .A(n14181), .ZN(n12571) );
  NAND4_X1 U11419 ( .A1(n15533), .A2(n12571), .A3(n13966), .A4(n8815), .ZN(
        n8816) );
  OAI211_X1 U11420 ( .C1(n11915), .C2(n8781), .A(n8816), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8817) );
  NOR2_X1 U11421 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8823) );
  NOR2_X1 U11422 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n8822) );
  NOR2_X1 U11423 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n8821) );
  INV_X1 U11424 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8825) );
  OR2_X1 U11425 ( .A1(n8859), .A2(n10453), .ZN(n8833) );
  NAND2_X1 U11426 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n15193), .ZN(n8830) );
  OR2_X1 U11427 ( .A1(n8843), .A2(n14654), .ZN(n8832) );
  NAND3_X2 U11428 ( .A1(n8834), .A2(n8833), .A3(n8832), .ZN(n11370) );
  INV_X1 U11429 ( .A(n15193), .ZN(n15293) );
  INV_X1 U11430 ( .A(SI_0_), .ZN(n8835) );
  INV_X1 U11431 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9751) );
  OAI21_X1 U11432 ( .B1(n10436), .B2(n8835), .A(n9751), .ZN(n8836) );
  NAND2_X1 U11433 ( .A1(n8837), .A2(n8836), .ZN(n15192) );
  MUX2_X1 U11434 ( .A(n15293), .B(n15192), .S(n8843), .Z(n11378) );
  INV_X1 U11435 ( .A(n11378), .ZN(n11453) );
  INV_X1 U11436 ( .A(n8845), .ZN(n8838) );
  NOR2_X2 U11437 ( .A1(n15332), .A2(n15330), .ZN(n11375) );
  OR2_X1 U11438 ( .A1(n8845), .A2(n8827), .ZN(n8840) );
  OR2_X1 U11439 ( .A1(n8859), .A2(n10442), .ZN(n8842) );
  OR2_X1 U11440 ( .A1(n8949), .A2(n10443), .ZN(n8841) );
  INV_X1 U11441 ( .A(n8859), .ZN(n8856) );
  NAND2_X1 U11442 ( .A1(n8856), .A2(n10408), .ZN(n8850) );
  NAND2_X1 U11443 ( .A1(n8845), .A2(n8844), .ZN(n8905) );
  NAND2_X1 U11444 ( .A1(n8905), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8846) );
  MUX2_X1 U11445 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8846), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n8847) );
  NAND2_X1 U11446 ( .A1(n8847), .A2(n8853), .ZN(n10617) );
  OR2_X1 U11447 ( .A1(n8843), .A2(n10617), .ZN(n8849) );
  INV_X1 U11448 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10447) );
  OR2_X1 U11449 ( .A1(n8949), .A2(n10447), .ZN(n8848) );
  NAND2_X1 U11450 ( .A1(n8853), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8852) );
  MUX2_X1 U11451 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8852), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n8855) );
  INV_X1 U11452 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U11453 ( .A1(n8855), .A2(n8863), .ZN(n10696) );
  INV_X1 U11454 ( .A(n10696), .ZN(n10611) );
  AOI22_X1 U11455 ( .A1(n8925), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10456), 
        .B2(n10611), .ZN(n8858) );
  NAND2_X1 U11456 ( .A1(n10410), .A2(n8856), .ZN(n8857) );
  NAND2_X1 U11457 ( .A1(n10417), .A2(n8856), .ZN(n8862) );
  NAND2_X1 U11458 ( .A1(n8863), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8860) );
  XNOR2_X1 U11459 ( .A(n8860), .B(P1_IR_REG_6__SCAN_IN), .ZN(n14724) );
  AOI22_X1 U11460 ( .A1(n8925), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10456), 
        .B2(n14724), .ZN(n8861) );
  NAND2_X1 U11461 ( .A1(n8862), .A2(n8861), .ZN(n14413) );
  INV_X1 U11462 ( .A(n14413), .ZN(n15364) );
  NAND2_X1 U11463 ( .A1(n10432), .A2(n8948), .ZN(n8868) );
  INV_X1 U11464 ( .A(n8863), .ZN(n8865) );
  INV_X1 U11465 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8864) );
  NAND2_X1 U11466 ( .A1(n8865), .A2(n8864), .ZN(n8869) );
  NAND2_X1 U11467 ( .A1(n8869), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8866) );
  XNOR2_X1 U11468 ( .A(n8866), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U11469 ( .A1(n8925), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10456), 
        .B2(n10697), .ZN(n8867) );
  INV_X1 U11470 ( .A(n14419), .ZN(n11689) );
  NAND2_X1 U11471 ( .A1(n11644), .A2(n11689), .ZN(n11686) );
  NAND2_X1 U11472 ( .A1(n10448), .A2(n8948), .ZN(n8871) );
  XNOR2_X1 U11473 ( .A(n8873), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U11474 ( .A1(n8925), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10456), 
        .B2(n10874), .ZN(n8870) );
  OR2_X2 U11475 ( .A1(n11686), .A2(n14424), .ZN(n12222) );
  NAND2_X1 U11476 ( .A1(n10469), .A2(n8948), .ZN(n8876) );
  INV_X1 U11477 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U11478 ( .A1(n8873), .A2(n8872), .ZN(n8874) );
  XNOR2_X1 U11479 ( .A(n8884), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U11480 ( .A1(n8925), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11102), 
        .B2(n10456), .ZN(n8875) );
  NAND2_X1 U11481 ( .A1(n10472), .A2(n8948), .ZN(n8881) );
  INV_X1 U11482 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U11483 ( .A1(n8884), .A2(n8877), .ZN(n8878) );
  NAND2_X1 U11484 ( .A1(n8878), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8879) );
  XNOR2_X1 U11485 ( .A(n8879), .B(P1_IR_REG_10__SCAN_IN), .ZN(n14739) );
  AOI22_X1 U11486 ( .A1(n14739), .A2(n10456), .B1(n8925), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11487 ( .A1(n10486), .A2(n8948), .ZN(n8887) );
  OR2_X1 U11488 ( .A1(n8882), .A2(n8827), .ZN(n8883) );
  NAND2_X1 U11489 ( .A1(n8884), .A2(n8883), .ZN(n8888) );
  XNOR2_X1 U11490 ( .A(n8888), .B(n8885), .ZN(n11289) );
  AOI22_X1 U11491 ( .A1(n11289), .A2(n10456), .B1(n8925), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U11492 ( .A1(n10578), .A2(n8948), .ZN(n8891) );
  XNOR2_X1 U11493 ( .A(n8893), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U11494 ( .A1(n11441), .A2(n10456), .B1(n8925), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11495 ( .A1(n10678), .A2(n8948), .ZN(n8898) );
  INV_X1 U11496 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U11497 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  NAND2_X1 U11498 ( .A1(n8894), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U11499 ( .A1(n8895), .A2(n7239), .ZN(n8899) );
  OR2_X1 U11500 ( .A1(n8895), .A2(n7239), .ZN(n8896) );
  AOI22_X1 U11501 ( .A1(n11711), .A2(n10456), .B1(n8925), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8897) );
  NAND2_X1 U11502 ( .A1(n11198), .A2(n8948), .ZN(n8902) );
  NAND2_X1 U11503 ( .A1(n8899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8900) );
  XNOR2_X1 U11504 ( .A(n8900), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U11505 ( .A1(n12347), .A2(n10456), .B1(n8925), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U11506 ( .A1(n8903), .A2(n8904), .ZN(n8906) );
  OR2_X1 U11507 ( .A1(n8906), .A2(n8905), .ZN(n8910) );
  NAND2_X1 U11508 ( .A1(n8910), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8907) );
  XNOR2_X1 U11509 ( .A(n8907), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U11510 ( .A1(n8925), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10456), 
        .B2(n12350), .ZN(n8908) );
  INV_X1 U11511 ( .A(n15146), .ZN(n14995) );
  NAND2_X1 U11512 ( .A1(n11297), .A2(n8948), .ZN(n8914) );
  OAI21_X1 U11513 ( .B1(n8910), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8911) );
  MUX2_X1 U11514 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8911), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8912) );
  NAND2_X1 U11515 ( .A1(n8912), .A2(n8916), .ZN(n12352) );
  INV_X1 U11516 ( .A(n12352), .ZN(n14749) );
  AOI22_X1 U11517 ( .A1(n8925), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10456), 
        .B2(n14749), .ZN(n8913) );
  NAND2_X1 U11518 ( .A1(n11365), .A2(n8948), .ZN(n8919) );
  NAND2_X1 U11519 ( .A1(n8916), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8915) );
  MUX2_X1 U11520 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8915), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n8917) );
  NAND2_X1 U11521 ( .A1(n8917), .A2(n6603), .ZN(n14762) );
  INV_X1 U11522 ( .A(n14762), .ZN(n14765) );
  AOI22_X1 U11523 ( .A1(n8925), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10456), 
        .B2(n14765), .ZN(n8918) );
  NAND2_X1 U11524 ( .A1(n11525), .A2(n8948), .ZN(n8922) );
  NAND2_X1 U11525 ( .A1(n6603), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8920) );
  XNOR2_X1 U11526 ( .A(n8920), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14779) );
  AOI22_X1 U11527 ( .A1(n8925), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10456), 
        .B2(n14779), .ZN(n8921) );
  XNOR2_X2 U11528 ( .A(n8924), .B(n8955), .ZN(n14958) );
  AOI22_X1 U11529 ( .A1(n8925), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14381), 
        .B2(n10456), .ZN(n8926) );
  INV_X1 U11530 ( .A(n15128), .ZN(n14931) );
  OR2_X1 U11531 ( .A1(n6952), .A2(n11710), .ZN(n8927) );
  NAND2_X1 U11532 ( .A1(n11769), .A2(n8948), .ZN(n8930) );
  INV_X1 U11533 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12566) );
  OR2_X1 U11534 ( .A1(n6952), .A2(n12566), .ZN(n8929) );
  OR2_X1 U11535 ( .A1(n6952), .A2(n12136), .ZN(n8933) );
  INV_X1 U11536 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12209) );
  OR2_X1 U11537 ( .A1(n6952), .A2(n12209), .ZN(n8935) );
  NAND2_X1 U11538 ( .A1(n12318), .A2(n8948), .ZN(n8938) );
  OR2_X1 U11539 ( .A1(n6952), .A2(n12320), .ZN(n8937) );
  NOR2_X4 U11540 ( .A1(n14839), .A2(n14829), .ZN(n14825) );
  NAND2_X1 U11541 ( .A1(n14183), .A2(n8948), .ZN(n8940) );
  OR2_X1 U11542 ( .A1(n6952), .A2(n15186), .ZN(n8939) );
  OR2_X1 U11543 ( .A1(n6952), .A2(n15184), .ZN(n8941) );
  OR2_X1 U11544 ( .A1(n6952), .A2(n12609), .ZN(n8943) );
  NAND2_X1 U11545 ( .A1(n14172), .A2(n8948), .ZN(n8946) );
  OR2_X1 U11546 ( .A1(n6952), .A2(n15182), .ZN(n8945) );
  INV_X1 U11547 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12584) );
  NOR2_X1 U11548 ( .A1(n6952), .A2(n12584), .ZN(n8947) );
  NAND2_X1 U11549 ( .A1(n14164), .A2(n8948), .ZN(n8951) );
  INV_X1 U11550 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15175) );
  OR2_X1 U11551 ( .A1(n6952), .A2(n15175), .ZN(n8950) );
  XNOR2_X1 U11552 ( .A(n14795), .B(n14624), .ZN(n8960) );
  INV_X1 U11553 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8956) );
  INV_X1 U11554 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10744) );
  INV_X1 U11555 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8952) );
  INV_X1 U11556 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8953) );
  AND2_X1 U11557 ( .A1(n14575), .A2(n11709), .ZN(n14535) );
  NAND2_X1 U11558 ( .A1(n8960), .A2(n15333), .ZN(n14794) );
  NAND2_X1 U11559 ( .A1(n14544), .A2(n14575), .ZN(n10721) );
  NAND2_X1 U11560 ( .A1(n11709), .A2(n14958), .ZN(n8987) );
  INV_X1 U11561 ( .A(n8987), .ZN(n8961) );
  INV_X1 U11562 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n15173) );
  INV_X1 U11563 ( .A(n8964), .ZN(n9220) );
  NAND2_X4 U11564 ( .A1(n9220), .A2(n15181), .ZN(n12508) );
  INV_X1 U11565 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14791) );
  AND2_X4 U11566 ( .A1(n12468), .A2(n8965), .ZN(n9638) );
  NAND2_X1 U11567 ( .A1(n9638), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8968) );
  NAND2_X2 U11568 ( .A1(n15181), .A2(n12468), .ZN(n12510) );
  INV_X1 U11569 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8966) );
  OR2_X1 U11570 ( .A1(n6440), .A2(n8966), .ZN(n8967) );
  OAI211_X1 U11571 ( .C1(n12508), .C2(n14791), .A(n8968), .B(n8967), .ZN(
        n14634) );
  AND2_X1 U11572 ( .A1(n9219), .A2(n15190), .ZN(n10458) );
  NAND2_X1 U11573 ( .A1(n10458), .A2(n14671), .ZN(n15052) );
  INV_X1 U11574 ( .A(P1_B_REG_SCAN_IN), .ZN(n14574) );
  NOR2_X1 U11575 ( .A1(n15291), .A2(n14574), .ZN(n8970) );
  NOR2_X1 U11576 ( .A1(n15052), .A2(n8970), .ZN(n12514) );
  NAND2_X1 U11577 ( .A1(n14634), .A2(n12514), .ZN(n15064) );
  INV_X1 U11578 ( .A(n8985), .ZN(n8974) );
  INV_X1 U11579 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8973) );
  INV_X1 U11580 ( .A(n8984), .ZN(n12319) );
  NAND2_X1 U11581 ( .A1(n8976), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8977) );
  INV_X1 U11582 ( .A(n8983), .ZN(n12208) );
  NAND3_X1 U11583 ( .A1(n12319), .A2(P1_B_REG_SCAN_IN), .A3(n12208), .ZN(n8981) );
  NAND2_X1 U11584 ( .A1(n8978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8979) );
  XNOR2_X1 U11585 ( .A(n8979), .B(P1_IR_REG_26__SCAN_IN), .ZN(n8982) );
  INV_X1 U11586 ( .A(n8982), .ZN(n15189) );
  AOI21_X1 U11587 ( .B1(n8983), .B2(n14574), .A(n15189), .ZN(n8980) );
  NOR2_X1 U11588 ( .A1(n10460), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9000) );
  AND2_X1 U11589 ( .A1(n12319), .A2(n15189), .ZN(n10461) );
  NAND2_X1 U11590 ( .A1(n8985), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8986) );
  XNOR2_X1 U11591 ( .A(n8986), .B(n8973), .ZN(n10457) );
  NAND2_X1 U11592 ( .A1(n10458), .A2(n8987), .ZN(n9667) );
  NOR4_X1 U11593 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8991) );
  NOR4_X1 U11594 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n8990) );
  NOR4_X1 U11595 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8989) );
  NOR4_X1 U11596 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n8988) );
  NAND4_X1 U11597 ( .A1(n8991), .A2(n8990), .A3(n8989), .A4(n8988), .ZN(n8997)
         );
  NOR2_X1 U11598 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n8995) );
  NOR4_X1 U11599 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n8994) );
  NOR4_X1 U11600 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n8993) );
  NOR4_X1 U11601 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n8992) );
  NAND4_X1 U11602 ( .A1(n8995), .A2(n8994), .A3(n8993), .A4(n8992), .ZN(n8996)
         );
  NOR2_X1 U11603 ( .A1(n8997), .A2(n8996), .ZN(n9629) );
  NAND2_X1 U11604 ( .A1(n15333), .A2(n14381), .ZN(n11264) );
  OAI21_X1 U11605 ( .B1(n10460), .B2(n9629), .A(n11264), .ZN(n8998) );
  INV_X1 U11606 ( .A(n8998), .ZN(n8999) );
  OAI211_X1 U11607 ( .C1(n9000), .C2(n10461), .A(n14577), .B(n8999), .ZN(
        n10718) );
  OR2_X1 U11608 ( .A1(n10460), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9001) );
  NAND2_X1 U11609 ( .A1(n12208), .A2(n15189), .ZN(n10463) );
  INV_X2 U11610 ( .A(n15406), .ZN(n15408) );
  NAND2_X1 U11611 ( .A1(n15406), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U11612 ( .A1(n13673), .A2(n10637), .ZN(n11348) );
  NAND2_X1 U11613 ( .A1(n11251), .A2(n15537), .ZN(n11242) );
  NAND2_X1 U11614 ( .A1(n12120), .A2(n8567), .ZN(n11240) );
  NAND2_X1 U11615 ( .A1(n11241), .A2(n11242), .ZN(n9004) );
  INV_X1 U11616 ( .A(n13671), .ZN(n12119) );
  NAND2_X1 U11617 ( .A1(n12119), .A2(n12056), .ZN(n9007) );
  INV_X1 U11618 ( .A(n11307), .ZN(n11328) );
  INV_X1 U11619 ( .A(n13670), .ZN(n11181) );
  INV_X1 U11620 ( .A(n6432), .ZN(n12029) );
  NAND2_X1 U11621 ( .A1(n11181), .A2(n12029), .ZN(n9008) );
  NAND2_X1 U11622 ( .A1(n12046), .A2(n11312), .ZN(n9009) );
  OAI21_X1 U11623 ( .B1(n12038), .B2(n13669), .A(n9009), .ZN(n9014) );
  NAND2_X1 U11624 ( .A1(n13669), .A2(n12038), .ZN(n9010) );
  NAND2_X1 U11625 ( .A1(n9010), .A2(n11312), .ZN(n9012) );
  INV_X1 U11626 ( .A(n9010), .ZN(n9011) );
  AOI22_X1 U11627 ( .A1(n15543), .A2(n9012), .B1(n13668), .B2(n9011), .ZN(
        n9013) );
  INV_X1 U11628 ( .A(n11992), .ZN(n11988) );
  OR2_X1 U11629 ( .A1(n11999), .A2(n11475), .ZN(n9015) );
  OR2_X1 U11630 ( .A1(n12015), .A2(n11702), .ZN(n9016) );
  AOI22_X1 U11631 ( .A1(n12110), .A2(n12168), .B1(n11754), .B2(n11984), .ZN(
        n9017) );
  OR2_X1 U11632 ( .A1(n11984), .A2(n11754), .ZN(n11967) );
  NAND2_X1 U11633 ( .A1(n11967), .A2(n12168), .ZN(n9019) );
  NOR2_X1 U11634 ( .A1(n11754), .A2(n12168), .ZN(n9018) );
  AOI22_X1 U11635 ( .A1(n9020), .A2(n9019), .B1(n9018), .B2(n14106), .ZN(n9021) );
  NAND2_X1 U11636 ( .A1(n14161), .A2(n12195), .ZN(n9022) );
  INV_X1 U11637 ( .A(n9023), .ZN(n9025) );
  NOR2_X1 U11638 ( .A1(n14089), .A2(n13967), .ZN(n9027) );
  NAND2_X1 U11639 ( .A1(n14089), .A2(n13967), .ZN(n9026) );
  NOR2_X1 U11640 ( .A1(n13941), .A2(n13641), .ZN(n13911) );
  NAND2_X1 U11641 ( .A1(n13901), .A2(n13549), .ZN(n9030) );
  OR2_X1 U11642 ( .A1(n13882), .A2(n13859), .ZN(n9031) );
  NAND2_X1 U11643 ( .A1(n13882), .A2(n13859), .ZN(n9032) );
  NAND2_X1 U11644 ( .A1(n14140), .A2(n13656), .ZN(n9033) );
  OR2_X1 U11645 ( .A1(n14133), .A2(n13843), .ZN(n9035) );
  NAND2_X1 U11646 ( .A1(n14036), .A2(n13810), .ZN(n9037) );
  NAND3_X1 U11647 ( .A1(n9039), .A2(n13705), .A3(n12562), .ZN(n15546) );
  NAND2_X1 U11648 ( .A1(n13896), .A2(n15546), .ZN(n15541) );
  INV_X1 U11649 ( .A(n15541), .ZN(n15557) );
  INV_X1 U11650 ( .A(n11355), .ZN(n9040) );
  NAND2_X1 U11651 ( .A1(n12120), .A2(n6645), .ZN(n12116) );
  NAND2_X1 U11652 ( .A1(n9041), .A2(n11241), .ZN(n11247) );
  AOI22_X1 U11653 ( .A1(n12056), .A2(n13671), .B1(n13670), .B2(n12029), .ZN(
        n9042) );
  NAND2_X1 U11654 ( .A1(n11327), .A2(n13670), .ZN(n9045) );
  NOR2_X1 U11655 ( .A1(n13671), .A2(n13670), .ZN(n9044) );
  AOI22_X1 U11656 ( .A1(n9045), .A2(n6432), .B1(n9044), .B2(n8571), .ZN(n9046)
         );
  OR2_X1 U11657 ( .A1(n13668), .A2(n12046), .ZN(n9050) );
  NAND2_X1 U11658 ( .A1(n11999), .A2(n13666), .ZN(n9051) );
  NAND2_X1 U11659 ( .A1(n11993), .A2(n9051), .ZN(n9053) );
  OR2_X1 U11660 ( .A1(n11999), .A2(n13666), .ZN(n9052) );
  INV_X1 U11661 ( .A(n12004), .ZN(n12007) );
  OR2_X1 U11662 ( .A1(n12015), .A2(n13665), .ZN(n9054) );
  NOR2_X1 U11663 ( .A1(n11984), .A2(n13664), .ZN(n9057) );
  NAND2_X1 U11664 ( .A1(n11984), .A2(n13664), .ZN(n9056) );
  OR2_X1 U11665 ( .A1(n12110), .A2(n13663), .ZN(n12162) );
  OR2_X1 U11666 ( .A1(n14161), .A2(n13662), .ZN(n9059) );
  NAND2_X1 U11667 ( .A1(n12282), .A2(n13661), .ZN(n9060) );
  OR2_X1 U11668 ( .A1(n12282), .A2(n13661), .ZN(n9061) );
  AND2_X1 U11669 ( .A1(n14089), .A2(n13530), .ZN(n9062) );
  OR2_X1 U11670 ( .A1(n13955), .A2(n13931), .ZN(n9064) );
  NAND2_X1 U11671 ( .A1(n13955), .A2(n13931), .ZN(n9065) );
  INV_X1 U11672 ( .A(n13893), .ZN(n13933) );
  OR2_X1 U11673 ( .A1(n13920), .A2(n13933), .ZN(n9067) );
  AND2_X1 U11674 ( .A1(n13901), .A2(n13657), .ZN(n9070) );
  OR2_X1 U11675 ( .A1(n13901), .A2(n13657), .ZN(n9069) );
  NOR2_X1 U11676 ( .A1(n13882), .A2(n13894), .ZN(n9071) );
  INV_X1 U11677 ( .A(n13794), .ZN(n13595) );
  NAND2_X1 U11678 ( .A1(n13541), .A2(n13595), .ZN(n13791) );
  INV_X1 U11679 ( .A(n13791), .ZN(n9074) );
  OR2_X1 U11680 ( .A1(n14137), .A2(n13655), .ZN(n13789) );
  AND2_X1 U11681 ( .A1(n13790), .A2(n13595), .ZN(n9076) );
  OAI22_X1 U11682 ( .A1(n9076), .A2(n13541), .B1(n13595), .B2(n13790), .ZN(
        n9077) );
  NOR2_X1 U11683 ( .A1(n9077), .A2(n13802), .ZN(n9078) );
  NAND2_X1 U11684 ( .A1(n13751), .A2(n13635), .ZN(n9085) );
  OR2_X1 U11685 ( .A1(n11770), .A2(n12562), .ZN(n9083) );
  AOI21_X1 U11686 ( .B1(n13741), .B2(n9085), .A(n14008), .ZN(n9087) );
  AOI22_X1 U11687 ( .A1(n13653), .A2(n13968), .B1(n13760), .B2(n13966), .ZN(
        n9086) );
  NAND2_X1 U11688 ( .A1(n12123), .A2(n15537), .ZN(n12122) );
  NOR2_X2 U11689 ( .A1(n12122), .A2(n8571), .ZN(n11335) );
  NAND2_X1 U11690 ( .A1(n11335), .A2(n12029), .ZN(n11336) );
  NOR2_X4 U11691 ( .A1(n13878), .A2(n14140), .ZN(n13865) );
  AOI211_X1 U11692 ( .C1(n13720), .C2(n13747), .A(n13974), .B(n6431), .ZN(
        n9199) );
  INV_X1 U11693 ( .A(n9199), .ZN(n9089) );
  INV_X1 U11694 ( .A(n13720), .ZN(n9088) );
  NAND4_X1 U11695 ( .A1(n9192), .A2(n15532), .A3(n9092), .A4(n9091), .ZN(n9214) );
  NOR2_X1 U11696 ( .A1(n9214), .A2(n15529), .ZN(n15569) );
  NAND2_X1 U11697 ( .A1(n9095), .A2(n9094), .ZN(P2_U3527) );
  INV_X1 U11698 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15507) );
  INV_X1 U11699 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15280) );
  INV_X1 U11700 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9166) );
  XNOR2_X1 U11701 ( .A(n6946), .B(n9166), .ZN(n9164) );
  INV_X1 U11702 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9121) );
  XNOR2_X1 U11703 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9124) );
  INV_X1 U11704 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11817) );
  XNOR2_X1 U11705 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9159) );
  INV_X1 U11706 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9115) );
  XNOR2_X1 U11707 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9127) );
  INV_X1 U11708 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n9113) );
  XNOR2_X1 U11709 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9157) );
  INV_X1 U11710 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10839) );
  XNOR2_X1 U11711 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n9150) );
  NAND2_X1 U11712 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n9102), .ZN(n9103) );
  NAND2_X1 U11713 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n9104), .ZN(n9105) );
  NAND2_X1 U11714 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n9106), .ZN(n9108) );
  NAND2_X1 U11715 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n9110), .ZN(n9111) );
  NAND2_X1 U11716 ( .A1(n9127), .A2(n9126), .ZN(n9114) );
  NAND2_X1 U11717 ( .A1(n9115), .A2(n9116), .ZN(n9117) );
  NAND2_X1 U11718 ( .A1(n9124), .A2(n9125), .ZN(n9119) );
  INV_X1 U11719 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U11720 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n10837), .ZN(n9120) );
  XOR2_X1 U11721 ( .A(n9164), .B(n9163), .Z(n15278) );
  INV_X1 U11722 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15275) );
  XNOR2_X1 U11723 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9123) );
  XNOR2_X1 U11724 ( .A(n9123), .B(n9122), .ZN(n15273) );
  XNOR2_X1 U11725 ( .A(n9125), .B(n9124), .ZN(n9161) );
  INV_X1 U11726 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15269) );
  XNOR2_X1 U11727 ( .A(n9127), .B(n9126), .ZN(n15210) );
  XNOR2_X1 U11728 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9128), .ZN(n15658) );
  NOR2_X1 U11729 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9143), .ZN(n9145) );
  INV_X1 U11730 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15201) );
  XNOR2_X1 U11731 ( .A(n9131), .B(n9130), .ZN(n9139) );
  XNOR2_X1 U11732 ( .A(n9132), .B(n9135), .ZN(n9134) );
  NAND2_X1 U11733 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9134), .ZN(n9137) );
  AOI21_X1 U11734 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n11425), .A(n9135), .ZN(
        n15657) );
  INV_X1 U11735 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15656) );
  NOR2_X1 U11736 ( .A1(n15657), .A2(n15656), .ZN(n15665) );
  NAND2_X1 U11737 ( .A1(n9137), .A2(n9136), .ZN(n9138) );
  NAND2_X1 U11738 ( .A1(n9139), .A2(n9138), .ZN(n15198) );
  NOR2_X1 U11739 ( .A1(n9139), .A2(n9138), .ZN(n15199) );
  XNOR2_X1 U11740 ( .A(n9141), .B(n9140), .ZN(n15662) );
  NOR2_X1 U11741 ( .A1(n15661), .A2(n15662), .ZN(n9142) );
  INV_X1 U11742 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15456) );
  NAND2_X1 U11743 ( .A1(n15661), .A2(n15662), .ZN(n15660) );
  OAI21_X1 U11744 ( .B1(n9142), .B2(n15456), .A(n15660), .ZN(n15654) );
  XNOR2_X1 U11745 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n9143), .ZN(n15653) );
  XNOR2_X1 U11746 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9146), .ZN(n9147) );
  XNOR2_X1 U11747 ( .A(n9151), .B(n9150), .ZN(n15203) );
  NAND2_X1 U11748 ( .A1(n15202), .A2(n15203), .ZN(n9154) );
  NAND2_X1 U11749 ( .A1(n9152), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9153) );
  XNOR2_X1 U11750 ( .A(n9157), .B(n9156), .ZN(n15206) );
  INV_X1 U11751 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15495) );
  NAND2_X1 U11752 ( .A1(n15210), .A2(n15209), .ZN(n15208) );
  XNOR2_X1 U11753 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n9158), .ZN(n15214) );
  INV_X1 U11754 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15215) );
  XNOR2_X1 U11755 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n9167) );
  NAND2_X1 U11756 ( .A1(n9164), .A2(n9163), .ZN(n9165) );
  XOR2_X1 U11757 ( .A(n9167), .B(n9169), .Z(n9168) );
  INV_X1 U11758 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n13073) );
  NAND2_X1 U11759 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n13073), .ZN(n9173) );
  OAI21_X1 U11760 ( .B1(n13073), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9173), .ZN(
        n9171) );
  INV_X1 U11761 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13038) );
  INV_X1 U11762 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15320) );
  NOR2_X1 U11763 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15320), .ZN(n9170) );
  XOR2_X1 U11764 ( .A(n9171), .B(n9174), .Z(n15287) );
  NOR2_X1 U11765 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n13073), .ZN(n9175) );
  XOR2_X1 U11766 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9176), .Z(n9177) );
  INV_X1 U11767 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15523) );
  NOR2_X1 U11768 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9176), .ZN(n9179) );
  XOR2_X1 U11769 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n9182) );
  XNOR2_X1 U11770 ( .A(n9183), .B(n9182), .ZN(n9180) );
  INV_X1 U11771 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9185) );
  NOR2_X1 U11772 ( .A1(n9183), .A2(n9182), .ZN(n9184) );
  AOI21_X1 U11773 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n9185), .A(n9184), .ZN(
        n9186) );
  XNOR2_X1 U11774 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9187) );
  INV_X1 U11775 ( .A(n13956), .ZN(n13990) );
  INV_X1 U11776 ( .A(n9191), .ZN(n9193) );
  NAND3_X1 U11777 ( .A1(n9193), .A2(n9192), .A3(n15529), .ZN(n9194) );
  INV_X1 U11778 ( .A(n13896), .ZN(n15550) );
  AND2_X2 U11779 ( .A1(n13987), .A2(n11614), .ZN(n13995) );
  INV_X1 U11780 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9197) );
  OAI22_X1 U11781 ( .A1(n9088), .A2(n13979), .B1(n13987), .B2(n9197), .ZN(
        n9198) );
  OAI211_X1 U11782 ( .C1(n9205), .C2(n9204), .A(n9203), .B(n13610), .ZN(n9212)
         );
  INV_X1 U11783 ( .A(n13749), .ZN(n9206) );
  AOI22_X1 U11784 ( .A1(n9206), .A2(n13631), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9207) );
  OAI21_X1 U11785 ( .B1(n13744), .B2(n13623), .A(n9207), .ZN(n9208) );
  AOI21_X1 U11786 ( .B1(n13568), .B2(n13742), .A(n9208), .ZN(n9209) );
  OAI21_X1 U11787 ( .B1(n14121), .B2(n13620), .A(n9209), .ZN(n9210) );
  NAND2_X1 U11788 ( .A1(n9212), .A2(n9211), .ZN(P2_U3186) );
  INV_X1 U11789 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9215) );
  NOR2_X1 U11790 ( .A1(n15561), .A2(n9215), .ZN(n9216) );
  INV_X1 U11791 ( .A(n9218), .ZN(P2_U3495) );
  INV_X4 U11792 ( .A(n12510), .ZN(n9658) );
  NAND2_X1 U11793 ( .A1(n9658), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9227) );
  INV_X1 U11794 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10873) );
  OR2_X1 U11795 ( .A1(n9288), .A2(n10873), .ZN(n9226) );
  NAND2_X1 U11796 ( .A1(n9331), .A2(n10871), .ZN(n9223) );
  NAND2_X1 U11797 ( .A1(n9353), .A2(n9223), .ZN(n12260) );
  OR2_X1 U11798 ( .A1(n6433), .A2(n12260), .ZN(n9225) );
  INV_X1 U11799 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n12221) );
  OR2_X1 U11800 ( .A1(n12508), .A2(n12221), .ZN(n9224) );
  AOI22_X1 U11801 ( .A1(n14428), .A2(n9649), .B1(n9648), .B2(n15048), .ZN(
        n9340) );
  AOI22_X1 U11802 ( .A1(n14428), .A2(n9634), .B1(n9649), .B2(n15048), .ZN(
        n9228) );
  XNOR2_X1 U11803 ( .A(n9228), .B(n10720), .ZN(n9339) );
  NAND2_X1 U11804 ( .A1(n9658), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9234) );
  INV_X1 U11805 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9229) );
  OR2_X1 U11806 ( .A1(n9288), .A2(n9229), .ZN(n9233) );
  NAND2_X1 U11807 ( .A1(n9314), .A2(n10708), .ZN(n9230) );
  NAND2_X1 U11808 ( .A1(n9329), .A2(n9230), .ZN(n11743) );
  OR2_X1 U11809 ( .A1(n6433), .A2(n11743), .ZN(n9232) );
  INV_X1 U11810 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11685) );
  OR2_X1 U11811 ( .A1(n12508), .A2(n11685), .ZN(n9231) );
  OAI22_X1 U11812 ( .A1(n11689), .A2(n9284), .B1(n11948), .B2(n9621), .ZN(
        n9327) );
  NAND2_X1 U11813 ( .A1(n14419), .A2(n9634), .ZN(n9236) );
  OR2_X1 U11814 ( .A1(n11948), .A2(n9284), .ZN(n9235) );
  NAND2_X1 U11815 ( .A1(n9236), .A2(n9235), .ZN(n9237) );
  XNOR2_X1 U11816 ( .A(n9237), .B(n10720), .ZN(n9326) );
  INV_X1 U11817 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n14655) );
  INV_X1 U11818 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11271) );
  OR2_X1 U11819 ( .A1(n9463), .A2(n11271), .ZN(n9240) );
  INV_X1 U11820 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9238) );
  OR2_X1 U11821 ( .A1(n6439), .A2(n9238), .ZN(n9239) );
  NAND2_X1 U11822 ( .A1(n11380), .A2(n9644), .ZN(n9244) );
  NAND2_X1 U11823 ( .A1(n11370), .A2(n9634), .ZN(n9243) );
  NAND2_X1 U11824 ( .A1(n9244), .A2(n9243), .ZN(n9245) );
  XNOR2_X1 U11825 ( .A(n9245), .B(n9619), .ZN(n9247) );
  INV_X1 U11826 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11449) );
  OR2_X1 U11827 ( .A1(n6434), .A2(n11449), .ZN(n9249) );
  INV_X1 U11828 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U11829 ( .A1(n9638), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9250) );
  NAND3_X2 U11830 ( .A1(n6430), .A2(n9251), .A3(n9250), .ZN(n11377) );
  NAND2_X1 U11831 ( .A1(n11377), .A2(n9648), .ZN(n9253) );
  INV_X1 U11832 ( .A(n10393), .ZN(n9254) );
  AOI22_X1 U11833 ( .A1(n11453), .A2(n9649), .B1(n15193), .B2(n9254), .ZN(
        n9252) );
  NAND2_X1 U11834 ( .A1(n11377), .A2(n9649), .ZN(n9256) );
  AOI22_X1 U11835 ( .A1(n11453), .A2(n9634), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n9254), .ZN(n9255) );
  NAND2_X1 U11836 ( .A1(n9638), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9262) );
  INV_X1 U11837 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9257) );
  OR2_X1 U11838 ( .A1(n6434), .A2(n9257), .ZN(n9261) );
  INV_X1 U11839 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n14676) );
  INV_X1 U11840 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9258) );
  OR2_X1 U11841 ( .A1(n6440), .A2(n9258), .ZN(n9259) );
  NAND2_X1 U11842 ( .A1(n11381), .A2(n9644), .ZN(n9264) );
  NAND2_X1 U11843 ( .A1(n9634), .A2(n15330), .ZN(n9263) );
  NAND2_X1 U11844 ( .A1(n9264), .A2(n9263), .ZN(n9265) );
  XNOR2_X1 U11845 ( .A(n9265), .B(n10720), .ZN(n9273) );
  AOI22_X1 U11846 ( .A1(n11381), .A2(n9648), .B1(n9649), .B2(n15330), .ZN(
        n9274) );
  XNOR2_X1 U11847 ( .A(n9273), .B(n9274), .ZN(n11154) );
  INV_X1 U11848 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10615) );
  INV_X1 U11849 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U11850 ( .A1(n9638), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U11851 ( .A1(n14652), .A2(n9644), .ZN(n9269) );
  NAND2_X1 U11852 ( .A1(n9634), .A2(n11629), .ZN(n9268) );
  NAND2_X1 U11853 ( .A1(n9269), .A2(n9268), .ZN(n9270) );
  XNOR2_X1 U11854 ( .A(n9270), .B(n10720), .ZN(n10397) );
  NAND2_X1 U11855 ( .A1(n14652), .A2(n9648), .ZN(n9272) );
  NAND2_X1 U11856 ( .A1(n9649), .A2(n11629), .ZN(n9271) );
  NAND2_X1 U11857 ( .A1(n9272), .A2(n9271), .ZN(n10396) );
  INV_X1 U11858 ( .A(n9273), .ZN(n9275) );
  NAND2_X1 U11859 ( .A1(n9275), .A2(n9274), .ZN(n10398) );
  NAND2_X1 U11860 ( .A1(n9638), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9280) );
  INV_X1 U11861 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9276) );
  OR2_X1 U11862 ( .A1(n12510), .A2(n9276), .ZN(n9279) );
  OAI21_X1 U11863 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9289), .ZN(n11553) );
  OR2_X1 U11864 ( .A1(n6434), .A2(n11553), .ZN(n9278) );
  INV_X1 U11865 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11552) );
  OR2_X1 U11866 ( .A1(n12508), .A2(n11552), .ZN(n9277) );
  NAND2_X1 U11867 ( .A1(n14651), .A2(n9644), .ZN(n9282) );
  OR2_X1 U11868 ( .A1(n11622), .A2(n9604), .ZN(n9281) );
  NAND2_X1 U11869 ( .A1(n9282), .A2(n9281), .ZN(n9283) );
  XNOR2_X1 U11870 ( .A(n9283), .B(n9619), .ZN(n9303) );
  NAND2_X1 U11871 ( .A1(n14651), .A2(n9648), .ZN(n9286) );
  OR2_X1 U11872 ( .A1(n11622), .A2(n9284), .ZN(n9285) );
  INV_X1 U11873 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10684) );
  OR2_X1 U11874 ( .A1(n9288), .A2(n10684), .ZN(n9293) );
  INV_X1 U11875 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10743) );
  NAND2_X1 U11876 ( .A1(n9289), .A2(n10743), .ZN(n9290) );
  NAND2_X1 U11877 ( .A1(n9312), .A2(n9290), .ZN(n11609) );
  OR2_X1 U11878 ( .A1(n6433), .A2(n11609), .ZN(n9292) );
  INV_X1 U11879 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11594) );
  OR2_X1 U11880 ( .A1(n12508), .A2(n11594), .ZN(n9291) );
  NAND2_X1 U11881 ( .A1(n14650), .A2(n9644), .ZN(n9296) );
  OR2_X1 U11882 ( .A1(n11635), .A2(n9604), .ZN(n9295) );
  NAND2_X1 U11883 ( .A1(n9296), .A2(n9295), .ZN(n9297) );
  XNOR2_X1 U11884 ( .A(n9297), .B(n9619), .ZN(n11603) );
  NAND2_X1 U11885 ( .A1(n14650), .A2(n9648), .ZN(n9299) );
  OR2_X1 U11886 ( .A1(n11635), .A2(n9284), .ZN(n9298) );
  AND2_X1 U11887 ( .A1(n9299), .A2(n9298), .ZN(n11602) );
  NAND2_X1 U11888 ( .A1(n11603), .A2(n11602), .ZN(n11601) );
  NOR2_X1 U11889 ( .A1(n9301), .A2(n9300), .ZN(n9302) );
  OAI21_X1 U11890 ( .B1(n11153), .B2(n11516), .A(n9302), .ZN(n9309) );
  INV_X1 U11891 ( .A(n9303), .ZN(n11599) );
  INV_X1 U11892 ( .A(n11519), .ZN(n11598) );
  INV_X1 U11893 ( .A(n11602), .ZN(n9304) );
  AOI21_X1 U11894 ( .B1(n11599), .B2(n11598), .A(n9304), .ZN(n9306) );
  NAND3_X1 U11895 ( .A1(n11599), .A2(n9304), .A3(n11598), .ZN(n9305) );
  NAND2_X1 U11896 ( .A1(n9638), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9318) );
  INV_X1 U11897 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9310) );
  OR2_X1 U11898 ( .A1(n12510), .A2(n9310), .ZN(n9317) );
  INV_X1 U11899 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U11900 ( .A1(n9312), .A2(n9311), .ZN(n9313) );
  NAND2_X1 U11901 ( .A1(n9314), .A2(n9313), .ZN(n11544) );
  OR2_X1 U11902 ( .A1(n6433), .A2(n11544), .ZN(n9316) );
  INV_X1 U11903 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11643) );
  OR2_X1 U11904 ( .A1(n12508), .A2(n11643), .ZN(n9315) );
  NAND4_X1 U11905 ( .A1(n9318), .A2(n9317), .A3(n9316), .A4(n9315), .ZN(n14649) );
  NAND2_X1 U11906 ( .A1(n14649), .A2(n9644), .ZN(n9320) );
  NAND2_X1 U11907 ( .A1(n14413), .A2(n9634), .ZN(n9319) );
  NAND2_X1 U11908 ( .A1(n9320), .A2(n9319), .ZN(n9321) );
  XNOR2_X1 U11909 ( .A(n9321), .B(n10720), .ZN(n9322) );
  AOI22_X1 U11910 ( .A1(n9648), .A2(n14649), .B1(n14413), .B2(n9644), .ZN(
        n9323) );
  XNOR2_X1 U11911 ( .A(n9322), .B(n9323), .ZN(n11542) );
  INV_X1 U11912 ( .A(n9323), .ZN(n9324) );
  NAND2_X1 U11913 ( .A1(n9322), .A2(n9324), .ZN(n9325) );
  XOR2_X1 U11914 ( .A(n9327), .B(n9326), .Z(n11741) );
  NAND2_X1 U11915 ( .A1(n9658), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9335) );
  INV_X1 U11916 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9328) );
  OR2_X1 U11917 ( .A1(n9288), .A2(n9328), .ZN(n9334) );
  NAND2_X1 U11918 ( .A1(n9329), .A2(n11952), .ZN(n9330) );
  NAND2_X1 U11919 ( .A1(n9331), .A2(n9330), .ZN(n12185) );
  OR2_X1 U11920 ( .A1(n6433), .A2(n12185), .ZN(n9333) );
  INV_X1 U11921 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10698) );
  OR2_X1 U11922 ( .A1(n12508), .A2(n10698), .ZN(n9332) );
  NAND4_X1 U11923 ( .A1(n9335), .A2(n9334), .A3(n9333), .A4(n9332), .ZN(n14648) );
  AOI22_X1 U11924 ( .A1(n14424), .A2(n9634), .B1(n9649), .B2(n14648), .ZN(
        n9336) );
  XNOR2_X1 U11925 ( .A(n9336), .B(n10720), .ZN(n9338) );
  AOI22_X1 U11926 ( .A1(n14424), .A2(n9649), .B1(n9648), .B2(n14648), .ZN(
        n9337) );
  XNOR2_X1 U11927 ( .A(n9338), .B(n9337), .ZN(n11947) );
  XOR2_X1 U11928 ( .A(n9340), .B(n9339), .Z(n12258) );
  NAND2_X1 U11929 ( .A1(n9658), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9345) );
  INV_X1 U11930 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9341) );
  OR2_X1 U11931 ( .A1(n9288), .A2(n9341), .ZN(n9344) );
  INV_X1 U11932 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9352) );
  XNOR2_X1 U11933 ( .A(n9353), .B(n9352), .ZN(n15056) );
  OR2_X1 U11934 ( .A1(n6434), .A2(n15056), .ZN(n9343) );
  INV_X1 U11935 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n15050) );
  OR2_X1 U11936 ( .A1(n12508), .A2(n15050), .ZN(n9342) );
  NOR2_X1 U11937 ( .A1(n14439), .A2(n9284), .ZN(n9346) );
  AOI21_X1 U11938 ( .B1(n15399), .B2(n9634), .A(n9346), .ZN(n9347) );
  XNOR2_X1 U11939 ( .A(n9347), .B(n10720), .ZN(n9349) );
  OAI22_X1 U11940 ( .A1(n15058), .A2(n9284), .B1(n14439), .B2(n9621), .ZN(
        n9348) );
  XNOR2_X1 U11941 ( .A(n9349), .B(n9348), .ZN(n14213) );
  INV_X1 U11942 ( .A(n9348), .ZN(n9350) );
  NAND2_X1 U11943 ( .A1(n9658), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9361) );
  INV_X1 U11944 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9351) );
  OAI21_X1 U11945 ( .B1(n9353), .B2(n9352), .A(n9351), .ZN(n9356) );
  NAND2_X1 U11946 ( .A1(n9356), .A2(n9368), .ZN(n14343) );
  OR2_X1 U11947 ( .A1(n6433), .A2(n14343), .ZN(n9360) );
  INV_X1 U11948 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9357) );
  OR2_X1 U11949 ( .A1(n9288), .A2(n9357), .ZN(n9359) );
  INV_X1 U11950 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11939) );
  OR2_X1 U11951 ( .A1(n12508), .A2(n11939), .ZN(n9358) );
  OAI22_X1 U11952 ( .A1(n15259), .A2(n9604), .B1(n15053), .B2(n9284), .ZN(
        n9362) );
  XNOR2_X1 U11953 ( .A(n9362), .B(n10720), .ZN(n9365) );
  OAI22_X1 U11954 ( .A1(n15259), .A2(n9284), .B1(n15053), .B2(n9621), .ZN(
        n9364) );
  XNOR2_X1 U11955 ( .A(n9365), .B(n9364), .ZN(n14342) );
  INV_X1 U11956 ( .A(n14342), .ZN(n9363) );
  OR2_X1 U11957 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  NAND2_X1 U11958 ( .A1(n9658), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9374) );
  INV_X1 U11959 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11288) );
  OR2_X1 U11960 ( .A1(n9288), .A2(n11288), .ZN(n9373) );
  NAND2_X1 U11961 ( .A1(n9368), .A2(n9367), .ZN(n9369) );
  NAND2_X1 U11962 ( .A1(n9387), .A2(n9369), .ZN(n15228) );
  OR2_X1 U11963 ( .A1(n6434), .A2(n15228), .ZN(n9372) );
  INV_X1 U11964 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9370) );
  OR2_X1 U11965 ( .A1(n12508), .A2(n9370), .ZN(n9371) );
  NAND4_X1 U11966 ( .A1(n9374), .A2(n9373), .A3(n9372), .A4(n9371), .ZN(n15027) );
  AND2_X1 U11967 ( .A1(n15027), .A2(n9648), .ZN(n9375) );
  AOI21_X1 U11968 ( .B1(n15230), .B2(n9649), .A(n9375), .ZN(n9381) );
  NAND2_X1 U11969 ( .A1(n15230), .A2(n9634), .ZN(n9377) );
  NAND2_X1 U11970 ( .A1(n15027), .A2(n9649), .ZN(n9376) );
  NAND2_X1 U11971 ( .A1(n9377), .A2(n9376), .ZN(n9378) );
  XNOR2_X1 U11972 ( .A(n9378), .B(n10720), .ZN(n9380) );
  XOR2_X1 U11973 ( .A(n9381), .B(n9380), .Z(n14250) );
  INV_X1 U11974 ( .A(n9381), .ZN(n9382) );
  NAND2_X1 U11975 ( .A1(n9380), .A2(n9382), .ZN(n9383) );
  INV_X1 U11976 ( .A(n15036), .ZN(n15252) );
  NAND2_X1 U11977 ( .A1(n9638), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9392) );
  INV_X1 U11978 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9384) );
  OR2_X1 U11979 ( .A1(n6440), .A2(n9384), .ZN(n9391) );
  INV_X1 U11980 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U11981 ( .A1(n9387), .A2(n9386), .ZN(n9388) );
  NAND2_X1 U11982 ( .A1(n9400), .A2(n9388), .ZN(n15033) );
  OR2_X1 U11983 ( .A1(n6433), .A2(n15033), .ZN(n9390) );
  INV_X1 U11984 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n15034) );
  OR2_X1 U11985 ( .A1(n12508), .A2(n15034), .ZN(n9389) );
  NAND4_X1 U11986 ( .A1(n9392), .A2(n9391), .A3(n9390), .A4(n9389), .ZN(n15221) );
  INV_X1 U11987 ( .A(n15221), .ZN(n14443) );
  OAI22_X1 U11988 ( .A1(n15252), .A2(n9604), .B1(n14443), .B2(n9284), .ZN(
        n9393) );
  XNOR2_X1 U11989 ( .A(n9393), .B(n10720), .ZN(n9395) );
  AND2_X1 U11990 ( .A1(n15221), .A2(n9648), .ZN(n9394) );
  AOI21_X1 U11991 ( .B1(n15036), .B2(n9649), .A(n9394), .ZN(n9396) );
  XNOR2_X1 U11992 ( .A(n9395), .B(n9396), .ZN(n14321) );
  INV_X1 U11993 ( .A(n9396), .ZN(n9397) );
  NAND2_X1 U11994 ( .A1(n9395), .A2(n9397), .ZN(n9398) );
  NAND2_X1 U11995 ( .A1(n15151), .A2(n9634), .ZN(n9407) );
  NAND2_X1 U11996 ( .A1(n9659), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9405) );
  INV_X1 U11997 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10755) );
  OR2_X1 U11998 ( .A1(n12510), .A2(n10755), .ZN(n9404) );
  INV_X1 U11999 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9399) );
  OR2_X1 U12000 ( .A1(n9288), .A2(n9399), .ZN(n9403) );
  INV_X1 U12001 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11725) );
  NAND2_X1 U12002 ( .A1(n9400), .A2(n11725), .ZN(n9401) );
  NAND2_X1 U12003 ( .A1(n9428), .A2(n9401), .ZN(n15007) );
  OR2_X1 U12004 ( .A1(n6434), .A2(n15007), .ZN(n9402) );
  NAND4_X1 U12005 ( .A1(n9405), .A2(n9404), .A3(n9403), .A4(n9402), .ZN(n15026) );
  NAND2_X1 U12006 ( .A1(n15026), .A2(n9649), .ZN(n9406) );
  NAND2_X1 U12007 ( .A1(n9407), .A2(n9406), .ZN(n9408) );
  XNOR2_X1 U12008 ( .A(n9408), .B(n10720), .ZN(n9411) );
  INV_X1 U12009 ( .A(n15151), .ZN(n15010) );
  INV_X1 U12010 ( .A(n15026), .ZN(n14324) );
  OAI22_X1 U12011 ( .A1(n15010), .A2(n9284), .B1(n14324), .B2(n9621), .ZN(
        n9410) );
  XNOR2_X1 U12012 ( .A(n9411), .B(n9410), .ZN(n14192) );
  OR2_X1 U12013 ( .A1(n9411), .A2(n9410), .ZN(n9412) );
  NAND2_X1 U12014 ( .A1(n15142), .A2(n9634), .ZN(n9422) );
  INV_X1 U12015 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U12016 ( .A1(n9638), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9413) );
  OAI21_X1 U12017 ( .B1(n6440), .B2(n9414), .A(n9413), .ZN(n9420) );
  INV_X1 U12018 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U12019 ( .A1(n9430), .A2(n9416), .ZN(n9417) );
  NAND2_X1 U12020 ( .A1(n9446), .A2(n9417), .ZN(n14979) );
  NAND2_X1 U12021 ( .A1(n9659), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9418) );
  OAI21_X1 U12022 ( .B1(n14979), .B2(n6434), .A(n9418), .ZN(n9419) );
  NAND2_X1 U12023 ( .A1(n14987), .A2(n9649), .ZN(n9421) );
  NAND2_X1 U12024 ( .A1(n9422), .A2(n9421), .ZN(n9423) );
  XNOR2_X1 U12025 ( .A(n9423), .B(n10720), .ZN(n14277) );
  NAND2_X1 U12026 ( .A1(n15142), .A2(n9649), .ZN(n9425) );
  NAND2_X1 U12027 ( .A1(n14987), .A2(n9648), .ZN(n9424) );
  NAND2_X1 U12028 ( .A1(n9425), .A2(n9424), .ZN(n14278) );
  NAND2_X1 U12029 ( .A1(n14277), .A2(n14278), .ZN(n9440) );
  NAND2_X1 U12030 ( .A1(n15146), .A2(n9634), .ZN(n9436) );
  NAND2_X1 U12031 ( .A1(n9658), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9434) );
  INV_X1 U12032 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15308) );
  OR2_X1 U12033 ( .A1(n9288), .A2(n15308), .ZN(n9433) );
  INV_X1 U12034 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9426) );
  OR2_X1 U12035 ( .A1(n12508), .A2(n9426), .ZN(n9432) );
  INV_X1 U12036 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U12037 ( .A1(n9428), .A2(n9427), .ZN(n9429) );
  NAND2_X1 U12038 ( .A1(n9430), .A2(n9429), .ZN(n14992) );
  OR2_X1 U12039 ( .A1(n6433), .A2(n14992), .ZN(n9431) );
  INV_X1 U12040 ( .A(n14975), .ZN(n14647) );
  NAND2_X1 U12041 ( .A1(n14647), .A2(n9649), .ZN(n9435) );
  NAND2_X1 U12042 ( .A1(n9436), .A2(n9435), .ZN(n9437) );
  XNOR2_X1 U12043 ( .A(n9437), .B(n9619), .ZN(n14276) );
  NOR2_X1 U12044 ( .A1(n14975), .A2(n9621), .ZN(n9438) );
  AOI21_X1 U12045 ( .B1(n15146), .B2(n9649), .A(n9438), .ZN(n14274) );
  NAND3_X1 U12046 ( .A1(n9440), .A2(n14276), .A3(n14274), .ZN(n9442) );
  NAND2_X1 U12047 ( .A1(n15137), .A2(n9634), .ZN(n9452) );
  INV_X1 U12048 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U12049 ( .A1(n9446), .A2(n9445), .ZN(n9447) );
  NAND2_X1 U12050 ( .A1(n9461), .A2(n9447), .ZN(n14959) );
  OR2_X1 U12051 ( .A1(n14959), .A2(n6433), .ZN(n9450) );
  AOI22_X1 U12052 ( .A1(n9658), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n9638), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n9449) );
  INV_X1 U12053 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14960) );
  OR2_X1 U12054 ( .A1(n12508), .A2(n14960), .ZN(n9448) );
  OR2_X1 U12055 ( .A1(n14974), .A2(n9284), .ZN(n9451) );
  NAND2_X1 U12056 ( .A1(n9452), .A2(n9451), .ZN(n9453) );
  XNOR2_X1 U12057 ( .A(n9453), .B(n10720), .ZN(n14288) );
  NAND2_X1 U12058 ( .A1(n15137), .A2(n9649), .ZN(n9455) );
  OR2_X1 U12059 ( .A1(n14974), .A2(n9621), .ZN(n9454) );
  NAND2_X1 U12060 ( .A1(n9455), .A2(n9454), .ZN(n14287) );
  NOR2_X1 U12061 ( .A1(n14288), .A2(n14287), .ZN(n9458) );
  INV_X1 U12062 ( .A(n14288), .ZN(n9457) );
  INV_X1 U12063 ( .A(n14287), .ZN(n9456) );
  INV_X1 U12064 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U12065 ( .A1(n9461), .A2(n9460), .ZN(n9462) );
  NAND2_X1 U12066 ( .A1(n9471), .A2(n9462), .ZN(n14938) );
  OR2_X1 U12067 ( .A1(n14938), .A2(n6434), .ZN(n9466) );
  AOI22_X1 U12068 ( .A1(n9658), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n9638), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U12069 ( .A1(n9659), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9464) );
  OAI22_X1 U12070 ( .A1(n14941), .A2(n9604), .B1(n14957), .B2(n9284), .ZN(
        n9467) );
  XNOR2_X1 U12071 ( .A(n9467), .B(n10720), .ZN(n14220) );
  INV_X1 U12072 ( .A(n14220), .ZN(n9496) );
  NAND2_X1 U12073 ( .A1(n15131), .A2(n9649), .ZN(n9469) );
  OR2_X1 U12074 ( .A1(n14957), .A2(n9621), .ZN(n9468) );
  NAND2_X1 U12075 ( .A1(n9469), .A2(n9468), .ZN(n14219) );
  INV_X1 U12076 ( .A(n14219), .ZN(n9494) );
  NAND2_X1 U12077 ( .A1(n15128), .A2(n9634), .ZN(n9480) );
  INV_X1 U12078 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U12079 ( .A1(n9471), .A2(n9470), .ZN(n9472) );
  NAND2_X1 U12080 ( .A1(n9484), .A2(n9472), .ZN(n14927) );
  OR2_X1 U12081 ( .A1(n14927), .A2(n6433), .ZN(n9478) );
  INV_X1 U12082 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U12083 ( .A1(n9638), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U12084 ( .A1(n9658), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9473) );
  OAI211_X1 U12085 ( .C1(n12508), .C2(n9475), .A(n9474), .B(n9473), .ZN(n9476)
         );
  INV_X1 U12086 ( .A(n9476), .ZN(n9477) );
  INV_X1 U12087 ( .A(n14944), .ZN(n14644) );
  NAND2_X1 U12088 ( .A1(n14644), .A2(n9649), .ZN(n9479) );
  NAND2_X1 U12089 ( .A1(n9480), .A2(n9479), .ZN(n9481) );
  XNOR2_X1 U12090 ( .A(n9481), .B(n9619), .ZN(n14223) );
  INV_X1 U12091 ( .A(n14223), .ZN(n9483) );
  NOR2_X1 U12092 ( .A1(n14944), .A2(n9621), .ZN(n9482) );
  AOI21_X1 U12093 ( .B1(n15128), .B2(n9649), .A(n9482), .ZN(n9495) );
  INV_X1 U12094 ( .A(n9495), .ZN(n14222) );
  NAND2_X1 U12095 ( .A1(n9483), .A2(n14222), .ZN(n14309) );
  OAI21_X1 U12096 ( .B1(n9496), .B2(n9494), .A(n14309), .ZN(n9500) );
  INV_X1 U12097 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14313) );
  NAND2_X1 U12098 ( .A1(n9484), .A2(n14313), .ZN(n9485) );
  NAND2_X1 U12099 ( .A1(n9507), .A2(n9485), .ZN(n14316) );
  INV_X1 U12100 ( .A(n14316), .ZN(n14912) );
  NAND2_X1 U12101 ( .A1(n14912), .A2(n9664), .ZN(n9491) );
  INV_X1 U12102 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U12103 ( .A1(n9658), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U12104 ( .A1(n9638), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9486) );
  OAI211_X1 U12105 ( .C1(n9488), .C2(n12508), .A(n9487), .B(n9486), .ZN(n9489)
         );
  INV_X1 U12106 ( .A(n9489), .ZN(n9490) );
  NOR2_X1 U12107 ( .A1(n14923), .A2(n9621), .ZN(n9492) );
  AOI21_X1 U12108 ( .B1(n15122), .B2(n9649), .A(n9492), .ZN(n9502) );
  AOI22_X1 U12109 ( .A1(n15122), .A2(n9634), .B1(n9649), .B2(n14643), .ZN(
        n9493) );
  XNOR2_X1 U12110 ( .A(n9493), .B(n10720), .ZN(n9501) );
  XOR2_X1 U12111 ( .A(n9502), .B(n9501), .Z(n14311) );
  NOR2_X1 U12112 ( .A1(n14220), .A2(n14219), .ZN(n14221) );
  OAI21_X1 U12113 ( .B1(n14221), .B2(n9495), .A(n14223), .ZN(n9498) );
  NAND3_X1 U12114 ( .A1(n9496), .A2(n9495), .A3(n9494), .ZN(n9497) );
  AND2_X1 U12115 ( .A1(n9498), .A2(n9497), .ZN(n9499) );
  INV_X1 U12116 ( .A(n9501), .ZN(n9504) );
  INV_X1 U12117 ( .A(n9502), .ZN(n9503) );
  NAND2_X1 U12118 ( .A1(n14889), .A2(n9634), .ZN(n9516) );
  INV_X1 U12119 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9506) );
  NAND2_X1 U12120 ( .A1(n9507), .A2(n9506), .ZN(n9508) );
  AND2_X1 U12121 ( .A1(n9523), .A2(n9508), .ZN(n14893) );
  NAND2_X1 U12122 ( .A1(n14893), .A2(n9664), .ZN(n9514) );
  INV_X1 U12123 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U12124 ( .A1(n9658), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9510) );
  NAND2_X1 U12125 ( .A1(n9638), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9509) );
  OAI211_X1 U12126 ( .C1(n9511), .C2(n12508), .A(n9510), .B(n9509), .ZN(n9512)
         );
  INV_X1 U12127 ( .A(n9512), .ZN(n9513) );
  NAND2_X1 U12128 ( .A1(n14870), .A2(n9649), .ZN(n9515) );
  NAND2_X1 U12129 ( .A1(n9516), .A2(n9515), .ZN(n9517) );
  XNOR2_X1 U12130 ( .A(n9517), .B(n9619), .ZN(n9520) );
  AND2_X1 U12131 ( .A1(n14870), .A2(n9648), .ZN(n9518) );
  AOI21_X1 U12132 ( .B1(n14889), .B2(n9649), .A(n9518), .ZN(n9519) );
  NAND2_X1 U12133 ( .A1(n9520), .A2(n9519), .ZN(n14329) );
  OAI21_X1 U12134 ( .B1(n9520), .B2(n9519), .A(n14329), .ZN(n14239) );
  NAND2_X1 U12135 ( .A1(n15111), .A2(n9634), .ZN(n9531) );
  INV_X1 U12136 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U12137 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  NAND2_X1 U12138 ( .A1(n9539), .A2(n9524), .ZN(n14875) );
  OR2_X1 U12139 ( .A1(n14875), .A2(n6433), .ZN(n9529) );
  INV_X1 U12140 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10816) );
  NAND2_X1 U12141 ( .A1(n9659), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U12142 ( .A1(n9638), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9525) );
  OAI211_X1 U12143 ( .C1(n12510), .C2(n10816), .A(n9526), .B(n9525), .ZN(n9527) );
  INV_X1 U12144 ( .A(n9527), .ZN(n9528) );
  NAND2_X1 U12145 ( .A1(n14642), .A2(n9649), .ZN(n9530) );
  NAND2_X1 U12146 ( .A1(n9531), .A2(n9530), .ZN(n9532) );
  XNOR2_X1 U12147 ( .A(n9532), .B(n9619), .ZN(n9534) );
  NOR2_X1 U12148 ( .A1(n14241), .A2(n9621), .ZN(n9533) );
  AOI21_X1 U12149 ( .B1(n15111), .B2(n9649), .A(n9533), .ZN(n9535) );
  NAND2_X1 U12150 ( .A1(n9534), .A2(n9535), .ZN(n14202) );
  INV_X1 U12151 ( .A(n9534), .ZN(n9537) );
  INV_X1 U12152 ( .A(n9535), .ZN(n9536) );
  NAND2_X1 U12153 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  NAND2_X1 U12154 ( .A1(n15104), .A2(n9634), .ZN(n9548) );
  INV_X1 U12155 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14206) );
  NAND2_X1 U12156 ( .A1(n9539), .A2(n14206), .ZN(n9540) );
  NAND2_X1 U12157 ( .A1(n14857), .A2(n9664), .ZN(n9546) );
  INV_X1 U12158 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U12159 ( .A1(n9638), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U12160 ( .A1(n9658), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9541) );
  OAI211_X1 U12161 ( .C1(n12508), .C2(n9543), .A(n9542), .B(n9541), .ZN(n9544)
         );
  INV_X1 U12162 ( .A(n9544), .ZN(n9545) );
  NAND2_X1 U12163 ( .A1(n14871), .A2(n9649), .ZN(n9547) );
  NAND2_X1 U12164 ( .A1(n9548), .A2(n9547), .ZN(n9549) );
  XNOR2_X1 U12165 ( .A(n9549), .B(n9619), .ZN(n9551) );
  AND2_X1 U12166 ( .A1(n14871), .A2(n9648), .ZN(n9550) );
  AOI21_X1 U12167 ( .B1(n15104), .B2(n9649), .A(n9550), .ZN(n9552) );
  NAND2_X1 U12168 ( .A1(n9551), .A2(n9552), .ZN(n14297) );
  INV_X1 U12169 ( .A(n9551), .ZN(n9554) );
  INV_X1 U12170 ( .A(n9552), .ZN(n9553) );
  NAND2_X1 U12171 ( .A1(n9554), .A2(n9553), .ZN(n9555) );
  AND2_X1 U12172 ( .A1(n14200), .A2(n14202), .ZN(n9558) );
  NAND2_X1 U12173 ( .A1(n14838), .A2(n9634), .ZN(n9570) );
  INV_X1 U12174 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14303) );
  NAND2_X1 U12175 ( .A1(n9561), .A2(n14303), .ZN(n9562) );
  NAND2_X1 U12176 ( .A1(n9578), .A2(n9562), .ZN(n14841) );
  INV_X1 U12177 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U12178 ( .A1(n9658), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9564) );
  NAND2_X1 U12179 ( .A1(n9638), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9563) );
  OAI211_X1 U12180 ( .C1(n9565), .C2(n12508), .A(n9564), .B(n9563), .ZN(n9566)
         );
  INV_X1 U12181 ( .A(n9566), .ZN(n9567) );
  AND2_X2 U12182 ( .A1(n9568), .A2(n9567), .ZN(n14266) );
  INV_X2 U12183 ( .A(n14266), .ZN(n14641) );
  NAND2_X1 U12184 ( .A1(n14641), .A2(n9644), .ZN(n9569) );
  NAND2_X1 U12185 ( .A1(n9570), .A2(n9569), .ZN(n9571) );
  XNOR2_X1 U12186 ( .A(n9571), .B(n9619), .ZN(n9573) );
  NOR2_X1 U12187 ( .A1(n14266), .A2(n9621), .ZN(n9572) );
  AOI21_X1 U12188 ( .B1(n14838), .B2(n9649), .A(n9572), .ZN(n9574) );
  NAND2_X1 U12189 ( .A1(n9573), .A2(n9574), .ZN(n14260) );
  INV_X1 U12190 ( .A(n9573), .ZN(n9576) );
  INV_X1 U12191 ( .A(n9574), .ZN(n9575) );
  NAND2_X1 U12192 ( .A1(n9576), .A2(n9575), .ZN(n9577) );
  INV_X1 U12193 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14269) );
  OR2_X2 U12194 ( .A1(n9578), .A2(n14269), .ZN(n9596) );
  NAND2_X1 U12195 ( .A1(n9578), .A2(n14269), .ZN(n9579) );
  NAND2_X1 U12196 ( .A1(n14268), .A2(n9664), .ZN(n9584) );
  INV_X1 U12197 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14822) );
  NAND2_X1 U12198 ( .A1(n9638), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U12199 ( .A1(n9658), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9580) );
  OAI211_X1 U12200 ( .C1(n12508), .C2(n14822), .A(n9581), .B(n9580), .ZN(n9582) );
  INV_X1 U12201 ( .A(n9582), .ZN(n9583) );
  INV_X1 U12202 ( .A(n14640), .ZN(n14802) );
  OAI22_X1 U12203 ( .A1(n14603), .A2(n9604), .B1(n14802), .B2(n9284), .ZN(
        n9585) );
  XNOR2_X1 U12204 ( .A(n9585), .B(n9619), .ZN(n9588) );
  NAND2_X1 U12205 ( .A1(n14640), .A2(n9648), .ZN(n9586) );
  NAND2_X1 U12206 ( .A1(n9588), .A2(n9589), .ZN(n9594) );
  INV_X1 U12207 ( .A(n9588), .ZN(n9591) );
  INV_X1 U12208 ( .A(n9589), .ZN(n9590) );
  NAND2_X1 U12209 ( .A1(n9591), .A2(n9590), .ZN(n9592) );
  INV_X1 U12210 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14366) );
  NAND2_X1 U12211 ( .A1(n9596), .A2(n14366), .ZN(n9597) );
  NAND2_X1 U12212 ( .A1(n9636), .A2(n9597), .ZN(n14808) );
  INV_X1 U12213 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9600) );
  NAND2_X1 U12214 ( .A1(n9658), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9599) );
  NAND2_X1 U12215 ( .A1(n9638), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9598) );
  OAI211_X1 U12216 ( .C1(n9600), .C2(n12508), .A(n9599), .B(n9598), .ZN(n9601)
         );
  INV_X1 U12217 ( .A(n9601), .ZN(n9602) );
  NAND2_X2 U12218 ( .A1(n9603), .A2(n9602), .ZN(n14639) );
  OAI22_X1 U12219 ( .A1(n14811), .A2(n9604), .B1(n14522), .B2(n9284), .ZN(
        n9605) );
  XNOR2_X1 U12220 ( .A(n9605), .B(n10720), .ZN(n9609) );
  NAND2_X1 U12221 ( .A1(n14639), .A2(n9648), .ZN(n9606) );
  NAND2_X1 U12222 ( .A1(n9607), .A2(n9606), .ZN(n9608) );
  NAND2_X1 U12223 ( .A1(n15082), .A2(n9634), .ZN(n9618) );
  NAND2_X1 U12224 ( .A1(n12437), .A2(n9664), .ZN(n9616) );
  INV_X1 U12225 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U12226 ( .A1(n9658), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9612) );
  NAND2_X1 U12227 ( .A1(n9638), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9611) );
  OAI211_X1 U12228 ( .C1(n9613), .C2(n12508), .A(n9612), .B(n9611), .ZN(n9614)
         );
  INV_X1 U12229 ( .A(n9614), .ZN(n9615) );
  AND2_X2 U12230 ( .A1(n9616), .A2(n9615), .ZN(n14365) );
  OR2_X1 U12231 ( .A1(n14365), .A2(n9284), .ZN(n9617) );
  NAND2_X1 U12232 ( .A1(n9618), .A2(n9617), .ZN(n9620) );
  XNOR2_X1 U12233 ( .A(n9620), .B(n9619), .ZN(n9624) );
  INV_X1 U12234 ( .A(n9624), .ZN(n9626) );
  NOR2_X1 U12235 ( .A1(n14365), .A2(n9621), .ZN(n9622) );
  AOI21_X1 U12236 ( .B1(n15082), .B2(n9649), .A(n9622), .ZN(n9623) );
  INV_X1 U12237 ( .A(n9623), .ZN(n9625) );
  INV_X1 U12238 ( .A(n10380), .ZN(n9652) );
  INV_X1 U12239 ( .A(n10458), .ZN(n14537) );
  AND2_X1 U12240 ( .A1(n15363), .A2(n14537), .ZN(n9627) );
  NAND2_X1 U12241 ( .A1(n11266), .A2(n9627), .ZN(n9628) );
  NOR2_X1 U12242 ( .A1(n11262), .A2(n9628), .ZN(n9633) );
  AND2_X1 U12243 ( .A1(n9629), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9630) );
  OR2_X1 U12244 ( .A1(n10460), .A2(n9630), .ZN(n9632) );
  INV_X1 U12245 ( .A(n10461), .ZN(n9631) );
  NAND2_X1 U12246 ( .A1(n15077), .A2(n9634), .ZN(n9646) );
  INV_X1 U12247 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10384) );
  INV_X1 U12248 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n10764) );
  OAI21_X1 U12249 ( .B1(n9636), .B2(n10384), .A(n10764), .ZN(n9637) );
  NAND2_X1 U12250 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9635) );
  NAND2_X1 U12251 ( .A1(n12597), .A2(n9664), .ZN(n9643) );
  INV_X1 U12252 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10756) );
  NAND2_X1 U12253 ( .A1(n9659), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12254 ( .A1(n9638), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9639) );
  OAI211_X1 U12255 ( .C1(n6440), .C2(n10756), .A(n9640), .B(n9639), .ZN(n9641)
         );
  INV_X1 U12256 ( .A(n9641), .ZN(n9642) );
  NAND2_X1 U12257 ( .A1(n14637), .A2(n9644), .ZN(n9645) );
  NAND2_X1 U12258 ( .A1(n9646), .A2(n9645), .ZN(n9647) );
  XNOR2_X1 U12259 ( .A(n9647), .B(n10720), .ZN(n9651) );
  AOI22_X1 U12260 ( .A1(n15077), .A2(n9649), .B1(n9648), .B2(n14637), .ZN(
        n9650) );
  XNOR2_X1 U12261 ( .A(n9651), .B(n9650), .ZN(n9656) );
  NAND3_X1 U12262 ( .A1(n9652), .A2(n14370), .A3(n9656), .ZN(n9677) );
  INV_X1 U12263 ( .A(n9656), .ZN(n9654) );
  INV_X1 U12264 ( .A(n9655), .ZN(n9653) );
  NAND3_X1 U12265 ( .A1(n9656), .A2(n9655), .A3(n14370), .ZN(n9674) );
  INV_X1 U12266 ( .A(n14671), .ZN(n10608) );
  AND2_X1 U12267 ( .A1(n14368), .A2(n15223), .ZN(n14377) );
  INV_X1 U12268 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9662) );
  NAND2_X1 U12269 ( .A1(n9658), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U12270 ( .A1(n9659), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9660) );
  OAI211_X1 U12271 ( .C1(n9662), .C2(n9288), .A(n9661), .B(n9660), .ZN(n9663)
         );
  NAND2_X1 U12272 ( .A1(n14368), .A2(n15222), .ZN(n14374) );
  NAND2_X1 U12273 ( .A1(n9665), .A2(n11263), .ZN(n9666) );
  NAND2_X1 U12274 ( .A1(n9666), .A2(n11264), .ZN(n10652) );
  AND2_X1 U12275 ( .A1(n9667), .A2(n10393), .ZN(n9668) );
  NAND2_X1 U12276 ( .A1(n10652), .A2(n9668), .ZN(n9669) );
  OR2_X1 U12277 ( .A1(n10457), .A2(n6428), .ZN(n14560) );
  AOI21_X1 U12278 ( .B1(n9669), .B2(P1_STATE_REG_SCAN_IN), .A(n14627), .ZN(
        n14353) );
  AOI22_X1 U12279 ( .A1(n12597), .A2(n14242), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(n6428), .ZN(n9670) );
  OAI21_X1 U12280 ( .B1(n14548), .B2(n14374), .A(n9670), .ZN(n9672) );
  INV_X1 U12281 ( .A(n15077), .ZN(n12504) );
  NAND2_X1 U12282 ( .A1(n10652), .A2(n11266), .ZN(n14308) );
  NOR2_X1 U12283 ( .A1(n12504), .A2(n14380), .ZN(n9671) );
  AOI211_X1 U12284 ( .C1(n14377), .C2(n14638), .A(n9672), .B(n9671), .ZN(n9673) );
  AOI21_X1 U12285 ( .B1(n10380), .B2(n7821), .A(n9675), .ZN(n9676) );
  NAND2_X1 U12286 ( .A1(n9677), .A2(n9676), .ZN(P1_U3220) );
  NOR2_X2 U12287 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n9685) );
  NAND2_X1 U12288 ( .A1(n10200), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9688) );
  NAND3_X1 U12289 ( .A1(n9705), .A2(n9704), .A3(n9683), .ZN(n9697) );
  NAND2_X1 U12290 ( .A1(n9697), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9696) );
  INV_X1 U12291 ( .A(n9697), .ZN(n9699) );
  INV_X1 U12292 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9698) );
  NAND2_X1 U12293 ( .A1(n9699), .A2(n9698), .ZN(n9701) );
  NAND2_X1 U12294 ( .A1(n9700), .A2(n9701), .ZN(n12091) );
  XNOR2_X1 U12295 ( .A(n12091), .B(P3_B_REG_SCAN_IN), .ZN(n9707) );
  NAND2_X1 U12296 ( .A1(n9701), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9702) );
  MUX2_X1 U12297 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9702), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9706) );
  NAND2_X1 U12298 ( .A1(n9706), .A2(n9719), .ZN(n12293) );
  NAND2_X1 U12299 ( .A1(n9719), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9709) );
  INV_X1 U12300 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9708) );
  XNOR2_X1 U12301 ( .A(n9709), .B(n9708), .ZN(n13523) );
  INV_X1 U12302 ( .A(n12091), .ZN(n9712) );
  NAND2_X1 U12303 ( .A1(n9713), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9714) );
  MUX2_X1 U12304 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9714), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n9715) );
  NAND2_X1 U12305 ( .A1(n9715), .A2(n10200), .ZN(n11540) );
  NOR2_X2 U12306 ( .A1(n10021), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n10039) );
  INV_X1 U12307 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n10058) );
  INV_X1 U12308 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9717) );
  NAND2_X4 U12309 ( .A1(n9718), .A2(n12800), .ZN(n11041) );
  INV_X1 U12310 ( .A(n10301), .ZN(n9804) );
  INV_X1 U12311 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15607) );
  OR2_X1 U12312 ( .A1(n9804), .A2(n15607), .ZN(n9731) );
  INV_X1 U12313 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9724) );
  INV_X1 U12314 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11050) );
  AND2_X1 U12315 ( .A1(n9727), .A2(n9726), .ZN(n9730) );
  INV_X1 U12316 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9736) );
  NAND2_X1 U12317 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9735) );
  XNOR2_X2 U12318 ( .A(n9735), .B(n9736), .ZN(n10978) );
  OR2_X1 U12319 ( .A1(n10911), .A2(n10978), .ZN(n9742) );
  NAND2_X1 U12320 ( .A1(n9738), .A2(n9753), .ZN(n9741) );
  INV_X1 U12321 ( .A(n9753), .ZN(n9739) );
  AND2_X1 U12322 ( .A1(n9741), .A2(n9760), .ZN(n10414) );
  OAI21_X1 U12323 ( .B1(n11041), .B2(n9757), .A(n12806), .ZN(n9744) );
  INV_X1 U12324 ( .A(n9745), .ZN(n9743) );
  NAND2_X1 U12325 ( .A1(n9745), .A2(n9757), .ZN(n9746) );
  NAND2_X1 U12326 ( .A1(n12093), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9750) );
  NAND2_X1 U12327 ( .A1(n10165), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9749) );
  INV_X1 U12328 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11428) );
  OR2_X1 U12329 ( .A1(n9804), .A2(n11428), .ZN(n9748) );
  INV_X1 U12330 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10918) );
  OR2_X1 U12331 ( .A1(n9828), .A2(n10918), .ZN(n9747) );
  INV_X1 U12332 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11429) );
  NAND2_X1 U12333 ( .A1(n9751), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9752) );
  AND2_X1 U12334 ( .A1(n9753), .A2(n9752), .ZN(n9754) );
  OAI21_X1 U12335 ( .B1(n9755), .B2(n9754), .A(n7891), .ZN(n13524) );
  INV_X1 U12336 ( .A(n13524), .ZN(n9756) );
  MUX2_X1 U12337 ( .A(n11429), .B(n9756), .S(n10911), .Z(n11423) );
  NAND2_X1 U12338 ( .A1(n10258), .A2(n11041), .ZN(n9758) );
  NAND2_X1 U12339 ( .A1(n15596), .A2(n7150), .ZN(n15594) );
  NAND2_X1 U12340 ( .A1(n10415), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9759) );
  OAI21_X1 U12341 ( .B1(n9762), .B2(n9761), .A(n9771), .ZN(n10428) );
  OR2_X1 U12342 ( .A1(n9877), .A2(n10428), .ZN(n9766) );
  OR2_X1 U12343 ( .A1(n10911), .A2(n7009), .ZN(n9764) );
  XNOR2_X1 U12344 ( .A(n11041), .B(n15573), .ZN(n9785) );
  NAND2_X1 U12345 ( .A1(n10165), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9770) );
  NAND2_X1 U12346 ( .A1(n12093), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9769) );
  INV_X1 U12347 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10919) );
  OR2_X1 U12348 ( .A1(n9828), .A2(n10919), .ZN(n9768) );
  INV_X1 U12349 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15592) );
  OR2_X1 U12350 ( .A1(n12269), .A2(n15592), .ZN(n9767) );
  XNOR2_X1 U12351 ( .A(n9785), .B(n10259), .ZN(n11096) );
  NAND2_X1 U12352 ( .A1(n11095), .A2(n11096), .ZN(n11094) );
  OR2_X1 U12353 ( .A1(n12761), .A2(SI_3_), .ZN(n9779) );
  OR2_X1 U12354 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  NAND2_X1 U12355 ( .A1(n9791), .A2(n9774), .ZN(n10424) );
  OR2_X1 U12356 ( .A1(n9877), .A2(n10424), .ZN(n9778) );
  INV_X1 U12357 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U12358 ( .A1(n9796), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9776) );
  OR2_X1 U12359 ( .A1(n10911), .A2(n10924), .ZN(n9777) );
  XNOR2_X1 U12360 ( .A(n11041), .B(n11498), .ZN(n9787) );
  NAND2_X1 U12361 ( .A1(n9854), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9784) );
  OR2_X1 U12362 ( .A1(n9826), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9783) );
  OR2_X1 U12363 ( .A1(n12269), .A2(n7511), .ZN(n9782) );
  INV_X1 U12364 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n9780) );
  OR2_X1 U12365 ( .A1(n9822), .A2(n9780), .ZN(n9781) );
  XNOR2_X1 U12366 ( .A(n9787), .B(n12979), .ZN(n11137) );
  NAND2_X1 U12367 ( .A1(n9785), .A2(n11494), .ZN(n11138) );
  AND2_X1 U12368 ( .A1(n11137), .A2(n11138), .ZN(n9786) );
  INV_X1 U12369 ( .A(n9787), .ZN(n9788) );
  NAND2_X1 U12370 ( .A1(n9788), .A2(n12979), .ZN(n9789) );
  OR2_X1 U12371 ( .A1(n12761), .A2(SI_4_), .ZN(n9800) );
  NAND2_X1 U12372 ( .A1(n10447), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9792) );
  OR2_X1 U12373 ( .A1(n9794), .A2(n9793), .ZN(n9795) );
  NAND2_X1 U12374 ( .A1(n9815), .A2(n9795), .ZN(n10430) );
  OR2_X1 U12375 ( .A1(n9877), .A2(n10430), .ZN(n9799) );
  NAND2_X1 U12376 ( .A1(n9817), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9797) );
  OR2_X1 U12377 ( .A1(n10911), .A2(n10979), .ZN(n9798) );
  XNOR2_X1 U12378 ( .A(n11041), .B(n15624), .ZN(n9809) );
  INV_X1 U12379 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n9801) );
  INV_X1 U12380 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10901) );
  OR2_X1 U12381 ( .A1(n9828), .A2(n10901), .ZN(n9807) );
  NAND2_X1 U12382 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9803) );
  AND2_X1 U12383 ( .A1(n9824), .A2(n9803), .ZN(n11731) );
  OR2_X1 U12384 ( .A1(n9826), .A2(n11731), .ZN(n9806) );
  INV_X1 U12385 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10945) );
  OR2_X1 U12386 ( .A1(n9804), .A2(n10945), .ZN(n9805) );
  NAND2_X1 U12387 ( .A1(n9809), .A2(n11784), .ZN(n9813) );
  INV_X1 U12388 ( .A(n9809), .ZN(n9810) );
  NAND2_X1 U12389 ( .A1(n9810), .A2(n12978), .ZN(n9811) );
  NAND2_X1 U12390 ( .A1(n9813), .A2(n9811), .ZN(n11406) );
  XNOR2_X1 U12391 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9816) );
  XNOR2_X1 U12392 ( .A(n9836), .B(n9816), .ZN(n10426) );
  OR2_X1 U12393 ( .A1(n9877), .A2(n10426), .ZN(n9821) );
  OR2_X1 U12394 ( .A1(n12761), .A2(SI_5_), .ZN(n9820) );
  OAI21_X1 U12395 ( .B1(n9817), .B2(P3_IR_REG_4__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9818) );
  XNOR2_X1 U12396 ( .A(n9818), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10934) );
  OR2_X1 U12397 ( .A1(n10911), .A2(n10934), .ZN(n9819) );
  XNOR2_X1 U12398 ( .A(n11041), .B(n11774), .ZN(n9871) );
  INV_X2 U12399 ( .A(n9822), .ZN(n12266) );
  NAND2_X1 U12400 ( .A1(n12266), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U12401 ( .A1(n9824), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9825) );
  AND2_X1 U12402 ( .A1(n9880), .A2(n9825), .ZN(n11775) );
  OR2_X1 U12403 ( .A1(n9826), .A2(n11775), .ZN(n9830) );
  INV_X1 U12404 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9827) );
  OR2_X1 U12405 ( .A1(n9828), .A2(n9827), .ZN(n9829) );
  INV_X1 U12406 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9832) );
  OR2_X1 U12407 ( .A1(n12269), .A2(n9832), .ZN(n9833) );
  XNOR2_X1 U12408 ( .A(n9871), .B(n12977), .ZN(n11561) );
  NAND2_X1 U12409 ( .A1(n10441), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9835) );
  NAND2_X1 U12410 ( .A1(n10439), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U12411 ( .A1(n10418), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U12412 ( .A1(n9838), .A2(n9837), .ZN(n9875) );
  NAND2_X1 U12413 ( .A1(n10445), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U12414 ( .A1(n10480), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9839) );
  NAND2_X1 U12415 ( .A1(n10451), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9901) );
  INV_X1 U12416 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10449) );
  NAND2_X1 U12417 ( .A1(n10449), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9841) );
  NAND2_X1 U12418 ( .A1(n9901), .A2(n9841), .ZN(n9898) );
  XNOR2_X1 U12419 ( .A(n9900), .B(n9898), .ZN(n10419) );
  INV_X1 U12420 ( .A(n9877), .ZN(n9903) );
  NAND2_X1 U12421 ( .A1(n10419), .A2(n9903), .ZN(n9846) );
  INV_X2 U12422 ( .A(n10911), .ZN(n10093) );
  OR2_X1 U12423 ( .A1(n9872), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n9866) );
  INV_X1 U12424 ( .A(n9866), .ZN(n9843) );
  NAND2_X1 U12425 ( .A1(n9843), .A2(n9842), .ZN(n9904) );
  NAND2_X1 U12426 ( .A1(n9904), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9844) );
  XNOR2_X1 U12427 ( .A(n11041), .B(n12842), .ZN(n9893) );
  NAND2_X1 U12428 ( .A1(n12266), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9853) );
  INV_X1 U12429 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n12080) );
  OR2_X1 U12430 ( .A1(n9828), .A2(n12080), .ZN(n9852) );
  NAND2_X1 U12431 ( .A1(n9856), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9849) );
  AND2_X1 U12432 ( .A1(n9912), .A2(n9849), .ZN(n12200) );
  OR2_X1 U12433 ( .A1(n6957), .A2(n12200), .ZN(n9851) );
  INV_X1 U12434 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11214) );
  OR2_X1 U12435 ( .A1(n12269), .A2(n11214), .ZN(n9850) );
  NAND2_X1 U12436 ( .A1(n9854), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9861) );
  NAND2_X1 U12437 ( .A1(n10301), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U12438 ( .A1(n9882), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9855) );
  AND2_X1 U12439 ( .A1(n9856), .A2(n9855), .ZN(n12082) );
  OR2_X1 U12440 ( .A1(n6957), .A2(n12082), .ZN(n9859) );
  INV_X1 U12441 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n9857) );
  OR2_X1 U12442 ( .A1(n9822), .A2(n9857), .ZN(n9858) );
  NAND4_X2 U12443 ( .A1(n9861), .A2(n9860), .A3(n9859), .A4(n9858), .ZN(n12837) );
  OR2_X1 U12444 ( .A1(n9863), .A2(n9862), .ZN(n9864) );
  NAND2_X1 U12445 ( .A1(n9865), .A2(n9864), .ZN(n10407) );
  NAND2_X1 U12446 ( .A1(n10407), .A2(n9903), .ZN(n9870) );
  OR2_X1 U12447 ( .A1(n12761), .A2(SI_7_), .ZN(n9869) );
  NAND2_X1 U12448 ( .A1(n9866), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9867) );
  XNOR2_X1 U12449 ( .A(n9867), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11063) );
  OR2_X1 U12450 ( .A1(n10911), .A2(n11063), .ZN(n9868) );
  XNOR2_X1 U12451 ( .A(n12835), .B(n11041), .ZN(n9892) );
  NAND2_X1 U12452 ( .A1(n9871), .A2(n10316), .ZN(n11831) );
  NAND2_X1 U12453 ( .A1(n9872), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9874) );
  INV_X1 U12454 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9873) );
  XNOR2_X1 U12455 ( .A(n9874), .B(n9873), .ZN(n11130) );
  OR2_X1 U12456 ( .A1(n12761), .A2(n6778), .ZN(n9879) );
  XNOR2_X1 U12457 ( .A(n9876), .B(n9875), .ZN(n10405) );
  OR2_X1 U12458 ( .A1(n9877), .A2(n10405), .ZN(n9878) );
  OAI211_X1 U12459 ( .C1(n6924), .C2(n11130), .A(n9879), .B(n9878), .ZN(n12721) );
  XNOR2_X1 U12460 ( .A(n11041), .B(n12721), .ZN(n11832) );
  NAND2_X1 U12461 ( .A1(n10165), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9886) );
  INV_X1 U12462 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10906) );
  OR2_X1 U12463 ( .A1(n9828), .A2(n10906), .ZN(n9885) );
  NAND2_X1 U12464 ( .A1(n9880), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9881) );
  AND2_X1 U12465 ( .A1(n9882), .A2(n9881), .ZN(n11512) );
  OR2_X1 U12466 ( .A1(n6957), .A2(n11512), .ZN(n9884) );
  INV_X1 U12467 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11511) );
  OR2_X1 U12468 ( .A1(n12269), .A2(n11511), .ZN(n9883) );
  NAND2_X1 U12469 ( .A1(n11832), .A2(n11785), .ZN(n9887) );
  NAND3_X1 U12470 ( .A1(n9892), .A2(n11831), .A3(n9887), .ZN(n9888) );
  NOR2_X1 U12471 ( .A1(n12139), .A2(n9888), .ZN(n9889) );
  INV_X1 U12472 ( .A(n12837), .ZN(n9890) );
  INV_X1 U12473 ( .A(n9892), .ZN(n12137) );
  OAI21_X1 U12474 ( .B1(n12139), .B2(n9890), .A(n12137), .ZN(n9896) );
  INV_X1 U12475 ( .A(n11832), .ZN(n9891) );
  NAND2_X1 U12476 ( .A1(n9891), .A2(n12976), .ZN(n11833) );
  OAI21_X1 U12477 ( .B1(n12139), .B2(n11833), .A(n9892), .ZN(n9895) );
  INV_X1 U12478 ( .A(n9893), .ZN(n9894) );
  INV_X1 U12479 ( .A(n12843), .ZN(n11855) );
  INV_X1 U12480 ( .A(n9898), .ZN(n9899) );
  INV_X1 U12481 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10471) );
  NAND2_X1 U12482 ( .A1(n10471), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9921) );
  INV_X1 U12483 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10484) );
  NAND2_X1 U12484 ( .A1(n10484), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9902) );
  XNOR2_X1 U12485 ( .A(n9920), .B(n9919), .ZN(n10423) );
  NAND2_X1 U12486 ( .A1(n10423), .A2(n12758), .ZN(n9910) );
  INV_X1 U12487 ( .A(SI_9_), .ZN(n10422) );
  INV_X1 U12488 ( .A(n9904), .ZN(n9906) );
  INV_X1 U12489 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U12490 ( .A1(n9906), .A2(n9905), .ZN(n9923) );
  NAND2_X1 U12491 ( .A1(n9923), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9908) );
  XNOR2_X1 U12492 ( .A(n9908), .B(n9907), .ZN(n11229) );
  AOI22_X1 U12493 ( .A1(n10074), .A2(n10422), .B1(n10093), .B2(n11229), .ZN(
        n9909) );
  XNOR2_X1 U12494 ( .A(n12069), .B(n11041), .ZN(n9934) );
  NAND2_X1 U12495 ( .A1(n10165), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9918) );
  NAND2_X1 U12496 ( .A1(n9854), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U12497 ( .A1(n9912), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9913) );
  AND2_X1 U12498 ( .A1(n9928), .A2(n9913), .ZN(n11856) );
  OR2_X1 U12499 ( .A1(n6957), .A2(n11856), .ZN(n9916) );
  INV_X1 U12500 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n9914) );
  OR2_X1 U12501 ( .A1(n12269), .A2(n9914), .ZN(n9915) );
  NAND4_X1 U12502 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(n12975) );
  XNOR2_X1 U12503 ( .A(n9934), .B(n12975), .ZN(n11863) );
  INV_X1 U12504 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10476) );
  NAND2_X1 U12505 ( .A1(n10476), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9941) );
  INV_X1 U12506 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10773) );
  NAND2_X1 U12507 ( .A1(n10773), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9922) );
  XNOR2_X1 U12508 ( .A(n9940), .B(n9939), .ZN(n10435) );
  NAND2_X1 U12509 ( .A1(n10435), .A2(n12758), .ZN(n9927) );
  INV_X1 U12510 ( .A(SI_10_), .ZN(n10434) );
  NAND2_X1 U12511 ( .A1(n9944), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9925) );
  INV_X1 U12512 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9924) );
  XNOR2_X1 U12513 ( .A(n9925), .B(n9924), .ZN(n11808) );
  AOI22_X1 U12514 ( .A1(n10074), .A2(n10434), .B1(n10093), .B2(n11808), .ZN(
        n9926) );
  XNOR2_X1 U12515 ( .A(n12852), .B(n12496), .ZN(n9937) );
  NAND2_X1 U12516 ( .A1(n12266), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9933) );
  INV_X1 U12517 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11656) );
  OR2_X1 U12518 ( .A1(n9828), .A2(n11656), .ZN(n9932) );
  NAND2_X1 U12519 ( .A1(n9928), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9929) );
  AND2_X1 U12520 ( .A1(n9949), .A2(n9929), .ZN(n12156) );
  OR2_X1 U12521 ( .A1(n6957), .A2(n12156), .ZN(n9931) );
  INV_X1 U12522 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11657) );
  OR2_X1 U12523 ( .A1(n12269), .A2(n11657), .ZN(n9930) );
  XNOR2_X1 U12524 ( .A(n9937), .B(n12369), .ZN(n11907) );
  INV_X1 U12525 ( .A(n9934), .ZN(n9935) );
  INV_X1 U12526 ( .A(n12975), .ZN(n11910) );
  NAND2_X1 U12527 ( .A1(n9935), .A2(n11910), .ZN(n11905) );
  AND2_X1 U12528 ( .A1(n11907), .A2(n11905), .ZN(n9936) );
  NAND2_X1 U12529 ( .A1(n9937), .A2(n12974), .ZN(n9938) );
  NAND2_X1 U12530 ( .A1(n9940), .A2(n9939), .ZN(n9942) );
  NAND2_X1 U12531 ( .A1(n10489), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U12532 ( .A1(n10487), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9943) );
  XNOR2_X1 U12533 ( .A(n9956), .B(n9955), .ZN(n10455) );
  NAND2_X1 U12534 ( .A1(n10455), .A2(n12758), .ZN(n9948) );
  OAI21_X1 U12535 ( .B1(n9944), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9946) );
  INV_X1 U12536 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9945) );
  XNOR2_X1 U12537 ( .A(n9946), .B(n9945), .ZN(n11875) );
  AOI22_X1 U12538 ( .A1(n10074), .A2(n10454), .B1(n10093), .B2(n11875), .ZN(
        n9947) );
  XNOR2_X1 U12539 ( .A(n12252), .B(n12496), .ZN(n12363) );
  NAND2_X1 U12540 ( .A1(n12266), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9954) );
  NAND2_X1 U12541 ( .A1(n9854), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U12542 ( .A1(n9949), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9950) );
  AND2_X1 U12543 ( .A1(n9966), .A2(n9950), .ZN(n12372) );
  OR2_X1 U12544 ( .A1(n6957), .A2(n12372), .ZN(n9952) );
  INV_X1 U12545 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12251) );
  OR2_X1 U12546 ( .A1(n12269), .A2(n12251), .ZN(n9951) );
  NAND4_X1 U12547 ( .A1(n9954), .A2(n9953), .A3(n9952), .A4(n9951), .ZN(n12973) );
  AND2_X1 U12548 ( .A1(n12363), .A2(n12973), .ZN(n9974) );
  NAND2_X1 U12549 ( .A1(n10581), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U12550 ( .A1(n10579), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U12551 ( .A1(n9980), .A2(n9958), .ZN(n9977) );
  XNOR2_X1 U12552 ( .A(n9979), .B(n9977), .ZN(n10477) );
  NAND2_X1 U12553 ( .A1(n10477), .A2(n12758), .ZN(n9964) );
  NAND2_X1 U12554 ( .A1(n9959), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9960) );
  MUX2_X1 U12555 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9960), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9961) );
  INV_X1 U12556 ( .A(n9961), .ZN(n9962) );
  NOR2_X1 U12557 ( .A1(n9962), .A2(n9982), .ZN(n12980) );
  AOI22_X1 U12558 ( .A1(n10074), .A2(SI_12_), .B1(n10093), .B2(n12980), .ZN(
        n9963) );
  XNOR2_X1 U12559 ( .A(n12665), .B(n12496), .ZN(n9975) );
  NAND2_X1 U12560 ( .A1(n9854), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9971) );
  INV_X1 U12561 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n9965) );
  OR2_X1 U12562 ( .A1(n9822), .A2(n9965), .ZN(n9970) );
  INV_X1 U12563 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n10829) );
  NAND2_X1 U12564 ( .A1(n9966), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9967) );
  AND2_X1 U12565 ( .A1(n9989), .A2(n9967), .ZN(n12663) );
  OR2_X1 U12566 ( .A1(n6957), .A2(n12663), .ZN(n9969) );
  INV_X1 U12567 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12338) );
  OR2_X1 U12568 ( .A1(n12269), .A2(n12338), .ZN(n9968) );
  NAND2_X1 U12569 ( .A1(n9975), .A2(n12383), .ZN(n12651) );
  OAI21_X1 U12570 ( .B1(n12363), .B2(n12973), .A(n12651), .ZN(n9972) );
  INV_X1 U12571 ( .A(n9972), .ZN(n9973) );
  INV_X1 U12572 ( .A(n9975), .ZN(n9976) );
  INV_X1 U12573 ( .A(n12383), .ZN(n12972) );
  NAND2_X1 U12574 ( .A1(n9976), .A2(n12972), .ZN(n12652) );
  INV_X1 U12575 ( .A(n9977), .ZN(n9978) );
  NAND2_X1 U12576 ( .A1(n10018), .A2(n10681), .ZN(n9997) );
  XNOR2_X1 U12577 ( .A(n9998), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10625) );
  NAND2_X1 U12578 ( .A1(n10625), .A2(n12758), .ZN(n9986) );
  INV_X1 U12579 ( .A(n9982), .ZN(n9983) );
  NAND2_X1 U12580 ( .A1(n9983), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9984) );
  XNOR2_X1 U12581 ( .A(n9984), .B(P3_IR_REG_13__SCAN_IN), .ZN(n13018) );
  AOI22_X1 U12582 ( .A1(n10074), .A2(SI_13_), .B1(n10093), .B2(n13018), .ZN(
        n9985) );
  XNOR2_X1 U12583 ( .A(n13492), .B(n12496), .ZN(n12324) );
  NAND2_X1 U12584 ( .A1(n12266), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9994) );
  INV_X1 U12585 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12984) );
  OR2_X1 U12586 ( .A1(n9828), .A2(n12984), .ZN(n9993) );
  INV_X1 U12587 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U12588 ( .A1(n9989), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9990) );
  AND2_X1 U12589 ( .A1(n10005), .A2(n9990), .ZN(n12379) );
  OR2_X1 U12590 ( .A1(n6957), .A2(n12379), .ZN(n9992) );
  INV_X1 U12591 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12385) );
  OR2_X1 U12592 ( .A1(n12269), .A2(n12385), .ZN(n9991) );
  NAND2_X1 U12593 ( .A1(n12324), .A2(n13354), .ZN(n9996) );
  INV_X1 U12594 ( .A(n12324), .ZN(n9995) );
  INV_X1 U12595 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11199) );
  NAND2_X1 U12596 ( .A1(n11199), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n10019) );
  INV_X1 U12597 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11201) );
  NAND2_X1 U12598 ( .A1(n11201), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U12599 ( .A1(n10019), .A2(n9999), .ZN(n10015) );
  XNOR2_X1 U12600 ( .A(n10000), .B(n10015), .ZN(n10674) );
  NAND2_X1 U12601 ( .A1(n10674), .A2(n12758), .ZN(n10004) );
  NAND2_X1 U12602 ( .A1(n10001), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10002) );
  XNOR2_X1 U12603 ( .A(n10002), .B(P3_IR_REG_14__SCAN_IN), .ZN(n13028) );
  AOI22_X1 U12604 ( .A1(n10074), .A2(SI_14_), .B1(n10093), .B2(n13028), .ZN(
        n10003) );
  XNOR2_X1 U12605 ( .A(n13487), .B(n12487), .ZN(n10011) );
  NAND2_X1 U12606 ( .A1(n10005), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n10006) );
  NAND2_X1 U12607 ( .A1(n10028), .A2(n10006), .ZN(n13346) );
  NAND2_X1 U12608 ( .A1(n13346), .A2(n12093), .ZN(n10010) );
  NAND2_X1 U12609 ( .A1(n10165), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n10009) );
  INV_X1 U12610 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13006) );
  OR2_X1 U12611 ( .A1(n9828), .A2(n13006), .ZN(n10008) );
  INV_X1 U12612 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13359) );
  OR2_X1 U12613 ( .A1(n12269), .A2(n13359), .ZN(n10007) );
  NAND4_X1 U12614 ( .A1(n10010), .A2(n10009), .A3(n10008), .A4(n10007), .ZN(
        n12970) );
  NOR2_X1 U12615 ( .A1(n10011), .A2(n12970), .ZN(n10012) );
  AOI21_X1 U12616 ( .B1(n10011), .B2(n12970), .A(n10012), .ZN(n12620) );
  INV_X1 U12617 ( .A(n10012), .ZN(n10013) );
  AND2_X1 U12618 ( .A1(n10681), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n10017) );
  AND2_X1 U12619 ( .A1(n10679), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n10014) );
  NOR2_X1 U12620 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  NAND2_X1 U12621 ( .A1(n11303), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U12622 ( .A1(n11305), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n10020) );
  NAND2_X1 U12623 ( .A1(n10037), .A2(n10020), .ZN(n10035) );
  XNOR2_X1 U12624 ( .A(n10036), .B(n10035), .ZN(n10628) );
  NAND2_X1 U12625 ( .A1(n10628), .A2(n12758), .ZN(n10025) );
  NAND2_X1 U12626 ( .A1(n10021), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10023) );
  INV_X1 U12627 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n10022) );
  XNOR2_X1 U12628 ( .A(n10023), .B(n10022), .ZN(n13058) );
  INV_X1 U12629 ( .A(n13058), .ZN(n13066) );
  AOI22_X1 U12630 ( .A1(n10074), .A2(SI_15_), .B1(n10093), .B2(n13066), .ZN(
        n10024) );
  XNOR2_X1 U12631 ( .A(n13410), .B(n12496), .ZN(n12738) );
  INV_X1 U12632 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n10026) );
  NAND2_X1 U12633 ( .A1(n10028), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U12634 ( .A1(n10044), .A2(n10029), .ZN(n13338) );
  NAND2_X1 U12635 ( .A1(n13338), .A2(n12093), .ZN(n10032) );
  AOI22_X1 U12636 ( .A1(n10165), .A2(P3_REG0_REG_15__SCAN_IN), .B1(n9854), 
        .B2(P3_REG1_REG_15__SCAN_IN), .ZN(n10031) );
  INV_X1 U12637 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13036) );
  OR2_X1 U12638 ( .A1(n12269), .A2(n13036), .ZN(n10030) );
  INV_X1 U12639 ( .A(n13355), .ZN(n12969) );
  NAND2_X1 U12640 ( .A1(n12738), .A2(n13355), .ZN(n10034) );
  NAND2_X1 U12641 ( .A1(n11298), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U12642 ( .A1(n11301), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U12643 ( .A1(n10055), .A2(n10038), .ZN(n10052) );
  XNOR2_X1 U12644 ( .A(n10054), .B(n10052), .ZN(n10732) );
  NAND2_X1 U12645 ( .A1(n10732), .A2(n12758), .ZN(n10043) );
  INV_X1 U12646 ( .A(n10039), .ZN(n10040) );
  NAND2_X1 U12647 ( .A1(n10040), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10041) );
  XNOR2_X1 U12648 ( .A(n10041), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U12649 ( .A1(n10074), .A2(SI_16_), .B1(n10093), .B2(n13091), .ZN(
        n10042) );
  XNOR2_X1 U12650 ( .A(n13406), .B(n11041), .ZN(n12678) );
  NAND2_X1 U12651 ( .A1(n10044), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n10045) );
  NAND2_X1 U12652 ( .A1(n10062), .A2(n10045), .ZN(n13327) );
  NAND2_X1 U12653 ( .A1(n13327), .A2(n12093), .ZN(n10048) );
  AOI22_X1 U12654 ( .A1(n10165), .A2(P3_REG0_REG_16__SCAN_IN), .B1(n9854), 
        .B2(P3_REG1_REG_16__SCAN_IN), .ZN(n10047) );
  NAND2_X1 U12655 ( .A1(n10301), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n10046) );
  INV_X1 U12656 ( .A(n12678), .ZN(n10050) );
  INV_X1 U12657 ( .A(n13337), .ZN(n12968) );
  NAND2_X1 U12658 ( .A1(n10050), .A2(n12968), .ZN(n10051) );
  INV_X1 U12659 ( .A(n10052), .ZN(n10053) );
  NAND2_X1 U12660 ( .A1(n10054), .A2(n10053), .ZN(n10056) );
  NAND2_X1 U12661 ( .A1(n11366), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n10070) );
  NAND2_X1 U12662 ( .A1(n11369), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n10057) );
  AND2_X1 U12663 ( .A1(n10070), .A2(n10057), .ZN(n10068) );
  XNOR2_X1 U12664 ( .A(n10069), .B(n10068), .ZN(n10683) );
  NAND2_X1 U12665 ( .A1(n10683), .A2(n12758), .ZN(n10061) );
  NAND2_X1 U12666 ( .A1(n6615), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10059) );
  XNOR2_X1 U12667 ( .A(n10059), .B(n10058), .ZN(n13104) );
  AOI22_X1 U12668 ( .A1(n10074), .A2(n10682), .B1(n13104), .B2(n10093), .ZN(
        n10060) );
  XNOR2_X1 U12669 ( .A(n13400), .B(n12496), .ZN(n10066) );
  INV_X1 U12670 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13089) );
  NAND2_X1 U12671 ( .A1(n10062), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U12672 ( .A1(n10077), .A2(n10063), .ZN(n13317) );
  NAND2_X1 U12673 ( .A1(n13317), .A2(n12093), .ZN(n10065) );
  AOI22_X1 U12674 ( .A1(n10165), .A2(P3_REG0_REG_17__SCAN_IN), .B1(n9854), 
        .B2(P3_REG1_REG_17__SCAN_IN), .ZN(n10064) );
  OAI211_X1 U12675 ( .C1(n12269), .C2(n13089), .A(n10065), .B(n10064), .ZN(
        n12681) );
  XNOR2_X1 U12676 ( .A(n10066), .B(n12681), .ZN(n12688) );
  INV_X1 U12677 ( .A(n12681), .ZN(n13326) );
  INV_X1 U12678 ( .A(n10066), .ZN(n10067) );
  NAND2_X1 U12679 ( .A1(n11528), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U12680 ( .A1(n11526), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U12681 ( .A1(n10089), .A2(n10071), .ZN(n10086) );
  XNOR2_X1 U12682 ( .A(n10088), .B(n10086), .ZN(n11051) );
  NAND2_X1 U12683 ( .A1(n11051), .A2(n12758), .ZN(n10076) );
  NAND2_X1 U12684 ( .A1(n10072), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10073) );
  XNOR2_X1 U12685 ( .A(n10073), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U12686 ( .A1(n13131), .A2(n10093), .B1(SI_18_), .B2(n10074), .ZN(
        n10075) );
  XNOR2_X1 U12687 ( .A(n13470), .B(n12496), .ZN(n10084) );
  NAND2_X1 U12688 ( .A1(n10077), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n10078) );
  NAND2_X1 U12689 ( .A1(n10098), .A2(n10078), .ZN(n13303) );
  NAND2_X1 U12690 ( .A1(n13303), .A2(n12093), .ZN(n10083) );
  INV_X1 U12691 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13309) );
  NAND2_X1 U12692 ( .A1(n12266), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n10080) );
  NAND2_X1 U12693 ( .A1(n9854), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n10079) );
  OAI211_X1 U12694 ( .C1(n13309), .C2(n12101), .A(n10080), .B(n10079), .ZN(
        n10081) );
  INV_X1 U12695 ( .A(n10081), .ZN(n10082) );
  XNOR2_X1 U12696 ( .A(n10084), .B(n12967), .ZN(n12708) );
  INV_X1 U12697 ( .A(n10084), .ZN(n10085) );
  AOI21_X2 U12698 ( .B1(n12709), .B2(n12708), .A(n7816), .ZN(n12636) );
  INV_X1 U12699 ( .A(n10086), .ZN(n10087) );
  NAND2_X1 U12700 ( .A1(n10090), .A2(n10089), .ZN(n10108) );
  INV_X1 U12701 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U12702 ( .A1(n12406), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n10109) );
  INV_X1 U12703 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11615) );
  NAND2_X1 U12704 ( .A1(n11615), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n10091) );
  AND2_X1 U12705 ( .A1(n10109), .A2(n10091), .ZN(n10107) );
  XNOR2_X1 U12706 ( .A(n10108), .B(n10107), .ZN(n12568) );
  NAND2_X1 U12707 ( .A1(n12568), .A2(n12758), .ZN(n10095) );
  NOR2_X1 U12708 ( .A1(n12761), .A2(SI_19_), .ZN(n10092) );
  AOI21_X1 U12709 ( .B1(n13146), .B2(n10093), .A(n10092), .ZN(n10094) );
  XNOR2_X1 U12710 ( .A(n13299), .B(n12496), .ZN(n10105) );
  INV_X1 U12711 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U12712 ( .A1(n10098), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n10099) );
  NAND2_X1 U12713 ( .A1(n10113), .A2(n10099), .ZN(n13297) );
  NAND2_X1 U12714 ( .A1(n13297), .A2(n12093), .ZN(n10104) );
  INV_X1 U12715 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U12716 ( .A1(n10165), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n10101) );
  NAND2_X1 U12717 ( .A1(n9854), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n10100) );
  OAI211_X1 U12718 ( .C1(n13129), .C2(n12101), .A(n10101), .B(n10100), .ZN(
        n10102) );
  INV_X1 U12719 ( .A(n10102), .ZN(n10103) );
  XNOR2_X1 U12720 ( .A(n10105), .B(n12710), .ZN(n12635) );
  INV_X1 U12721 ( .A(n10105), .ZN(n10106) );
  NAND2_X1 U12722 ( .A1(n10108), .A2(n10107), .ZN(n10110) );
  XNOR2_X1 U12723 ( .A(n10139), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n10122) );
  XNOR2_X1 U12724 ( .A(n10122), .B(n11710), .ZN(n11537) );
  NAND2_X1 U12725 ( .A1(n11537), .A2(n12758), .ZN(n10112) );
  OR2_X1 U12726 ( .A1(n12761), .A2(n11539), .ZN(n10111) );
  XNOR2_X1 U12727 ( .A(n13391), .B(n12496), .ZN(n10120) );
  NAND2_X1 U12728 ( .A1(n10113), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n10114) );
  NAND2_X1 U12729 ( .A1(n10129), .A2(n10114), .ZN(n13273) );
  NAND2_X1 U12730 ( .A1(n13273), .A2(n12093), .ZN(n10119) );
  INV_X1 U12731 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U12732 ( .A1(n12266), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n10116) );
  NAND2_X1 U12733 ( .A1(n9854), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n10115) );
  OAI211_X1 U12734 ( .C1(n13274), .C2(n12101), .A(n10116), .B(n10115), .ZN(
        n10117) );
  INV_X1 U12735 ( .A(n10117), .ZN(n10118) );
  XNOR2_X1 U12736 ( .A(n10120), .B(n13294), .ZN(n12694) );
  INV_X1 U12737 ( .A(n10120), .ZN(n10121) );
  NAND2_X1 U12738 ( .A1(n10139), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U12739 ( .A1(n10124), .A2(n10123), .ZN(n10126) );
  NAND2_X1 U12740 ( .A1(n11771), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n10140) );
  NAND2_X1 U12741 ( .A1(n12566), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n10141) );
  NAND2_X1 U12742 ( .A1(n10140), .A2(n10141), .ZN(n10125) );
  INV_X1 U12743 ( .A(SI_21_), .ZN(n11651) );
  OR2_X1 U12744 ( .A1(n12761), .A2(n11651), .ZN(n10127) );
  XNOR2_X1 U12745 ( .A(n13457), .B(n12487), .ZN(n10134) );
  NAND2_X1 U12746 ( .A1(n10129), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n10130) );
  NAND2_X1 U12747 ( .A1(n10147), .A2(n10130), .ZN(n13258) );
  INV_X1 U12748 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13267) );
  NAND2_X1 U12749 ( .A1(n12266), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U12750 ( .A1(n9854), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n10131) );
  OAI211_X1 U12751 ( .C1(n13267), .C2(n12101), .A(n10132), .B(n10131), .ZN(
        n10133) );
  AOI21_X1 U12752 ( .B1(n10134), .B2(n13252), .A(n10135), .ZN(n12644) );
  NAND2_X1 U12753 ( .A1(n12643), .A2(n12644), .ZN(n12642) );
  INV_X1 U12754 ( .A(n10135), .ZN(n10136) );
  NAND3_X1 U12755 ( .A1(n10140), .A2(P1_DATAO_REG_20__SCAN_IN), .A3(n11710), 
        .ZN(n10142) );
  AND2_X1 U12756 ( .A1(n10142), .A2(n10141), .ZN(n10143) );
  INV_X1 U12757 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10158) );
  XNOR2_X1 U12758 ( .A(n10158), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n10157) );
  XNOR2_X1 U12759 ( .A(n10156), .B(n10157), .ZN(n11456) );
  NAND2_X1 U12760 ( .A1(n11456), .A2(n12758), .ZN(n10146) );
  OR2_X1 U12761 ( .A1(n12761), .A2(n10144), .ZN(n10145) );
  XNOR2_X1 U12762 ( .A(n13451), .B(n11041), .ZN(n10192) );
  NAND2_X1 U12763 ( .A1(n10191), .A2(n10192), .ZN(n10154) );
  OAI21_X1 U12764 ( .B1(n10191), .B2(n10192), .A(n10154), .ZN(n12702) );
  NAND2_X1 U12765 ( .A1(n10147), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n10148) );
  NAND2_X1 U12766 ( .A1(n10163), .A2(n10148), .ZN(n13248) );
  NAND2_X1 U12767 ( .A1(n13248), .A2(n12093), .ZN(n10153) );
  INV_X1 U12768 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13254) );
  NAND2_X1 U12769 ( .A1(n12266), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n10150) );
  NAND2_X1 U12770 ( .A1(n9854), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n10149) );
  OAI211_X1 U12771 ( .C1(n13254), .C2(n12101), .A(n10150), .B(n10149), .ZN(
        n10151) );
  INV_X1 U12772 ( .A(n10151), .ZN(n10152) );
  INV_X1 U12773 ( .A(n10154), .ZN(n10155) );
  NAND2_X1 U12774 ( .A1(n10158), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n10159) );
  XNOR2_X1 U12775 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n10173) );
  XNOR2_X1 U12776 ( .A(n10174), .B(n10173), .ZN(n11616) );
  NAND2_X1 U12777 ( .A1(n11616), .A2(n12758), .ZN(n10161) );
  OR2_X1 U12778 ( .A1(n12761), .A2(n11618), .ZN(n10160) );
  XNOR2_X1 U12779 ( .A(n12918), .B(n12496), .ZN(n10193) );
  INV_X1 U12780 ( .A(n10193), .ZN(n10162) );
  NAND2_X1 U12781 ( .A1(n10163), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U12782 ( .A1(n10182), .A2(n10164), .ZN(n12630) );
  NAND2_X1 U12783 ( .A1(n12630), .A2(n12093), .ZN(n10171) );
  INV_X1 U12784 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n10168) );
  NAND2_X1 U12785 ( .A1(n10165), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n10167) );
  NAND2_X1 U12786 ( .A1(n9854), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n10166) );
  OAI211_X1 U12787 ( .C1(n10168), .C2(n12101), .A(n10167), .B(n10166), .ZN(
        n10169) );
  INV_X1 U12788 ( .A(n10169), .ZN(n10170) );
  NAND2_X1 U12789 ( .A1(n12628), .A2(n13227), .ZN(n12627) );
  INV_X1 U12790 ( .A(n10172), .ZN(n10190) );
  NAND2_X1 U12791 ( .A1(n10174), .A2(n10173), .ZN(n10177) );
  NAND2_X1 U12792 ( .A1(n10175), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n10176) );
  INV_X1 U12793 ( .A(n10179), .ZN(n10178) );
  XNOR2_X1 U12794 ( .A(n10266), .B(n12209), .ZN(n12088) );
  NAND2_X1 U12795 ( .A1(n12088), .A2(n12758), .ZN(n10181) );
  OR2_X1 U12796 ( .A1(n12761), .A2(n12089), .ZN(n10180) );
  XNOR2_X1 U12797 ( .A(n13223), .B(n12496), .ZN(n10189) );
  INV_X1 U12798 ( .A(n10232), .ZN(n10233) );
  NAND2_X1 U12799 ( .A1(n10182), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n10183) );
  NAND2_X1 U12800 ( .A1(n10233), .A2(n10183), .ZN(n13222) );
  NAND2_X1 U12801 ( .A1(n13222), .A2(n12093), .ZN(n10188) );
  INV_X1 U12802 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13230) );
  NAND2_X1 U12803 ( .A1(n12266), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n10185) );
  NAND2_X1 U12804 ( .A1(n9854), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n10184) );
  OAI211_X1 U12805 ( .C1(n13230), .C2(n12101), .A(n10185), .B(n10184), .ZN(
        n10186) );
  INV_X1 U12806 ( .A(n10186), .ZN(n10187) );
  NAND2_X1 U12807 ( .A1(n10189), .A2(n13238), .ZN(n12479) );
  OAI21_X1 U12808 ( .B1(n10189), .B2(n13238), .A(n12479), .ZN(n10195) );
  NAND2_X1 U12809 ( .A1(n12627), .A2(n7823), .ZN(n10199) );
  AOI22_X1 U12810 ( .A1(n10193), .A2(n13227), .B1(n13264), .B2(n10192), .ZN(
        n10197) );
  NOR2_X1 U12811 ( .A1(n10193), .A2(n13227), .ZN(n10194) );
  INV_X1 U12812 ( .A(n12671), .ZN(n10198) );
  NAND2_X1 U12813 ( .A1(n10199), .A2(n10198), .ZN(n10228) );
  NAND2_X1 U12814 ( .A1(n13146), .A2(n6928), .ZN(n10203) );
  NAND2_X1 U12815 ( .A1(n10222), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10201) );
  AND2_X1 U12816 ( .A1(n6928), .A2(n11540), .ZN(n10373) );
  XNOR2_X1 U12817 ( .A(n12801), .B(n10373), .ZN(n10202) );
  NAND2_X1 U12818 ( .A1(n10203), .A2(n10202), .ZN(n10363) );
  AND2_X1 U12819 ( .A1(n10363), .A2(n15638), .ZN(n10256) );
  INV_X1 U12820 ( .A(n10369), .ZN(n13499) );
  INV_X1 U12821 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10205) );
  NAND2_X1 U12822 ( .A1(n10545), .A2(n10205), .ZN(n10207) );
  NAND2_X1 U12823 ( .A1(n12293), .A2(n13523), .ZN(n10206) );
  NOR2_X1 U12824 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .ZN(
        n10211) );
  NOR4_X1 U12825 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n10210) );
  NOR4_X1 U12826 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n10209) );
  NOR4_X1 U12827 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n10208) );
  NAND4_X1 U12828 ( .A1(n10211), .A2(n10210), .A3(n10209), .A4(n10208), .ZN(
        n10217) );
  NOR4_X1 U12829 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n10215) );
  NOR4_X1 U12830 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n10214) );
  NOR4_X1 U12831 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n10213) );
  NOR4_X1 U12832 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n10212) );
  NAND4_X1 U12833 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n10216) );
  OAI21_X1 U12834 ( .B1(n10217), .B2(n10216), .A(n10545), .ZN(n10370) );
  NAND2_X1 U12835 ( .A1(n10256), .A2(n10365), .ZN(n10221) );
  NAND3_X1 U12836 ( .A1(n12957), .A2(n6928), .A3(n12952), .ZN(n10218) );
  NAND2_X1 U12837 ( .A1(n10369), .A2(n10370), .ZN(n10219) );
  NOR2_X1 U12838 ( .A1(n10219), .A2(n13497), .ZN(n10362) );
  NAND2_X1 U12839 ( .A1(n6602), .A2(n10362), .ZN(n10220) );
  NAND2_X1 U12840 ( .A1(n10221), .A2(n10220), .ZN(n10227) );
  OAI21_X1 U12841 ( .B1(n10222), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n10224) );
  XNOR2_X1 U12842 ( .A(n10224), .B(n10223), .ZN(n10910) );
  INV_X1 U12843 ( .A(n12293), .ZN(n10226) );
  NOR2_X1 U12844 ( .A1(n12091), .A2(n13523), .ZN(n10225) );
  NAND2_X1 U12845 ( .A1(n10226), .A2(n10225), .ZN(n10394) );
  NAND2_X1 U12846 ( .A1(n10227), .A2(n10909), .ZN(n12749) );
  NAND2_X1 U12847 ( .A1(n10228), .A2(n12730), .ZN(n10255) );
  INV_X1 U12848 ( .A(n13223), .ZN(n13438) );
  NAND2_X1 U12849 ( .A1(n10909), .A2(n15623), .ZN(n10229) );
  OR2_X1 U12850 ( .A1(n13146), .A2(n12952), .ZN(n15603) );
  INV_X1 U12851 ( .A(n10365), .ZN(n10242) );
  OR2_X1 U12852 ( .A1(n10229), .A2(n10242), .ZN(n10230) );
  INV_X1 U12853 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n10231) );
  INV_X1 U12854 ( .A(n10280), .ZN(n10281) );
  NAND2_X1 U12855 ( .A1(n10233), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n10234) );
  NAND2_X1 U12856 ( .A1(n10281), .A2(n10234), .ZN(n13213) );
  NAND2_X1 U12857 ( .A1(n13213), .A2(n12093), .ZN(n10240) );
  INV_X1 U12858 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U12859 ( .A1(n12266), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n10236) );
  NAND2_X1 U12860 ( .A1(n9854), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n10235) );
  OAI211_X1 U12861 ( .C1(n10237), .C2(n12101), .A(n10236), .B(n10235), .ZN(
        n10238) );
  INV_X1 U12862 ( .A(n10238), .ZN(n10239) );
  NOR2_X1 U12863 ( .A1(n12800), .A2(n12946), .ZN(n11158) );
  NAND2_X1 U12864 ( .A1(n11158), .A2(n10909), .ZN(n12953) );
  INV_X1 U12865 ( .A(n13513), .ZN(n12954) );
  NAND2_X1 U12866 ( .A1(n12954), .A2(n13134), .ZN(n10951) );
  NAND2_X1 U12867 ( .A1(n6924), .A2(n10951), .ZN(n10356) );
  INV_X1 U12868 ( .A(n10356), .ZN(n10241) );
  INV_X1 U12869 ( .A(n10362), .ZN(n10243) );
  OR2_X1 U12870 ( .A1(n12953), .A2(n10362), .ZN(n10249) );
  NAND2_X1 U12871 ( .A1(n10242), .A2(n10363), .ZN(n10246) );
  NAND2_X1 U12872 ( .A1(n10243), .A2(n6602), .ZN(n10245) );
  AND2_X1 U12873 ( .A1(n10910), .A2(n10394), .ZN(n10244) );
  NAND2_X1 U12874 ( .A1(n12800), .A2(n12930), .ZN(n10368) );
  NAND4_X1 U12875 ( .A1(n10246), .A2(n10245), .A3(n10244), .A4(n10368), .ZN(
        n10247) );
  NAND2_X1 U12876 ( .A1(n10247), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10248) );
  AOI22_X1 U12877 ( .A1(n13222), .A2(n12747), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10250) );
  OAI21_X1 U12878 ( .B1(n13227), .B2(n12733), .A(n10250), .ZN(n10251) );
  AOI21_X1 U12879 ( .B1(n12963), .B2(n12735), .A(n10251), .ZN(n10252) );
  OAI21_X1 U12880 ( .B1(n13438), .B2(n12744), .A(n10252), .ZN(n10253) );
  INV_X1 U12881 ( .A(n10253), .ZN(n10254) );
  INV_X1 U12882 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n10830) );
  MUX2_X1 U12883 ( .A(n10256), .B(n12957), .S(n12952), .Z(n10257) );
  NAND2_X1 U12884 ( .A1(n10257), .A2(n13146), .ZN(n15588) );
  OR2_X1 U12885 ( .A1(n15603), .A2(n12957), .ZN(n15627) );
  NAND2_X1 U12886 ( .A1(n15588), .A2(n15627), .ZN(n13372) );
  NAND2_X1 U12887 ( .A1(n10258), .A2(n12806), .ZN(n15572) );
  NAND2_X1 U12888 ( .A1(n11494), .A2(n15573), .ZN(n12811) );
  NAND2_X1 U12889 ( .A1(n10260), .A2(n12811), .ZN(n11493) );
  NAND2_X1 U12890 ( .A1(n15581), .A2(n11498), .ZN(n12820) );
  INV_X1 U12891 ( .A(n11498), .ZN(n10261) );
  NAND2_X1 U12892 ( .A1(n12979), .A2(n10261), .ZN(n12818) );
  AND2_X2 U12893 ( .A1(n12820), .A2(n12818), .ZN(n12767) );
  NAND2_X1 U12894 ( .A1(n11784), .A2(n15624), .ZN(n12821) );
  INV_X1 U12895 ( .A(n15624), .ZN(n11732) );
  NAND2_X1 U12896 ( .A1(n12978), .A2(n11732), .ZN(n12822) );
  AND2_X2 U12897 ( .A1(n12821), .A2(n12822), .ZN(n12819) );
  NAND2_X1 U12898 ( .A1(n10316), .A2(n11774), .ZN(n12827) );
  INV_X1 U12899 ( .A(n11774), .ZN(n11563) );
  NAND2_X1 U12900 ( .A1(n11563), .A2(n12977), .ZN(n12826) );
  NAND2_X1 U12901 ( .A1(n11785), .A2(n12721), .ZN(n12832) );
  INV_X1 U12902 ( .A(n12721), .ZN(n15639) );
  NAND2_X1 U12903 ( .A1(n12976), .A2(n15639), .ZN(n12833) );
  NAND2_X1 U12904 ( .A1(n11505), .A2(n12771), .ZN(n11504) );
  INV_X1 U12905 ( .A(n11767), .ZN(n12838) );
  NOR2_X1 U12906 ( .A1(n12069), .A2(n12975), .ZN(n12849) );
  XNOR2_X1 U12907 ( .A(n12852), .B(n12369), .ZN(n12851) );
  AND2_X1 U12908 ( .A1(n12852), .A2(n12974), .ZN(n12853) );
  NAND2_X1 U12909 ( .A1(n12252), .A2(n12973), .ZN(n12863) );
  NAND2_X1 U12910 ( .A1(n12241), .A2(n12858), .ZN(n12240) );
  NAND2_X1 U12911 ( .A1(n12665), .A2(n12383), .ZN(n12866) );
  INV_X1 U12912 ( .A(n12866), .ZN(n10262) );
  NOR2_X1 U12913 ( .A1(n13492), .A2(n13354), .ZN(n12870) );
  NAND2_X1 U12914 ( .A1(n13492), .A2(n13354), .ZN(n12377) );
  NAND2_X1 U12915 ( .A1(n13487), .A2(n12970), .ZN(n10330) );
  OR2_X1 U12916 ( .A1(n13487), .A2(n12970), .ZN(n10263) );
  INV_X1 U12917 ( .A(n12970), .ZN(n13336) );
  AND2_X1 U12918 ( .A1(n13487), .A2(n13336), .ZN(n12874) );
  OR2_X1 U12919 ( .A1(n13410), .A2(n13355), .ZN(n12878) );
  NAND2_X1 U12920 ( .A1(n13410), .A2(n13355), .ZN(n12881) );
  NAND2_X1 U12921 ( .A1(n12878), .A2(n12881), .ZN(n13334) );
  INV_X1 U12922 ( .A(n12881), .ZN(n10264) );
  OR2_X1 U12923 ( .A1(n13406), .A2(n13337), .ZN(n12879) );
  NAND2_X1 U12924 ( .A1(n13406), .A2(n13337), .ZN(n12882) );
  NAND2_X1 U12925 ( .A1(n12879), .A2(n12882), .ZN(n13324) );
  OR2_X1 U12926 ( .A1(n13400), .A2(n12681), .ZN(n10265) );
  NAND2_X1 U12927 ( .A1(n13400), .A2(n12681), .ZN(n12893) );
  INV_X1 U12928 ( .A(n10265), .ZN(n12889) );
  NAND2_X1 U12929 ( .A1(n13470), .A2(n13316), .ZN(n12894) );
  NAND2_X1 U12930 ( .A1(n13299), .A2(n12710), .ZN(n12901) );
  INV_X1 U12931 ( .A(n13299), .ZN(n13395) );
  INV_X1 U12932 ( .A(n13294), .ZN(n13265) );
  NAND2_X1 U12933 ( .A1(n13457), .A2(n13283), .ZN(n12909) );
  NOR2_X1 U12934 ( .A1(n13457), .A2(n13283), .ZN(n12911) );
  XNOR2_X1 U12935 ( .A(n12323), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n10268) );
  XNOR2_X1 U12936 ( .A(n10274), .B(n10268), .ZN(n12290) );
  NAND2_X1 U12937 ( .A1(n12290), .A2(n12758), .ZN(n10270) );
  OR2_X1 U12938 ( .A1(n12761), .A2(n12292), .ZN(n10269) );
  OR2_X1 U12939 ( .A1(n13223), .A2(n13238), .ZN(n12921) );
  NAND2_X1 U12940 ( .A1(n12921), .A2(n13218), .ZN(n10271) );
  NAND2_X1 U12941 ( .A1(n13223), .A2(n13238), .ZN(n12920) );
  AND2_X1 U12942 ( .A1(n10271), .A2(n12920), .ZN(n10272) );
  NAND2_X1 U12943 ( .A1(n12918), .A2(n13227), .ZN(n10344) );
  AND2_X1 U12944 ( .A1(n12920), .A2(n10344), .ZN(n13195) );
  NAND2_X1 U12945 ( .A1(n12323), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U12946 ( .A1(n12320), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n10275) );
  XNOR2_X1 U12947 ( .A(n14185), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n10276) );
  XNOR2_X1 U12948 ( .A(n10292), .B(n10276), .ZN(n13518) );
  NAND2_X1 U12949 ( .A1(n13518), .A2(n12758), .ZN(n10278) );
  OR2_X1 U12950 ( .A1(n12761), .A2(n13521), .ZN(n10277) );
  INV_X1 U12951 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n10279) );
  INV_X1 U12952 ( .A(n10298), .ZN(n10299) );
  NAND2_X1 U12953 ( .A1(n10281), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U12954 ( .A1(n10299), .A2(n10282), .ZN(n13201) );
  NAND2_X1 U12955 ( .A1(n13201), .A2(n12093), .ZN(n10288) );
  INV_X1 U12956 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U12957 ( .A1(n12266), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n10284) );
  NAND2_X1 U12958 ( .A1(n9854), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n10283) );
  OAI211_X1 U12959 ( .C1(n10285), .C2(n12101), .A(n10284), .B(n10283), .ZN(
        n10286) );
  INV_X1 U12960 ( .A(n10286), .ZN(n10287) );
  NAND2_X1 U12961 ( .A1(n12483), .A2(n13212), .ZN(n12932) );
  AND2_X1 U12962 ( .A1(n12932), .A2(n13196), .ZN(n10289) );
  NAND2_X1 U12963 ( .A1(n10290), .A2(n10289), .ZN(n10309) );
  INV_X1 U12964 ( .A(n10309), .ZN(n10310) );
  OAI21_X1 U12965 ( .B1(n10311), .B2(n13194), .A(n10310), .ZN(n10307) );
  AND2_X1 U12966 ( .A1(n15186), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U12967 ( .A1(n14185), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n10293) );
  XNOR2_X1 U12968 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n10294) );
  XNOR2_X1 U12969 ( .A(n12491), .B(n10294), .ZN(n13514) );
  NAND2_X1 U12970 ( .A1(n13514), .A2(n12758), .ZN(n10296) );
  OR2_X1 U12971 ( .A1(n12761), .A2(n13515), .ZN(n10295) );
  INV_X1 U12972 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n10297) );
  NAND2_X1 U12973 ( .A1(n10299), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U12974 ( .A1(n10351), .A2(n10300), .ZN(n13185) );
  NAND2_X1 U12975 ( .A1(n13185), .A2(n12093), .ZN(n10306) );
  NAND2_X1 U12976 ( .A1(n9854), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U12977 ( .A1(n10301), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n10302) );
  OAI211_X1 U12978 ( .C1(n9822), .C2(n10830), .A(n10303), .B(n10302), .ZN(
        n10304) );
  INV_X1 U12979 ( .A(n10304), .ZN(n10305) );
  AOI21_X1 U12980 ( .B1(n10307), .B2(n12931), .A(n12934), .ZN(n10312) );
  INV_X1 U12981 ( .A(n13194), .ZN(n10308) );
  OR2_X1 U12982 ( .A1(n10312), .A2(n12544), .ZN(n13189) );
  NAND2_X1 U12983 ( .A1(n11040), .A2(n15594), .ZN(n10314) );
  NAND2_X1 U12984 ( .A1(n15583), .A2(n15593), .ZN(n10313) );
  NAND2_X1 U12985 ( .A1(n10314), .A2(n10313), .ZN(n15579) );
  INV_X1 U12986 ( .A(n15573), .ZN(n12815) );
  NAND2_X1 U12987 ( .A1(n11494), .A2(n12815), .ZN(n10315) );
  AND2_X1 U12988 ( .A1(n10316), .A2(n11563), .ZN(n10318) );
  OR2_X1 U12989 ( .A1(n12819), .A2(n10318), .ZN(n10319) );
  NAND2_X1 U12990 ( .A1(n12978), .A2(n15624), .ZN(n11777) );
  INV_X1 U12991 ( .A(n12771), .ZN(n11507) );
  NAND2_X1 U12992 ( .A1(n12976), .A2(n12721), .ZN(n10320) );
  NAND2_X1 U12993 ( .A1(n12842), .A2(n11855), .ZN(n10321) );
  NAND2_X1 U12994 ( .A1(n12837), .A2(n11767), .ZN(n11794) );
  AND2_X1 U12995 ( .A1(n10321), .A2(n11794), .ZN(n10322) );
  XNOR2_X1 U12996 ( .A(n12069), .B(n12975), .ZN(n12846) );
  INV_X1 U12997 ( .A(n12842), .ZN(n12201) );
  NAND2_X1 U12998 ( .A1(n12201), .A2(n12843), .ZN(n11796) );
  AND2_X1 U12999 ( .A1(n12846), .A2(n11796), .ZN(n10323) );
  OR2_X1 U13000 ( .A1(n12069), .A2(n11910), .ZN(n12151) );
  OR2_X1 U13001 ( .A1(n12852), .A2(n12369), .ZN(n12235) );
  INV_X1 U13002 ( .A(n12973), .ZN(n12659) );
  AOI22_X1 U13003 ( .A1(n12252), .A2(n12659), .B1(n12369), .B2(n12852), .ZN(
        n10324) );
  OR2_X1 U13004 ( .A1(n12252), .A2(n12659), .ZN(n10326) );
  NAND2_X1 U13005 ( .A1(n12665), .A2(n12972), .ZN(n10327) );
  NAND2_X1 U13006 ( .A1(n10328), .A2(n10327), .ZN(n12381) );
  OR2_X1 U13007 ( .A1(n13492), .A2(n12971), .ZN(n13348) );
  NAND2_X1 U13008 ( .A1(n13410), .A2(n12969), .ZN(n10331) );
  NAND2_X1 U13009 ( .A1(n13406), .A2(n12968), .ZN(n10332) );
  NAND2_X1 U13010 ( .A1(n10333), .A2(n10332), .ZN(n13313) );
  NAND2_X1 U13011 ( .A1(n13313), .A2(n13314), .ZN(n10335) );
  OR2_X1 U13012 ( .A1(n13400), .A2(n13326), .ZN(n10334) );
  NAND2_X1 U13013 ( .A1(n10335), .A2(n10334), .ZN(n13277) );
  OR2_X1 U13014 ( .A1(n13299), .A2(n13307), .ZN(n13279) );
  INV_X1 U13015 ( .A(n13305), .ZN(n10336) );
  NAND2_X1 U13016 ( .A1(n13279), .A2(n10336), .ZN(n10338) );
  INV_X1 U13017 ( .A(n13271), .ZN(n13280) );
  INV_X1 U13018 ( .A(n12888), .ZN(n12900) );
  NAND2_X1 U13019 ( .A1(n12900), .A2(n12901), .ZN(n13292) );
  OR2_X1 U13020 ( .A1(n13470), .A2(n12967), .ZN(n13289) );
  NAND2_X1 U13021 ( .A1(n13292), .A2(n13289), .ZN(n13278) );
  NAND2_X1 U13022 ( .A1(n13278), .A2(n13279), .ZN(n10337) );
  NAND2_X1 U13023 ( .A1(n13391), .A2(n13294), .ZN(n10339) );
  OR2_X1 U13024 ( .A1(n13457), .A2(n13252), .ZN(n10341) );
  NAND2_X1 U13025 ( .A1(n13451), .A2(n12966), .ZN(n10343) );
  NOR2_X1 U13026 ( .A1(n13451), .A2(n12966), .ZN(n10342) );
  INV_X1 U13027 ( .A(n13238), .ZN(n12964) );
  INV_X1 U13028 ( .A(n13376), .ZN(n13215) );
  NOR2_X1 U13029 ( .A1(n13433), .A2(n13212), .ZN(n10345) );
  INV_X1 U13030 ( .A(n13146), .ZN(n12799) );
  NAND2_X1 U13031 ( .A1(n12799), .A2(n12957), .ZN(n10348) );
  NAND2_X1 U13032 ( .A1(n12797), .A2(n12952), .ZN(n10347) );
  NAND2_X1 U13033 ( .A1(n10350), .A2(n10349), .ZN(n10360) );
  NAND2_X1 U13034 ( .A1(n10351), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U13035 ( .A1(n12092), .A2(n10352), .ZN(n13181) );
  INV_X1 U13036 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n13180) );
  NAND2_X1 U13037 ( .A1(n12266), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U13038 ( .A1(n9854), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n10353) );
  OAI211_X1 U13039 ( .C1(n13180), .C2(n12101), .A(n10354), .B(n10353), .ZN(
        n10355) );
  AOI21_X1 U13040 ( .B1(n13372), .B2(n13189), .A(n13184), .ZN(n10378) );
  NAND2_X1 U13041 ( .A1(n6602), .A2(n10909), .ZN(n10361) );
  NAND2_X1 U13042 ( .A1(n12953), .A2(n10361), .ZN(n10366) );
  AND3_X1 U13043 ( .A1(n10363), .A2(n10909), .A3(n10362), .ZN(n10364) );
  INV_X1 U13044 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n10379) );
  NAND3_X1 U13045 ( .A1(n13146), .A2(n12952), .A3(n12957), .ZN(n10367) );
  NAND2_X1 U13046 ( .A1(n10367), .A2(n12946), .ZN(n10372) );
  NAND2_X1 U13047 ( .A1(n10368), .A2(n10372), .ZN(n11414) );
  NAND2_X1 U13048 ( .A1(n11414), .A2(n13497), .ZN(n10377) );
  XNOR2_X1 U13049 ( .A(n13497), .B(n10369), .ZN(n10371) );
  INV_X1 U13050 ( .A(n10372), .ZN(n11418) );
  NAND3_X1 U13051 ( .A1(n12800), .A2(n10373), .A3(n12801), .ZN(n10374) );
  NAND2_X1 U13052 ( .A1(n11418), .A2(n10374), .ZN(n10375) );
  INV_X1 U13053 ( .A(n13497), .ZN(n11417) );
  NAND2_X1 U13054 ( .A1(n10375), .A2(n11417), .ZN(n10376) );
  NAND2_X1 U13055 ( .A1(n10382), .A2(n14370), .ZN(n10390) );
  INV_X1 U13056 ( .A(n15082), .ZN(n12439) );
  INV_X1 U13057 ( .A(n14637), .ZN(n10383) );
  OAI22_X1 U13058 ( .A1(n10383), .A2(n15052), .B1(n14522), .B2(n14976), .ZN(
        n12433) );
  INV_X1 U13059 ( .A(n12437), .ZN(n10385) );
  OAI22_X1 U13060 ( .A1(n10385), .A2(n14291), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10384), .ZN(n10386) );
  AOI21_X1 U13061 ( .B1(n12433), .B2(n14368), .A(n10386), .ZN(n10387) );
  NAND2_X1 U13062 ( .A1(n10390), .A2(n10389), .ZN(P1_U3214) );
  NAND2_X1 U13063 ( .A1(n10490), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10391) );
  NOR2_X1 U13064 ( .A1(n10496), .A2(n10391), .ZN(P2_U3947) );
  INV_X1 U13065 ( .A(n10464), .ZN(n10392) );
  OR2_X2 U13066 ( .A1(n10393), .A2(n10392), .ZN(n14653) );
  INV_X1 U13067 ( .A(n10394), .ZN(n10395) );
  NAND2_X1 U13068 ( .A1(n13498), .A2(n10395), .ZN(n12965) );
  INV_X2 U13069 ( .A(n12965), .ZN(P3_U3897) );
  XNOR2_X1 U13070 ( .A(n10397), .B(n10396), .ZN(n10401) );
  NAND2_X1 U13071 ( .A1(n11153), .A2(n10398), .ZN(n10400) );
  OR2_X1 U13072 ( .A1(n10400), .A2(n10401), .ZN(n11518) );
  INV_X1 U13073 ( .A(n11518), .ZN(n10399) );
  AOI211_X1 U13074 ( .C1(n10401), .C2(n10400), .A(n14359), .B(n10399), .ZN(
        n10404) );
  MUX2_X1 U13075 ( .A(n14242), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n10403) );
  AOI22_X1 U13076 ( .A1(n15223), .A2(n11381), .B1(n14651), .B2(n15222), .ZN(
        n11384) );
  INV_X1 U13077 ( .A(n14368), .ZN(n14244) );
  OAI22_X1 U13078 ( .A1(n14380), .A2(n14399), .B1(n11384), .B2(n14244), .ZN(
        n10402) );
  OR3_X1 U13079 ( .A1(n10404), .A2(n10403), .A3(n10402), .ZN(P1_U3218) );
  NOR2_X1 U13080 ( .A1(n10436), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13500) );
  INV_X1 U13081 ( .A(n13500), .ZN(n13520) );
  NAND2_X2 U13082 ( .A1(n10436), .A2(P3_U3151), .ZN(n13522) );
  OAI222_X1 U13083 ( .A1(n13520), .A2(n10405), .B1(n13522), .B2(n6778), .C1(
        n11130), .C2(P3_U3151), .ZN(P3_U3289) );
  INV_X1 U13084 ( .A(SI_7_), .ZN(n10406) );
  INV_X1 U13085 ( .A(n11063), .ZN(n11056) );
  OAI222_X1 U13086 ( .A1(n13520), .A2(n10407), .B1(n13522), .B2(n10406), .C1(
        n11056), .C2(P3_U3151), .ZN(P3_U3288) );
  NOR2_X1 U13087 ( .A1(n10436), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14169) );
  INV_X2 U13088 ( .A(n14169), .ZN(n14184) );
  AND2_X1 U13089 ( .A1(n10436), .A2(P2_U3088), .ZN(n14175) );
  OAI222_X1 U13090 ( .A1(n14184), .A2(n10738), .B1(n6438), .B2(n10442), .C1(
        P2_U3088), .C2(n6667), .ZN(P2_U3324) );
  INV_X1 U13091 ( .A(n10408), .ZN(n10446) );
  OAI222_X1 U13092 ( .A1(n14184), .A2(n10409), .B1(n6438), .B2(n10446), .C1(
        P2_U3088), .C2(n10507), .ZN(P2_U3323) );
  INV_X1 U13093 ( .A(n10410), .ZN(n10440) );
  INV_X1 U13094 ( .A(n15466), .ZN(n10411) );
  OAI222_X1 U13095 ( .A1(n14184), .A2(n10412), .B1(n6438), .B2(n10440), .C1(
        P2_U3088), .C2(n10411), .ZN(P2_U3322) );
  OAI222_X1 U13096 ( .A1(n10978), .A2(P3_U3151), .B1(n13520), .B2(n10414), 
        .C1(n10413), .C2(n13522), .ZN(P3_U3294) );
  OAI222_X1 U13097 ( .A1(n15427), .A2(P2_U3088), .B1(n6438), .B2(n10453), .C1(
        n10415), .C2(n14184), .ZN(P2_U3326) );
  OAI222_X1 U13098 ( .A1(n10598), .A2(P2_U3088), .B1(n6438), .B2(n10468), .C1(
        n10416), .C2(n14184), .ZN(P2_U3325) );
  INV_X1 U13099 ( .A(n10417), .ZN(n10438) );
  INV_X1 U13100 ( .A(n10538), .ZN(n15479) );
  OAI222_X1 U13101 ( .A1(n14184), .A2(n10418), .B1(n6438), .B2(n10438), .C1(
        P2_U3088), .C2(n15479), .ZN(P2_U3321) );
  INV_X1 U13102 ( .A(n11225), .ZN(n11068) );
  INV_X1 U13103 ( .A(n10419), .ZN(n10421) );
  INV_X1 U13104 ( .A(SI_8_), .ZN(n10420) );
  OAI222_X1 U13105 ( .A1(n11068), .A2(P3_U3151), .B1(n13520), .B2(n10421), 
        .C1(n10420), .C2(n13522), .ZN(P3_U3287) );
  OAI222_X1 U13106 ( .A1(n11229), .A2(P3_U3151), .B1(n13520), .B2(n10423), 
        .C1(n10422), .C2(n13522), .ZN(P3_U3286) );
  INV_X1 U13107 ( .A(n13522), .ZN(n10731) );
  AOI222_X1 U13108 ( .A1(n10424), .A2(n13500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10924), .C1(SI_3_), .C2(n10731), .ZN(n10425) );
  INV_X1 U13109 ( .A(n10425), .ZN(P3_U3292) );
  AOI222_X1 U13110 ( .A1(n10426), .A2(n13500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10934), .C1(SI_5_), .C2(n10731), .ZN(n10427) );
  INV_X1 U13111 ( .A(n10427), .ZN(P3_U3290) );
  AOI222_X1 U13112 ( .A1(n10428), .A2(n13500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n7009), .C1(SI_2_), .C2(n10731), .ZN(n10429) );
  INV_X1 U13113 ( .A(n10429), .ZN(P3_U3293) );
  AOI222_X1 U13114 ( .A1(n10430), .A2(n13500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10979), .C1(SI_4_), .C2(n10731), .ZN(n10431) );
  INV_X1 U13115 ( .A(n10431), .ZN(P3_U3291) );
  INV_X1 U13116 ( .A(n10432), .ZN(n10444) );
  INV_X1 U13117 ( .A(n10664), .ZN(n10433) );
  OAI222_X1 U13118 ( .A1(n14184), .A2(n10480), .B1(n6438), .B2(n10444), .C1(
        P2_U3088), .C2(n10433), .ZN(P2_U3320) );
  OAI222_X1 U13119 ( .A1(n11808), .A2(P3_U3151), .B1(n13520), .B2(n10435), 
        .C1(n10434), .C2(n13522), .ZN(P3_U3285) );
  NAND2_X1 U13120 ( .A1(n10436), .A2(P1_U3086), .ZN(n15185) );
  CLKBUF_X1 U13121 ( .A(n15185), .Z(n15174) );
  NOR2_X1 U13122 ( .A1(n10436), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15178) );
  INV_X2 U13123 ( .A(n15178), .ZN(n15188) );
  INV_X1 U13124 ( .A(n14724), .ZN(n10437) );
  OAI222_X1 U13125 ( .A1(n15174), .A2(n10439), .B1(n15188), .B2(n10438), .C1(
        n6428), .C2(n10437), .ZN(P1_U3349) );
  OAI222_X1 U13126 ( .A1(n15174), .A2(n10441), .B1(n15188), .B2(n10440), .C1(
        P1_U3086), .C2(n10696), .ZN(P1_U3350) );
  OAI222_X1 U13127 ( .A1(n15174), .A2(n10443), .B1(n15188), .B2(n10442), .C1(
        n6428), .C2(n10616), .ZN(P1_U3352) );
  INV_X1 U13128 ( .A(n10697), .ZN(n10709) );
  OAI222_X1 U13129 ( .A1(n15185), .A2(n10445), .B1(n15188), .B2(n10444), .C1(
        P1_U3086), .C2(n10709), .ZN(P1_U3348) );
  OAI222_X1 U13130 ( .A1(n15174), .A2(n10447), .B1(n15188), .B2(n10446), .C1(
        n6428), .C2(n10617), .ZN(P1_U3351) );
  INV_X1 U13131 ( .A(n10448), .ZN(n10450) );
  OAI222_X1 U13132 ( .A1(n14184), .A2(n10449), .B1(n6438), .B2(n10450), .C1(
        P2_U3088), .C2(n15489), .ZN(P2_U3319) );
  INV_X1 U13133 ( .A(n10874), .ZN(n10693) );
  OAI222_X1 U13134 ( .A1(n15174), .A2(n10451), .B1(n15188), .B2(n10450), .C1(
        P1_U3086), .C2(n10693), .ZN(P1_U3347) );
  OAI222_X1 U13135 ( .A1(n14654), .A2(P1_U3086), .B1(n15188), .B2(n10453), 
        .C1(n10452), .C2(n15174), .ZN(P1_U3354) );
  OAI222_X1 U13136 ( .A1(n11875), .A2(P3_U3151), .B1(n13520), .B2(n10455), 
        .C1(n10454), .C2(n13522), .ZN(P3_U3284) );
  OR2_X1 U13137 ( .A1(n11266), .A2(n14627), .ZN(n10607) );
  AOI21_X1 U13138 ( .B1(n10458), .B2(n10457), .A(n10456), .ZN(n10606) );
  INV_X1 U13139 ( .A(n10606), .ZN(n10459) );
  AND2_X1 U13140 ( .A1(n10607), .A2(n10459), .ZN(n15299) );
  NOR2_X1 U13141 ( .A1(n15299), .A2(P1_U4016), .ZN(P1_U3085) );
  NAND2_X1 U13142 ( .A1(n11266), .A2(n10460), .ZN(n15341) );
  INV_X1 U13143 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13144 ( .A1(n15341), .A2(n10462), .B1(n10464), .B2(n10461), .ZN(
        P1_U3446) );
  INV_X1 U13145 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10466) );
  INV_X1 U13146 ( .A(n10463), .ZN(n10465) );
  AOI22_X1 U13147 ( .A1(n15341), .A2(n10466), .B1(n10465), .B2(n10464), .ZN(
        P1_U3445) );
  OAI222_X1 U13148 ( .A1(n14675), .A2(n6428), .B1(n15188), .B2(n10468), .C1(
        n10467), .C2(n15174), .ZN(P1_U3353) );
  INV_X1 U13149 ( .A(n10469), .ZN(n10470) );
  OAI222_X1 U13150 ( .A1(n14184), .A2(n10484), .B1(n6438), .B2(n10470), .C1(
        P2_U3088), .C2(n6676), .ZN(P2_U3318) );
  INV_X1 U13151 ( .A(n11102), .ZN(n11109) );
  OAI222_X1 U13152 ( .A1(n15174), .A2(n10471), .B1(n15188), .B2(n10470), .C1(
        n6428), .C2(n11109), .ZN(P1_U3346) );
  INV_X1 U13153 ( .A(n10472), .ZN(n10475) );
  INV_X1 U13154 ( .A(n11465), .ZN(n10473) );
  OAI222_X1 U13155 ( .A1(n14184), .A2(n10773), .B1(n6438), .B2(n10475), .C1(
        P2_U3088), .C2(n10473), .ZN(P2_U3317) );
  INV_X1 U13156 ( .A(n14739), .ZN(n10474) );
  OAI222_X1 U13157 ( .A1(n15174), .A2(n10476), .B1(n15188), .B2(n10475), .C1(
        P1_U3086), .C2(n10474), .ZN(P1_U3345) );
  INV_X1 U13158 ( .A(n12980), .ZN(n12988) );
  INV_X1 U13159 ( .A(n10477), .ZN(n10479) );
  OAI222_X1 U13160 ( .A1(n12988), .A2(P3_U3151), .B1(n13520), .B2(n10479), 
        .C1(n10478), .C2(n13522), .ZN(P3_U3283) );
  MUX2_X1 U13161 ( .A(n10480), .B(n11948), .S(P1_U4016), .Z(n10481) );
  INV_X1 U13162 ( .A(n10481), .ZN(P1_U3567) );
  MUX2_X1 U13163 ( .A(n10773), .B(n14439), .S(P1_U4016), .Z(n10482) );
  INV_X1 U13164 ( .A(n10482), .ZN(P1_U3570) );
  MUX2_X1 U13165 ( .A(n10487), .B(n15053), .S(P1_U4016), .Z(n10483) );
  INV_X1 U13166 ( .A(n10483), .ZN(P1_U3571) );
  MUX2_X1 U13167 ( .A(n10484), .B(n11949), .S(P1_U4016), .Z(n10485) );
  INV_X1 U13168 ( .A(n10485), .ZN(P1_U3569) );
  INV_X1 U13169 ( .A(n10486), .ZN(n10488) );
  OAI222_X1 U13170 ( .A1(n14184), .A2(n10487), .B1(n6438), .B2(n10488), .C1(
        P2_U3088), .C2(n11568), .ZN(P2_U3316) );
  INV_X1 U13171 ( .A(n11289), .ZN(n11113) );
  OAI222_X1 U13172 ( .A1(n10489), .A2(n15185), .B1(P1_U3086), .B2(n11113), 
        .C1(n15188), .C2(n10488), .ZN(P1_U3344) );
  NAND2_X1 U13173 ( .A1(n10491), .A2(n10490), .ZN(n10493) );
  NAND2_X1 U13174 ( .A1(n10493), .A2(n10492), .ZN(n10494) );
  OAI21_X1 U13175 ( .B1(n10496), .B2(n10495), .A(n10494), .ZN(n10515) );
  NAND2_X1 U13176 ( .A1(n10515), .A2(n8541), .ZN(n15428) );
  NOR2_X2 U13177 ( .A1(n15428), .A2(P2_U3088), .ZN(n15519) );
  INV_X1 U13178 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10506) );
  INV_X1 U13179 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n11339) );
  MUX2_X1 U13180 ( .A(n11339), .B(P2_REG1_REG_4__SCAN_IN), .S(n10507), .Z(
        n10504) );
  INV_X1 U13181 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10497) );
  MUX2_X1 U13182 ( .A(n10497), .B(P2_REG1_REG_1__SCAN_IN), .S(n15427), .Z(
        n15434) );
  NAND2_X1 U13183 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15438) );
  INV_X1 U13184 ( .A(n15438), .ZN(n10498) );
  NAND2_X1 U13185 ( .A1(n15434), .A2(n10498), .ZN(n15435) );
  NAND2_X1 U13186 ( .A1(n10508), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10499) );
  NAND2_X1 U13187 ( .A1(n15435), .A2(n10499), .ZN(n10588) );
  INV_X1 U13188 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n15562) );
  MUX2_X1 U13189 ( .A(n15562), .B(P2_REG1_REG_2__SCAN_IN), .S(n10598), .Z(
        n10589) );
  NAND2_X1 U13190 ( .A1(n10588), .A2(n10589), .ZN(n10587) );
  NAND2_X1 U13191 ( .A1(n10510), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10500) );
  NAND2_X1 U13192 ( .A1(n10587), .A2(n10500), .ZN(n15448) );
  INV_X1 U13193 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11256) );
  NAND2_X1 U13194 ( .A1(n15448), .A2(n15449), .ZN(n15447) );
  NAND2_X1 U13195 ( .A1(n15453), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10501) );
  NAND2_X1 U13196 ( .A1(n15447), .A2(n10501), .ZN(n10503) );
  OR2_X1 U13197 ( .A1(n8541), .A2(P2_U3088), .ZN(n14177) );
  NOR2_X1 U13198 ( .A1(n14177), .A2(n12571), .ZN(n10502) );
  AND2_X1 U13199 ( .A1(n10515), .A2(n10502), .ZN(n15471) );
  NAND2_X1 U13200 ( .A1(n10503), .A2(n10504), .ZN(n10524) );
  OAI211_X1 U13201 ( .C1(n10504), .C2(n10503), .A(n15471), .B(n10524), .ZN(
        n10505) );
  OAI21_X1 U13202 ( .B1(n10506), .B2(n15522), .A(n10505), .ZN(n10521) );
  MUX2_X1 U13203 ( .A(n12027), .B(P2_REG2_REG_4__SCAN_IN), .S(n10507), .Z(
        n10517) );
  MUX2_X1 U13204 ( .A(n13989), .B(P2_REG2_REG_1__SCAN_IN), .S(n15427), .Z(
        n15432) );
  AND2_X1 U13205 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15431) );
  NAND2_X1 U13206 ( .A1(n15432), .A2(n15431), .ZN(n15430) );
  NAND2_X1 U13207 ( .A1(n10508), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10509) );
  NAND2_X1 U13208 ( .A1(n15430), .A2(n10509), .ZN(n10592) );
  MUX2_X1 U13209 ( .A(n7899), .B(P2_REG2_REG_2__SCAN_IN), .S(n10598), .Z(
        n10593) );
  NAND2_X1 U13210 ( .A1(n10592), .A2(n10593), .ZN(n10591) );
  NAND2_X1 U13211 ( .A1(n10510), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U13212 ( .A1(n10591), .A2(n10511), .ZN(n15445) );
  INV_X1 U13213 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10512) );
  MUX2_X1 U13214 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10512), .S(n15453), .Z(
        n15446) );
  NAND2_X1 U13215 ( .A1(n15445), .A2(n15446), .ZN(n15444) );
  NAND2_X1 U13216 ( .A1(n15453), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10513) );
  NAND2_X1 U13217 ( .A1(n15444), .A2(n10513), .ZN(n10516) );
  NOR2_X1 U13218 ( .A1(n14177), .A2(n14181), .ZN(n10514) );
  NAND2_X1 U13219 ( .A1(n10515), .A2(n10514), .ZN(n15421) );
  NAND2_X1 U13220 ( .A1(n10516), .A2(n10517), .ZN(n10534) );
  OAI211_X1 U13221 ( .C1(n10517), .C2(n10516), .A(n15508), .B(n10534), .ZN(
        n10519) );
  NAND2_X1 U13222 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10518) );
  NAND2_X1 U13223 ( .A1(n10519), .A2(n10518), .ZN(n10520) );
  AOI211_X1 U13224 ( .C1(n10532), .C2(n15519), .A(n10521), .B(n10520), .ZN(
        n10522) );
  INV_X1 U13225 ( .A(n10522), .ZN(P2_U3218) );
  NAND2_X1 U13226 ( .A1(n10532), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10523) );
  NAND2_X1 U13227 ( .A1(n10524), .A2(n10523), .ZN(n15461) );
  INV_X1 U13228 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11319) );
  MUX2_X1 U13229 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n11319), .S(n15466), .Z(
        n15462) );
  NAND2_X1 U13230 ( .A1(n15461), .A2(n15462), .ZN(n15460) );
  NAND2_X1 U13231 ( .A1(n15466), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10525) );
  NAND2_X1 U13232 ( .A1(n15460), .A2(n10525), .ZN(n15472) );
  INV_X1 U13233 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15565) );
  MUX2_X1 U13234 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n15565), .S(n10538), .Z(
        n15473) );
  NAND2_X1 U13235 ( .A1(n15472), .A2(n15473), .ZN(n15470) );
  NAND2_X1 U13236 ( .A1(n10538), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10526) );
  MUX2_X1 U13237 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8019), .S(n10664), .Z(
        n10528) );
  OAI21_X1 U13238 ( .B1(n10528), .B2(n10527), .A(n15471), .ZN(n10544) );
  INV_X1 U13239 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10530) );
  NAND2_X1 U13240 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n10529) );
  OAI21_X1 U13241 ( .B1(n15522), .B2(n10530), .A(n10529), .ZN(n10531) );
  AOI21_X1 U13242 ( .B1(n15519), .B2(n10664), .A(n10531), .ZN(n10543) );
  MUX2_X1 U13243 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11997), .S(n10664), .Z(
        n10541) );
  NAND2_X1 U13244 ( .A1(n10532), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U13245 ( .A1(n10534), .A2(n10533), .ZN(n15458) );
  INV_X1 U13246 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10535) );
  MUX2_X1 U13247 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10535), .S(n15466), .Z(
        n15459) );
  NAND2_X1 U13248 ( .A1(n15458), .A2(n15459), .ZN(n15457) );
  NAND2_X1 U13249 ( .A1(n15466), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10536) );
  NAND2_X1 U13250 ( .A1(n15457), .A2(n10536), .ZN(n15475) );
  XNOR2_X1 U13251 ( .A(n10538), .B(n10537), .ZN(n15476) );
  NAND2_X1 U13252 ( .A1(n15475), .A2(n15476), .ZN(n15474) );
  NAND2_X1 U13253 ( .A1(n10538), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10539) );
  NAND2_X1 U13254 ( .A1(n15474), .A2(n10539), .ZN(n10540) );
  NAND2_X1 U13255 ( .A1(n10540), .A2(n10541), .ZN(n10658) );
  OAI211_X1 U13256 ( .C1(n10541), .C2(n10540), .A(n15508), .B(n10658), .ZN(
        n10542) );
  OAI211_X1 U13257 ( .C1(n10663), .C2(n10544), .A(n10543), .B(n10542), .ZN(
        P2_U3221) );
  INV_X1 U13258 ( .A(n13498), .ZN(n10546) );
  NOR2_X1 U13259 ( .A1(n10546), .A2(n10545), .ZN(n10548) );
  CLKBUF_X1 U13260 ( .A(n10548), .Z(n10565) );
  INV_X1 U13261 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10547) );
  NOR2_X1 U13262 ( .A1(n10565), .A2(n10547), .ZN(P3_U3263) );
  INV_X1 U13263 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10549) );
  NOR2_X1 U13264 ( .A1(n10565), .A2(n10549), .ZN(P3_U3260) );
  INV_X1 U13265 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10550) );
  NOR2_X1 U13266 ( .A1(n10565), .A2(n10550), .ZN(P3_U3259) );
  INV_X1 U13267 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10551) );
  NOR2_X1 U13268 ( .A1(n10548), .A2(n10551), .ZN(P3_U3258) );
  INV_X1 U13269 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10788) );
  NOR2_X1 U13270 ( .A1(n10565), .A2(n10788), .ZN(P3_U3261) );
  INV_X1 U13271 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10552) );
  NOR2_X1 U13272 ( .A1(n10548), .A2(n10552), .ZN(P3_U3262) );
  INV_X1 U13273 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10553) );
  NOR2_X1 U13274 ( .A1(n10565), .A2(n10553), .ZN(P3_U3257) );
  INV_X1 U13275 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10554) );
  NOR2_X1 U13276 ( .A1(n10565), .A2(n10554), .ZN(P3_U3253) );
  INV_X1 U13277 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10555) );
  NOR2_X1 U13278 ( .A1(n10565), .A2(n10555), .ZN(P3_U3256) );
  INV_X1 U13279 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10556) );
  NOR2_X1 U13280 ( .A1(n10565), .A2(n10556), .ZN(P3_U3255) );
  INV_X1 U13281 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10557) );
  NOR2_X1 U13282 ( .A1(n10565), .A2(n10557), .ZN(P3_U3252) );
  INV_X1 U13283 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10558) );
  NOR2_X1 U13284 ( .A1(n10565), .A2(n10558), .ZN(P3_U3251) );
  INV_X1 U13285 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10559) );
  NOR2_X1 U13286 ( .A1(n10565), .A2(n10559), .ZN(P3_U3250) );
  INV_X1 U13287 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10560) );
  NOR2_X1 U13288 ( .A1(n10565), .A2(n10560), .ZN(P3_U3249) );
  INV_X1 U13289 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10561) );
  NOR2_X1 U13290 ( .A1(n10565), .A2(n10561), .ZN(P3_U3248) );
  INV_X1 U13291 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10562) );
  NOR2_X1 U13292 ( .A1(n10565), .A2(n10562), .ZN(P3_U3247) );
  INV_X1 U13293 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10563) );
  NOR2_X1 U13294 ( .A1(n10565), .A2(n10563), .ZN(P3_U3246) );
  INV_X1 U13295 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10564) );
  NOR2_X1 U13296 ( .A1(n10565), .A2(n10564), .ZN(P3_U3254) );
  INV_X1 U13297 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10566) );
  NOR2_X1 U13298 ( .A1(n10548), .A2(n10566), .ZN(P3_U3245) );
  INV_X1 U13299 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10567) );
  NOR2_X1 U13300 ( .A1(n10548), .A2(n10567), .ZN(P3_U3244) );
  INV_X1 U13301 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10568) );
  NOR2_X1 U13302 ( .A1(n10548), .A2(n10568), .ZN(P3_U3243) );
  INV_X1 U13303 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10569) );
  NOR2_X1 U13304 ( .A1(n10548), .A2(n10569), .ZN(P3_U3242) );
  INV_X1 U13305 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10570) );
  NOR2_X1 U13306 ( .A1(n10548), .A2(n10570), .ZN(P3_U3238) );
  INV_X1 U13307 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10571) );
  NOR2_X1 U13308 ( .A1(n10548), .A2(n10571), .ZN(P3_U3241) );
  INV_X1 U13309 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10572) );
  NOR2_X1 U13310 ( .A1(n10548), .A2(n10572), .ZN(P3_U3240) );
  INV_X1 U13311 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10573) );
  NOR2_X1 U13312 ( .A1(n10548), .A2(n10573), .ZN(P3_U3239) );
  INV_X1 U13313 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10574) );
  NOR2_X1 U13314 ( .A1(n10548), .A2(n10574), .ZN(P3_U3237) );
  INV_X1 U13315 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10575) );
  NOR2_X1 U13316 ( .A1(n10565), .A2(n10575), .ZN(P3_U3236) );
  INV_X1 U13317 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10576) );
  NOR2_X1 U13318 ( .A1(n10565), .A2(n10576), .ZN(P3_U3235) );
  INV_X1 U13319 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10577) );
  NOR2_X1 U13320 ( .A1(n10565), .A2(n10577), .ZN(P3_U3234) );
  INV_X1 U13321 ( .A(n10578), .ZN(n10580) );
  INV_X1 U13322 ( .A(n11842), .ZN(n11578) );
  OAI222_X1 U13323 ( .A1(n14184), .A2(n10579), .B1(n6438), .B2(n10580), .C1(
        P2_U3088), .C2(n11578), .ZN(P2_U3315) );
  INV_X1 U13324 ( .A(n11441), .ZN(n11285) );
  OAI222_X1 U13325 ( .A1(n15174), .A2(n10581), .B1(n15188), .B2(n10580), .C1(
        n6428), .C2(n11285), .ZN(P1_U3343) );
  INV_X1 U13326 ( .A(n10582), .ZN(n11824) );
  NAND2_X1 U13327 ( .A1(n13896), .A2(n13951), .ZN(n10583) );
  NOR2_X1 U13328 ( .A1(n12120), .A2(n13932), .ZN(n10635) );
  AOI21_X1 U13329 ( .B1(n11824), .B2(n10583), .A(n10635), .ZN(n11826) );
  INV_X1 U13330 ( .A(n15546), .ZN(n11362) );
  NOR2_X1 U13331 ( .A1(n11353), .A2(n10584), .ZN(n11825) );
  AOI21_X1 U13332 ( .B1(n11824), .B2(n11362), .A(n11825), .ZN(n10585) );
  AND2_X1 U13333 ( .A1(n11826), .A2(n10585), .ZN(n15534) );
  NAND2_X1 U13334 ( .A1(n15567), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10586) );
  OAI21_X1 U13335 ( .B1(n15534), .B2(n15567), .A(n10586), .ZN(P2_U3499) );
  INV_X1 U13336 ( .A(n15519), .ZN(n15490) );
  INV_X1 U13337 ( .A(n15522), .ZN(n15441) );
  OAI211_X1 U13338 ( .C1(n10589), .C2(n10588), .A(n15471), .B(n10587), .ZN(
        n10590) );
  OAI21_X1 U13339 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n12121), .A(n10590), .ZN(
        n10596) );
  OAI211_X1 U13340 ( .C1(n10593), .C2(n10592), .A(n15508), .B(n10591), .ZN(
        n10594) );
  INV_X1 U13341 ( .A(n10594), .ZN(n10595) );
  AOI211_X1 U13342 ( .C1(n15441), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10596), .B(
        n10595), .ZN(n10597) );
  OAI21_X1 U13343 ( .B1(n10598), .B2(n15490), .A(n10597), .ZN(P2_U3216) );
  MUX2_X1 U13344 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10684), .S(n10696), .Z(
        n10605) );
  INV_X1 U13345 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15411) );
  MUX2_X1 U13346 ( .A(n15411), .B(P1_REG1_REG_2__SCAN_IN), .S(n14675), .Z(
        n14682) );
  INV_X1 U13347 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15409) );
  AND2_X1 U13348 ( .A1(n15193), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n14662) );
  INV_X1 U13349 ( .A(n14654), .ZN(n14660) );
  NAND2_X1 U13350 ( .A1(n14660), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U13351 ( .A1(n14661), .A2(n10599), .ZN(n14681) );
  NAND2_X1 U13352 ( .A1(n14682), .A2(n14681), .ZN(n14680) );
  OR2_X1 U13353 ( .A1(n14675), .A2(n15411), .ZN(n10600) );
  NAND2_X1 U13354 ( .A1(n14680), .A2(n10600), .ZN(n14693) );
  XNOR2_X1 U13355 ( .A(n10616), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n14694) );
  NAND2_X1 U13356 ( .A1(n14693), .A2(n14694), .ZN(n14692) );
  INV_X1 U13357 ( .A(n10616), .ZN(n14691) );
  NAND2_X1 U13358 ( .A1(n14691), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13359 ( .A1(n14692), .A2(n10601), .ZN(n14704) );
  XNOR2_X1 U13360 ( .A(n10617), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n14705) );
  NAND2_X1 U13361 ( .A1(n14704), .A2(n14705), .ZN(n14703) );
  INV_X1 U13362 ( .A(n10617), .ZN(n14702) );
  NAND2_X1 U13363 ( .A1(n14702), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10602) );
  INV_X1 U13364 ( .A(n10686), .ZN(n10603) );
  AOI21_X1 U13365 ( .B1(n10605), .B2(n10604), .A(n10603), .ZN(n10624) );
  NAND2_X1 U13366 ( .A1(n10607), .A2(n10606), .ZN(n15302) );
  INV_X1 U13367 ( .A(n15291), .ZN(n14576) );
  NOR2_X2 U13368 ( .A1(n15302), .A2(n14576), .ZN(n15310) );
  NOR2_X2 U13369 ( .A1(n15302), .A2(n10608), .ZN(n14783) );
  INV_X1 U13370 ( .A(n15299), .ZN(n15319) );
  INV_X1 U13371 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U13372 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11608) );
  OAI21_X1 U13373 ( .B1(n15319), .B2(n10609), .A(n11608), .ZN(n10610) );
  AOI21_X1 U13374 ( .B1(n10611), .B2(n14783), .A(n10610), .ZN(n10623) );
  INV_X1 U13375 ( .A(n15302), .ZN(n10613) );
  NOR2_X1 U13376 ( .A1(n14671), .A2(n15291), .ZN(n10612) );
  NAND2_X1 U13377 ( .A1(n10613), .A2(n10612), .ZN(n15305) );
  AOI21_X1 U13378 ( .B1(n14660), .B2(P1_REG2_REG_1__SCAN_IN), .A(n14656), .ZN(
        n14677) );
  MUX2_X1 U13379 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n14676), .S(n14675), .Z(
        n10614) );
  OR2_X1 U13380 ( .A1(n14677), .A2(n10614), .ZN(n14688) );
  INV_X1 U13381 ( .A(n14675), .ZN(n14674) );
  NAND2_X1 U13382 ( .A1(n14674), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14687) );
  MUX2_X1 U13383 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10615), .S(n10616), .Z(
        n14686) );
  AOI21_X1 U13384 ( .B1(n14688), .B2(n14687), .A(n14686), .ZN(n14708) );
  NOR2_X1 U13385 ( .A1(n10616), .A2(n10615), .ZN(n14707) );
  MUX2_X1 U13386 ( .A(n11552), .B(P1_REG2_REG_4__SCAN_IN), .S(n10617), .Z(
        n14706) );
  NAND2_X1 U13387 ( .A1(n14702), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10619) );
  MUX2_X1 U13388 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11594), .S(n10696), .Z(
        n10618) );
  INV_X1 U13389 ( .A(n14717), .ZN(n10621) );
  NAND3_X1 U13390 ( .A1(n14710), .A2(n10619), .A3(n10618), .ZN(n10620) );
  NAND3_X1 U13391 ( .A1(n14785), .A2(n10621), .A3(n10620), .ZN(n10622) );
  OAI211_X1 U13392 ( .C1(n10624), .C2(n6633), .A(n10623), .B(n10622), .ZN(
        P1_U3248) );
  INV_X1 U13393 ( .A(n10625), .ZN(n10627) );
  INV_X1 U13394 ( .A(n13018), .ZN(n13004) );
  OAI222_X1 U13395 ( .A1(n13520), .A2(n10627), .B1(n13522), .B2(n10626), .C1(
        n13004), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U13396 ( .A(n10628), .ZN(n10630) );
  OAI222_X1 U13397 ( .A1(n13058), .A2(P3_U3151), .B1(n13520), .B2(n10630), 
        .C1(n10629), .C2(n13522), .ZN(P3_U3280) );
  NOR2_X1 U13398 ( .A1(n10631), .A2(P2_U3088), .ZN(n11190) );
  INV_X1 U13399 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10640) );
  OAI21_X1 U13400 ( .B1(n10634), .B2(n12569), .A(n10633), .ZN(n10636) );
  AOI22_X1 U13401 ( .A1(n13610), .A2(n10636), .B1(n13643), .B2(n10635), .ZN(
        n10639) );
  NAND2_X1 U13402 ( .A1(n13647), .A2(n10637), .ZN(n10638) );
  OAI211_X1 U13403 ( .C1(n11190), .C2(n10640), .A(n10639), .B(n10638), .ZN(
        P2_U3204) );
  INV_X1 U13404 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n10848) );
  NAND2_X1 U13405 ( .A1(P3_U3897), .A2(n12837), .ZN(n10641) );
  OAI21_X1 U13406 ( .B1(P3_U3897), .B2(n10848), .A(n10641), .ZN(P3_U3498) );
  OAI22_X1 U13407 ( .A1(n10642), .A2(n13930), .B1(n11251), .B2(n13932), .ZN(
        n11360) );
  AOI22_X1 U13408 ( .A1(n6645), .A2(n13647), .B1(n13643), .B2(n11360), .ZN(
        n10648) );
  OAI21_X1 U13409 ( .B1(n10645), .B2(n10644), .A(n10643), .ZN(n10646) );
  NAND2_X1 U13410 ( .A1(n13610), .A2(n10646), .ZN(n10647) );
  OAI211_X1 U13411 ( .C1(n11190), .C2(n10649), .A(n10648), .B(n10647), .ZN(
        P2_U3194) );
  INV_X1 U13412 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n10762) );
  NAND2_X1 U13413 ( .A1(n11855), .A2(P3_U3897), .ZN(n10650) );
  OAI21_X1 U13414 ( .B1(P3_U3897), .B2(n10762), .A(n10650), .ZN(P3_U3499) );
  INV_X1 U13415 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n10805) );
  NAND2_X1 U13416 ( .A1(n12681), .A2(P3_U3897), .ZN(n10651) );
  OAI21_X1 U13417 ( .B1(P3_U3897), .B2(n10805), .A(n10651), .ZN(P3_U3508) );
  INV_X1 U13418 ( .A(n14374), .ZN(n14336) );
  NAND2_X1 U13419 ( .A1(n10652), .A2(n14577), .ZN(n14234) );
  AOI22_X1 U13420 ( .A1(n14336), .A2(n11380), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n14234), .ZN(n10656) );
  XNOR2_X1 U13421 ( .A(n10654), .B(n10653), .ZN(n14668) );
  NAND2_X1 U13422 ( .A1(n14668), .A2(n14370), .ZN(n10655) );
  OAI211_X1 U13423 ( .C1(n14380), .C2(n11378), .A(n10656), .B(n10655), .ZN(
        P1_U3232) );
  MUX2_X1 U13424 ( .A(n11979), .B(P2_REG2_REG_9__SCAN_IN), .S(n11168), .Z(
        n10662) );
  NAND2_X1 U13425 ( .A1(n10664), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10657) );
  NAND2_X1 U13426 ( .A1(n10658), .A2(n10657), .ZN(n15486) );
  MUX2_X1 U13427 ( .A(n12010), .B(P2_REG2_REG_8__SCAN_IN), .S(n15489), .Z(
        n15487) );
  NAND2_X1 U13428 ( .A1(n15486), .A2(n15487), .ZN(n15485) );
  NAND2_X1 U13429 ( .A1(n10665), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10659) );
  NAND2_X1 U13430 ( .A1(n15485), .A2(n10659), .ZN(n10661) );
  INV_X1 U13431 ( .A(n11170), .ZN(n10660) );
  AOI21_X1 U13432 ( .B1(n10662), .B2(n10661), .A(n10660), .ZN(n10673) );
  XNOR2_X1 U13433 ( .A(n11168), .B(n6675), .ZN(n10667) );
  XNOR2_X1 U13434 ( .A(n10665), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n15483) );
  AOI21_X1 U13435 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n10665), .A(n6502), .ZN(
        n10666) );
  OAI21_X1 U13436 ( .B1(n10667), .B2(n10666), .A(n11164), .ZN(n10668) );
  NAND2_X1 U13437 ( .A1(n10668), .A2(n15471), .ZN(n10672) );
  NOR2_X1 U13438 ( .A1(n10669), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11703) );
  NOR2_X1 U13439 ( .A1(n15490), .A2(n6676), .ZN(n10670) );
  AOI211_X1 U13440 ( .C1(n15441), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n11703), .B(
        n10670), .ZN(n10671) );
  OAI211_X1 U13441 ( .C1(n10673), .C2(n15421), .A(n10672), .B(n10671), .ZN(
        P2_U3223) );
  INV_X1 U13442 ( .A(n13028), .ZN(n10677) );
  INV_X1 U13443 ( .A(n10674), .ZN(n10676) );
  OAI222_X1 U13444 ( .A1(n10677), .A2(P3_U3151), .B1(n13520), .B2(n10676), 
        .C1(n10675), .C2(n13522), .ZN(P3_U3281) );
  INV_X1 U13445 ( .A(n10678), .ZN(n10680) );
  INV_X1 U13446 ( .A(n12392), .ZN(n11852) );
  OAI222_X1 U13447 ( .A1(n14184), .A2(n10679), .B1(n6438), .B2(n10680), .C1(
        P2_U3088), .C2(n11852), .ZN(P2_U3314) );
  INV_X1 U13448 ( .A(n11711), .ZN(n11718) );
  OAI222_X1 U13449 ( .A1(n15174), .A2(n10681), .B1(n15188), .B2(n10680), .C1(
        P1_U3086), .C2(n11718), .ZN(P1_U3342) );
  OAI222_X1 U13450 ( .A1(n13104), .A2(P3_U3151), .B1(n13520), .B2(n10683), 
        .C1(n10682), .C2(n13522), .ZN(P3_U3278) );
  MUX2_X1 U13451 ( .A(n9328), .B(P1_REG1_REG_8__SCAN_IN), .S(n10874), .Z(
        n10692) );
  NAND2_X1 U13452 ( .A1(n10696), .A2(n10684), .ZN(n10685) );
  INV_X1 U13453 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10687) );
  XNOR2_X1 U13454 ( .A(n14724), .B(n10687), .ZN(n14723) );
  NAND2_X1 U13455 ( .A1(n14722), .A2(n14723), .ZN(n14721) );
  NAND2_X1 U13456 ( .A1(n14724), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10688) );
  NAND2_X1 U13457 ( .A1(n14721), .A2(n10688), .ZN(n10712) );
  MUX2_X1 U13458 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9229), .S(n10697), .Z(
        n10713) );
  NAND2_X1 U13459 ( .A1(n10712), .A2(n10713), .ZN(n10711) );
  NAND2_X1 U13460 ( .A1(n10697), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10689) );
  NAND2_X1 U13461 ( .A1(n10711), .A2(n10689), .ZN(n10691) );
  INV_X1 U13462 ( .A(n10876), .ZN(n10690) );
  AOI21_X1 U13463 ( .B1(n10692), .B2(n10691), .A(n10690), .ZN(n10704) );
  AND2_X1 U13464 ( .A1(n6428), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10695) );
  INV_X1 U13465 ( .A(n14783), .ZN(n15315) );
  NOR2_X1 U13466 ( .A1(n15315), .A2(n10693), .ZN(n10694) );
  AOI211_X1 U13467 ( .C1(n15299), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10695), .B(
        n10694), .ZN(n10703) );
  NOR2_X1 U13468 ( .A1(n10696), .A2(n11594), .ZN(n14716) );
  MUX2_X1 U13469 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11643), .S(n14724), .Z(
        n14715) );
  NAND2_X1 U13470 ( .A1(n14724), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10706) );
  MUX2_X1 U13471 ( .A(n11685), .B(P1_REG2_REG_7__SCAN_IN), .S(n10697), .Z(
        n10705) );
  NOR2_X1 U13472 ( .A1(n10709), .A2(n11685), .ZN(n10700) );
  MUX2_X1 U13473 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10698), .S(n10874), .Z(
        n10699) );
  OAI21_X1 U13474 ( .B1(n10717), .B2(n10700), .A(n10699), .ZN(n10869) );
  OR3_X1 U13475 ( .A1(n10717), .A2(n10700), .A3(n10699), .ZN(n10701) );
  NAND3_X1 U13476 ( .A1(n10869), .A2(n14785), .A3(n10701), .ZN(n10702) );
  OAI211_X1 U13477 ( .C1(n10704), .C2(n6633), .A(n10703), .B(n10702), .ZN(
        P1_U3251) );
  NAND3_X1 U13478 ( .A1(n14719), .A2(n10706), .A3(n10705), .ZN(n10707) );
  NAND2_X1 U13479 ( .A1(n10707), .A2(n14785), .ZN(n10716) );
  NOR2_X1 U13480 ( .A1(n10708), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11745) );
  NOR2_X1 U13481 ( .A1(n15315), .A2(n10709), .ZN(n10710) );
  AOI211_X1 U13482 ( .C1(n15299), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n11745), .B(
        n10710), .ZN(n10715) );
  OAI211_X1 U13483 ( .C1(n10713), .C2(n10712), .A(n15310), .B(n10711), .ZN(
        n10714) );
  OAI211_X1 U13484 ( .C1(n10717), .C2(n10716), .A(n10715), .B(n10714), .ZN(
        P1_U3250) );
  INV_X2 U13485 ( .A(n15418), .ZN(n15420) );
  INV_X1 U13486 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15290) );
  OR2_X1 U13487 ( .A1(n11377), .A2(n11453), .ZN(n10719) );
  NAND2_X1 U13488 ( .A1(n11377), .A2(n11453), .ZN(n11260) );
  AND2_X1 U13489 ( .A1(n10719), .A2(n11260), .ZN(n14388) );
  INV_X1 U13490 ( .A(n14388), .ZN(n14581) );
  OAI21_X1 U13491 ( .B1(n14387), .B2(n14383), .A(n10720), .ZN(n11448) );
  OR2_X1 U13492 ( .A1(n11448), .A2(n14381), .ZN(n15375) );
  NAND2_X1 U13493 ( .A1(n14535), .A2(n14381), .ZN(n15374) );
  NAND2_X1 U13494 ( .A1(n15375), .A2(n15374), .ZN(n15395) );
  OAI22_X1 U13495 ( .A1(n14581), .A2(n15404), .B1(n11378), .B2(n10721), .ZN(
        n10726) );
  INV_X1 U13496 ( .A(n11709), .ZN(n14384) );
  NAND2_X1 U13497 ( .A1(n9219), .A2(n14384), .ZN(n10723) );
  NAND2_X1 U13498 ( .A1(n15190), .A2(n14381), .ZN(n10722) );
  NAND2_X1 U13499 ( .A1(n14388), .A2(n15024), .ZN(n10725) );
  NAND2_X1 U13500 ( .A1(n11380), .A2(n15222), .ZN(n10724) );
  NAND2_X1 U13501 ( .A1(n10725), .A2(n10724), .ZN(n11452) );
  OR2_X1 U13502 ( .A1(n10726), .A2(n11452), .ZN(n10728) );
  NAND2_X1 U13503 ( .A1(n10728), .A2(n15420), .ZN(n10727) );
  OAI21_X1 U13504 ( .B1(n15420), .B2(n15290), .A(n10727), .ZN(P1_U3528) );
  INV_X1 U13505 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10730) );
  NAND2_X1 U13506 ( .A1(n10728), .A2(n15408), .ZN(n10729) );
  OAI21_X1 U13507 ( .B1(n15408), .B2(n10730), .A(n10729), .ZN(P1_U3459) );
  AOI222_X1 U13508 ( .A1(n10732), .A2(n13500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13091), .C1(SI_16_), .C2(n10731), .ZN(n10866) );
  NAND4_X1 U13509 ( .A1(P2_REG0_REG_11__SCAN_IN), .A2(P3_DATAO_REG_19__SCAN_IN), .A3(n10825), .A4(n10615), .ZN(n10754) );
  NOR3_X1 U13510 ( .A1(P2_REG2_REG_31__SCAN_IN), .A2(P3_DATAO_REG_17__SCAN_IN), 
        .A3(n10918), .ZN(n10736) );
  NOR4_X1 U13511 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_REG0_REG_27__SCAN_IN), 
        .A3(n13903), .A4(n12221), .ZN(n10733) );
  NAND4_X1 U13512 ( .A1(n12121), .A2(P2_REG1_REG_0__SCAN_IN), .A3(
        P2_IR_REG_7__SCAN_IN), .A4(n10733), .ZN(n10734) );
  NOR3_X1 U13513 ( .A1(n10734), .A2(P3_IR_REG_29__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .ZN(n10735) );
  NAND2_X1 U13514 ( .A1(n10736), .A2(n10735), .ZN(n10753) );
  NOR4_X1 U13515 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .A3(n15656), .A4(n15456), .ZN(n10751) );
  NAND4_X1 U13516 ( .A1(P3_REG2_REG_28__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .A3(P1_REG2_REG_6__SCAN_IN), .A4(P3_DATAO_REG_8__SCAN_IN), .ZN(n10741)
         );
  INV_X1 U13517 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n10737) );
  NAND4_X1 U13518 ( .A1(n10738), .A2(n10737), .A3(P1_DATAO_REG_12__SCAN_IN), 
        .A4(P1_DATAO_REG_10__SCAN_IN), .ZN(n10740) );
  NAND4_X1 U13519 ( .A1(n10798), .A2(n13502), .A3(P3_IR_REG_8__SCAN_IN), .A4(
        P2_ADDR_REG_5__SCAN_IN), .ZN(n10739) );
  NOR3_X1 U13520 ( .A1(n10741), .A2(n10740), .A3(n10739), .ZN(n10750) );
  NOR4_X1 U13521 ( .A1(SI_0_), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P3_ADDR_REG_13__SCAN_IN), .A4(P3_DATAO_REG_7__SCAN_IN), .ZN(n10749) );
  NAND4_X1 U13522 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_REG0_REG_22__SCAN_IN), 
        .A3(P1_REG0_REG_13__SCAN_IN), .A4(P3_DATAO_REG_30__SCAN_IN), .ZN(
        n10747) );
  NAND4_X1 U13523 ( .A1(n12984), .A2(n10742), .A3(P2_REG2_REG_7__SCAN_IN), 
        .A4(n13989), .ZN(n10746) );
  NAND4_X1 U13524 ( .A1(n10744), .A2(n10743), .A3(P3_REG0_REG_31__SCAN_IN), 
        .A4(P3_REG3_REG_20__SCAN_IN), .ZN(n10745) );
  NOR3_X1 U13525 ( .A1(n10747), .A2(n10746), .A3(n10745), .ZN(n10748) );
  NAND4_X1 U13526 ( .A1(n10751), .A2(n10750), .A3(n10749), .A4(n10748), .ZN(
        n10752) );
  NOR3_X1 U13527 ( .A1(n10754), .A2(n10753), .A3(n10752), .ZN(n10864) );
  INV_X1 U13528 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11424) );
  NAND4_X1 U13529 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_WR_REG_SCAN_IN), .A3(
        n11424), .A4(n10755), .ZN(n10760) );
  NAND4_X1 U13530 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(P3_REG3_REG_28__SCAN_IN), 
        .A3(P1_IR_REG_20__SCAN_IN), .A4(n15409), .ZN(n10758) );
  NAND4_X1 U13531 ( .A1(P3_B_REG_SCAN_IN), .A2(P2_REG1_REG_6__SCAN_IN), .A3(
        n11528), .A4(n10756), .ZN(n10757) );
  OR4_X1 U13532 ( .A1(n10788), .A2(P3_REG2_REG_15__SCAN_IN), .A3(n10758), .A4(
        n10757), .ZN(n10759) );
  INV_X1 U13533 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10787) );
  NOR4_X1 U13534 ( .A1(n10760), .A2(n10759), .A3(P1_IR_REG_8__SCAN_IN), .A4(
        n10787), .ZN(n10863) );
  AOI22_X1 U13535 ( .A1(n13180), .A2(keyinput11), .B1(keyinput38), .B2(n10762), 
        .ZN(n10761) );
  OAI221_X1 U13536 ( .B1(n13180), .B2(keyinput11), .C1(n10762), .C2(keyinput38), .A(n10761), .ZN(n10771) );
  AOI22_X1 U13537 ( .A1(n11424), .A2(keyinput7), .B1(keyinput57), .B2(n10764), 
        .ZN(n10763) );
  OAI221_X1 U13538 ( .B1(n11424), .B2(keyinput7), .C1(n10764), .C2(keyinput57), 
        .A(n10763), .ZN(n10770) );
  XNOR2_X1 U13539 ( .A(keyinput24), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n10768) );
  XNOR2_X1 U13540 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput22), .ZN(n10767) );
  XNOR2_X1 U13541 ( .A(P1_REG0_REG_14__SCAN_IN), .B(keyinput48), .ZN(n10766)
         );
  XNOR2_X1 U13542 ( .A(P3_IR_REG_4__SCAN_IN), .B(keyinput4), .ZN(n10765) );
  NAND4_X1 U13543 ( .A1(n10768), .A2(n10767), .A3(n10766), .A4(n10765), .ZN(
        n10769) );
  NOR3_X1 U13544 ( .A1(n10771), .A2(n10770), .A3(n10769), .ZN(n10812) );
  AOI22_X1 U13545 ( .A1(n11528), .A2(keyinput59), .B1(keyinput32), .B2(n9098), 
        .ZN(n10772) );
  OAI221_X1 U13546 ( .B1(n11528), .B2(keyinput59), .C1(n9098), .C2(keyinput32), 
        .A(n10772), .ZN(n10783) );
  XNOR2_X1 U13547 ( .A(keyinput5), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n10779) );
  XNOR2_X1 U13548 ( .A(keyinput26), .B(n10773), .ZN(n10775) );
  XOR2_X1 U13549 ( .A(P1_REG0_REG_28__SCAN_IN), .B(keyinput43), .Z(n10774) );
  NOR2_X1 U13550 ( .A1(n10775), .A2(n10774), .ZN(n10778) );
  XNOR2_X1 U13551 ( .A(P3_B_REG_SCAN_IN), .B(keyinput14), .ZN(n10777) );
  XNOR2_X1 U13552 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput27), .ZN(n10776) );
  NAND4_X1 U13553 ( .A1(n10779), .A2(n10778), .A3(n10777), .A4(n10776), .ZN(
        n10782) );
  INV_X1 U13554 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10780) );
  XNOR2_X1 U13555 ( .A(n10780), .B(keyinput49), .ZN(n10781) );
  NOR3_X1 U13556 ( .A1(n10783), .A2(n10782), .A3(n10781), .ZN(n10811) );
  INV_X1 U13557 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U13558 ( .A1(n15409), .A2(keyinput63), .B1(n10785), .B2(keyinput29), 
        .ZN(n10784) );
  OAI221_X1 U13559 ( .B1(n15409), .B2(keyinput63), .C1(n10785), .C2(keyinput29), .A(n10784), .ZN(n10795) );
  AOI22_X1 U13560 ( .A1(n13036), .A2(keyinput61), .B1(keyinput15), .B2(n10787), 
        .ZN(n10786) );
  OAI221_X1 U13561 ( .B1(n13036), .B2(keyinput61), .C1(n10787), .C2(keyinput15), .A(n10786), .ZN(n10794) );
  XOR2_X1 U13562 ( .A(n10788), .B(keyinput8), .Z(n10792) );
  XNOR2_X1 U13563 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput23), .ZN(n10791) );
  XNOR2_X1 U13564 ( .A(P3_REG1_REG_12__SCAN_IN), .B(keyinput35), .ZN(n10790)
         );
  XNOR2_X1 U13565 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput34), .ZN(n10789) );
  NAND4_X1 U13566 ( .A1(n10792), .A2(n10791), .A3(n10790), .A4(n10789), .ZN(
        n10793) );
  NOR3_X1 U13567 ( .A1(n10795), .A2(n10794), .A3(n10793), .ZN(n10810) );
  INV_X1 U13568 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U13569 ( .A1(n10797), .A2(keyinput56), .B1(n7152), .B2(keyinput45), 
        .ZN(n10796) );
  OAI221_X1 U13570 ( .B1(n10797), .B2(keyinput56), .C1(n7152), .C2(keyinput45), 
        .A(n10796), .ZN(n10808) );
  XOR2_X1 U13571 ( .A(n12121), .B(keyinput39), .Z(n10804) );
  XNOR2_X1 U13572 ( .A(keyinput50), .B(n10798), .ZN(n10801) );
  XOR2_X1 U13573 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput60), .Z(n10800) );
  XNOR2_X1 U13574 ( .A(n10918), .B(keyinput44), .ZN(n10799) );
  NOR3_X1 U13575 ( .A1(n10801), .A2(n10800), .A3(n10799), .ZN(n10803) );
  XNOR2_X1 U13576 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput12), .ZN(n10802) );
  NAND3_X1 U13577 ( .A1(n10804), .A2(n10803), .A3(n10802), .ZN(n10807) );
  XNOR2_X1 U13578 ( .A(n10805), .B(keyinput10), .ZN(n10806) );
  NOR3_X1 U13579 ( .A1(n10808), .A2(n10807), .A3(n10806), .ZN(n10809) );
  NAND4_X1 U13580 ( .A1(n10812), .A2(n10811), .A3(n10810), .A4(n10809), .ZN(
        n10862) );
  INV_X1 U13581 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13582 ( .A1(n7161), .A2(keyinput47), .B1(keyinput52), .B2(n10814), 
        .ZN(n10813) );
  OAI221_X1 U13583 ( .B1(n7161), .B2(keyinput47), .C1(n10814), .C2(keyinput52), 
        .A(n10813), .ZN(n10823) );
  INV_X1 U13584 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U13585 ( .A1(n12274), .A2(keyinput25), .B1(n10816), .B2(keyinput37), 
        .ZN(n10815) );
  OAI221_X1 U13586 ( .B1(n12274), .B2(keyinput25), .C1(n10816), .C2(keyinput37), .A(n10815), .ZN(n10822) );
  INV_X1 U13587 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13421) );
  AOI22_X1 U13588 ( .A1(n12984), .A2(keyinput36), .B1(keyinput54), .B2(n13421), 
        .ZN(n10817) );
  OAI221_X1 U13589 ( .B1(n12984), .B2(keyinput36), .C1(n13421), .C2(keyinput54), .A(n10817), .ZN(n10821) );
  XOR2_X1 U13590 ( .A(n12221), .B(keyinput6), .Z(n10819) );
  XNOR2_X1 U13591 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput33), .ZN(n10818) );
  NAND2_X1 U13592 ( .A1(n10819), .A2(n10818), .ZN(n10820) );
  NOR4_X1 U13593 ( .A1(n10823), .A2(n10822), .A3(n10821), .A4(n10820), .ZN(
        n10860) );
  AOI22_X1 U13594 ( .A1(n10825), .A2(keyinput51), .B1(keyinput21), .B2(n10615), 
        .ZN(n10824) );
  OAI221_X1 U13595 ( .B1(n10825), .B2(keyinput51), .C1(n10615), .C2(keyinput21), .A(n10824), .ZN(n10835) );
  AOI22_X1 U13596 ( .A1(n10827), .A2(keyinput62), .B1(n14158), .B2(keyinput41), 
        .ZN(n10826) );
  OAI221_X1 U13597 ( .B1(n10827), .B2(keyinput62), .C1(n14158), .C2(keyinput41), .A(n10826), .ZN(n10834) );
  AOI22_X1 U13598 ( .A1(n10830), .A2(keyinput53), .B1(n10829), .B2(keyinput42), 
        .ZN(n10828) );
  OAI221_X1 U13599 ( .B1(n10830), .B2(keyinput53), .C1(n10829), .C2(keyinput42), .A(n10828), .ZN(n10833) );
  INV_X1 U13600 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U13601 ( .A1(n10884), .A2(keyinput46), .B1(n13903), .B2(keyinput40), 
        .ZN(n10831) );
  OAI221_X1 U13602 ( .B1(n10884), .B2(keyinput46), .C1(n13903), .C2(keyinput40), .A(n10831), .ZN(n10832) );
  NOR4_X1 U13603 ( .A1(n10835), .A2(n10834), .A3(n10833), .A4(n10832), .ZN(
        n10859) );
  AOI22_X1 U13604 ( .A1(n15656), .A2(keyinput18), .B1(n10837), .B2(keyinput3), 
        .ZN(n10836) );
  OAI221_X1 U13605 ( .B1(n15656), .B2(keyinput18), .C1(n10837), .C2(keyinput3), 
        .A(n10836), .ZN(n10846) );
  INV_X1 U13606 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15525) );
  AOI22_X1 U13607 ( .A1(n15456), .A2(keyinput1), .B1(n15525), .B2(keyinput58), 
        .ZN(n10838) );
  OAI221_X1 U13608 ( .B1(n15456), .B2(keyinput1), .C1(n15525), .C2(keyinput58), 
        .A(n10838), .ZN(n10845) );
  XOR2_X1 U13609 ( .A(n10839), .B(keyinput13), .Z(n10843) );
  XNOR2_X1 U13610 ( .A(SI_0_), .B(keyinput17), .ZN(n10842) );
  XNOR2_X1 U13611 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput28), .ZN(n10841)
         );
  XNOR2_X1 U13612 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(keyinput16), .ZN(n10840)
         );
  NAND4_X1 U13613 ( .A1(n10843), .A2(n10842), .A3(n10841), .A4(n10840), .ZN(
        n10844) );
  NOR3_X1 U13614 ( .A1(n10846), .A2(n10845), .A3(n10844), .ZN(n10858) );
  AOI22_X1 U13615 ( .A1(n13989), .A2(keyinput30), .B1(keyinput9), .B2(n10848), 
        .ZN(n10847) );
  OAI221_X1 U13616 ( .B1(n13989), .B2(keyinput30), .C1(n10848), .C2(keyinput9), 
        .A(n10847), .ZN(n10856) );
  XNOR2_X1 U13617 ( .A(keyinput31), .B(n9384), .ZN(n10855) );
  INV_X1 U13618 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15469) );
  XNOR2_X1 U13619 ( .A(keyinput0), .B(n15469), .ZN(n10854) );
  XNOR2_X1 U13620 ( .A(P3_IR_REG_31__SCAN_IN), .B(keyinput55), .ZN(n10852) );
  XNOR2_X1 U13621 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput2), .ZN(n10851) );
  XNOR2_X1 U13622 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput20), .ZN(n10850) );
  XNOR2_X1 U13623 ( .A(keyinput19), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n10849) );
  NAND4_X1 U13624 ( .A1(n10852), .A2(n10851), .A3(n10850), .A4(n10849), .ZN(
        n10853) );
  NOR4_X1 U13625 ( .A1(n10856), .A2(n10855), .A3(n10854), .A4(n10853), .ZN(
        n10857) );
  NAND4_X1 U13626 ( .A1(n10860), .A2(n10859), .A3(n10858), .A4(n10857), .ZN(
        n10861) );
  AOI211_X1 U13627 ( .C1(n10864), .C2(n10863), .A(n10862), .B(n10861), .ZN(
        n10865) );
  XNOR2_X1 U13628 ( .A(n10866), .B(n10865), .ZN(P3_U3279) );
  NAND2_X1 U13629 ( .A1(n10874), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10868) );
  MUX2_X1 U13630 ( .A(n12221), .B(P1_REG2_REG_9__SCAN_IN), .S(n11102), .Z(
        n10867) );
  AOI21_X1 U13631 ( .B1(n10869), .B2(n10868), .A(n10867), .ZN(n14731) );
  NAND3_X1 U13632 ( .A1(n10869), .A2(n10868), .A3(n10867), .ZN(n10870) );
  NAND2_X1 U13633 ( .A1(n10870), .A2(n14785), .ZN(n10882) );
  NOR2_X1 U13634 ( .A1(n10871), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12262) );
  NOR2_X1 U13635 ( .A1(n15315), .A2(n11109), .ZN(n10872) );
  AOI211_X1 U13636 ( .C1(n15299), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n12262), .B(
        n10872), .ZN(n10881) );
  MUX2_X1 U13637 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10873), .S(n11102), .Z(
        n10878) );
  OR2_X1 U13638 ( .A1(n10874), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10875) );
  OAI21_X1 U13639 ( .B1(n10878), .B2(n10877), .A(n11104), .ZN(n10879) );
  NAND2_X1 U13640 ( .A1(n10879), .A2(n15310), .ZN(n10880) );
  OAI211_X1 U13641 ( .C1(n14731), .C2(n10882), .A(n10881), .B(n10880), .ZN(
        P1_U3252) );
  NAND2_X1 U13642 ( .A1(n12710), .A2(P3_U3897), .ZN(n10883) );
  OAI21_X1 U13643 ( .B1(P3_U3897), .B2(n10884), .A(n10883), .ZN(P3_U3510) );
  INV_X1 U13644 ( .A(n10885), .ZN(n10886) );
  AOI21_X1 U13645 ( .B1(n10888), .B2(n10887), .A(n10886), .ZN(n10895) );
  INV_X1 U13646 ( .A(n12028), .ZN(n10893) );
  NAND2_X1 U13647 ( .A1(n13669), .A2(n13968), .ZN(n10890) );
  NAND2_X1 U13648 ( .A1(n13671), .A2(n13966), .ZN(n10889) );
  NAND2_X1 U13649 ( .A1(n10890), .A2(n10889), .ZN(n11325) );
  AOI22_X1 U13650 ( .A1(n13643), .A2(n11325), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10891) );
  OAI21_X1 U13651 ( .B1(n13620), .B2(n12029), .A(n10891), .ZN(n10892) );
  AOI21_X1 U13652 ( .B1(n10893), .B2(n13631), .A(n10892), .ZN(n10894) );
  OAI21_X1 U13653 ( .B1(n10895), .B2(n13649), .A(n10894), .ZN(P2_U3202) );
  OR2_X1 U13654 ( .A1(n10918), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10896) );
  INV_X1 U13655 ( .A(n10896), .ZN(n11434) );
  INV_X1 U13656 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U13657 ( .A1(n10965), .A2(n10897), .ZN(n11024) );
  OR2_X1 U13658 ( .A1(n10943), .A2(n10919), .ZN(n10898) );
  XNOR2_X1 U13659 ( .A(n10899), .B(n10924), .ZN(n11004) );
  NAND2_X1 U13660 ( .A1(n10899), .A2(n11018), .ZN(n10900) );
  MUX2_X1 U13661 ( .A(n10901), .B(P3_REG1_REG_4__SCAN_IN), .S(n10979), .Z(
        n10982) );
  OR2_X1 U13662 ( .A1(n10979), .A2(n10901), .ZN(n10902) );
  XNOR2_X1 U13663 ( .A(n10903), .B(n10934), .ZN(n11084) );
  NAND2_X1 U13664 ( .A1(n11084), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10905) );
  NAND2_X1 U13665 ( .A1(n10903), .A2(n11089), .ZN(n10904) );
  NAND2_X1 U13666 ( .A1(n10905), .A2(n10904), .ZN(n11122) );
  MUX2_X1 U13667 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10906), .S(n11130), .Z(
        n11123) );
  NAND2_X1 U13668 ( .A1(n11122), .A2(n11123), .ZN(n11121) );
  NAND2_X1 U13669 ( .A1(n11130), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U13670 ( .A1(n11121), .A2(n10907), .ZN(n11057) );
  XNOR2_X1 U13671 ( .A(n11057), .B(n11063), .ZN(n11055) );
  INV_X1 U13672 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11871) );
  XNOR2_X1 U13673 ( .A(n11055), .B(n11871), .ZN(n10962) );
  OR2_X1 U13674 ( .A1(n10910), .A2(P3_U3151), .ZN(n12959) );
  INV_X1 U13675 ( .A(n12959), .ZN(n10908) );
  OR2_X1 U13676 ( .A1(n10909), .A2(n10908), .ZN(n10956) );
  NAND2_X1 U13677 ( .A1(n12930), .A2(n10910), .ZN(n10912) );
  NAND2_X1 U13678 ( .A1(n10912), .A2(n6924), .ZN(n10955) );
  INV_X1 U13679 ( .A(n10955), .ZN(n10913) );
  NAND2_X1 U13680 ( .A1(n10953), .A2(n7029), .ZN(n13143) );
  INV_X1 U13681 ( .A(n10978), .ZN(n10914) );
  NAND2_X1 U13682 ( .A1(n10915), .A2(n10914), .ZN(n11031) );
  INV_X1 U13683 ( .A(n10915), .ZN(n10916) );
  NAND2_X1 U13684 ( .A1(n10916), .A2(n10978), .ZN(n10917) );
  NAND2_X1 U13685 ( .A1(n11030), .A2(n11031), .ZN(n10923) );
  MUX2_X1 U13686 ( .A(n15592), .B(n10919), .S(n13039), .Z(n10920) );
  NAND2_X1 U13687 ( .A1(n10920), .A2(n7009), .ZN(n11010) );
  INV_X1 U13688 ( .A(n10920), .ZN(n10921) );
  INV_X1 U13689 ( .A(n7009), .ZN(n11039) );
  NAND2_X1 U13690 ( .A1(n10921), .A2(n11039), .ZN(n10922) );
  AND2_X1 U13691 ( .A1(n11010), .A2(n10922), .ZN(n11032) );
  NAND2_X1 U13692 ( .A1(n10923), .A2(n11032), .ZN(n11009) );
  NAND2_X1 U13693 ( .A1(n11009), .A2(n11010), .ZN(n10928) );
  INV_X1 U13694 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11003) );
  MUX2_X1 U13695 ( .A(n7511), .B(n11003), .S(n13039), .Z(n10925) );
  NAND2_X1 U13696 ( .A1(n10925), .A2(n10924), .ZN(n10929) );
  INV_X1 U13697 ( .A(n10925), .ZN(n10926) );
  NAND2_X1 U13698 ( .A1(n10926), .A2(n11018), .ZN(n10927) );
  AND2_X1 U13699 ( .A1(n10929), .A2(n10927), .ZN(n11011) );
  MUX2_X1 U13700 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n7029), .Z(n10930) );
  XNOR2_X1 U13701 ( .A(n10930), .B(n10979), .ZN(n10992) );
  INV_X1 U13702 ( .A(n10930), .ZN(n10931) );
  NAND2_X1 U13703 ( .A1(n10931), .A2(n10979), .ZN(n10932) );
  MUX2_X1 U13704 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n7029), .Z(n10933) );
  NAND2_X1 U13705 ( .A1(n10933), .A2(n11089), .ZN(n11080) );
  NAND2_X1 U13706 ( .A1(n11083), .A2(n11080), .ZN(n10936) );
  INV_X1 U13707 ( .A(n10933), .ZN(n10935) );
  NAND2_X1 U13708 ( .A1(n10935), .A2(n10934), .ZN(n11081) );
  MUX2_X1 U13709 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n7029), .Z(n10937) );
  INV_X1 U13710 ( .A(n11130), .ZN(n10938) );
  XNOR2_X1 U13711 ( .A(n10937), .B(n10938), .ZN(n11120) );
  INV_X1 U13712 ( .A(n10937), .ZN(n10939) );
  MUX2_X1 U13713 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n7029), .Z(n11062) );
  XNOR2_X1 U13714 ( .A(n11062), .B(n11063), .ZN(n11060) );
  XNOR2_X1 U13715 ( .A(n11061), .B(n11060), .ZN(n10960) );
  AND2_X1 U13716 ( .A1(P3_U3897), .A2(n13513), .ZN(n13149) );
  INV_X1 U13717 ( .A(n10953), .ZN(n10940) );
  MUX2_X1 U13718 ( .A(n10940), .B(n12965), .S(n12954), .Z(n13147) );
  XNOR2_X1 U13719 ( .A(n10943), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n11021) );
  NOR2_X1 U13720 ( .A1(n11428), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10941) );
  OAI21_X1 U13721 ( .B1(n10978), .B2(n10941), .A(n10942), .ZN(n10971) );
  OR2_X1 U13722 ( .A1(n10971), .A2(n15607), .ZN(n10969) );
  NAND2_X1 U13723 ( .A1(n10969), .A2(n10942), .ZN(n11020) );
  NAND2_X1 U13724 ( .A1(n11021), .A2(n11020), .ZN(n11019) );
  OR2_X1 U13725 ( .A1(n10943), .A2(n15592), .ZN(n10944) );
  XNOR2_X1 U13726 ( .A(n10979), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n10983) );
  OR2_X1 U13727 ( .A1(n10979), .A2(n10945), .ZN(n10946) );
  XNOR2_X1 U13728 ( .A(n11130), .B(n11511), .ZN(n11124) );
  NAND2_X1 U13729 ( .A1(n11130), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10947) );
  OAI21_X1 U13730 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n10950), .A(n11073), .ZN(
        n10954) );
  INV_X1 U13731 ( .A(n10951), .ZN(n10952) );
  NAND2_X1 U13732 ( .A1(n10953), .A2(n10952), .ZN(n13151) );
  NAND2_X1 U13733 ( .A1(n10954), .A2(n13112), .ZN(n10958) );
  AND2_X1 U13734 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11836) );
  AOI21_X1 U13735 ( .B1(n15570), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11836), .ZN(
        n10957) );
  OAI211_X1 U13736 ( .C1(n13147), .C2(n11056), .A(n10958), .B(n10957), .ZN(
        n10959) );
  AOI21_X1 U13737 ( .B1(n10960), .B2(n13149), .A(n10959), .ZN(n10961) );
  OAI21_X1 U13738 ( .B1(n10962), .B2(n13143), .A(n10961), .ZN(P3_U3189) );
  OAI21_X1 U13739 ( .B1(n10964), .B2(n10963), .A(n11030), .ZN(n10976) );
  INV_X1 U13740 ( .A(n15570), .ZN(n13074) );
  OAI22_X1 U13741 ( .A1(n13074), .A2(n9097), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11050), .ZN(n10975) );
  INV_X1 U13742 ( .A(n10965), .ZN(n10966) );
  AOI21_X1 U13743 ( .B1(n10968), .B2(n10967), .A(n10966), .ZN(n10973) );
  INV_X1 U13744 ( .A(n10969), .ZN(n10970) );
  AOI21_X1 U13745 ( .B1(n15607), .B2(n10971), .A(n10970), .ZN(n10972) );
  OAI22_X1 U13746 ( .A1(n10973), .A2(n13143), .B1(n13151), .B2(n10972), .ZN(
        n10974) );
  AOI211_X1 U13747 ( .C1(n13149), .C2(n10976), .A(n10975), .B(n10974), .ZN(
        n10977) );
  OAI21_X1 U13748 ( .B1(n10978), .B2(n13147), .A(n10977), .ZN(P3_U3183) );
  INV_X1 U13749 ( .A(n10979), .ZN(n10997) );
  INV_X1 U13750 ( .A(n13143), .ZN(n13122) );
  OAI21_X1 U13751 ( .B1(n10982), .B2(n10981), .A(n10980), .ZN(n10990) );
  NAND2_X1 U13752 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11408) );
  OAI21_X1 U13753 ( .B1(n13074), .B2(n7599), .A(n11408), .ZN(n10989) );
  INV_X1 U13754 ( .A(n10983), .ZN(n10985) );
  NAND3_X1 U13755 ( .A1(n11001), .A2(n10985), .A3(n10984), .ZN(n10986) );
  AOI21_X1 U13756 ( .B1(n10987), .B2(n10986), .A(n13151), .ZN(n10988) );
  AOI211_X1 U13757 ( .C1(n13122), .C2(n10990), .A(n10989), .B(n10988), .ZN(
        n10996) );
  OAI21_X1 U13758 ( .B1(n10993), .B2(n10992), .A(n10991), .ZN(n10994) );
  NAND2_X1 U13759 ( .A1(n10994), .A2(n13149), .ZN(n10995) );
  OAI211_X1 U13760 ( .C1(n13147), .C2(n10997), .A(n10996), .B(n10995), .ZN(
        P3_U3186) );
  NOR2_X1 U13761 ( .A1(n12747), .A2(P3_U3151), .ZN(n11101) );
  NAND2_X1 U13762 ( .A1(n15596), .A2(n11423), .ZN(n12803) );
  NAND2_X1 U13763 ( .A1(n15598), .A2(n12803), .ZN(n12769) );
  OAI22_X1 U13764 ( .A1(n12744), .A2(n11423), .B1(n12743), .B2(n15583), .ZN(
        n10999) );
  AOI21_X1 U13765 ( .B1(n12730), .B2(n12769), .A(n10999), .ZN(n11000) );
  OAI21_X1 U13766 ( .B1(n11101), .B2(n11424), .A(n11000), .ZN(P3_U3172) );
  OAI21_X1 U13767 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n11002), .A(n11001), .ZN(
        n11008) );
  XNOR2_X1 U13768 ( .A(n11004), .B(n11003), .ZN(n11006) );
  AOI22_X1 U13769 ( .A1(n15570), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n11005) );
  OAI21_X1 U13770 ( .B1(n11006), .B2(n13143), .A(n11005), .ZN(n11007) );
  AOI21_X1 U13771 ( .B1(n13112), .B2(n11008), .A(n11007), .ZN(n11017) );
  INV_X1 U13772 ( .A(n11009), .ZN(n11035) );
  INV_X1 U13773 ( .A(n11010), .ZN(n11012) );
  NOR3_X1 U13774 ( .A1(n11035), .A2(n11012), .A3(n11011), .ZN(n11015) );
  INV_X1 U13775 ( .A(n11013), .ZN(n11014) );
  OAI21_X1 U13776 ( .B1(n11015), .B2(n11014), .A(n13149), .ZN(n11016) );
  OAI211_X1 U13777 ( .C1(n13147), .C2(n11018), .A(n11017), .B(n11016), .ZN(
        P3_U3185) );
  OAI21_X1 U13778 ( .B1(n11021), .B2(n11020), .A(n11019), .ZN(n11029) );
  INV_X1 U13779 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15576) );
  OAI22_X1 U13780 ( .A1(n13074), .A2(n11022), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15576), .ZN(n11028) );
  OAI21_X1 U13781 ( .B1(n11025), .B2(n11024), .A(n11023), .ZN(n11026) );
  AND2_X1 U13782 ( .A1(n13122), .A2(n11026), .ZN(n11027) );
  AOI211_X1 U13783 ( .C1(n13112), .C2(n11029), .A(n11028), .B(n11027), .ZN(
        n11038) );
  INV_X1 U13784 ( .A(n11030), .ZN(n11034) );
  INV_X1 U13785 ( .A(n11031), .ZN(n11033) );
  NOR3_X1 U13786 ( .A1(n11034), .A2(n11033), .A3(n11032), .ZN(n11036) );
  OAI21_X1 U13787 ( .B1(n11036), .B2(n11035), .A(n13149), .ZN(n11037) );
  OAI211_X1 U13788 ( .C1(n13147), .C2(n11039), .A(n11038), .B(n11037), .ZN(
        P3_U3184) );
  NAND3_X1 U13789 ( .A1(n15598), .A2(n11040), .A3(n12496), .ZN(n11042) );
  OAI211_X1 U13790 ( .C1(n6623), .C2(n15594), .A(n11043), .B(n11042), .ZN(
        n11044) );
  NAND2_X1 U13791 ( .A1(n11044), .A2(n12730), .ZN(n11049) );
  INV_X1 U13792 ( .A(n15596), .ZN(n11045) );
  OAI22_X1 U13793 ( .A1(n11494), .A2(n12743), .B1(n12733), .B2(n11045), .ZN(
        n11046) );
  AOI21_X1 U13794 ( .B1(n11047), .B2(n12720), .A(n11046), .ZN(n11048) );
  OAI211_X1 U13795 ( .C1(n11101), .C2(n11050), .A(n11049), .B(n11048), .ZN(
        P3_U3162) );
  INV_X1 U13796 ( .A(n13131), .ZN(n13138) );
  INV_X1 U13797 ( .A(n11051), .ZN(n11053) );
  OAI222_X1 U13798 ( .A1(n13138), .A2(P3_U3151), .B1(n13520), .B2(n11053), 
        .C1(n11052), .C2(n13522), .ZN(P3_U3277) );
  XNOR2_X1 U13799 ( .A(n11225), .B(P3_REG1_REG_8__SCAN_IN), .ZN(n11212) );
  NAND2_X1 U13800 ( .A1(n11055), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n11059) );
  NAND2_X1 U13801 ( .A1(n11057), .A2(n11056), .ZN(n11058) );
  XOR2_X1 U13802 ( .A(n11212), .B(n11213), .Z(n11079) );
  INV_X1 U13803 ( .A(n11062), .ZN(n11064) );
  NAND2_X1 U13804 ( .A1(n11064), .A2(n11063), .ZN(n11065) );
  NAND2_X1 U13805 ( .A1(n11066), .A2(n11065), .ZN(n11223) );
  MUX2_X1 U13806 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n7029), .Z(n11224) );
  XNOR2_X1 U13807 ( .A(n11224), .B(n11225), .ZN(n11222) );
  XNOR2_X1 U13808 ( .A(n11223), .B(n11222), .ZN(n11077) );
  AND2_X1 U13809 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n12141) );
  AOI21_X1 U13810 ( .B1(n15570), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12141), .ZN(
        n11067) );
  OAI21_X1 U13811 ( .B1(n13147), .B2(n11068), .A(n11067), .ZN(n11076) );
  XNOR2_X1 U13812 ( .A(n11225), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n11070) );
  INV_X1 U13813 ( .A(n11070), .ZN(n11072) );
  NAND3_X1 U13814 ( .A1(n11073), .A2(n11072), .A3(n11071), .ZN(n11074) );
  AOI21_X1 U13815 ( .B1(n11216), .B2(n11074), .A(n13151), .ZN(n11075) );
  AOI211_X1 U13816 ( .C1(n11077), .C2(n13149), .A(n11076), .B(n11075), .ZN(
        n11078) );
  OAI21_X1 U13817 ( .B1(n11079), .B2(n13143), .A(n11078), .ZN(P3_U3190) );
  INV_X1 U13818 ( .A(n13149), .ZN(n13125) );
  NAND2_X1 U13819 ( .A1(n11081), .A2(n11080), .ZN(n11082) );
  XNOR2_X1 U13820 ( .A(n11083), .B(n11082), .ZN(n11093) );
  XNOR2_X1 U13821 ( .A(n11084), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n11091) );
  OAI21_X1 U13822 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11085), .A(n11126), .ZN(
        n11086) );
  NAND2_X1 U13823 ( .A1(n13112), .A2(n11086), .ZN(n11088) );
  AND2_X1 U13824 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11565) );
  AOI21_X1 U13825 ( .B1(n15570), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11565), .ZN(
        n11087) );
  OAI211_X1 U13826 ( .C1(n13147), .C2(n11089), .A(n11088), .B(n11087), .ZN(
        n11090) );
  AOI21_X1 U13827 ( .B1(n13122), .B2(n11091), .A(n11090), .ZN(n11092) );
  OAI21_X1 U13828 ( .B1(n13125), .B2(n11093), .A(n11092), .ZN(P3_U3187) );
  OAI21_X1 U13829 ( .B1(n11096), .B2(n11095), .A(n11094), .ZN(n11097) );
  NAND2_X1 U13830 ( .A1(n11097), .A2(n12730), .ZN(n11100) );
  OAI22_X1 U13831 ( .A1(n15583), .A2(n12733), .B1(n12743), .B2(n15581), .ZN(
        n11098) );
  AOI21_X1 U13832 ( .B1(n15573), .B2(n12720), .A(n11098), .ZN(n11099) );
  OAI211_X1 U13833 ( .C1(n11101), .C2(n15576), .A(n11100), .B(n11099), .ZN(
        P3_U3177) );
  MUX2_X1 U13834 ( .A(n9357), .B(P1_REG1_REG_11__SCAN_IN), .S(n11289), .Z(
        n11108) );
  OR2_X1 U13835 ( .A1(n11102), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11103) );
  MUX2_X1 U13836 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9341), .S(n14739), .Z(
        n14737) );
  NAND2_X1 U13837 ( .A1(n14739), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U13838 ( .A1(n14736), .A2(n11105), .ZN(n11107) );
  INV_X1 U13839 ( .A(n11291), .ZN(n11106) );
  AOI21_X1 U13840 ( .B1(n11108), .B2(n11107), .A(n11106), .ZN(n11118) );
  NOR2_X1 U13841 ( .A1(n11109), .A2(n12221), .ZN(n14730) );
  MUX2_X1 U13842 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n15050), .S(n14739), .Z(
        n14729) );
  NAND2_X1 U13843 ( .A1(n14739), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11111) );
  MUX2_X1 U13844 ( .A(n11939), .B(P1_REG2_REG_11__SCAN_IN), .S(n11289), .Z(
        n11110) );
  NAND3_X1 U13845 ( .A1(n14733), .A2(n11111), .A3(n11110), .ZN(n11112) );
  NAND3_X1 U13846 ( .A1(n6625), .A2(n14785), .A3(n11112), .ZN(n11117) );
  NAND2_X1 U13847 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(n6428), .ZN(n14344) );
  INV_X1 U13848 ( .A(n14344), .ZN(n11115) );
  NOR2_X1 U13849 ( .A1(n15315), .A2(n11113), .ZN(n11114) );
  AOI211_X1 U13850 ( .C1(n15299), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n11115), 
        .B(n11114), .ZN(n11116) );
  OAI211_X1 U13851 ( .C1(n11118), .C2(n6633), .A(n11117), .B(n11116), .ZN(
        P1_U3254) );
  XOR2_X1 U13852 ( .A(n11119), .B(n11120), .Z(n11135) );
  OAI21_X1 U13853 ( .B1(n11123), .B2(n11122), .A(n11121), .ZN(n11133) );
  NAND3_X1 U13854 ( .A1(n11126), .A2(n7519), .A3(n11125), .ZN(n11127) );
  AOI21_X1 U13855 ( .B1(n11128), .B2(n11127), .A(n13151), .ZN(n11132) );
  AND2_X1 U13856 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n12719) );
  AOI21_X1 U13857 ( .B1(n15570), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n12719), .ZN(
        n11129) );
  OAI21_X1 U13858 ( .B1(n13147), .B2(n11130), .A(n11129), .ZN(n11131) );
  AOI211_X1 U13859 ( .C1(n13122), .C2(n11133), .A(n11132), .B(n11131), .ZN(
        n11134) );
  OAI21_X1 U13860 ( .B1(n11135), .B2(n13125), .A(n11134), .ZN(P3_U3188) );
  NAND2_X1 U13861 ( .A1(n11136), .A2(n12730), .ZN(n11143) );
  AOI21_X1 U13862 ( .B1(n11094), .B2(n11138), .A(n11137), .ZN(n11142) );
  OAI22_X1 U13863 ( .A1(n11494), .A2(n12733), .B1(n12743), .B2(n11784), .ZN(
        n11140) );
  MUX2_X1 U13864 ( .A(n12747), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n11139) );
  AOI211_X1 U13865 ( .C1(n11498), .C2(n12720), .A(n11140), .B(n11139), .ZN(
        n11141) );
  OAI21_X1 U13866 ( .B1(n11143), .B2(n11142), .A(n11141), .ZN(P3_U3158) );
  XNOR2_X1 U13867 ( .A(n11145), .B(n11144), .ZN(n11151) );
  INV_X1 U13868 ( .A(n11146), .ZN(n12044) );
  NAND2_X1 U13869 ( .A1(n13669), .A2(n13966), .ZN(n11147) );
  OAI21_X1 U13870 ( .B1(n11475), .B2(n13932), .A(n11147), .ZN(n12050) );
  AOI22_X1 U13871 ( .A1(n13643), .A2(n12050), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11148) );
  OAI21_X1 U13872 ( .B1(n13620), .B2(n12046), .A(n11148), .ZN(n11149) );
  AOI21_X1 U13873 ( .B1(n12044), .B2(n13631), .A(n11149), .ZN(n11150) );
  OAI21_X1 U13874 ( .B1(n11151), .B2(n13649), .A(n11150), .ZN(P2_U3211) );
  INV_X1 U13875 ( .A(n15330), .ZN(n15348) );
  OAI21_X1 U13876 ( .B1(n11154), .B2(n11152), .A(n11153), .ZN(n11155) );
  NAND2_X1 U13877 ( .A1(n11155), .A2(n14370), .ZN(n11157) );
  INV_X1 U13878 ( .A(n11380), .ZN(n11275) );
  INV_X1 U13879 ( .A(n14652), .ZN(n14398) );
  OAI22_X1 U13880 ( .A1(n11275), .A2(n14976), .B1(n14398), .B2(n15052), .ZN(
        n15328) );
  AOI22_X1 U13881 ( .A1(n15328), .A2(n14368), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n14234), .ZN(n11156) );
  OAI211_X1 U13882 ( .C1(n15348), .C2(n14380), .A(n11157), .B(n11156), .ZN(
        P1_U3237) );
  NOR2_X1 U13883 ( .A1(n11158), .A2(n15623), .ZN(n11159) );
  NAND2_X1 U13884 ( .A1(n12769), .A2(n11159), .ZN(n11161) );
  NAND2_X1 U13885 ( .A1(n9757), .A2(n15597), .ZN(n11160) );
  NAND2_X1 U13886 ( .A1(n11161), .A2(n11160), .ZN(n11419) );
  NOR2_X1 U13887 ( .A1(n15652), .A2(n10918), .ZN(n11162) );
  AOI21_X1 U13888 ( .B1(n15652), .B2(n11419), .A(n11162), .ZN(n11163) );
  OAI21_X1 U13889 ( .B1(n11423), .B2(n13382), .A(n11163), .ZN(P3_U3459) );
  XNOR2_X1 U13890 ( .A(n11465), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n11166) );
  INV_X1 U13891 ( .A(n15471), .ZN(n15513) );
  AOI211_X1 U13892 ( .C1(n11166), .C2(n11165), .A(n15513), .B(n11464), .ZN(
        n11178) );
  MUX2_X1 U13893 ( .A(n11167), .B(P2_REG2_REG_10__SCAN_IN), .S(n11465), .Z(
        n11173) );
  OR2_X1 U13894 ( .A1(n11168), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n11169) );
  NAND2_X1 U13895 ( .A1(n11170), .A2(n11169), .ZN(n11172) );
  INV_X1 U13896 ( .A(n11460), .ZN(n11171) );
  AOI211_X1 U13897 ( .C1(n11173), .C2(n11172), .A(n15421), .B(n11171), .ZN(
        n11177) );
  NAND2_X1 U13898 ( .A1(n15519), .A2(n11465), .ZN(n11175) );
  NAND2_X1 U13899 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11174)
         );
  OAI211_X1 U13900 ( .C1(n15215), .C2(n15522), .A(n11175), .B(n11174), .ZN(
        n11176) );
  OR3_X1 U13901 ( .A1(n11178), .A2(n11177), .A3(n11176), .ZN(P2_U3224) );
  XNOR2_X1 U13902 ( .A(n11180), .B(n11179), .ZN(n11186) );
  INV_X1 U13903 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11184) );
  OAI22_X1 U13904 ( .A1(n13620), .A2(n12056), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11184), .ZN(n11183) );
  OAI22_X1 U13905 ( .A1(n13634), .A2(n11181), .B1(n11251), .B2(n13623), .ZN(
        n11182) );
  AOI211_X1 U13906 ( .C1(n13631), .C2(n11184), .A(n11183), .B(n11182), .ZN(
        n11185) );
  OAI21_X1 U13907 ( .B1(n11186), .B2(n13649), .A(n11185), .ZN(P2_U3190) );
  OAI21_X1 U13908 ( .B1(n11189), .B2(n11188), .A(n11187), .ZN(n11193) );
  OAI22_X1 U13909 ( .A1(n11190), .A2(n12121), .B1(n13623), .B2(n12120), .ZN(
        n11192) );
  OAI22_X1 U13910 ( .A1(n13634), .A2(n12119), .B1(n15537), .B2(n13620), .ZN(
        n11191) );
  AOI211_X1 U13911 ( .C1(n13610), .C2(n11193), .A(n11192), .B(n11191), .ZN(
        n11194) );
  INV_X1 U13912 ( .A(n11194), .ZN(P2_U3209) );
  INV_X1 U13913 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11195) );
  NOR2_X1 U13914 ( .A1(n15645), .A2(n11195), .ZN(n11196) );
  AOI21_X1 U13915 ( .B1(n15645), .B2(n11419), .A(n11196), .ZN(n11197) );
  OAI21_X1 U13916 ( .B1(n11423), .B2(n13443), .A(n11197), .ZN(P3_U3390) );
  INV_X1 U13917 ( .A(n11198), .ZN(n11200) );
  INV_X1 U13918 ( .A(n12347), .ZN(n12342) );
  OAI222_X1 U13919 ( .A1(n15174), .A2(n11199), .B1(n15188), .B2(n11200), .C1(
        n12342), .C2(n6428), .ZN(P1_U3341) );
  INV_X1 U13920 ( .A(n12474), .ZN(n12395) );
  OAI222_X1 U13921 ( .A1(n14184), .A2(n11201), .B1(n6438), .B2(n11200), .C1(
        n12395), .C2(P2_U3088), .ZN(P2_U3313) );
  OAI21_X1 U13922 ( .B1(n11204), .B2(n11203), .A(n11202), .ZN(n11209) );
  INV_X1 U13923 ( .A(n13623), .ZN(n13630) );
  AOI22_X1 U13924 ( .A1(n13630), .A2(n13670), .B1(n13568), .B2(n13668), .ZN(
        n11207) );
  NAND2_X1 U13925 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n15467) );
  INV_X1 U13926 ( .A(n15467), .ZN(n11205) );
  AOI21_X1 U13927 ( .B1(n13647), .B2(n12038), .A(n11205), .ZN(n11206) );
  OAI211_X1 U13928 ( .C1(n12020), .C2(n13645), .A(n11207), .B(n11206), .ZN(
        n11208) );
  AOI21_X1 U13929 ( .B1(n11209), .B2(n13610), .A(n11208), .ZN(n11210) );
  INV_X1 U13930 ( .A(n11210), .ZN(P2_U3199) );
  NOR2_X1 U13931 ( .A1(n11225), .A2(n12080), .ZN(n11211) );
  INV_X1 U13932 ( .A(n11229), .ZN(n11654) );
  XNOR2_X1 U13933 ( .A(n11655), .B(P3_REG1_REG_9__SCAN_IN), .ZN(n11239) );
  OR2_X1 U13934 ( .A1(n11225), .A2(n11214), .ZN(n11215) );
  OAI21_X1 U13935 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11217), .A(n11670), .ZN(
        n11221) );
  NAND2_X1 U13936 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11858) );
  INV_X1 U13937 ( .A(n11858), .ZN(n11218) );
  AOI21_X1 U13938 ( .B1(n15570), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11218), .ZN(
        n11219) );
  OAI21_X1 U13939 ( .B1(n13147), .B2(n11229), .A(n11219), .ZN(n11220) );
  AOI21_X1 U13940 ( .B1(n11221), .B2(n13112), .A(n11220), .ZN(n11238) );
  NAND2_X1 U13941 ( .A1(n11223), .A2(n11222), .ZN(n11228) );
  INV_X1 U13942 ( .A(n11224), .ZN(n11226) );
  NAND2_X1 U13943 ( .A1(n11226), .A2(n11225), .ZN(n11227) );
  NAND2_X1 U13944 ( .A1(n11228), .A2(n11227), .ZN(n11233) );
  MUX2_X1 U13945 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n7029), .Z(n11230) );
  NAND2_X1 U13946 ( .A1(n11230), .A2(n11229), .ZN(n11234) );
  INV_X1 U13947 ( .A(n11230), .ZN(n11231) );
  NAND2_X1 U13948 ( .A1(n11231), .A2(n11654), .ZN(n11664) );
  INV_X1 U13949 ( .A(n11664), .ZN(n11232) );
  NOR2_X1 U13950 ( .A1(n11665), .A2(n11232), .ZN(n11236) );
  AOI21_X1 U13951 ( .B1(n11664), .B2(n11234), .A(n11233), .ZN(n11235) );
  OAI21_X1 U13952 ( .B1(n11236), .B2(n11235), .A(n13149), .ZN(n11237) );
  OAI211_X1 U13953 ( .C1(n11239), .C2(n13143), .A(n11238), .B(n11237), .ZN(
        P3_U3191) );
  NAND2_X1 U13954 ( .A1(n11352), .A2(n11240), .ZN(n12129) );
  INV_X1 U13955 ( .A(n11241), .ZN(n12128) );
  NAND2_X1 U13956 ( .A1(n12129), .A2(n12128), .ZN(n12127) );
  INV_X1 U13957 ( .A(n11249), .ZN(n11245) );
  NAND3_X1 U13958 ( .A1(n12127), .A2(n11242), .A3(n11245), .ZN(n11244) );
  AND2_X1 U13959 ( .A1(n11243), .A2(n11244), .ZN(n12061) );
  NAND2_X1 U13960 ( .A1(n11246), .A2(n11245), .ZN(n11329) );
  NAND3_X1 U13961 ( .A1(n11247), .A2(n11249), .A3(n11248), .ZN(n11250) );
  NAND2_X1 U13962 ( .A1(n11329), .A2(n11250), .ZN(n11252) );
  AOI222_X1 U13963 ( .A1(n13971), .A2(n11252), .B1(n13670), .B2(n13968), .C1(
        n8790), .C2(n13966), .ZN(n12055) );
  NAND2_X1 U13964 ( .A1(n12122), .A2(n8571), .ZN(n11253) );
  NAND2_X1 U13965 ( .A1(n11253), .A2(n12569), .ZN(n11254) );
  NOR2_X1 U13966 ( .A1(n11335), .A2(n11254), .ZN(n12058) );
  INV_X1 U13967 ( .A(n12058), .ZN(n11255) );
  OAI211_X1 U13968 ( .C1(n15557), .C2(n12061), .A(n12055), .B(n11255), .ZN(
        n11398) );
  NAND2_X1 U13969 ( .A1(n15564), .A2(n15553), .ZN(n14104) );
  OAI22_X1 U13970 ( .A1(n14104), .A2(n12056), .B1(n15564), .B2(n11256), .ZN(
        n11257) );
  AOI21_X1 U13971 ( .B1(n11398), .B2(n15564), .A(n11257), .ZN(n11258) );
  INV_X1 U13972 ( .A(n11258), .ZN(P2_U3502) );
  NAND2_X1 U13973 ( .A1(n11259), .A2(n11260), .ZN(n11372) );
  OR2_X1 U13974 ( .A1(n11259), .A2(n11260), .ZN(n11261) );
  NAND2_X1 U13975 ( .A1(n11372), .A2(n11261), .ZN(n15346) );
  INV_X1 U13976 ( .A(n15346), .ZN(n11282) );
  NAND3_X1 U13977 ( .A1(n14577), .A2(n11263), .A3(n11262), .ZN(n12506) );
  INV_X1 U13978 ( .A(n11264), .ZN(n11265) );
  OR2_X1 U13979 ( .A1(n14387), .A2(n14958), .ZN(n14538) );
  INV_X1 U13980 ( .A(n14538), .ZN(n11267) );
  NAND2_X1 U13981 ( .A1(n15049), .A2(n11267), .ZN(n15231) );
  OR2_X1 U13982 ( .A1(n9219), .A2(n11709), .ZN(n14614) );
  OR2_X1 U13983 ( .A1(n14614), .A2(n15190), .ZN(n11268) );
  NOR2_X2 U13984 ( .A1(n15340), .A2(n11268), .ZN(n15329) );
  NOR2_X1 U13985 ( .A1(n15049), .A2(n14655), .ZN(n11273) );
  INV_X1 U13986 ( .A(n15235), .ZN(n14860) );
  OR2_X1 U13987 ( .A1(n15343), .A2(n11378), .ZN(n11269) );
  NAND2_X1 U13988 ( .A1(n11269), .A2(n15332), .ZN(n11274) );
  INV_X1 U13989 ( .A(n11274), .ZN(n11270) );
  NAND2_X1 U13990 ( .A1(n11270), .A2(n15333), .ZN(n15342) );
  OAI22_X1 U13991 ( .A1(n14860), .A2(n15342), .B1(n11271), .B2(n15055), .ZN(
        n11272) );
  AOI211_X1 U13992 ( .C1(n15329), .C2(n11370), .A(n11273), .B(n11272), .ZN(
        n11281) );
  XNOR2_X1 U13993 ( .A(n11275), .B(n11274), .ZN(n11276) );
  INV_X1 U13994 ( .A(n11259), .ZN(n14583) );
  MUX2_X1 U13995 ( .A(n11276), .B(n14583), .S(n11377), .Z(n11279) );
  AOI22_X1 U13996 ( .A1(n15223), .A2(n11377), .B1(n11381), .B2(n15222), .ZN(
        n11278) );
  INV_X1 U13997 ( .A(n15375), .ZN(n15361) );
  NAND2_X1 U13998 ( .A1(n15346), .A2(n15361), .ZN(n11277) );
  OAI211_X1 U13999 ( .C1(n11279), .C2(n15325), .A(n11278), .B(n11277), .ZN(
        n15344) );
  NAND2_X1 U14000 ( .A1(n15344), .A2(n15049), .ZN(n11280) );
  OAI211_X1 U14001 ( .C1(n11282), .C2(n15231), .A(n11281), .B(n11280), .ZN(
        P1_U3292) );
  MUX2_X1 U14002 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9370), .S(n11441), .Z(
        n11283) );
  OAI21_X1 U14003 ( .B1(n11283), .B2(n6624), .A(n11436), .ZN(n11287) );
  NAND2_X1 U14004 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14254)
         );
  NAND2_X1 U14005 ( .A1(n15299), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n11284) );
  OAI211_X1 U14006 ( .C1(n15315), .C2(n11285), .A(n14254), .B(n11284), .ZN(
        n11286) );
  AOI21_X1 U14007 ( .B1(n11287), .B2(n14785), .A(n11286), .ZN(n11296) );
  MUX2_X1 U14008 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n11288), .S(n11441), .Z(
        n11293) );
  OR2_X1 U14009 ( .A1(n11289), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11290) );
  OAI21_X1 U14010 ( .B1(n11293), .B2(n11292), .A(n11443), .ZN(n11294) );
  NAND2_X1 U14011 ( .A1(n11294), .A2(n15310), .ZN(n11295) );
  NAND2_X1 U14012 ( .A1(n11296), .A2(n11295), .ZN(P1_U3255) );
  INV_X1 U14013 ( .A(n11297), .ZN(n11300) );
  OAI222_X1 U14014 ( .A1(n15174), .A2(n11298), .B1(n15188), .B2(n11300), .C1(
        n12352), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U14015 ( .A(n15504), .ZN(n11299) );
  OAI222_X1 U14016 ( .A1(n14184), .A2(n11301), .B1(n6438), .B2(n11300), .C1(
        n11299), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U14017 ( .A(n11302), .ZN(n11304) );
  INV_X1 U14018 ( .A(n12350), .ZN(n15314) );
  OAI222_X1 U14019 ( .A1(n15174), .A2(n11303), .B1(n15188), .B2(n11304), .C1(
        n15314), .C2(n6428), .ZN(P1_U3340) );
  INV_X1 U14020 ( .A(n13685), .ZN(n12398) );
  OAI222_X1 U14021 ( .A1(n14184), .A2(n11305), .B1(n6438), .B2(n11304), .C1(
        n12398), .C2(P2_U3088), .ZN(P2_U3312) );
  XNOR2_X1 U14022 ( .A(n6949), .B(n11309), .ZN(n11306) );
  INV_X1 U14023 ( .A(n11306), .ZN(n12025) );
  NAND2_X1 U14024 ( .A1(n11306), .A2(n15550), .ZN(n11316) );
  NAND2_X1 U14025 ( .A1(n11329), .A2(n11327), .ZN(n11308) );
  NAND2_X1 U14026 ( .A1(n11308), .A2(n11307), .ZN(n11331) );
  OAI211_X1 U14027 ( .C1(n12029), .C2(n13670), .A(n11331), .B(n11309), .ZN(
        n11310) );
  NAND2_X1 U14028 ( .A1(n11310), .A2(n7833), .ZN(n11314) );
  NAND2_X1 U14029 ( .A1(n13670), .A2(n13966), .ZN(n11311) );
  OAI21_X1 U14030 ( .B1(n11312), .B2(n13932), .A(n11311), .ZN(n11313) );
  AOI21_X1 U14031 ( .B1(n11314), .B2(n13971), .A(n11313), .ZN(n11315) );
  AND2_X1 U14032 ( .A1(n11316), .A2(n11315), .ZN(n12019) );
  AOI211_X1 U14033 ( .C1(n12038), .C2(n11336), .A(n13974), .B(n6435), .ZN(
        n12022) );
  INV_X1 U14034 ( .A(n12022), .ZN(n11317) );
  OAI211_X1 U14035 ( .C1(n12025), .C2(n15546), .A(n12019), .B(n11317), .ZN(
        n11402) );
  OAI22_X1 U14036 ( .A1(n14104), .A2(n11318), .B1(n15564), .B2(n11319), .ZN(
        n11320) );
  AOI21_X1 U14037 ( .B1(n11402), .B2(n15564), .A(n11320), .ZN(n11321) );
  INV_X1 U14038 ( .A(n11321), .ZN(P2_U3504) );
  OR2_X1 U14039 ( .A1(n11323), .A2(n11328), .ZN(n11324) );
  NAND2_X1 U14040 ( .A1(n11322), .A2(n11324), .ZN(n11326) );
  INV_X1 U14041 ( .A(n11326), .ZN(n12035) );
  AOI21_X1 U14042 ( .B1(n11326), .B2(n15550), .A(n11325), .ZN(n11334) );
  NAND3_X1 U14043 ( .A1(n11329), .A2(n11328), .A3(n11327), .ZN(n11330) );
  NAND2_X1 U14044 ( .A1(n11331), .A2(n11330), .ZN(n11332) );
  NAND2_X1 U14045 ( .A1(n11332), .A2(n13971), .ZN(n11333) );
  AND2_X1 U14046 ( .A1(n11334), .A2(n11333), .ZN(n12026) );
  INV_X1 U14047 ( .A(n11335), .ZN(n11337) );
  AOI211_X1 U14048 ( .C1(n6432), .C2(n11337), .A(n13974), .B(n6436), .ZN(
        n12031) );
  INV_X1 U14049 ( .A(n12031), .ZN(n11338) );
  OAI211_X1 U14050 ( .C1(n12035), .C2(n15546), .A(n12026), .B(n11338), .ZN(
        n11394) );
  OAI22_X1 U14051 ( .A1(n14104), .A2(n12029), .B1(n15564), .B2(n11339), .ZN(
        n11340) );
  AOI21_X1 U14052 ( .B1(n11394), .B2(n15564), .A(n11340), .ZN(n11341) );
  INV_X1 U14053 ( .A(n11341), .ZN(P2_U3503) );
  XNOR2_X1 U14054 ( .A(n11343), .B(n11342), .ZN(n11347) );
  AOI22_X1 U14055 ( .A1(n13966), .A2(n13668), .B1(n13665), .B2(n13968), .ZN(
        n11994) );
  OAI22_X1 U14056 ( .A1(n13616), .A2(n11994), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8020), .ZN(n11345) );
  NOR2_X1 U14057 ( .A1(n13645), .A2(n11998), .ZN(n11344) );
  AOI211_X1 U14058 ( .C1(n15552), .C2(n13647), .A(n11345), .B(n11344), .ZN(
        n11346) );
  OAI21_X1 U14059 ( .B1(n11347), .B2(n13649), .A(n11346), .ZN(P2_U3185) );
  INV_X1 U14060 ( .A(n11348), .ZN(n11349) );
  NAND2_X1 U14061 ( .A1(n11350), .A2(n11349), .ZN(n11351) );
  NAND2_X1 U14062 ( .A1(n11352), .A2(n11351), .ZN(n13992) );
  OAI21_X1 U14063 ( .B1(n8567), .B2(n11353), .A(n12569), .ZN(n11354) );
  NOR2_X1 U14064 ( .A1(n11354), .A2(n12123), .ZN(n13994) );
  NAND2_X1 U14065 ( .A1(n11356), .A2(n11355), .ZN(n11358) );
  AOI21_X1 U14066 ( .B1(n11358), .B2(n11357), .A(n13951), .ZN(n11359) );
  AOI211_X1 U14067 ( .C1(n15550), .C2(n13992), .A(n11360), .B(n11359), .ZN(
        n13988) );
  INV_X1 U14068 ( .A(n13988), .ZN(n11361) );
  AOI211_X1 U14069 ( .C1(n11362), .C2(n13992), .A(n13994), .B(n11361), .ZN(
        n11392) );
  NAND2_X1 U14070 ( .A1(n15561), .A2(n15553), .ZN(n14160) );
  OAI22_X1 U14071 ( .A1(n14160), .A2(n8567), .B1(n15561), .B2(n7881), .ZN(
        n11363) );
  INV_X1 U14072 ( .A(n11363), .ZN(n11364) );
  OAI21_X1 U14073 ( .B1(n11392), .B2(n15559), .A(n11364), .ZN(P2_U3433) );
  INV_X1 U14074 ( .A(n11365), .ZN(n11368) );
  OAI222_X1 U14075 ( .A1(n15174), .A2(n11366), .B1(n15188), .B2(n11368), .C1(
        n14762), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U14076 ( .A(n15518), .ZN(n11367) );
  OAI222_X1 U14077 ( .A1(n14184), .A2(n11369), .B1(n6438), .B2(n11368), .C1(
        n11367), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U14078 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n11388) );
  OR2_X1 U14079 ( .A1(n11380), .A2(n11370), .ZN(n11371) );
  NAND2_X1 U14080 ( .A1(n11372), .A2(n11371), .ZN(n15322) );
  NAND2_X1 U14081 ( .A1(n15322), .A2(n15323), .ZN(n15321) );
  OR2_X1 U14082 ( .A1(n11381), .A2(n15330), .ZN(n11373) );
  NAND2_X1 U14083 ( .A1(n11633), .A2(n7435), .ZN(n11480) );
  INV_X1 U14084 ( .A(n11480), .ZN(n11374) );
  AOI21_X1 U14085 ( .B1(n7059), .B2(n14584), .A(n11374), .ZN(n11536) );
  INV_X1 U14086 ( .A(n11375), .ZN(n15334) );
  AOI211_X1 U14087 ( .C1(n11629), .C2(n15334), .A(n15365), .B(n8851), .ZN(
        n11532) );
  INV_X1 U14088 ( .A(n11377), .ZN(n11379) );
  NAND2_X1 U14089 ( .A1(n11379), .A2(n11453), .ZN(n14385) );
  AND2_X1 U14090 ( .A1(n11380), .A2(n15343), .ZN(n14389) );
  INV_X1 U14091 ( .A(n11381), .ZN(n11382) );
  NAND2_X1 U14092 ( .A1(n11382), .A2(n15330), .ZN(n11383) );
  XNOR2_X1 U14093 ( .A(n11482), .B(n7435), .ZN(n11385) );
  OAI21_X1 U14094 ( .B1(n11385), .B2(n15325), .A(n11384), .ZN(n11533) );
  AOI211_X1 U14095 ( .C1(n15400), .C2(n11629), .A(n11532), .B(n11533), .ZN(
        n11386) );
  OAI21_X1 U14096 ( .B1(n15404), .B2(n11536), .A(n11386), .ZN(n11389) );
  NAND2_X1 U14097 ( .A1(n11389), .A2(n15420), .ZN(n11387) );
  OAI21_X1 U14098 ( .B1(n15420), .B2(n11388), .A(n11387), .ZN(P1_U3531) );
  NAND2_X1 U14099 ( .A1(n11389), .A2(n15408), .ZN(n11390) );
  OAI21_X1 U14100 ( .B1(n15408), .B2(n9266), .A(n11390), .ZN(P1_U3468) );
  INV_X1 U14101 ( .A(n14104), .ZN(n14096) );
  AOI22_X1 U14102 ( .A1(n14096), .A2(n6645), .B1(n15567), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n11391) );
  OAI21_X1 U14103 ( .B1(n11392), .B2(n15567), .A(n11391), .ZN(P2_U3500) );
  OAI22_X1 U14104 ( .A1(n14160), .A2(n12029), .B1(n15561), .B2(n7020), .ZN(
        n11393) );
  AOI21_X1 U14105 ( .B1(n11394), .B2(n15561), .A(n11393), .ZN(n11395) );
  INV_X1 U14106 ( .A(n11395), .ZN(P2_U3442) );
  INV_X1 U14107 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11396) );
  OAI22_X1 U14108 ( .A1(n14160), .A2(n12056), .B1(n15561), .B2(n11396), .ZN(
        n11397) );
  AOI21_X1 U14109 ( .B1(n11398), .B2(n15561), .A(n11397), .ZN(n11399) );
  INV_X1 U14110 ( .A(n11399), .ZN(P2_U3439) );
  INV_X1 U14111 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11400) );
  OAI22_X1 U14112 ( .A1(n14160), .A2(n11318), .B1(n15561), .B2(n11400), .ZN(
        n11401) );
  AOI21_X1 U14113 ( .B1(n11402), .B2(n15561), .A(n11401), .ZN(n11403) );
  INV_X1 U14114 ( .A(n11403), .ZN(P2_U3445) );
  INV_X1 U14115 ( .A(n11404), .ZN(n11405) );
  AOI21_X1 U14116 ( .B1(n11407), .B2(n11406), .A(n11405), .ZN(n11413) );
  INV_X1 U14117 ( .A(n11731), .ZN(n11411) );
  AOI22_X1 U14118 ( .A1(n12735), .A2(n12977), .B1(n15624), .B2(n12720), .ZN(
        n11409) );
  OAI211_X1 U14119 ( .C1(n15581), .C2(n12733), .A(n11409), .B(n11408), .ZN(
        n11410) );
  AOI21_X1 U14120 ( .B1(n11411), .B2(n12747), .A(n11410), .ZN(n11412) );
  OAI21_X1 U14121 ( .B1(n11413), .B2(n12749), .A(n11412), .ZN(P3_U3170) );
  NAND2_X1 U14122 ( .A1(n11414), .A2(n11417), .ZN(n11415) );
  OAI211_X1 U14123 ( .C1(n11418), .C2(n11417), .A(n11416), .B(n11415), .ZN(
        n11420) );
  INV_X1 U14124 ( .A(n15603), .ZN(n15575) );
  OR2_X1 U14125 ( .A1(n11420), .A2(n15575), .ZN(n11776) );
  AOI21_X1 U14126 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15604), .A(n11419), .ZN(
        n11421) );
  AND2_X2 U14127 ( .A1(n11420), .A2(n15577), .ZN(n15610) );
  INV_X2 U14128 ( .A(n15610), .ZN(n15608) );
  MUX2_X1 U14129 ( .A(n11428), .B(n11421), .S(n15608), .Z(n11422) );
  OAI21_X1 U14130 ( .B1(n13340), .B2(n11423), .A(n11422), .ZN(P3_U3233) );
  OAI22_X1 U14131 ( .A1(n13074), .A2(n11425), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11424), .ZN(n11433) );
  NOR3_X1 U14132 ( .A1(n13112), .A2(n13122), .A3(n13149), .ZN(n11427) );
  OAI21_X1 U14133 ( .B1(n11427), .B2(n11426), .A(n13147), .ZN(n11431) );
  MUX2_X1 U14134 ( .A(n11431), .B(n11430), .S(n11429), .Z(n11432) );
  AOI211_X1 U14135 ( .C1(n13122), .C2(n11434), .A(n11433), .B(n11432), .ZN(
        n11435) );
  INV_X1 U14136 ( .A(n11435), .ZN(P3_U3182) );
  NAND2_X1 U14137 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14323)
         );
  OAI21_X1 U14138 ( .B1(n15319), .B2(n9121), .A(n14323), .ZN(n11440) );
  OAI21_X1 U14139 ( .B1(n11441), .B2(P1_REG2_REG_12__SCAN_IN), .A(n11436), 
        .ZN(n11438) );
  MUX2_X1 U14140 ( .A(n15034), .B(P1_REG2_REG_13__SCAN_IN), .S(n11711), .Z(
        n11437) );
  AOI211_X1 U14141 ( .C1(n11438), .C2(n11437), .A(n15305), .B(n11724), .ZN(
        n11439) );
  AOI211_X1 U14142 ( .C1(n14783), .C2(n11711), .A(n11440), .B(n11439), .ZN(
        n11447) );
  OR2_X1 U14143 ( .A1(n11441), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11442) );
  INV_X1 U14144 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n15256) );
  MUX2_X1 U14145 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15256), .S(n11711), .Z(
        n11444) );
  OAI211_X1 U14146 ( .C1(n11445), .C2(n11444), .A(n11713), .B(n15310), .ZN(
        n11446) );
  NAND2_X1 U14147 ( .A1(n11447), .A2(n11446), .ZN(P1_U3256) );
  NOR2_X1 U14148 ( .A1(n15340), .A2(n11448), .ZN(n14865) );
  OAI22_X1 U14149 ( .A1(n15049), .A2(n11450), .B1(n11449), .B2(n15055), .ZN(
        n11451) );
  AOI21_X1 U14150 ( .B1(n15049), .B2(n11452), .A(n11451), .ZN(n11455) );
  AND2_X1 U14151 ( .A1(n15235), .A2(n15333), .ZN(n14950) );
  OAI21_X1 U14152 ( .B1(n15329), .B2(n14950), .A(n11453), .ZN(n11454) );
  OAI211_X1 U14153 ( .C1(n15062), .C2(n14581), .A(n11455), .B(n11454), .ZN(
        P1_U3293) );
  INV_X1 U14154 ( .A(n11456), .ZN(n11458) );
  OAI22_X1 U14155 ( .A1(n12957), .A2(P3_U3151), .B1(SI_22_), .B2(n13522), .ZN(
        n11457) );
  AOI21_X1 U14156 ( .B1(n11458), .B2(n13500), .A(n11457), .ZN(P3_U3273) );
  XNOR2_X1 U14157 ( .A(n11568), .B(n12173), .ZN(n11463) );
  NAND2_X1 U14158 ( .A1(n11465), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11459) );
  NAND2_X1 U14159 ( .A1(n11460), .A2(n11459), .ZN(n11462) );
  INV_X1 U14160 ( .A(n11570), .ZN(n11461) );
  AOI21_X1 U14161 ( .B1(n11463), .B2(n11462), .A(n11461), .ZN(n11471) );
  NAND2_X1 U14162 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11900)
         );
  OAI21_X1 U14163 ( .B1(n15522), .B2(n15269), .A(n11900), .ZN(n11469) );
  XNOR2_X1 U14164 ( .A(n11573), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n11466) );
  AOI211_X1 U14165 ( .C1(n11467), .C2(n11466), .A(n15513), .B(n11572), .ZN(
        n11468) );
  AOI211_X1 U14166 ( .C1(n15519), .C2(n11573), .A(n11469), .B(n11468), .ZN(
        n11470) );
  OAI21_X1 U14167 ( .B1(n11471), .B2(n15421), .A(n11470), .ZN(P2_U3225) );
  XNOR2_X1 U14168 ( .A(n11694), .B(n11473), .ZN(n11474) );
  XNOR2_X1 U14169 ( .A(n11472), .B(n11474), .ZN(n11479) );
  OAI22_X1 U14170 ( .A1(n11754), .A2(n13932), .B1(n11475), .B2(n13930), .ZN(
        n12008) );
  AOI22_X1 U14171 ( .A1(n13643), .A2(n12008), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11476) );
  OAI21_X1 U14172 ( .B1(n13645), .B2(n12014), .A(n11476), .ZN(n11477) );
  AOI21_X1 U14173 ( .B1(n14111), .B2(n13647), .A(n11477), .ZN(n11478) );
  OAI21_X1 U14174 ( .B1(n11479), .B2(n13649), .A(n11478), .ZN(P2_U3193) );
  INV_X1 U14175 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n11489) );
  NAND2_X1 U14176 ( .A1(n11480), .A2(n11627), .ZN(n11583) );
  XNOR2_X1 U14177 ( .A(n14651), .B(n14404), .ZN(n14582) );
  XNOR2_X1 U14178 ( .A(n11583), .B(n14582), .ZN(n11558) );
  INV_X1 U14179 ( .A(n11587), .ZN(n11481) );
  AOI211_X1 U14180 ( .C1(n14404), .C2(n11376), .A(n15365), .B(n11481), .ZN(
        n11555) );
  OR2_X1 U14181 ( .A1(n14652), .A2(n14399), .ZN(n11483) );
  XOR2_X1 U14182 ( .A(n11589), .B(n14582), .Z(n11486) );
  NAND2_X1 U14183 ( .A1(n14652), .A2(n15223), .ZN(n11485) );
  NAND2_X1 U14184 ( .A1(n14650), .A2(n15222), .ZN(n11484) );
  AND2_X1 U14185 ( .A1(n11485), .A2(n11484), .ZN(n11520) );
  OAI21_X1 U14186 ( .B1(n11486), .B2(n15325), .A(n11520), .ZN(n11550) );
  AOI211_X1 U14187 ( .C1(n15400), .C2(n14404), .A(n11555), .B(n11550), .ZN(
        n11487) );
  OAI21_X1 U14188 ( .B1(n15404), .B2(n11558), .A(n11487), .ZN(n11490) );
  NAND2_X1 U14189 ( .A1(n11490), .A2(n15420), .ZN(n11488) );
  OAI21_X1 U14190 ( .B1(n15420), .B2(n11489), .A(n11488), .ZN(P1_U3532) );
  NAND2_X1 U14191 ( .A1(n11490), .A2(n15408), .ZN(n11491) );
  OAI21_X1 U14192 ( .B1(n15408), .B2(n9276), .A(n11491), .ZN(P1_U3471) );
  OAI21_X1 U14193 ( .B1(n11493), .B2(n12767), .A(n11492), .ZN(n15621) );
  INV_X1 U14194 ( .A(n15621), .ZN(n11502) );
  OR2_X1 U14195 ( .A1(n15603), .A2(n6928), .ZN(n15571) );
  INV_X1 U14196 ( .A(n15588), .ZN(n15642) );
  OAI22_X1 U14197 ( .A1(n11494), .A2(n15582), .B1(n11784), .B2(n15580), .ZN(
        n11497) );
  AOI211_X1 U14198 ( .C1(n12767), .C2(n11495), .A(n15601), .B(n7196), .ZN(
        n11496) );
  AOI211_X1 U14199 ( .C1(n15642), .C2(n15621), .A(n11497), .B(n11496), .ZN(
        n15618) );
  MUX2_X1 U14200 ( .A(n7511), .B(n15618), .S(n15608), .Z(n11501) );
  INV_X1 U14201 ( .A(n11776), .ZN(n13165) );
  AND2_X1 U14202 ( .A1(n11498), .A2(n15623), .ZN(n15620) );
  AOI22_X1 U14203 ( .A1(n13165), .A2(n15620), .B1(n15604), .B2(n11499), .ZN(
        n11500) );
  OAI211_X1 U14204 ( .C1(n11502), .C2(n11773), .A(n11501), .B(n11500), .ZN(
        P3_U3230) );
  OR2_X1 U14205 ( .A1(n15588), .A2(n15610), .ZN(n11503) );
  OAI21_X1 U14206 ( .B1(n11505), .B2(n12771), .A(n11504), .ZN(n15641) );
  INV_X1 U14207 ( .A(n15641), .ZN(n11515) );
  OAI211_X1 U14208 ( .C1(n11508), .C2(n11507), .A(n11506), .B(n10349), .ZN(
        n11510) );
  INV_X1 U14209 ( .A(n15582), .ZN(n15595) );
  AOI22_X1 U14210 ( .A1(n12977), .A2(n15595), .B1(n15597), .B2(n12837), .ZN(
        n11509) );
  AND2_X1 U14211 ( .A1(n11510), .A2(n11509), .ZN(n15637) );
  MUX2_X1 U14212 ( .A(n15637), .B(n11511), .S(n15610), .Z(n11514) );
  INV_X1 U14213 ( .A(n11512), .ZN(n12722) );
  AOI22_X1 U14214 ( .A1(n13347), .A2(n12721), .B1(n15604), .B2(n12722), .ZN(
        n11513) );
  OAI211_X1 U14215 ( .C1(n13363), .C2(n11515), .A(n11514), .B(n11513), .ZN(
        P3_U3227) );
  INV_X1 U14216 ( .A(n11516), .ZN(n11517) );
  NAND2_X1 U14217 ( .A1(n11518), .A2(n11517), .ZN(n11597) );
  XNOR2_X1 U14218 ( .A(n11597), .B(n11519), .ZN(n11600) );
  XNOR2_X1 U14219 ( .A(n11600), .B(n11599), .ZN(n11524) );
  INV_X1 U14220 ( .A(n14380), .ZN(n14357) );
  NAND2_X1 U14221 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14699) );
  OAI21_X1 U14222 ( .B1(n14244), .B2(n11520), .A(n14699), .ZN(n11522) );
  NOR2_X1 U14223 ( .A1(n14291), .A2(n11553), .ZN(n11521) );
  AOI211_X1 U14224 ( .C1(n14357), .C2(n14404), .A(n11522), .B(n11521), .ZN(
        n11523) );
  OAI21_X1 U14225 ( .B1(n11524), .B2(n14359), .A(n11523), .ZN(P1_U3230) );
  INV_X1 U14226 ( .A(n11525), .ZN(n11527) );
  OAI222_X1 U14227 ( .A1(P2_U3088), .A2(n7381), .B1(n6438), .B2(n11527), .C1(
        n11526), .C2(n14184), .ZN(P2_U3309) );
  INV_X1 U14228 ( .A(n14779), .ZN(n14773) );
  OAI222_X1 U14229 ( .A1(n15185), .A2(n11528), .B1(n15188), .B2(n11527), .C1(
        n14773), .C2(n6428), .ZN(P1_U3337) );
  NAND2_X1 U14230 ( .A1(n15049), .A2(n15361), .ZN(n11529) );
  OAI22_X1 U14231 ( .A1(n15049), .A2(n10615), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15055), .ZN(n11531) );
  NOR2_X1 U14232 ( .A1(n15057), .A2(n14399), .ZN(n11530) );
  AOI211_X1 U14233 ( .C1(n11532), .C2(n15235), .A(n11531), .B(n11530), .ZN(
        n11535) );
  NAND2_X1 U14234 ( .A1(n11533), .A2(n15049), .ZN(n11534) );
  OAI211_X1 U14235 ( .C1(n11536), .C2(n14952), .A(n11535), .B(n11534), .ZN(
        P1_U3290) );
  INV_X1 U14236 ( .A(n11537), .ZN(n11538) );
  OAI222_X1 U14237 ( .A1(P3_U3151), .A2(n11540), .B1(n13522), .B2(n11539), 
        .C1(n13520), .C2(n11538), .ZN(P3_U3275) );
  OAI211_X1 U14238 ( .C1(n11543), .C2(n11542), .A(n11541), .B(n14370), .ZN(
        n11549) );
  INV_X1 U14239 ( .A(n11544), .ZN(n11641) );
  OR2_X1 U14240 ( .A1(n11948), .A2(n15052), .ZN(n11546) );
  NAND2_X1 U14241 ( .A1(n14650), .A2(n15223), .ZN(n11545) );
  AND2_X1 U14242 ( .A1(n11546), .A2(n11545), .ZN(n11639) );
  OAI22_X1 U14243 ( .A1(n11639), .A2(n14244), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9311), .ZN(n11547) );
  AOI21_X1 U14244 ( .B1(n14242), .B2(n11641), .A(n11547), .ZN(n11548) );
  OAI211_X1 U14245 ( .C1(n15364), .C2(n14380), .A(n11549), .B(n11548), .ZN(
        P1_U3239) );
  INV_X1 U14246 ( .A(n11550), .ZN(n11551) );
  MUX2_X1 U14247 ( .A(n11552), .B(n11551), .S(n15049), .Z(n11557) );
  OAI22_X1 U14248 ( .A1(n15057), .A2(n11622), .B1(n15055), .B2(n11553), .ZN(
        n11554) );
  AOI21_X1 U14249 ( .B1(n11555), .B2(n15235), .A(n11554), .ZN(n11556) );
  OAI211_X1 U14250 ( .C1(n11558), .C2(n15062), .A(n11557), .B(n11556), .ZN(
        P1_U3289) );
  OAI21_X1 U14251 ( .B1(n11561), .B2(n11560), .A(n11559), .ZN(n11562) );
  NAND2_X1 U14252 ( .A1(n11562), .A2(n12730), .ZN(n11567) );
  OAI22_X1 U14253 ( .A1(n12744), .A2(n11563), .B1(n12743), .B2(n11785), .ZN(
        n11564) );
  AOI211_X1 U14254 ( .C1(n12741), .C2(n12978), .A(n11565), .B(n11564), .ZN(
        n11566) );
  OAI211_X1 U14255 ( .C1(n11775), .C2(n12662), .A(n11567), .B(n11566), .ZN(
        P3_U3167) );
  XNOR2_X1 U14256 ( .A(n11842), .B(n12284), .ZN(n11844) );
  NAND2_X1 U14257 ( .A1(n11568), .A2(n12173), .ZN(n11569) );
  NAND2_X1 U14258 ( .A1(n11570), .A2(n11569), .ZN(n11845) );
  XOR2_X1 U14259 ( .A(n11844), .B(n11845), .Z(n11582) );
  XNOR2_X1 U14260 ( .A(n11842), .B(n11571), .ZN(n11575) );
  OAI21_X1 U14261 ( .B1(n11575), .B2(n11574), .A(n11839), .ZN(n11580) );
  NAND2_X1 U14262 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11577)
         );
  NAND2_X1 U14263 ( .A1(n15441), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n11576) );
  OAI211_X1 U14264 ( .C1(n15490), .C2(n11578), .A(n11577), .B(n11576), .ZN(
        n11579) );
  AOI21_X1 U14265 ( .B1(n11580), .B2(n15471), .A(n11579), .ZN(n11581) );
  OAI21_X1 U14266 ( .B1(n15421), .B2(n11582), .A(n11581), .ZN(P2_U3226) );
  XNOR2_X1 U14267 ( .A(n14650), .B(n11635), .ZN(n14586) );
  INV_X1 U14268 ( .A(n11583), .ZN(n11585) );
  INV_X1 U14269 ( .A(n14651), .ZN(n11623) );
  OAI21_X1 U14270 ( .B1(n11583), .B2(n11623), .A(n11622), .ZN(n11584) );
  OAI21_X1 U14271 ( .B1(n11585), .B2(n14651), .A(n11584), .ZN(n11586) );
  XOR2_X1 U14272 ( .A(n14586), .B(n11586), .Z(n15358) );
  AOI211_X1 U14273 ( .C1(n15355), .C2(n11587), .A(n15365), .B(n11645), .ZN(
        n15354) );
  OAI22_X1 U14274 ( .A1(n15057), .A2(n11635), .B1(n15055), .B2(n11609), .ZN(
        n11588) );
  AOI21_X1 U14275 ( .B1(n15354), .B2(n15235), .A(n11588), .ZN(n11596) );
  NAND2_X1 U14276 ( .A1(n14651), .A2(n11622), .ZN(n11590) );
  XNOR2_X1 U14277 ( .A(n11637), .B(n14586), .ZN(n11593) );
  NAND2_X1 U14278 ( .A1(n14651), .A2(n15223), .ZN(n11592) );
  NAND2_X1 U14279 ( .A1(n14649), .A2(n15222), .ZN(n11591) );
  NAND2_X1 U14280 ( .A1(n11592), .A2(n11591), .ZN(n11606) );
  AOI21_X1 U14281 ( .B1(n11593), .B2(n15024), .A(n11606), .ZN(n15357) );
  MUX2_X1 U14282 ( .A(n11594), .B(n15357), .S(n15049), .Z(n11595) );
  OAI211_X1 U14283 ( .C1(n15358), .C2(n14952), .A(n11596), .B(n11595), .ZN(
        P1_U3288) );
  AOI22_X1 U14284 ( .A1(n11600), .A2(n11599), .B1(n11598), .B2(n11597), .ZN(
        n11605) );
  OAI21_X1 U14285 ( .B1(n11603), .B2(n11602), .A(n11601), .ZN(n11604) );
  XNOR2_X1 U14286 ( .A(n11605), .B(n11604), .ZN(n11612) );
  NAND2_X1 U14287 ( .A1(n14368), .A2(n11606), .ZN(n11607) );
  OAI211_X1 U14288 ( .C1(n14291), .C2(n11609), .A(n11608), .B(n11607), .ZN(
        n11610) );
  AOI21_X1 U14289 ( .B1(n14357), .B2(n15355), .A(n11610), .ZN(n11611) );
  OAI21_X1 U14290 ( .B1(n11612), .B2(n14359), .A(n11611), .ZN(P1_U3227) );
  INV_X1 U14291 ( .A(n11613), .ZN(n12405) );
  OAI222_X1 U14292 ( .A1(n14184), .A2(n11615), .B1(n6438), .B2(n12405), .C1(
        P2_U3088), .C2(n11614), .ZN(P2_U3308) );
  NAND2_X1 U14293 ( .A1(n11616), .A2(n13500), .ZN(n11617) );
  OAI211_X1 U14294 ( .C1(n11618), .C2(n13522), .A(n11617), .B(n12959), .ZN(
        P3_U3272) );
  NAND2_X1 U14295 ( .A1(n14651), .A2(n14404), .ZN(n11620) );
  NAND2_X1 U14296 ( .A1(n14650), .A2(n15355), .ZN(n11619) );
  NAND2_X1 U14297 ( .A1(n11620), .A2(n11619), .ZN(n11631) );
  OAI21_X1 U14298 ( .B1(n14651), .B2(n14404), .A(n14650), .ZN(n11621) );
  NAND2_X1 U14299 ( .A1(n11621), .A2(n11635), .ZN(n11626) );
  INV_X1 U14300 ( .A(n14650), .ZN(n11624) );
  NAND3_X1 U14301 ( .A1(n11624), .A2(n11623), .A3(n11622), .ZN(n11625) );
  OAI211_X1 U14302 ( .C1(n11631), .C2(n11627), .A(n11626), .B(n11625), .ZN(
        n11628) );
  INV_X1 U14303 ( .A(n11628), .ZN(n11634) );
  AND2_X1 U14304 ( .A1(n14652), .A2(n11629), .ZN(n11630) );
  NOR2_X1 U14305 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  XNOR2_X1 U14306 ( .A(n14649), .B(n14413), .ZN(n14589) );
  XNOR2_X1 U14307 ( .A(n11680), .B(n14589), .ZN(n15369) );
  INV_X1 U14308 ( .A(n15055), .ZN(n15331) );
  AND2_X1 U14309 ( .A1(n14650), .A2(n11635), .ZN(n11636) );
  XNOR2_X1 U14310 ( .A(n11681), .B(n14589), .ZN(n11638) );
  NAND2_X1 U14311 ( .A1(n11638), .A2(n15024), .ZN(n11640) );
  NAND2_X1 U14312 ( .A1(n11640), .A2(n11639), .ZN(n15372) );
  AOI21_X1 U14313 ( .B1(n11641), .B2(n15331), .A(n15372), .ZN(n11642) );
  MUX2_X1 U14314 ( .A(n11643), .B(n11642), .S(n15049), .Z(n11649) );
  NOR2_X1 U14315 ( .A1(n11645), .A2(n15364), .ZN(n11646) );
  OR2_X1 U14316 ( .A1(n11644), .A2(n11646), .ZN(n15366) );
  INV_X1 U14317 ( .A(n15366), .ZN(n11647) );
  AOI22_X1 U14318 ( .A1(n11647), .A2(n14950), .B1(n15329), .B2(n14413), .ZN(
        n11648) );
  OAI211_X1 U14319 ( .C1(n14952), .C2(n15369), .A(n11649), .B(n11648), .ZN(
        P1_U3287) );
  INV_X1 U14320 ( .A(n11650), .ZN(n11652) );
  OAI222_X1 U14321 ( .A1(n6928), .A2(P3_U3151), .B1(n13520), .B2(n11652), .C1(
        n11651), .C2(n13522), .ZN(P3_U3274) );
  INV_X1 U14322 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12064) );
  XNOR2_X1 U14323 ( .A(n11808), .B(n11656), .ZN(n11806) );
  XNOR2_X1 U14324 ( .A(n6626), .B(n11806), .ZN(n11677) );
  MUX2_X1 U14325 ( .A(n11657), .B(n11656), .S(n7029), .Z(n11659) );
  INV_X1 U14326 ( .A(n11808), .ZN(n11658) );
  NAND2_X1 U14327 ( .A1(n11659), .A2(n11658), .ZN(n11812) );
  INV_X1 U14328 ( .A(n11659), .ZN(n11660) );
  NAND2_X1 U14329 ( .A1(n11660), .A2(n11808), .ZN(n11661) );
  AND2_X1 U14330 ( .A1(n11812), .A2(n11661), .ZN(n11662) );
  INV_X1 U14331 ( .A(n11662), .ZN(n11663) );
  NAND3_X1 U14332 ( .A1(n11665), .A2(n11664), .A3(n11663), .ZN(n11666) );
  AOI21_X1 U14333 ( .B1(n11813), .B2(n11666), .A(n13125), .ZN(n11676) );
  INV_X1 U14334 ( .A(n11667), .ZN(n11668) );
  XNOR2_X1 U14335 ( .A(n11808), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n11669) );
  AND3_X1 U14336 ( .A1(n11670), .A2(n11669), .A3(n11668), .ZN(n11671) );
  OAI21_X1 U14337 ( .B1(n11807), .B2(n11671), .A(n13112), .ZN(n11674) );
  NAND2_X1 U14338 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11909)
         );
  INV_X1 U14339 ( .A(n11909), .ZN(n11672) );
  AOI21_X1 U14340 ( .B1(n15570), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11672), 
        .ZN(n11673) );
  OAI211_X1 U14341 ( .C1(n13147), .C2(n11808), .A(n11674), .B(n11673), .ZN(
        n11675) );
  AOI211_X1 U14342 ( .C1(n13122), .C2(n11677), .A(n11676), .B(n11675), .ZN(
        n11678) );
  INV_X1 U14343 ( .A(n11678), .ZN(P3_U3192) );
  INV_X1 U14344 ( .A(n14589), .ZN(n11679) );
  XNOR2_X1 U14345 ( .A(n14419), .B(n11948), .ZN(n11918) );
  INV_X1 U14346 ( .A(n11918), .ZN(n14588) );
  XNOR2_X1 U14347 ( .A(n11919), .B(n14588), .ZN(n15376) );
  OR2_X1 U14348 ( .A1(n14649), .A2(n15364), .ZN(n11682) );
  XNOR2_X1 U14349 ( .A(n11926), .B(n14588), .ZN(n11684) );
  INV_X1 U14350 ( .A(n14649), .ZN(n11683) );
  INV_X1 U14351 ( .A(n14648), .ZN(n11927) );
  OAI22_X1 U14352 ( .A1(n11683), .A2(n14976), .B1(n11927), .B2(n15052), .ZN(
        n11746) );
  AOI21_X1 U14353 ( .B1(n11684), .B2(n15024), .A(n11746), .ZN(n15373) );
  MUX2_X1 U14354 ( .A(n11685), .B(n15373), .S(n15049), .Z(n11692) );
  INV_X1 U14355 ( .A(n11644), .ZN(n11688) );
  INV_X1 U14356 ( .A(n11686), .ZN(n11687) );
  AOI211_X1 U14357 ( .C1(n14419), .C2(n11688), .A(n15365), .B(n11687), .ZN(
        n15379) );
  OAI22_X1 U14358 ( .A1(n15057), .A2(n11689), .B1(n15055), .B2(n11743), .ZN(
        n11690) );
  AOI21_X1 U14359 ( .B1(n15379), .B2(n15235), .A(n11690), .ZN(n11691) );
  OAI211_X1 U14360 ( .C1(n14952), .C2(n15376), .A(n11692), .B(n11691), .ZN(
        P1_U3286) );
  OAI21_X1 U14361 ( .B1(n11695), .B2(n11694), .A(n11693), .ZN(n11696) );
  OAI21_X1 U14362 ( .B1(n11697), .B2(n11472), .A(n11696), .ZN(n11701) );
  XNOR2_X1 U14363 ( .A(n11699), .B(n11698), .ZN(n11700) );
  XNOR2_X1 U14364 ( .A(n11701), .B(n11700), .ZN(n11707) );
  OAI22_X1 U14365 ( .A1(n12168), .A2(n13932), .B1(n11702), .B2(n13930), .ZN(
        n11977) );
  AOI21_X1 U14366 ( .B1(n13643), .B2(n11977), .A(n11703), .ZN(n11704) );
  OAI21_X1 U14367 ( .B1(n13645), .B2(n11983), .A(n11704), .ZN(n11705) );
  AOI21_X1 U14368 ( .B1(n14106), .B2(n13647), .A(n11705), .ZN(n11706) );
  OAI21_X1 U14369 ( .B1(n11707), .B2(n13649), .A(n11706), .ZN(P2_U3203) );
  INV_X1 U14370 ( .A(n11708), .ZN(n12563) );
  OAI222_X1 U14371 ( .A1(n15174), .A2(n11710), .B1(n6428), .B2(n11709), .C1(
        n15188), .C2(n12563), .ZN(P1_U3335) );
  XNOR2_X1 U14372 ( .A(n12347), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n11716) );
  NAND2_X1 U14373 ( .A1(n11711), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11712) );
  NAND2_X1 U14374 ( .A1(n11713), .A2(n11712), .ZN(n11715) );
  INV_X1 U14375 ( .A(n12349), .ZN(n11714) );
  AOI21_X1 U14376 ( .B1(n11716), .B2(n11715), .A(n11714), .ZN(n11729) );
  INV_X1 U14377 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11717) );
  MUX2_X1 U14378 ( .A(n11717), .B(P1_REG2_REG_14__SCAN_IN), .S(n12347), .Z(
        n11720) );
  NOR2_X1 U14379 ( .A1(n11718), .A2(n15034), .ZN(n11722) );
  INV_X1 U14380 ( .A(n11722), .ZN(n11719) );
  NAND2_X1 U14381 ( .A1(n11720), .A2(n11719), .ZN(n11723) );
  MUX2_X1 U14382 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11717), .S(n12347), .Z(
        n11721) );
  OAI21_X1 U14383 ( .B1(n11724), .B2(n11722), .A(n11721), .ZN(n12341) );
  OAI211_X1 U14384 ( .C1(n11724), .C2(n11723), .A(n12341), .B(n14785), .ZN(
        n11728) );
  NOR2_X1 U14385 ( .A1(n11725), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14194) );
  NOR2_X1 U14386 ( .A1(n15315), .A2(n12342), .ZN(n11726) );
  AOI211_X1 U14387 ( .C1(n15299), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n14194), 
        .B(n11726), .ZN(n11727) );
  OAI211_X1 U14388 ( .C1(n11729), .C2(n6633), .A(n11728), .B(n11727), .ZN(
        P1_U3257) );
  XNOR2_X1 U14389 ( .A(n11730), .B(n11733), .ZN(n15626) );
  INV_X1 U14390 ( .A(n15626), .ZN(n15629) );
  INV_X1 U14391 ( .A(n13363), .ZN(n13245) );
  OAI22_X1 U14392 ( .A1(n13340), .A2(n11732), .B1(n11731), .B2(n15577), .ZN(
        n11738) );
  NAND2_X1 U14393 ( .A1(n11779), .A2(n7839), .ZN(n11734) );
  NAND2_X1 U14394 ( .A1(n11734), .A2(n11733), .ZN(n11778) );
  OAI211_X1 U14395 ( .C1(n11734), .C2(n11733), .A(n11778), .B(n10349), .ZN(
        n11736) );
  NAND2_X1 U14396 ( .A1(n12977), .A2(n15597), .ZN(n11735) );
  OAI211_X1 U14397 ( .C1(n15581), .C2(n15582), .A(n11736), .B(n11735), .ZN(
        n15622) );
  MUX2_X1 U14398 ( .A(n15622), .B(P3_REG2_REG_4__SCAN_IN), .S(n15610), .Z(
        n11737) );
  AOI211_X1 U14399 ( .C1(n15629), .C2(n13245), .A(n11738), .B(n11737), .ZN(
        n11739) );
  INV_X1 U14400 ( .A(n11739), .ZN(P3_U3229) );
  AND2_X1 U14401 ( .A1(n14419), .A2(n15400), .ZN(n15378) );
  INV_X1 U14402 ( .A(n15378), .ZN(n11749) );
  OAI211_X1 U14403 ( .C1(n11742), .C2(n11741), .A(n11740), .B(n14370), .ZN(
        n11748) );
  NOR2_X1 U14404 ( .A1(n14291), .A2(n11743), .ZN(n11744) );
  AOI211_X1 U14405 ( .C1(n14368), .C2(n11746), .A(n11745), .B(n11744), .ZN(
        n11747) );
  OAI211_X1 U14406 ( .C1(n14308), .C2(n11749), .A(n11748), .B(n11747), .ZN(
        P1_U3213) );
  OAI211_X1 U14407 ( .C1(n6469), .C2(n11751), .A(n11750), .B(n13610), .ZN(
        n11759) );
  INV_X1 U14408 ( .A(n11752), .ZN(n11963) );
  OR2_X1 U14409 ( .A1(n12195), .A2(n13932), .ZN(n11753) );
  OAI21_X1 U14410 ( .B1(n11754), .B2(n13930), .A(n11753), .ZN(n11960) );
  INV_X1 U14411 ( .A(n11960), .ZN(n11756) );
  OAI22_X1 U14412 ( .A1(n13616), .A2(n11756), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11755), .ZN(n11757) );
  AOI21_X1 U14413 ( .B1(n11963), .B2(n13631), .A(n11757), .ZN(n11758) );
  OAI211_X1 U14414 ( .C1(n12110), .C2(n13620), .A(n11759), .B(n11758), .ZN(
        P2_U3189) );
  INV_X1 U14415 ( .A(n15627), .ZN(n15635) );
  XNOR2_X1 U14416 ( .A(n7014), .B(n12835), .ZN(n12086) );
  NAND2_X1 U14417 ( .A1(n12086), .A2(n15642), .ZN(n11766) );
  OAI211_X1 U14418 ( .C1(n11761), .C2(n7717), .A(n11795), .B(n10349), .ZN(
        n11764) );
  OAI22_X1 U14419 ( .A1(n11785), .A2(n15582), .B1(n12843), .B2(n15580), .ZN(
        n11762) );
  INV_X1 U14420 ( .A(n11762), .ZN(n11763) );
  AND2_X1 U14421 ( .A1(n11764), .A2(n11763), .ZN(n11765) );
  NAND2_X1 U14422 ( .A1(n11766), .A2(n11765), .ZN(n12083) );
  AOI21_X1 U14423 ( .B1(n15635), .B2(n12086), .A(n12083), .ZN(n11870) );
  AOI22_X1 U14424 ( .A1(n13493), .A2(n11767), .B1(P3_REG0_REG_7__SCAN_IN), 
        .B2(n15643), .ZN(n11768) );
  OAI21_X1 U14425 ( .B1(n11870), .B2(n15643), .A(n11768), .ZN(P3_U3411) );
  INV_X1 U14426 ( .A(n11769), .ZN(n12565) );
  OAI222_X1 U14427 ( .A1(n14184), .A2(n11771), .B1(n6438), .B2(n12565), .C1(
        P2_U3088), .C2(n11770), .ZN(P2_U3306) );
  XNOR2_X1 U14428 ( .A(n11772), .B(n12824), .ZN(n15633) );
  INV_X1 U14429 ( .A(n11773), .ZN(n15605) );
  NAND2_X1 U14430 ( .A1(n11774), .A2(n15623), .ZN(n15630) );
  OAI22_X1 U14431 ( .A1(n11776), .A2(n15630), .B1(n11775), .B2(n15577), .ZN(
        n11791) );
  NAND2_X1 U14432 ( .A1(n15633), .A2(n15642), .ZN(n11789) );
  AOI21_X1 U14433 ( .B1(n11778), .B2(n11777), .A(n12768), .ZN(n11783) );
  OR2_X1 U14434 ( .A1(n11779), .A2(n12819), .ZN(n11781) );
  AND2_X1 U14435 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  OAI21_X1 U14436 ( .B1(n11783), .B2(n11782), .A(n10349), .ZN(n11788) );
  OAI22_X1 U14437 ( .A1(n11785), .A2(n15580), .B1(n11784), .B2(n15582), .ZN(
        n11786) );
  INV_X1 U14438 ( .A(n11786), .ZN(n11787) );
  NAND3_X1 U14439 ( .A1(n11789), .A2(n11788), .A3(n11787), .ZN(n15631) );
  MUX2_X1 U14440 ( .A(n15631), .B(P3_REG2_REG_5__SCAN_IN), .S(n15610), .Z(
        n11790) );
  AOI211_X1 U14441 ( .C1(n15633), .C2(n15605), .A(n11791), .B(n11790), .ZN(
        n11792) );
  INV_X1 U14442 ( .A(n11792), .ZN(P3_U3228) );
  XOR2_X1 U14443 ( .A(n12846), .B(n11793), .Z(n12063) );
  INV_X1 U14444 ( .A(n12063), .ZN(n11805) );
  NAND2_X1 U14445 ( .A1(n11795), .A2(n11794), .ZN(n12071) );
  OR2_X1 U14446 ( .A1(n12071), .A2(n6437), .ZN(n12073) );
  AOI21_X1 U14447 ( .B1(n12073), .B2(n11796), .A(n12846), .ZN(n11800) );
  NAND2_X1 U14448 ( .A1(n11797), .A2(n10349), .ZN(n11799) );
  AOI22_X1 U14449 ( .A1(n15595), .A2(n11855), .B1(n12974), .B2(n15597), .ZN(
        n11798) );
  OAI21_X1 U14450 ( .B1(n11800), .B2(n11799), .A(n11798), .ZN(n12062) );
  NOR2_X1 U14451 ( .A1(n15577), .A2(n11856), .ZN(n11801) );
  AOI21_X1 U14452 ( .B1(n15610), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11801), .ZN(
        n11802) );
  OAI21_X1 U14453 ( .B1(n13340), .B2(n12069), .A(n11802), .ZN(n11803) );
  AOI21_X1 U14454 ( .B1(n12062), .B2(n15608), .A(n11803), .ZN(n11804) );
  OAI21_X1 U14455 ( .B1(n11805), .B2(n13363), .A(n11804), .ZN(P3_U3224) );
  INV_X1 U14456 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n12245) );
  XNOR2_X1 U14457 ( .A(n11876), .B(n12245), .ZN(n11822) );
  AOI21_X1 U14458 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11808), .A(n11807), 
        .ZN(n11809) );
  INV_X1 U14459 ( .A(n11875), .ZN(n11884) );
  OAI21_X1 U14460 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n11810), .A(n11880), 
        .ZN(n11811) );
  NAND2_X1 U14461 ( .A1(n11811), .A2(n13112), .ZN(n11821) );
  MUX2_X1 U14462 ( .A(n12251), .B(n12245), .S(n7029), .Z(n11883) );
  XNOR2_X1 U14463 ( .A(n11883), .B(n11875), .ZN(n11814) );
  OAI21_X1 U14464 ( .B1(n11815), .B2(n11814), .A(n11888), .ZN(n11819) );
  INV_X1 U14465 ( .A(n13147), .ZN(n13100) );
  NAND2_X1 U14466 ( .A1(n13100), .A2(n11884), .ZN(n11816) );
  NAND2_X1 U14467 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12368)
         );
  OAI211_X1 U14468 ( .C1(n11817), .C2(n13074), .A(n11816), .B(n12368), .ZN(
        n11818) );
  AOI21_X1 U14469 ( .B1(n11819), .B2(n13149), .A(n11818), .ZN(n11820) );
  OAI211_X1 U14470 ( .C1(n11822), .C2(n13143), .A(n11821), .B(n11820), .ZN(
        P3_U3193) );
  AND2_X1 U14471 ( .A1(n11823), .A2(n13987), .ZN(n13993) );
  AOI22_X1 U14472 ( .A1(n11825), .A2(n13995), .B1(n13993), .B2(n11824), .ZN(
        n11830) );
  INV_X1 U14473 ( .A(n11825), .ZN(n11827) );
  OAI21_X1 U14474 ( .B1(n12562), .B2(n11827), .A(n11826), .ZN(n11828) );
  AOI22_X1 U14475 ( .A1(n11828), .A2(n13987), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13990), .ZN(n11829) );
  OAI211_X1 U14476 ( .C1(n7622), .C2(n13987), .A(n11830), .B(n11829), .ZN(
        P2_U3265) );
  AND2_X1 U14477 ( .A1(n11559), .A2(n11831), .ZN(n12718) );
  XNOR2_X1 U14478 ( .A(n11832), .B(n12976), .ZN(n12717) );
  NAND2_X1 U14479 ( .A1(n12718), .A2(n12717), .ZN(n12716) );
  NAND2_X1 U14480 ( .A1(n12716), .A2(n11833), .ZN(n12138) );
  XNOR2_X1 U14481 ( .A(n12138), .B(n12137), .ZN(n11834) );
  NAND2_X1 U14482 ( .A1(n11834), .A2(n12730), .ZN(n11838) );
  OAI22_X1 U14483 ( .A1(n12744), .A2(n12838), .B1(n12743), .B2(n12843), .ZN(
        n11835) );
  AOI211_X1 U14484 ( .C1(n12741), .C2(n12976), .A(n11836), .B(n11835), .ZN(
        n11837) );
  OAI211_X1 U14485 ( .C1(n12082), .C2(n12662), .A(n11838), .B(n11837), .ZN(
        P3_U3153) );
  XNOR2_X1 U14486 ( .A(n12392), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n11841) );
  AOI211_X1 U14487 ( .C1(n11841), .C2(n11840), .A(n15513), .B(n12388), .ZN(
        n11854) );
  NOR2_X1 U14488 ( .A1(n11842), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11843) );
  AOI21_X1 U14489 ( .B1(n11845), .B2(n11844), .A(n11843), .ZN(n11848) );
  INV_X1 U14490 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11846) );
  XNOR2_X1 U14491 ( .A(n12392), .B(n11846), .ZN(n11847) );
  NAND2_X1 U14492 ( .A1(n11848), .A2(n11847), .ZN(n12394) );
  OAI211_X1 U14493 ( .C1(n11848), .C2(n11847), .A(n12394), .B(n15508), .ZN(
        n11851) );
  NOR2_X1 U14494 ( .A1(n11849), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12311) );
  AOI21_X1 U14495 ( .B1(n15441), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n12311), 
        .ZN(n11850) );
  OAI211_X1 U14496 ( .C1(n15490), .C2(n11852), .A(n11851), .B(n11850), .ZN(
        n11853) );
  OR2_X1 U14497 ( .A1(n11854), .A2(n11853), .ZN(P2_U3227) );
  INV_X1 U14498 ( .A(n12069), .ZN(n11868) );
  NAND2_X1 U14499 ( .A1(n12741), .A2(n11855), .ZN(n11861) );
  NAND2_X1 U14500 ( .A1(n12735), .A2(n12974), .ZN(n11860) );
  INV_X1 U14501 ( .A(n11856), .ZN(n11857) );
  NAND2_X1 U14502 ( .A1(n12747), .A2(n11857), .ZN(n11859) );
  NAND4_X1 U14503 ( .A1(n11861), .A2(n11860), .A3(n11859), .A4(n11858), .ZN(
        n11867) );
  NAND2_X1 U14504 ( .A1(n11864), .A2(n11863), .ZN(n11865) );
  AOI21_X1 U14505 ( .B1(n11862), .B2(n11865), .A(n12749), .ZN(n11866) );
  AOI211_X1 U14506 ( .C1(n11868), .C2(n12720), .A(n11867), .B(n11866), .ZN(
        n11869) );
  INV_X1 U14507 ( .A(n11869), .ZN(P3_U3171) );
  MUX2_X1 U14508 ( .A(n11871), .B(n11870), .S(n15652), .Z(n11872) );
  OAI21_X1 U14509 ( .B1(n13382), .B2(n12838), .A(n11872), .ZN(P3_U3466) );
  XNOR2_X1 U14510 ( .A(n12988), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n12981) );
  INV_X1 U14511 ( .A(n11873), .ZN(n11874) );
  XOR2_X1 U14512 ( .A(n12982), .B(n12981), .Z(n11895) );
  XNOR2_X1 U14513 ( .A(n12980), .B(n12338), .ZN(n11879) );
  AND3_X1 U14514 ( .A1(n11880), .A2(n11879), .A3(n11878), .ZN(n11881) );
  OAI21_X1 U14515 ( .B1(n12986), .B2(n11881), .A(n13112), .ZN(n11894) );
  NAND2_X1 U14516 ( .A1(n15570), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n11882) );
  NAND2_X1 U14517 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12658)
         );
  NAND2_X1 U14518 ( .A1(n11882), .A2(n12658), .ZN(n11892) );
  MUX2_X1 U14519 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n7029), .Z(n12989) );
  XNOR2_X1 U14520 ( .A(n12989), .B(n12980), .ZN(n11886) );
  NAND2_X1 U14521 ( .A1(n11884), .A2(n11883), .ZN(n11887) );
  AND2_X1 U14522 ( .A1(n11886), .A2(n11887), .ZN(n11885) );
  INV_X1 U14523 ( .A(n12993), .ZN(n11890) );
  AOI21_X1 U14524 ( .B1(n11888), .B2(n11887), .A(n11886), .ZN(n11889) );
  NOR3_X1 U14525 ( .A1(n11890), .A2(n11889), .A3(n13125), .ZN(n11891) );
  AOI211_X1 U14526 ( .C1(n13100), .C2(n12980), .A(n11892), .B(n11891), .ZN(
        n11893) );
  OAI211_X1 U14527 ( .C1(n11895), .C2(n13143), .A(n11894), .B(n11893), .ZN(
        P3_U3194) );
  NAND2_X1 U14528 ( .A1(n11897), .A2(n11896), .ZN(n11899) );
  XOR2_X1 U14529 ( .A(n11899), .B(n11898), .Z(n11904) );
  OAI21_X1 U14530 ( .B1(n13623), .B2(n12168), .A(n11900), .ZN(n11902) );
  OAI22_X1 U14531 ( .A1(n13634), .A2(n12295), .B1(n13645), .B2(n12172), .ZN(
        n11901) );
  AOI211_X1 U14532 ( .C1(n12171), .C2(n13647), .A(n11902), .B(n11901), .ZN(
        n11903) );
  OAI21_X1 U14533 ( .B1(n11904), .B2(n13649), .A(n11903), .ZN(P2_U3208) );
  AND2_X1 U14534 ( .A1(n11862), .A2(n11905), .ZN(n11908) );
  OAI211_X1 U14535 ( .C1(n11908), .C2(n11907), .A(n12730), .B(n11906), .ZN(
        n11914) );
  OAI21_X1 U14536 ( .B1(n12733), .B2(n11910), .A(n11909), .ZN(n11912) );
  NOR2_X1 U14537 ( .A1(n12662), .A2(n12156), .ZN(n11911) );
  AOI211_X1 U14538 ( .C1(n12735), .C2(n12973), .A(n11912), .B(n11911), .ZN(
        n11913) );
  OAI211_X1 U14539 ( .C1(n12744), .C2(n12852), .A(n11914), .B(n11913), .ZN(
        P3_U3157) );
  AOI222_X1 U14540 ( .A1(n11916), .A2(n14175), .B1(P1_DATAO_REG_22__SCAN_IN), 
        .B2(n14169), .C1(n11915), .C2(P2_STATE_REG_SCAN_IN), .ZN(n11917) );
  INV_X1 U14541 ( .A(n11917), .ZN(P2_U3305) );
  NAND2_X1 U14542 ( .A1(n11919), .A2(n11918), .ZN(n11921) );
  INV_X1 U14543 ( .A(n11948), .ZN(n14418) );
  OR2_X1 U14544 ( .A1(n14419), .A2(n14418), .ZN(n11920) );
  NAND2_X2 U14545 ( .A1(n11921), .A2(n11920), .ZN(n12179) );
  XNOR2_X1 U14546 ( .A(n14424), .B(n14648), .ZN(n14590) );
  INV_X1 U14547 ( .A(n14590), .ZN(n12183) );
  OR2_X1 U14548 ( .A1(n14424), .A2(n14648), .ZN(n11922) );
  OR2_X1 U14549 ( .A1(n15399), .A2(n14439), .ZN(n11931) );
  NAND2_X1 U14550 ( .A1(n15399), .A2(n14439), .ZN(n11930) );
  NAND2_X1 U14551 ( .A1(n11931), .A2(n11930), .ZN(n15046) );
  INV_X1 U14552 ( .A(n14439), .ZN(n14437) );
  OR2_X1 U14553 ( .A1(n15399), .A2(n14437), .ZN(n11923) );
  XNOR2_X1 U14554 ( .A(n14438), .B(n15053), .ZN(n14593) );
  XNOR2_X1 U14555 ( .A(n12440), .B(n14593), .ZN(n15257) );
  INV_X1 U14556 ( .A(n15257), .ZN(n11944) );
  AND2_X1 U14557 ( .A1(n14419), .A2(n11948), .ZN(n11925) );
  OR2_X1 U14558 ( .A1(n14419), .A2(n11948), .ZN(n11924) );
  OR2_X1 U14559 ( .A1(n14424), .A2(n11927), .ZN(n12214) );
  OAI211_X1 U14560 ( .C1(n11949), .C2(n14428), .A(n11931), .B(n12214), .ZN(
        n11928) );
  NAND2_X1 U14561 ( .A1(n14428), .A2(n11949), .ZN(n15041) );
  NAND2_X1 U14562 ( .A1(n11930), .A2(n15041), .ZN(n11932) );
  INV_X1 U14563 ( .A(n14593), .ZN(n11933) );
  XNOR2_X1 U14564 ( .A(n12409), .B(n11933), .ZN(n11934) );
  NAND2_X1 U14565 ( .A1(n11934), .A2(n15024), .ZN(n11936) );
  AOI22_X1 U14566 ( .A1(n14437), .A2(n15223), .B1(n15222), .B2(n15027), .ZN(
        n11935) );
  NAND2_X1 U14567 ( .A1(n11936), .A2(n11935), .ZN(n15262) );
  OAI211_X1 U14568 ( .C1(n11937), .C2(n15259), .A(n15333), .B(n11938), .ZN(
        n15258) );
  OAI22_X1 U14569 ( .A1(n15049), .A2(n11939), .B1(n14343), .B2(n15055), .ZN(
        n11940) );
  AOI21_X1 U14570 ( .B1(n14438), .B2(n15329), .A(n11940), .ZN(n11941) );
  OAI21_X1 U14571 ( .B1(n15258), .B2(n14860), .A(n11941), .ZN(n11942) );
  AOI21_X1 U14572 ( .B1(n15262), .B2(n15049), .A(n11942), .ZN(n11943) );
  OAI21_X1 U14573 ( .B1(n15062), .B2(n11944), .A(n11943), .ZN(P1_U3282) );
  AOI21_X1 U14574 ( .B1(n11947), .B2(n11946), .A(n11945), .ZN(n11957) );
  INV_X1 U14575 ( .A(n12185), .ZN(n11955) );
  OR2_X1 U14576 ( .A1(n11948), .A2(n14976), .ZN(n11951) );
  OR2_X1 U14577 ( .A1(n11949), .A2(n15052), .ZN(n11950) );
  AND2_X1 U14578 ( .A1(n11951), .A2(n11950), .ZN(n15384) );
  OAI22_X1 U14579 ( .A1(n15384), .A2(n14244), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11952), .ZN(n11954) );
  NAND2_X1 U14580 ( .A1(n14424), .A2(n15400), .ZN(n15382) );
  NOR2_X1 U14581 ( .A1(n15382), .A2(n14308), .ZN(n11953) );
  AOI211_X1 U14582 ( .C1(n11955), .C2(n14242), .A(n11954), .B(n11953), .ZN(
        n11956) );
  OAI21_X1 U14583 ( .B1(n11957), .B2(n14359), .A(n11956), .ZN(P1_U3221) );
  INV_X1 U14584 ( .A(n11969), .ZN(n11959) );
  OAI21_X1 U14585 ( .B1(n6611), .B2(n11959), .A(n12164), .ZN(n11961) );
  AOI21_X1 U14586 ( .B1(n11961), .B2(n13971), .A(n11960), .ZN(n12109) );
  OAI211_X1 U14587 ( .C1(n11981), .C2(n12110), .A(n12569), .B(n12170), .ZN(
        n12108) );
  INV_X1 U14588 ( .A(n12108), .ZN(n11966) );
  AOI22_X1 U14589 ( .A1(n13909), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11963), 
        .B2(n13990), .ZN(n11964) );
  OAI21_X1 U14590 ( .B1(n12110), .B2(n13979), .A(n11964), .ZN(n11965) );
  AOI21_X1 U14591 ( .B1(n11966), .B2(n13995), .A(n11965), .ZN(n11971) );
  INV_X1 U14592 ( .A(n11976), .ZN(n11973) );
  NAND2_X1 U14593 ( .A1(n7031), .A2(n11973), .ZN(n11972) );
  NAND2_X1 U14594 ( .A1(n11972), .A2(n11967), .ZN(n11968) );
  XOR2_X1 U14595 ( .A(n11969), .B(n11968), .Z(n12112) );
  INV_X1 U14596 ( .A(n13983), .ZN(n12130) );
  NAND2_X1 U14597 ( .A1(n12112), .A2(n12130), .ZN(n11970) );
  OAI211_X1 U14598 ( .C1(n12109), .C2(n13909), .A(n11971), .B(n11970), .ZN(
        P2_U3255) );
  OAI21_X1 U14599 ( .B1(n7031), .B2(n11973), .A(n11972), .ZN(n14109) );
  XNOR2_X1 U14600 ( .A(n11975), .B(n11976), .ZN(n11978) );
  AOI21_X1 U14601 ( .B1(n11978), .B2(n13971), .A(n11977), .ZN(n14107) );
  MUX2_X1 U14602 ( .A(n11979), .B(n14107), .S(n13987), .Z(n11987) );
  INV_X1 U14603 ( .A(n12012), .ZN(n11982) );
  AOI211_X1 U14604 ( .C1(n14106), .C2(n11982), .A(n13974), .B(n11981), .ZN(
        n14105) );
  OAI22_X1 U14605 ( .A1(n13979), .A2(n11984), .B1(n11983), .B2(n13956), .ZN(
        n11985) );
  AOI21_X1 U14606 ( .B1(n14105), .B2(n13995), .A(n11985), .ZN(n11986) );
  OAI211_X1 U14607 ( .C1(n13983), .C2(n14109), .A(n11987), .B(n11986), .ZN(
        P2_U3256) );
  OR2_X1 U14608 ( .A1(n11989), .A2(n11988), .ZN(n11990) );
  NAND2_X1 U14609 ( .A1(n11991), .A2(n11990), .ZN(n15556) );
  XNOR2_X1 U14610 ( .A(n11993), .B(n11992), .ZN(n11996) );
  INV_X1 U14611 ( .A(n11994), .ZN(n11995) );
  AOI21_X1 U14612 ( .B1(n11996), .B2(n13971), .A(n11995), .ZN(n15554) );
  MUX2_X1 U14613 ( .A(n15554), .B(n11997), .S(n13909), .Z(n12002) );
  AOI211_X1 U14614 ( .C1(n15552), .C2(n12041), .A(n13974), .B(n12011), .ZN(
        n15551) );
  OAI22_X1 U14615 ( .A1(n13979), .A2(n11999), .B1(n13956), .B2(n11998), .ZN(
        n12000) );
  AOI21_X1 U14616 ( .B1(n15551), .B2(n13995), .A(n12000), .ZN(n12001) );
  OAI211_X1 U14617 ( .C1(n13983), .C2(n15556), .A(n12002), .B(n12001), .ZN(
        P2_U3258) );
  OAI21_X1 U14618 ( .B1(n12005), .B2(n12004), .A(n12003), .ZN(n14114) );
  XNOR2_X1 U14619 ( .A(n12006), .B(n12007), .ZN(n12009) );
  AOI21_X1 U14620 ( .B1(n12009), .B2(n13971), .A(n12008), .ZN(n14112) );
  MUX2_X1 U14621 ( .A(n12010), .B(n14112), .S(n13987), .Z(n12018) );
  INV_X1 U14622 ( .A(n12011), .ZN(n12013) );
  AOI211_X1 U14623 ( .C1(n14111), .C2(n12013), .A(n13974), .B(n12012), .ZN(
        n14110) );
  OAI22_X1 U14624 ( .A1(n13979), .A2(n12015), .B1(n13956), .B2(n12014), .ZN(
        n12016) );
  AOI21_X1 U14625 ( .B1(n14110), .B2(n13995), .A(n12016), .ZN(n12017) );
  OAI211_X1 U14626 ( .C1(n13983), .C2(n14114), .A(n12018), .B(n12017), .ZN(
        P2_U3257) );
  INV_X1 U14627 ( .A(n13993), .ZN(n12034) );
  MUX2_X1 U14628 ( .A(n10535), .B(n12019), .S(n13987), .Z(n12024) );
  OAI22_X1 U14629 ( .A1(n13979), .A2(n11318), .B1(n13956), .B2(n12020), .ZN(
        n12021) );
  AOI21_X1 U14630 ( .B1(n12022), .B2(n13995), .A(n12021), .ZN(n12023) );
  OAI211_X1 U14631 ( .C1(n12025), .C2(n12034), .A(n12024), .B(n12023), .ZN(
        P2_U3260) );
  MUX2_X1 U14632 ( .A(n12027), .B(n12026), .S(n13987), .Z(n12033) );
  OAI22_X1 U14633 ( .A1(n13979), .A2(n12029), .B1(n12028), .B2(n13956), .ZN(
        n12030) );
  AOI21_X1 U14634 ( .B1(n12031), .B2(n13995), .A(n12030), .ZN(n12032) );
  OAI211_X1 U14635 ( .C1(n12035), .C2(n12034), .A(n12033), .B(n12032), .ZN(
        P2_U3261) );
  INV_X1 U14636 ( .A(n6949), .ZN(n12039) );
  OAI21_X1 U14637 ( .B1(n6949), .B2(n11318), .A(n12036), .ZN(n12037) );
  OAI21_X1 U14638 ( .B1(n12039), .B2(n12038), .A(n12037), .ZN(n12040) );
  XNOR2_X1 U14639 ( .A(n12040), .B(n12048), .ZN(n15547) );
  INV_X1 U14640 ( .A(n12041), .ZN(n12042) );
  AOI211_X1 U14641 ( .C1(n15543), .C2(n12043), .A(n13974), .B(n12042), .ZN(
        n15542) );
  AOI22_X1 U14642 ( .A1(n13909), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n12044), 
        .B2(n13990), .ZN(n12045) );
  OAI21_X1 U14643 ( .B1(n12046), .B2(n13979), .A(n12045), .ZN(n12053) );
  OAI21_X1 U14644 ( .B1(n12049), .B2(n12048), .A(n12047), .ZN(n12051) );
  AOI21_X1 U14645 ( .B1(n12051), .B2(n13971), .A(n12050), .ZN(n15545) );
  NOR2_X1 U14646 ( .A1(n15545), .A2(n13909), .ZN(n12052) );
  AOI211_X1 U14647 ( .C1(n15542), .C2(n13995), .A(n12053), .B(n12052), .ZN(
        n12054) );
  OAI21_X1 U14648 ( .B1(n13983), .B2(n15547), .A(n12054), .ZN(P2_U3259) );
  MUX2_X1 U14649 ( .A(n10512), .B(n12055), .S(n13987), .Z(n12060) );
  OAI22_X1 U14650 ( .A1(n13979), .A2(n12056), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13956), .ZN(n12057) );
  AOI21_X1 U14651 ( .B1(n13995), .B2(n12058), .A(n12057), .ZN(n12059) );
  OAI211_X1 U14652 ( .C1(n12061), .C2(n13983), .A(n12060), .B(n12059), .ZN(
        P2_U3262) );
  AOI21_X1 U14653 ( .B1(n12063), .B2(n13372), .A(n12062), .ZN(n12066) );
  MUX2_X1 U14654 ( .A(n12064), .B(n12066), .S(n15652), .Z(n12065) );
  OAI21_X1 U14655 ( .B1(n13382), .B2(n12069), .A(n12065), .ZN(P3_U3468) );
  INV_X1 U14656 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n12067) );
  MUX2_X1 U14657 ( .A(n12067), .B(n12066), .S(n15645), .Z(n12068) );
  OAI21_X1 U14658 ( .B1(n13443), .B2(n12069), .A(n12068), .ZN(P3_U3417) );
  INV_X1 U14659 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n12077) );
  XNOR2_X1 U14660 ( .A(n12070), .B(n12773), .ZN(n12205) );
  NAND2_X1 U14661 ( .A1(n12071), .A2(n6437), .ZN(n12072) );
  AND2_X1 U14662 ( .A1(n12073), .A2(n12072), .ZN(n12076) );
  NAND2_X1 U14663 ( .A1(n12205), .A2(n15642), .ZN(n12075) );
  AOI22_X1 U14664 ( .A1(n15595), .A2(n12837), .B1(n12975), .B2(n15597), .ZN(
        n12074) );
  OAI211_X1 U14665 ( .C1(n15601), .C2(n12076), .A(n12075), .B(n12074), .ZN(
        n12202) );
  AOI21_X1 U14666 ( .B1(n15635), .B2(n12205), .A(n12202), .ZN(n12079) );
  MUX2_X1 U14667 ( .A(n12077), .B(n12079), .S(n15645), .Z(n12078) );
  OAI21_X1 U14668 ( .B1(n12201), .B2(n13443), .A(n12078), .ZN(P3_U3414) );
  MUX2_X1 U14669 ( .A(n12080), .B(n12079), .S(n15652), .Z(n12081) );
  OAI21_X1 U14670 ( .B1(n12201), .B2(n13382), .A(n12081), .ZN(P3_U3467) );
  OAI22_X1 U14671 ( .A1(n13340), .A2(n12838), .B1(n12082), .B2(n15577), .ZN(
        n12085) );
  MUX2_X1 U14672 ( .A(n12083), .B(P3_REG2_REG_7__SCAN_IN), .S(n15610), .Z(
        n12084) );
  AOI211_X1 U14673 ( .C1(n12086), .C2(n15605), .A(n12085), .B(n12084), .ZN(
        n12087) );
  INV_X1 U14674 ( .A(n12087), .ZN(P3_U3226) );
  INV_X1 U14675 ( .A(n12088), .ZN(n12090) );
  OAI222_X1 U14676 ( .A1(P3_U3151), .A2(n12091), .B1(n13520), .B2(n12090), 
        .C1(n12089), .C2(n13522), .ZN(P3_U3271) );
  INV_X1 U14677 ( .A(n12092), .ZN(n13154) );
  NAND2_X1 U14678 ( .A1(n13154), .A2(n12093), .ZN(n12272) );
  INV_X1 U14679 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n13163) );
  NAND2_X1 U14680 ( .A1(n9854), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n12095) );
  NAND2_X1 U14681 ( .A1(n12266), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n12094) );
  OAI211_X1 U14682 ( .C1(n12269), .C2(n13163), .A(n12095), .B(n12094), .ZN(
        n12096) );
  INV_X1 U14683 ( .A(n12096), .ZN(n12097) );
  NAND2_X1 U14684 ( .A1(n12965), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n12098) );
  OAI21_X1 U14685 ( .B1(n13176), .B2(n12965), .A(n12098), .ZN(P3_U3520) );
  INV_X1 U14686 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13157) );
  NAND2_X1 U14687 ( .A1(n12266), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12100) );
  INV_X1 U14688 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13365) );
  OR2_X1 U14689 ( .A1(n9828), .A2(n13365), .ZN(n12099) );
  OAI211_X1 U14690 ( .C1(n13157), .C2(n12101), .A(n12100), .B(n12099), .ZN(
        n12102) );
  INV_X1 U14691 ( .A(n12102), .ZN(n12103) );
  NAND2_X1 U14692 ( .A1(n12965), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(n12104) );
  OAI21_X1 U14693 ( .B1(n13153), .B2(n12965), .A(n12104), .ZN(P3_U3522) );
  INV_X1 U14694 ( .A(n12134), .ZN(n12107) );
  AOI21_X1 U14695 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14169), .A(n12105), 
        .ZN(n12106) );
  OAI21_X1 U14696 ( .B1(n12107), .B2(n6438), .A(n12106), .ZN(P2_U3304) );
  OAI211_X1 U14697 ( .C1(n12110), .C2(n15536), .A(n12109), .B(n12108), .ZN(
        n12111) );
  AOI21_X1 U14698 ( .B1(n15541), .B2(n12112), .A(n12111), .ZN(n12115) );
  NAND2_X1 U14699 ( .A1(n15567), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n12113) );
  OAI21_X1 U14700 ( .B1(n12115), .B2(n15567), .A(n12113), .ZN(P2_U3509) );
  NAND2_X1 U14701 ( .A1(n15559), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n12114) );
  OAI21_X1 U14702 ( .B1(n12115), .B2(n15559), .A(n12114), .ZN(P2_U3460) );
  NAND3_X1 U14703 ( .A1(n12128), .A2(n11357), .A3(n12116), .ZN(n12117) );
  AND2_X1 U14704 ( .A1(n11247), .A2(n12117), .ZN(n12118) );
  OAI222_X1 U14705 ( .A1(n13930), .A2(n12120), .B1(n13932), .B2(n12119), .C1(
        n13951), .C2(n12118), .ZN(n15538) );
  INV_X1 U14706 ( .A(n15538), .ZN(n12133) );
  INV_X1 U14707 ( .A(n13979), .ZN(n13991) );
  OAI22_X1 U14708 ( .A1(n13987), .A2(n7899), .B1(n12121), .B2(n13956), .ZN(
        n12125) );
  INV_X1 U14709 ( .A(n13995), .ZN(n13868) );
  OAI211_X1 U14710 ( .C1(n12123), .C2(n15537), .A(n12569), .B(n12122), .ZN(
        n15535) );
  NOR2_X1 U14711 ( .A1(n13868), .A2(n15535), .ZN(n12124) );
  AOI211_X1 U14712 ( .C1(n13991), .C2(n12126), .A(n12125), .B(n12124), .ZN(
        n12132) );
  OAI21_X1 U14713 ( .B1(n12129), .B2(n12128), .A(n12127), .ZN(n15540) );
  NAND2_X1 U14714 ( .A1(n12130), .A2(n15540), .ZN(n12131) );
  OAI211_X1 U14715 ( .C1(n13909), .C2(n12133), .A(n12132), .B(n12131), .ZN(
        P2_U3263) );
  NAND2_X1 U14716 ( .A1(n12134), .A2(n15178), .ZN(n12135) );
  OAI211_X1 U14717 ( .C1(n12136), .C2(n15174), .A(n12135), .B(n14560), .ZN(
        P1_U3332) );
  MUX2_X1 U14718 ( .A(n12138), .B(n12837), .S(n12137), .Z(n12140) );
  XNOR2_X1 U14719 ( .A(n12140), .B(n12139), .ZN(n12148) );
  AOI21_X1 U14720 ( .B1(n12741), .B2(n12837), .A(n12141), .ZN(n12146) );
  NAND2_X1 U14721 ( .A1(n12720), .A2(n12842), .ZN(n12145) );
  INV_X1 U14722 ( .A(n12200), .ZN(n12142) );
  NAND2_X1 U14723 ( .A1(n12747), .A2(n12142), .ZN(n12144) );
  NAND2_X1 U14724 ( .A1(n12735), .A2(n12975), .ZN(n12143) );
  NAND4_X1 U14725 ( .A1(n12146), .A2(n12145), .A3(n12144), .A4(n12143), .ZN(
        n12147) );
  AOI21_X1 U14726 ( .B1(n12148), .B2(n12730), .A(n12147), .ZN(n12149) );
  INV_X1 U14727 ( .A(n12149), .ZN(P3_U3161) );
  XNOR2_X1 U14728 ( .A(n12150), .B(n12851), .ZN(n12234) );
  NAND2_X1 U14729 ( .A1(n11797), .A2(n12151), .ZN(n12153) );
  INV_X1 U14730 ( .A(n12851), .ZN(n12152) );
  NAND2_X1 U14731 ( .A1(n12153), .A2(n12152), .ZN(n12236) );
  OAI211_X1 U14732 ( .C1(n12153), .C2(n12152), .A(n12236), .B(n10349), .ZN(
        n12155) );
  AOI22_X1 U14733 ( .A1(n15595), .A2(n12975), .B1(n12973), .B2(n15597), .ZN(
        n12154) );
  NAND2_X1 U14734 ( .A1(n12155), .A2(n12154), .ZN(n12230) );
  MUX2_X1 U14735 ( .A(n12230), .B(P3_REG2_REG_10__SCAN_IN), .S(n15610), .Z(
        n12158) );
  OAI22_X1 U14736 ( .A1(n13340), .A2(n12852), .B1(n12156), .B2(n15577), .ZN(
        n12157) );
  NOR2_X1 U14737 ( .A1(n12158), .A2(n12157), .ZN(n12159) );
  OAI21_X1 U14738 ( .B1(n12234), .B2(n13363), .A(n12159), .ZN(P3_U3223) );
  XNOR2_X1 U14739 ( .A(n12160), .B(n12161), .ZN(n14100) );
  INV_X1 U14740 ( .A(n14100), .ZN(n12178) );
  INV_X1 U14741 ( .A(n12161), .ZN(n12163) );
  NAND3_X1 U14742 ( .A1(n12164), .A2(n12163), .A3(n12162), .ZN(n12165) );
  AND2_X1 U14743 ( .A1(n12166), .A2(n12165), .ZN(n12167) );
  OAI222_X1 U14744 ( .A1(n13932), .A2(n12295), .B1(n13930), .B2(n12168), .C1(
        n13951), .C2(n12167), .ZN(n14098) );
  NAND2_X1 U14745 ( .A1(n14098), .A2(n13987), .ZN(n12177) );
  INV_X1 U14746 ( .A(n12281), .ZN(n12169) );
  AOI211_X1 U14747 ( .C1(n12171), .C2(n12170), .A(n13974), .B(n12169), .ZN(
        n14099) );
  NOR2_X1 U14748 ( .A1(n14161), .A2(n13979), .ZN(n12175) );
  OAI22_X1 U14749 ( .A1(n13987), .A2(n12173), .B1(n12172), .B2(n13956), .ZN(
        n12174) );
  AOI211_X1 U14750 ( .C1(n14099), .C2(n13995), .A(n12175), .B(n12174), .ZN(
        n12176) );
  OAI211_X1 U14751 ( .C1(n12178), .C2(n13983), .A(n12177), .B(n12176), .ZN(
        P2_U3254) );
  XNOR2_X1 U14752 ( .A(n12179), .B(n12183), .ZN(n15387) );
  AOI21_X1 U14753 ( .B1(n11686), .B2(n14424), .A(n15365), .ZN(n12180) );
  NAND2_X1 U14754 ( .A1(n12180), .A2(n12222), .ZN(n15383) );
  INV_X1 U14755 ( .A(n14424), .ZN(n12181) );
  OAI22_X1 U14756 ( .A1(n15383), .A2(n14860), .B1(n12181), .B2(n15057), .ZN(
        n12188) );
  XNOR2_X1 U14757 ( .A(n12182), .B(n12183), .ZN(n12184) );
  NAND2_X1 U14758 ( .A1(n12184), .A2(n15024), .ZN(n15385) );
  OAI211_X1 U14759 ( .C1(n15055), .C2(n12185), .A(n15385), .B(n15384), .ZN(
        n12186) );
  MUX2_X1 U14760 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n12186), .S(n15049), .Z(
        n12187) );
  AOI211_X1 U14761 ( .C1(n14865), .C2(n15387), .A(n12188), .B(n12187), .ZN(
        n12189) );
  INV_X1 U14762 ( .A(n12189), .ZN(P1_U3285) );
  INV_X1 U14763 ( .A(n12190), .ZN(n12191) );
  AOI21_X1 U14764 ( .B1(n12193), .B2(n12192), .A(n12191), .ZN(n12199) );
  NAND2_X1 U14765 ( .A1(n13967), .A2(n13968), .ZN(n12194) );
  OAI21_X1 U14766 ( .B1(n12195), .B2(n13930), .A(n12194), .ZN(n12278) );
  AOI22_X1 U14767 ( .A1(n13643), .A2(n12278), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12196) );
  OAI21_X1 U14768 ( .B1(n13645), .B2(n12283), .A(n12196), .ZN(n12197) );
  AOI21_X1 U14769 ( .B1(n14154), .B2(n13647), .A(n12197), .ZN(n12198) );
  OAI21_X1 U14770 ( .B1(n12199), .B2(n13649), .A(n12198), .ZN(P2_U3196) );
  OAI22_X1 U14771 ( .A1(n13340), .A2(n12201), .B1(n12200), .B2(n15577), .ZN(
        n12204) );
  MUX2_X1 U14772 ( .A(n12202), .B(P3_REG2_REG_8__SCAN_IN), .S(n15610), .Z(
        n12203) );
  AOI211_X1 U14773 ( .C1(n15605), .C2(n12205), .A(n12204), .B(n12203), .ZN(
        n12206) );
  INV_X1 U14774 ( .A(n12206), .ZN(P3_U3225) );
  INV_X1 U14775 ( .A(n12207), .ZN(n12211) );
  OAI222_X1 U14776 ( .A1(n15185), .A2(n12209), .B1(n15188), .B2(n12211), .C1(
        n6428), .C2(n12208), .ZN(P1_U3331) );
  OAI222_X1 U14777 ( .A1(n14184), .A2(n12212), .B1(n6438), .B2(n12211), .C1(
        P2_U3088), .C2(n12210), .ZN(P2_U3303) );
  XOR2_X1 U14778 ( .A(n12213), .B(n14592), .Z(n15389) );
  NAND2_X1 U14779 ( .A1(n12215), .A2(n12214), .ZN(n12216) );
  NOR2_X1 U14780 ( .A1(n12216), .A2(n14592), .ZN(n15043) );
  AOI21_X1 U14781 ( .B1(n14592), .B2(n12216), .A(n15043), .ZN(n12217) );
  NOR2_X1 U14782 ( .A1(n12217), .A2(n15325), .ZN(n15393) );
  OR2_X1 U14783 ( .A1(n14439), .A2(n15052), .ZN(n12219) );
  NAND2_X1 U14784 ( .A1(n14648), .A2(n15223), .ZN(n12218) );
  NAND2_X1 U14785 ( .A1(n12219), .A2(n12218), .ZN(n15390) );
  NOR2_X1 U14786 ( .A1(n15393), .A2(n15390), .ZN(n12220) );
  MUX2_X1 U14787 ( .A(n12221), .B(n12220), .S(n15049), .Z(n12227) );
  NAND2_X1 U14788 ( .A1(n12222), .A2(n14428), .ZN(n12223) );
  NAND2_X1 U14789 ( .A1(n12223), .A2(n15333), .ZN(n12224) );
  NOR2_X1 U14790 ( .A1(n15051), .A2(n12224), .ZN(n15391) );
  OAI22_X1 U14791 ( .A1(n15057), .A2(n7493), .B1(n12260), .B2(n15055), .ZN(
        n12225) );
  AOI21_X1 U14792 ( .B1(n15391), .B2(n15235), .A(n12225), .ZN(n12226) );
  OAI211_X1 U14793 ( .C1(n14952), .C2(n15389), .A(n12227), .B(n12226), .ZN(
        P1_U3284) );
  INV_X1 U14794 ( .A(n12852), .ZN(n12232) );
  MUX2_X1 U14795 ( .A(n12230), .B(P3_REG1_REG_10__SCAN_IN), .S(n7202), .Z(
        n12228) );
  AOI21_X1 U14796 ( .B1(n13416), .B2(n12232), .A(n12228), .ZN(n12229) );
  OAI21_X1 U14797 ( .B1(n12234), .B2(n13418), .A(n12229), .ZN(P3_U3469) );
  MUX2_X1 U14798 ( .A(n12230), .B(P3_REG0_REG_10__SCAN_IN), .S(n15643), .Z(
        n12231) );
  AOI21_X1 U14799 ( .B1(n13493), .B2(n12232), .A(n12231), .ZN(n12233) );
  OAI21_X1 U14800 ( .B1(n12234), .B2(n13495), .A(n12233), .ZN(P3_U3420) );
  INV_X1 U14801 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n12239) );
  NAND2_X1 U14802 ( .A1(n12236), .A2(n12235), .ZN(n12237) );
  XNOR2_X1 U14803 ( .A(n12237), .B(n12858), .ZN(n12238) );
  AOI222_X1 U14804 ( .A1(n10349), .A2(n12238), .B1(n12972), .B2(n15597), .C1(
        n12974), .C2(n15595), .ZN(n12250) );
  MUX2_X1 U14805 ( .A(n12239), .B(n12250), .S(n15645), .Z(n12244) );
  OAI21_X1 U14806 ( .B1(n12241), .B2(n12858), .A(n12240), .ZN(n12249) );
  INV_X1 U14807 ( .A(n13495), .ZN(n12242) );
  NAND2_X1 U14808 ( .A1(n12249), .A2(n12242), .ZN(n12243) );
  OAI211_X1 U14809 ( .C1(n13443), .C2(n12252), .A(n12244), .B(n12243), .ZN(
        P3_U3423) );
  MUX2_X1 U14810 ( .A(n12245), .B(n12250), .S(n15652), .Z(n12248) );
  INV_X1 U14811 ( .A(n13418), .ZN(n12246) );
  NAND2_X1 U14812 ( .A1(n12249), .A2(n12246), .ZN(n12247) );
  OAI211_X1 U14813 ( .C1(n13382), .C2(n12252), .A(n12248), .B(n12247), .ZN(
        P3_U3470) );
  INV_X1 U14814 ( .A(n12249), .ZN(n12256) );
  MUX2_X1 U14815 ( .A(n12251), .B(n12250), .S(n15608), .Z(n12255) );
  INV_X1 U14816 ( .A(n12252), .ZN(n12374) );
  INV_X1 U14817 ( .A(n12372), .ZN(n12253) );
  AOI22_X1 U14818 ( .A1(n13347), .A2(n12374), .B1(n15604), .B2(n12253), .ZN(
        n12254) );
  OAI211_X1 U14819 ( .C1(n13363), .C2(n12256), .A(n12255), .B(n12254), .ZN(
        P3_U3222) );
  AND2_X1 U14820 ( .A1(n14428), .A2(n15400), .ZN(n15392) );
  INV_X1 U14821 ( .A(n15392), .ZN(n12265) );
  OAI211_X1 U14822 ( .C1(n12259), .C2(n12258), .A(n12257), .B(n14370), .ZN(
        n12264) );
  NOR2_X1 U14823 ( .A1(n14353), .A2(n12260), .ZN(n12261) );
  AOI211_X1 U14824 ( .C1(n14368), .C2(n15390), .A(n12262), .B(n12261), .ZN(
        n12263) );
  OAI211_X1 U14825 ( .C1(n14308), .C2(n12265), .A(n12264), .B(n12263), .ZN(
        P1_U3231) );
  INV_X1 U14826 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n13161) );
  NAND2_X1 U14827 ( .A1(n12266), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n12268) );
  NAND2_X1 U14828 ( .A1(n9854), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12267) );
  OAI211_X1 U14829 ( .C1(n13161), .C2(n12269), .A(n12268), .B(n12267), .ZN(
        n12270) );
  INV_X1 U14830 ( .A(n12270), .ZN(n12271) );
  AND2_X1 U14831 ( .A1(n12272), .A2(n12271), .ZN(n12764) );
  INV_X1 U14832 ( .A(n12764), .ZN(n12785) );
  NAND2_X1 U14833 ( .A1(n12785), .A2(P3_U3897), .ZN(n12273) );
  OAI21_X1 U14834 ( .B1(P3_U3897), .B2(n12274), .A(n12273), .ZN(P3_U3521) );
  XNOR2_X1 U14835 ( .A(n12275), .B(n12276), .ZN(n14095) );
  INV_X1 U14836 ( .A(n14095), .ZN(n12289) );
  XOR2_X1 U14837 ( .A(n12277), .B(n12276), .Z(n12280) );
  INV_X1 U14838 ( .A(n12278), .ZN(n12279) );
  OAI21_X1 U14839 ( .B1(n12280), .B2(n13951), .A(n12279), .ZN(n14093) );
  NAND2_X1 U14840 ( .A1(n14093), .A2(n13987), .ZN(n12288) );
  AOI211_X1 U14841 ( .C1(n14154), .C2(n12281), .A(n13974), .B(n12298), .ZN(
        n14094) );
  NOR2_X1 U14842 ( .A1(n12282), .A2(n13979), .ZN(n12286) );
  OAI22_X1 U14843 ( .A1(n13987), .A2(n12284), .B1(n12283), .B2(n13956), .ZN(
        n12285) );
  AOI211_X1 U14844 ( .C1(n14094), .C2(n13995), .A(n12286), .B(n12285), .ZN(
        n12287) );
  OAI211_X1 U14845 ( .C1(n13983), .C2(n12289), .A(n12288), .B(n12287), .ZN(
        P2_U3253) );
  INV_X1 U14846 ( .A(n12290), .ZN(n12291) );
  OAI222_X1 U14847 ( .A1(n12293), .A2(P3_U3151), .B1(n13522), .B2(n12292), 
        .C1(n13520), .C2(n12291), .ZN(P3_U3270) );
  XOR2_X1 U14848 ( .A(n12294), .B(n12304), .Z(n12297) );
  OR2_X1 U14849 ( .A1(n12295), .A2(n13930), .ZN(n12296) );
  OAI21_X1 U14850 ( .B1(n13659), .B2(n13932), .A(n12296), .ZN(n12312) );
  AOI21_X1 U14851 ( .B1(n12297), .B2(n13971), .A(n12312), .ZN(n14091) );
  INV_X1 U14852 ( .A(n12298), .ZN(n12300) );
  AOI211_X1 U14853 ( .C1(n14089), .C2(n12300), .A(n13974), .B(n13972), .ZN(
        n14088) );
  INV_X1 U14854 ( .A(n12314), .ZN(n12301) );
  AOI22_X1 U14855 ( .A1(n13909), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12301), 
        .B2(n13990), .ZN(n12302) );
  OAI21_X1 U14856 ( .B1(n12303), .B2(n13979), .A(n12302), .ZN(n12307) );
  XOR2_X1 U14857 ( .A(n12305), .B(n12304), .Z(n14092) );
  NOR2_X1 U14858 ( .A1(n14092), .A2(n13983), .ZN(n12306) );
  AOI211_X1 U14859 ( .C1(n14088), .C2(n13995), .A(n12307), .B(n12306), .ZN(
        n12308) );
  OAI21_X1 U14860 ( .B1(n13909), .B2(n14091), .A(n12308), .ZN(P2_U3252) );
  XNOR2_X1 U14861 ( .A(n12310), .B(n12309), .ZN(n12317) );
  AOI21_X1 U14862 ( .B1(n13643), .B2(n12312), .A(n12311), .ZN(n12313) );
  OAI21_X1 U14863 ( .B1(n13645), .B2(n12314), .A(n12313), .ZN(n12315) );
  AOI21_X1 U14864 ( .B1(n14089), .B2(n13647), .A(n12315), .ZN(n12316) );
  OAI21_X1 U14865 ( .B1(n12317), .B2(n13649), .A(n12316), .ZN(P2_U3206) );
  INV_X1 U14866 ( .A(n12318), .ZN(n12322) );
  OAI222_X1 U14867 ( .A1(n15185), .A2(n12320), .B1(n15188), .B2(n12322), .C1(
        P1_U3086), .C2(n12319), .ZN(P1_U3330) );
  OAI222_X1 U14868 ( .A1(n14184), .A2(n12323), .B1(n6438), .B2(n12322), .C1(
        P2_U3088), .C2(n12321), .ZN(P2_U3302) );
  XNOR2_X1 U14869 ( .A(n12324), .B(n12971), .ZN(n12325) );
  XNOR2_X1 U14870 ( .A(n12326), .B(n12325), .ZN(n12331) );
  AND2_X1 U14871 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12996) );
  NOR2_X1 U14872 ( .A1(n12733), .A2(n12383), .ZN(n12327) );
  AOI211_X1 U14873 ( .C1(n12735), .C2(n12970), .A(n12996), .B(n12327), .ZN(
        n12328) );
  OAI21_X1 U14874 ( .B1(n12379), .B2(n12662), .A(n12328), .ZN(n12329) );
  AOI21_X1 U14875 ( .B1(n13492), .B2(n12720), .A(n12329), .ZN(n12330) );
  OAI21_X1 U14876 ( .B1(n12331), .B2(n12749), .A(n12330), .ZN(P3_U3174) );
  XNOR2_X1 U14877 ( .A(n12332), .B(n12335), .ZN(n12362) );
  INV_X1 U14878 ( .A(n12663), .ZN(n12333) );
  AOI22_X1 U14879 ( .A1(n12665), .A2(n13347), .B1(n15604), .B2(n12333), .ZN(
        n12340) );
  XNOR2_X1 U14880 ( .A(n12334), .B(n12335), .ZN(n12336) );
  OAI222_X1 U14881 ( .A1(n15580), .A2(n13354), .B1(n15582), .B2(n12659), .C1(
        n12336), .C2(n15601), .ZN(n12359) );
  INV_X1 U14882 ( .A(n12359), .ZN(n12337) );
  MUX2_X1 U14883 ( .A(n12338), .B(n12337), .S(n15608), .Z(n12339) );
  OAI211_X1 U14884 ( .C1(n12362), .C2(n13363), .A(n12340), .B(n12339), .ZN(
        P3_U3221) );
  NOR2_X1 U14885 ( .A1(n12350), .A2(n12343), .ZN(n12344) );
  XNOR2_X1 U14886 ( .A(n12352), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n14744) );
  XNOR2_X1 U14887 ( .A(n14745), .B(n14744), .ZN(n12356) );
  NAND2_X1 U14888 ( .A1(n15299), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n12345) );
  NAND2_X1 U14889 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14281)
         );
  NAND2_X1 U14890 ( .A1(n12345), .A2(n14281), .ZN(n12346) );
  AOI21_X1 U14891 ( .B1(n14749), .B2(n14783), .A(n12346), .ZN(n12355) );
  OR2_X1 U14892 ( .A1(n12347), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n12348) );
  XNOR2_X1 U14893 ( .A(n12351), .B(n12350), .ZN(n15309) );
  NAND2_X1 U14894 ( .A1(n15309), .A2(n15308), .ZN(n15307) );
  XNOR2_X1 U14895 ( .A(n12352), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12353) );
  OAI211_X1 U14896 ( .C1(n6473), .C2(n12353), .A(n14751), .B(n15310), .ZN(
        n12354) );
  OAI211_X1 U14897 ( .C1(n12356), .C2(n15305), .A(n12355), .B(n12354), .ZN(
        P1_U3259) );
  MUX2_X1 U14898 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n12359), .S(n15652), .Z(
        n12357) );
  AOI21_X1 U14899 ( .B1(n13416), .B2(n12665), .A(n12357), .ZN(n12358) );
  OAI21_X1 U14900 ( .B1(n13418), .B2(n12362), .A(n12358), .ZN(P3_U3471) );
  MUX2_X1 U14901 ( .A(P3_REG0_REG_12__SCAN_IN), .B(n12359), .S(n15645), .Z(
        n12360) );
  AOI21_X1 U14902 ( .B1(n13493), .B2(n12665), .A(n12360), .ZN(n12361) );
  OAI21_X1 U14903 ( .B1(n13495), .B2(n12362), .A(n12361), .ZN(P3_U3426) );
  INV_X1 U14904 ( .A(n12363), .ZN(n12366) );
  INV_X1 U14905 ( .A(n12364), .ZN(n12365) );
  OR2_X1 U14906 ( .A1(n12364), .A2(n12363), .ZN(n12653) );
  OAI21_X1 U14907 ( .B1(n12366), .B2(n12365), .A(n12653), .ZN(n12367) );
  NOR2_X1 U14908 ( .A1(n12367), .A2(n12973), .ZN(n12655) );
  AOI21_X1 U14909 ( .B1(n12973), .B2(n12367), .A(n12655), .ZN(n12376) );
  OAI21_X1 U14910 ( .B1(n12733), .B2(n12369), .A(n12368), .ZN(n12370) );
  AOI21_X1 U14911 ( .B1(n12735), .B2(n12972), .A(n12370), .ZN(n12371) );
  OAI21_X1 U14912 ( .B1(n12372), .B2(n12662), .A(n12371), .ZN(n12373) );
  AOI21_X1 U14913 ( .B1(n12374), .B2(n12720), .A(n12373), .ZN(n12375) );
  OAI21_X1 U14914 ( .B1(n12376), .B2(n12749), .A(n12375), .ZN(P3_U3176) );
  INV_X1 U14915 ( .A(n12377), .ZN(n12869) );
  OR2_X1 U14916 ( .A1(n12870), .A2(n12869), .ZN(n12867) );
  XOR2_X1 U14917 ( .A(n12378), .B(n12867), .Z(n13496) );
  INV_X1 U14918 ( .A(n12379), .ZN(n12380) );
  AOI22_X1 U14919 ( .A1(n13492), .A2(n13347), .B1(n15604), .B2(n12380), .ZN(
        n12387) );
  XNOR2_X1 U14920 ( .A(n12381), .B(n12867), .ZN(n12382) );
  OAI222_X1 U14921 ( .A1(n15580), .A2(n13336), .B1(n15582), .B2(n12383), .C1(
        n12382), .C2(n15601), .ZN(n13490) );
  INV_X1 U14922 ( .A(n13490), .ZN(n12384) );
  MUX2_X1 U14923 ( .A(n12385), .B(n12384), .S(n15608), .Z(n12386) );
  OAI211_X1 U14924 ( .C1(n13496), .C2(n13363), .A(n12387), .B(n12386), .ZN(
        P3_U3220) );
  XNOR2_X1 U14925 ( .A(n12474), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n12470) );
  OAI21_X1 U14926 ( .B1(n12389), .B2(P2_REG1_REG_15__SCAN_IN), .A(n15471), 
        .ZN(n12402) );
  NOR2_X1 U14927 ( .A1(n12390), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13642) );
  NOR2_X1 U14928 ( .A1(n15522), .A2(n7084), .ZN(n12391) );
  AOI211_X1 U14929 ( .C1(n15519), .C2(n13685), .A(n13642), .B(n12391), .ZN(
        n12401) );
  NAND2_X1 U14930 ( .A1(n12392), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12393) );
  NAND2_X1 U14931 ( .A1(n12394), .A2(n12393), .ZN(n12396) );
  XNOR2_X1 U14932 ( .A(n12396), .B(n12395), .ZN(n12476) );
  NAND2_X1 U14933 ( .A1(n12476), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n12475) );
  NAND2_X1 U14934 ( .A1(n12396), .A2(n12474), .ZN(n12397) );
  NAND2_X1 U14935 ( .A1(n12475), .A2(n12397), .ZN(n13674) );
  XNOR2_X1 U14936 ( .A(n13674), .B(n12398), .ZN(n12399) );
  NAND2_X1 U14937 ( .A1(n12399), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n13676) );
  OAI211_X1 U14938 ( .C1(n12399), .C2(P2_REG2_REG_15__SCAN_IN), .A(n13676), 
        .B(n15508), .ZN(n12400) );
  OAI211_X1 U14939 ( .C1(n12402), .C2(n13683), .A(n12401), .B(n12400), .ZN(
        P2_U3229) );
  INV_X1 U14940 ( .A(n12403), .ZN(n12467) );
  OAI222_X1 U14941 ( .A1(n14184), .A2(n12583), .B1(P2_U3088), .B2(n12404), 
        .C1(n6438), .C2(n12467), .ZN(P2_U3297) );
  OAI222_X1 U14942 ( .A1(n15185), .A2(n12406), .B1(n15188), .B2(n12405), .C1(
        n14958), .C2(P1_U3086), .ZN(P1_U3336) );
  OR2_X1 U14943 ( .A1(n14438), .A2(n15053), .ZN(n12408) );
  XNOR2_X1 U14944 ( .A(n15230), .B(n15027), .ZN(n15219) );
  INV_X1 U14945 ( .A(n15027), .ZN(n14445) );
  OR2_X1 U14946 ( .A1(n15230), .A2(n14445), .ZN(n15020) );
  OR2_X1 U14947 ( .A1(n15036), .A2(n14443), .ZN(n12410) );
  AND2_X1 U14948 ( .A1(n15020), .A2(n12410), .ZN(n12413) );
  INV_X1 U14949 ( .A(n12410), .ZN(n12411) );
  XNOR2_X1 U14950 ( .A(n15036), .B(n15221), .ZN(n15019) );
  OR2_X1 U14951 ( .A1(n15151), .A2(n14324), .ZN(n14442) );
  XNOR2_X1 U14952 ( .A(n15142), .B(n14956), .ZN(n14972) );
  NAND2_X1 U14953 ( .A1(n15142), .A2(n14956), .ZN(n12414) );
  OR2_X1 U14954 ( .A1(n15137), .A2(n14974), .ZN(n12415) );
  NAND2_X1 U14955 ( .A1(n15137), .A2(n14974), .ZN(n12416) );
  NAND2_X1 U14956 ( .A1(n15131), .A2(n14957), .ZN(n14496) );
  NAND2_X1 U14957 ( .A1(n14492), .A2(n14496), .ZN(n14942) );
  INV_X1 U14958 ( .A(n14942), .ZN(n12417) );
  INV_X1 U14959 ( .A(n14921), .ZN(n12418) );
  XNOR2_X1 U14960 ( .A(n15122), .B(n14923), .ZN(n14899) );
  OR2_X1 U14961 ( .A1(n15122), .A2(n14923), .ZN(n12419) );
  INV_X1 U14962 ( .A(n14870), .ZN(n14901) );
  NAND2_X1 U14963 ( .A1(n14878), .A2(n14642), .ZN(n12421) );
  XNOR2_X2 U14964 ( .A(n15104), .B(n14871), .ZN(n14863) );
  INV_X1 U14965 ( .A(n14871), .ZN(n12423) );
  NAND2_X1 U14966 ( .A1(n6476), .A2(n12424), .ZN(n12430) );
  INV_X1 U14967 ( .A(n14838), .ZN(n14844) );
  OAI21_X1 U14968 ( .B1(n14844), .B2(n14641), .A(n14640), .ZN(n12426) );
  NOR2_X1 U14969 ( .A1(n14640), .A2(n14641), .ZN(n12425) );
  AOI22_X1 U14970 ( .A1(n12426), .A2(n14829), .B1(n12425), .B2(n14838), .ZN(
        n12427) );
  OAI21_X1 U14971 ( .B1(n14811), .B2(n14639), .A(n12427), .ZN(n12428) );
  INV_X1 U14972 ( .A(n12428), .ZN(n12429) );
  INV_X1 U14973 ( .A(n12503), .ZN(n12432) );
  OAI21_X1 U14974 ( .B1(n14607), .B2(n6546), .A(n12432), .ZN(n12434) );
  AOI21_X2 U14975 ( .B1(n12434), .B2(n15024), .A(n12433), .ZN(n15084) );
  INV_X1 U14976 ( .A(n12593), .ZN(n12436) );
  AOI211_X1 U14977 ( .C1(n15082), .C2(n12435), .A(n15365), .B(n12436), .ZN(
        n15081) );
  AOI22_X1 U14978 ( .A1(n12437), .A2(n15331), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15340), .ZN(n12438) );
  OAI21_X1 U14979 ( .B1(n12439), .B2(n15057), .A(n12438), .ZN(n12465) );
  NAND2_X1 U14980 ( .A1(n12440), .A2(n14593), .ZN(n12442) );
  INV_X1 U14981 ( .A(n15053), .ZN(n15224) );
  OR2_X1 U14982 ( .A1(n14438), .A2(n15224), .ZN(n12441) );
  NAND2_X1 U14983 ( .A1(n12442), .A2(n12441), .ZN(n15217) );
  INV_X1 U14984 ( .A(n15219), .ZN(n15218) );
  NAND2_X1 U14985 ( .A1(n15217), .A2(n15218), .ZN(n12444) );
  OR2_X1 U14986 ( .A1(n15230), .A2(n15027), .ZN(n12443) );
  NAND2_X1 U14987 ( .A1(n12444), .A2(n12443), .ZN(n15018) );
  INV_X1 U14988 ( .A(n15019), .ZN(n15022) );
  OR2_X1 U14989 ( .A1(n15036), .A2(n15221), .ZN(n12445) );
  NAND2_X1 U14990 ( .A1(n15151), .A2(n15026), .ZN(n12447) );
  NAND2_X1 U14991 ( .A1(n15014), .A2(n12447), .ZN(n14996) );
  OR2_X1 U14992 ( .A1(n15146), .A2(n14647), .ZN(n12449) );
  OR2_X1 U14993 ( .A1(n15142), .A2(n14987), .ZN(n12450) );
  INV_X1 U14994 ( .A(n15137), .ZN(n12451) );
  INV_X1 U14995 ( .A(n14974), .ZN(n14646) );
  NAND2_X1 U14996 ( .A1(n15137), .A2(n14646), .ZN(n14596) );
  INV_X1 U14997 ( .A(n14957), .ZN(n14645) );
  AND2_X1 U14998 ( .A1(n15131), .A2(n14645), .ZN(n12453) );
  OR2_X1 U14999 ( .A1(n15131), .A2(n14645), .ZN(n12452) );
  OR2_X1 U15000 ( .A1(n15128), .A2(n14644), .ZN(n12454) );
  INV_X1 U15001 ( .A(n14899), .ZN(n14909) );
  NAND2_X1 U15002 ( .A1(n15122), .A2(n14643), .ZN(n14476) );
  INV_X1 U15003 ( .A(n14880), .ZN(n14601) );
  NAND2_X1 U15004 ( .A1(n14879), .A2(n14601), .ZN(n12456) );
  NAND2_X1 U15005 ( .A1(n14878), .A2(n14241), .ZN(n12455) );
  NAND2_X1 U15006 ( .A1(n15104), .A2(n14871), .ZN(n12457) );
  XNOR2_X2 U15007 ( .A(n14838), .B(n14641), .ZN(n14846) );
  OAI22_X1 U15008 ( .A1(n15087), .A2(n14639), .B1(n14640), .B2(n14829), .ZN(
        n12461) );
  NAND2_X1 U15009 ( .A1(n14829), .A2(n14640), .ZN(n14813) );
  NAND2_X1 U15010 ( .A1(n14813), .A2(n14522), .ZN(n12459) );
  AND2_X1 U15011 ( .A1(n14639), .A2(n14640), .ZN(n12458) );
  AOI22_X1 U15012 ( .A1(n15087), .A2(n12459), .B1(n12458), .B2(n14829), .ZN(
        n12460) );
  INV_X1 U15013 ( .A(n12463), .ZN(n15085) );
  NOR2_X1 U15014 ( .A1(n15085), .A2(n14952), .ZN(n12464) );
  OAI21_X1 U15015 ( .B1(n15084), .B2(n15340), .A(n12466), .ZN(P1_U3266) );
  OAI222_X1 U15016 ( .A1(n15174), .A2(n12584), .B1(P1_U3086), .B2(n12468), 
        .C1(n15188), .C2(n12467), .ZN(P1_U3325) );
  NAND2_X1 U15017 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n13529)
         );
  OAI21_X1 U15018 ( .B1(n15522), .B2(n15280), .A(n13529), .ZN(n12473) );
  AOI211_X1 U15019 ( .C1(n12471), .C2(n12470), .A(n15513), .B(n12469), .ZN(
        n12472) );
  AOI211_X1 U15020 ( .C1(n15519), .C2(n12474), .A(n12473), .B(n12472), .ZN(
        n12478) );
  OAI211_X1 U15021 ( .C1(n12476), .C2(P2_REG2_REG_14__SCAN_IN), .A(n12475), 
        .B(n15508), .ZN(n12477) );
  NAND2_X1 U15022 ( .A1(n12478), .A2(n12477), .ZN(P2_U3228) );
  INV_X1 U15023 ( .A(n12479), .ZN(n12670) );
  XNOR2_X1 U15024 ( .A(n13376), .B(n12487), .ZN(n12480) );
  AOI21_X1 U15025 ( .B1(n12480), .B2(n12963), .A(n12481), .ZN(n12669) );
  INV_X1 U15026 ( .A(n12481), .ZN(n12482) );
  XNOR2_X1 U15027 ( .A(n12483), .B(n12487), .ZN(n12484) );
  NOR2_X1 U15028 ( .A1(n12484), .A2(n12962), .ZN(n12485) );
  AOI21_X1 U15029 ( .B1(n12484), .B2(n12962), .A(n12485), .ZN(n12729) );
  NAND2_X1 U15030 ( .A1(n12728), .A2(n12729), .ZN(n12727) );
  INV_X1 U15031 ( .A(n12485), .ZN(n12486) );
  NOR2_X1 U15032 ( .A1(n12488), .A2(n12961), .ZN(n12489) );
  AOI21_X1 U15033 ( .B1(n12488), .B2(n12961), .A(n12489), .ZN(n12612) );
  AND2_X1 U15034 ( .A1(n14182), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12490) );
  NAND2_X1 U15035 ( .A1(n15184), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12492) );
  XNOR2_X1 U15036 ( .A(n14179), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n12493) );
  XNOR2_X1 U15037 ( .A(n12538), .B(n12493), .ZN(n13510) );
  NAND2_X1 U15038 ( .A1(n13510), .A2(n12758), .ZN(n12495) );
  OR2_X1 U15039 ( .A1(n12761), .A2(n13512), .ZN(n12494) );
  XNOR2_X1 U15040 ( .A(n13173), .B(n12496), .ZN(n12497) );
  NOR2_X1 U15041 ( .A1(n13176), .A2(n12743), .ZN(n12500) );
  AOI22_X1 U15042 ( .A1(n13181), .A2(n12747), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12498) );
  OAI21_X1 U15043 ( .B1(n13193), .B2(n12733), .A(n12498), .ZN(n12499) );
  AOI211_X1 U15044 ( .C1(n13427), .C2(n12720), .A(n12500), .B(n12499), .ZN(
        n12501) );
  OAI21_X1 U15045 ( .B1(n12502), .B2(n12749), .A(n12501), .ZN(P3_U3160) );
  NAND2_X1 U15046 ( .A1(n15049), .A2(n15024), .ZN(n12536) );
  INV_X1 U15047 ( .A(n12596), .ZN(n12505) );
  NAND2_X1 U15048 ( .A1(n14637), .A2(n15223), .ZN(n15068) );
  NAND2_X1 U15049 ( .A1(n14550), .A2(n15329), .ZN(n12520) );
  INV_X1 U15050 ( .A(n12506), .ZN(n12516) );
  INV_X1 U15051 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n12507) );
  NOR2_X1 U15052 ( .A1(n9288), .A2(n12507), .ZN(n12513) );
  INV_X1 U15053 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14797) );
  NOR2_X1 U15054 ( .A1(n12508), .A2(n14797), .ZN(n12512) );
  INV_X1 U15055 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n12509) );
  NOR2_X1 U15056 ( .A1(n12510), .A2(n12509), .ZN(n12511) );
  OR3_X1 U15057 ( .A1(n12513), .A2(n12512), .A3(n12511), .ZN(n14635) );
  NAND2_X1 U15058 ( .A1(n14635), .A2(n12514), .ZN(n15069) );
  AOI21_X1 U15059 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n15055), .A(n12516), 
        .ZN(n12515) );
  AOI21_X1 U15060 ( .B1(n12516), .B2(n15069), .A(n12515), .ZN(n12517) );
  AOI21_X1 U15061 ( .B1(n12518), .B2(n15331), .A(n12517), .ZN(n12519) );
  OAI211_X1 U15062 ( .C1(n15340), .C2(n15068), .A(n12520), .B(n12519), .ZN(
        n12521) );
  AOI21_X1 U15063 ( .B1(n15072), .B2(n15235), .A(n12521), .ZN(n12535) );
  NAND2_X1 U15064 ( .A1(n14610), .A2(n12526), .ZN(n12522) );
  NOR2_X1 U15065 ( .A1(n12602), .A2(n12522), .ZN(n12529) );
  OR2_X1 U15066 ( .A1(n15082), .A2(n14638), .ZN(n12601) );
  AND2_X1 U15067 ( .A1(n12523), .A2(n12601), .ZN(n12531) );
  INV_X1 U15068 ( .A(n12531), .ZN(n12524) );
  NAND2_X1 U15069 ( .A1(n12524), .A2(n12526), .ZN(n12525) );
  MUX2_X1 U15070 ( .A(n12526), .B(n12525), .S(n14610), .Z(n12527) );
  NOR2_X1 U15071 ( .A1(n12529), .A2(n12528), .ZN(n12533) );
  INV_X1 U15072 ( .A(n14610), .ZN(n12530) );
  NAND3_X1 U15073 ( .A1(n12602), .A2(n12531), .A3(n12530), .ZN(n12532) );
  NAND2_X1 U15074 ( .A1(n15067), .A2(n14865), .ZN(n12534) );
  OAI211_X1 U15075 ( .C1(n15073), .C2(n12536), .A(n12535), .B(n12534), .ZN(
        P1_U3356) );
  AND2_X1 U15076 ( .A1(n12609), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12537) );
  NAND2_X1 U15077 ( .A1(n14179), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12539) );
  XNOR2_X1 U15078 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12579) );
  XNOR2_X1 U15079 ( .A(n12581), .B(n12579), .ZN(n13506) );
  NAND2_X1 U15080 ( .A1(n13506), .A2(n12758), .ZN(n12542) );
  OR2_X1 U15081 ( .A1(n12761), .A2(n13509), .ZN(n12541) );
  NAND2_X1 U15082 ( .A1(n12556), .A2(n13176), .ZN(n12943) );
  INV_X1 U15083 ( .A(n12937), .ZN(n12543) );
  NOR2_X1 U15084 ( .A1(n12796), .A2(n12545), .ZN(n12546) );
  XOR2_X1 U15085 ( .A(n12784), .B(n12546), .Z(n13170) );
  INV_X1 U15086 ( .A(n13178), .ZN(n12547) );
  INV_X1 U15087 ( .A(n12551), .ZN(n12960) );
  INV_X1 U15088 ( .A(n13427), .ZN(n12549) );
  NOR4_X1 U15089 ( .A1(n12784), .A2(n12549), .A3(n12551), .A4(n15601), .ZN(
        n12553) );
  NAND2_X1 U15090 ( .A1(n12954), .A2(P3_B_REG_SCAN_IN), .ZN(n12550) );
  NAND2_X1 U15091 ( .A1(n15597), .A2(n12550), .ZN(n13152) );
  OAI22_X1 U15092 ( .A1(n12551), .A2(n15582), .B1(n12764), .B2(n13152), .ZN(
        n12552) );
  INV_X1 U15093 ( .A(n12556), .ZN(n12557) );
  NOR2_X1 U15094 ( .A1(n12557), .A2(n15638), .ZN(n13166) );
  NAND2_X1 U15095 ( .A1(n12561), .A2(n12560), .ZN(P3_U3456) );
  OAI222_X1 U15096 ( .A1(n14184), .A2(n12564), .B1(n6438), .B2(n12563), .C1(
        n12562), .C2(P2_U3088), .ZN(P2_U3307) );
  OAI222_X1 U15097 ( .A1(n15185), .A2(n12566), .B1(n15188), .B2(n12565), .C1(
        n14544), .C2(n6428), .ZN(P1_U3334) );
  OAI222_X1 U15098 ( .A1(n13146), .A2(P3_U3151), .B1(n13520), .B2(n12568), 
        .C1(n12567), .C2(n13522), .ZN(P3_U3276) );
  NAND2_X1 U15099 ( .A1(n12571), .A2(P2_B_REG_SCAN_IN), .ZN(n12572) );
  NAND2_X1 U15100 ( .A1(n13968), .A2(n12572), .ZN(n13721) );
  INV_X1 U15101 ( .A(n13721), .ZN(n12573) );
  NAND2_X1 U15102 ( .A1(n13651), .A2(n12573), .ZN(n14000) );
  OR2_X1 U15103 ( .A1(n15564), .A2(n8694), .ZN(n12574) );
  AOI21_X1 U15104 ( .B1(n14096), .B2(n12577), .A(n12576), .ZN(n12578) );
  INV_X1 U15105 ( .A(n12578), .ZN(P2_U3530) );
  INV_X1 U15106 ( .A(SI_30_), .ZN(n12760) );
  INV_X1 U15107 ( .A(n12579), .ZN(n12580) );
  NAND2_X1 U15108 ( .A1(n15182), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12582) );
  NAND2_X1 U15109 ( .A1(n12583), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U15110 ( .A1(n12584), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U15111 ( .A1(n12751), .A2(n12585), .ZN(n12752) );
  XNOR2_X1 U15112 ( .A(n12753), .B(n12752), .ZN(n12759) );
  INV_X1 U15113 ( .A(n12759), .ZN(n12586) );
  OAI222_X1 U15114 ( .A1(n13522), .A2(n12760), .B1(n13520), .B2(n12586), .C1(
        P3_U3151), .C2(n7790), .ZN(P3_U3265) );
  INV_X1 U15115 ( .A(n14605), .ZN(n12603) );
  NAND2_X1 U15116 ( .A1(n12603), .A2(n12587), .ZN(n12589) );
  OAI21_X1 U15117 ( .B1(n12503), .B2(n12589), .A(n12588), .ZN(n12590) );
  INV_X1 U15118 ( .A(n14548), .ZN(n14636) );
  NAND2_X1 U15119 ( .A1(n12593), .A2(n15077), .ZN(n12594) );
  NAND2_X1 U15120 ( .A1(n12594), .A2(n15333), .ZN(n12595) );
  NOR2_X1 U15121 ( .A1(n12596), .A2(n12595), .ZN(n15076) );
  NAND2_X1 U15122 ( .A1(n15077), .A2(n15329), .ZN(n12599) );
  AOI22_X1 U15123 ( .A1(n12597), .A2(n15331), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15340), .ZN(n12598) );
  NAND2_X1 U15124 ( .A1(n12599), .A2(n12598), .ZN(n12600) );
  AOI21_X1 U15125 ( .B1(n15076), .B2(n15235), .A(n12600), .ZN(n12607) );
  NAND2_X1 U15126 ( .A1(n12604), .A2(n12603), .ZN(n15074) );
  NAND2_X1 U15127 ( .A1(n12605), .A2(n14605), .ZN(n15075) );
  NAND3_X1 U15128 ( .A1(n15074), .A2(n14865), .A3(n15075), .ZN(n12606) );
  OAI211_X1 U15129 ( .C1(n15079), .C2(n15340), .A(n12607), .B(n12606), .ZN(
        P1_U3265) );
  INV_X1 U15130 ( .A(n14176), .ZN(n12608) );
  OAI222_X1 U15131 ( .A1(n15185), .A2(n12609), .B1(n15188), .B2(n12608), .C1(
        n14671), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI21_X1 U15132 ( .B1(n12612), .B2(n12610), .A(n12611), .ZN(n12613) );
  NAND2_X1 U15133 ( .A1(n12613), .A2(n12730), .ZN(n12617) );
  AOI22_X1 U15134 ( .A1(n13185), .A2(n12747), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12614) );
  OAI21_X1 U15135 ( .B1(n13212), .B2(n12733), .A(n12614), .ZN(n12615) );
  AOI21_X1 U15136 ( .B1(n12960), .B2(n12735), .A(n12615), .ZN(n12616) );
  OAI211_X1 U15137 ( .C1(n13187), .C2(n12744), .A(n12617), .B(n12616), .ZN(
        P3_U3154) );
  INV_X1 U15138 ( .A(n13487), .ZN(n12626) );
  OAI21_X1 U15139 ( .B1(n12620), .B2(n12619), .A(n12618), .ZN(n12621) );
  NAND2_X1 U15140 ( .A1(n12621), .A2(n12730), .ZN(n12625) );
  NAND2_X1 U15141 ( .A1(n12741), .A2(n12971), .ZN(n12622) );
  NAND2_X1 U15142 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13015)
         );
  OAI211_X1 U15143 ( .C1(n13355), .C2(n12743), .A(n12622), .B(n13015), .ZN(
        n12623) );
  AOI21_X1 U15144 ( .B1(n13346), .B2(n12747), .A(n12623), .ZN(n12624) );
  OAI211_X1 U15145 ( .C1(n12626), .C2(n12744), .A(n12625), .B(n12624), .ZN(
        P3_U3155) );
  INV_X1 U15146 ( .A(n12918), .ZN(n13444) );
  OAI21_X1 U15147 ( .B1(n13227), .B2(n12628), .A(n12627), .ZN(n12629) );
  NAND2_X1 U15148 ( .A1(n12629), .A2(n12730), .ZN(n12634) );
  INV_X1 U15149 ( .A(n12630), .ZN(n13242) );
  AOI22_X1 U15150 ( .A1(n12966), .A2(n12741), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12631) );
  OAI21_X1 U15151 ( .B1(n13242), .B2(n12662), .A(n12631), .ZN(n12632) );
  AOI21_X1 U15152 ( .B1(n12735), .B2(n12964), .A(n12632), .ZN(n12633) );
  OAI211_X1 U15153 ( .C1(n13444), .C2(n12744), .A(n12634), .B(n12633), .ZN(
        P3_U3156) );
  XNOR2_X1 U15154 ( .A(n12636), .B(n12635), .ZN(n12641) );
  NAND2_X1 U15155 ( .A1(n13294), .A2(n12735), .ZN(n12637) );
  NAND2_X1 U15156 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13145)
         );
  OAI211_X1 U15157 ( .C1(n13316), .C2(n12733), .A(n12637), .B(n13145), .ZN(
        n12639) );
  NOR2_X1 U15158 ( .A1(n13299), .A2(n12744), .ZN(n12638) );
  AOI211_X1 U15159 ( .C1(n13297), .C2(n12747), .A(n12639), .B(n12638), .ZN(
        n12640) );
  OAI21_X1 U15160 ( .B1(n12641), .B2(n12749), .A(n12640), .ZN(P3_U3159) );
  INV_X1 U15161 ( .A(n13457), .ZN(n12650) );
  OAI21_X1 U15162 ( .B1(n12644), .B2(n12643), .A(n12642), .ZN(n12645) );
  NAND2_X1 U15163 ( .A1(n12645), .A2(n12730), .ZN(n12649) );
  AOI22_X1 U15164 ( .A1(n13294), .A2(n12741), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12646) );
  OAI21_X1 U15165 ( .B1(n13264), .B2(n12743), .A(n12646), .ZN(n12647) );
  AOI21_X1 U15166 ( .B1(n13258), .B2(n12747), .A(n12647), .ZN(n12648) );
  OAI211_X1 U15167 ( .C1(n12650), .C2(n12744), .A(n12649), .B(n12648), .ZN(
        P3_U3163) );
  NAND2_X1 U15168 ( .A1(n12652), .A2(n12651), .ZN(n12657) );
  INV_X1 U15169 ( .A(n12653), .ZN(n12654) );
  NOR2_X1 U15170 ( .A1(n12655), .A2(n12654), .ZN(n12656) );
  XOR2_X1 U15171 ( .A(n12657), .B(n12656), .Z(n12667) );
  OAI21_X1 U15172 ( .B1(n12733), .B2(n12659), .A(n12658), .ZN(n12660) );
  AOI21_X1 U15173 ( .B1(n12735), .B2(n12971), .A(n12660), .ZN(n12661) );
  OAI21_X1 U15174 ( .B1(n12663), .B2(n12662), .A(n12661), .ZN(n12664) );
  AOI21_X1 U15175 ( .B1(n12665), .B2(n12720), .A(n12664), .ZN(n12666) );
  OAI21_X1 U15176 ( .B1(n12667), .B2(n12749), .A(n12666), .ZN(P3_U3164) );
  INV_X1 U15177 ( .A(n12668), .ZN(n12673) );
  NOR3_X1 U15178 ( .A1(n12671), .A2(n12670), .A3(n12669), .ZN(n12672) );
  OAI21_X1 U15179 ( .B1(n12673), .B2(n12672), .A(n12730), .ZN(n12677) );
  AOI22_X1 U15180 ( .A1(n13213), .A2(n12747), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12674) );
  OAI21_X1 U15181 ( .B1(n13238), .B2(n12733), .A(n12674), .ZN(n12675) );
  AOI21_X1 U15182 ( .B1(n12962), .B2(n12735), .A(n12675), .ZN(n12676) );
  OAI211_X1 U15183 ( .C1(n13215), .C2(n12744), .A(n12677), .B(n12676), .ZN(
        P3_U3165) );
  XNOR2_X1 U15184 ( .A(n12678), .B(n13337), .ZN(n12679) );
  XNOR2_X1 U15185 ( .A(n12680), .B(n12679), .ZN(n12686) );
  NAND2_X1 U15186 ( .A1(n12735), .A2(n12681), .ZN(n12682) );
  NAND2_X1 U15187 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13071)
         );
  OAI211_X1 U15188 ( .C1(n13355), .C2(n12733), .A(n12682), .B(n13071), .ZN(
        n12684) );
  INV_X1 U15189 ( .A(n13406), .ZN(n13329) );
  NOR2_X1 U15190 ( .A1(n13329), .A2(n12744), .ZN(n12683) );
  AOI211_X1 U15191 ( .C1(n13327), .C2(n12747), .A(n12684), .B(n12683), .ZN(
        n12685) );
  OAI21_X1 U15192 ( .B1(n12686), .B2(n12749), .A(n12685), .ZN(P3_U3166) );
  XNOR2_X1 U15193 ( .A(n12687), .B(n12688), .ZN(n12693) );
  NAND2_X1 U15194 ( .A1(n12741), .A2(n12968), .ZN(n12689) );
  NAND2_X1 U15195 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13093)
         );
  OAI211_X1 U15196 ( .C1(n13316), .C2(n12743), .A(n12689), .B(n13093), .ZN(
        n12691) );
  NOR2_X1 U15197 ( .A1(n13400), .A2(n12744), .ZN(n12690) );
  AOI211_X1 U15198 ( .C1(n13317), .C2(n12747), .A(n12691), .B(n12690), .ZN(
        n12692) );
  OAI21_X1 U15199 ( .B1(n12693), .B2(n12749), .A(n12692), .ZN(P3_U3168) );
  XNOR2_X1 U15200 ( .A(n12695), .B(n12694), .ZN(n12700) );
  AOI22_X1 U15201 ( .A1(n12710), .A2(n12741), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12697) );
  NAND2_X1 U15202 ( .A1(n13273), .A2(n12747), .ZN(n12696) );
  OAI211_X1 U15203 ( .C1(n13283), .C2(n12743), .A(n12697), .B(n12696), .ZN(
        n12698) );
  AOI21_X1 U15204 ( .B1(n13391), .B2(n12720), .A(n12698), .ZN(n12699) );
  OAI21_X1 U15205 ( .B1(n12700), .B2(n12749), .A(n12699), .ZN(P3_U3173) );
  AOI21_X1 U15206 ( .B1(n12966), .B2(n12702), .A(n12701), .ZN(n12707) );
  AOI22_X1 U15207 ( .A1(n13252), .A2(n12741), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12704) );
  NAND2_X1 U15208 ( .A1(n13248), .A2(n12747), .ZN(n12703) );
  OAI211_X1 U15209 ( .C1(n13227), .C2(n12743), .A(n12704), .B(n12703), .ZN(
        n12705) );
  AOI21_X1 U15210 ( .B1(n13451), .B2(n12720), .A(n12705), .ZN(n12706) );
  OAI21_X1 U15211 ( .B1(n12707), .B2(n12749), .A(n12706), .ZN(P3_U3175) );
  XNOR2_X1 U15212 ( .A(n12709), .B(n12708), .ZN(n12715) );
  NAND2_X1 U15213 ( .A1(n12710), .A2(n12735), .ZN(n12711) );
  NAND2_X1 U15214 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13119)
         );
  OAI211_X1 U15215 ( .C1(n13326), .C2(n12733), .A(n12711), .B(n13119), .ZN(
        n12712) );
  AOI21_X1 U15216 ( .B1(n13303), .B2(n12747), .A(n12712), .ZN(n12714) );
  NAND2_X1 U15217 ( .A1(n13470), .A2(n12720), .ZN(n12713) );
  OAI211_X1 U15218 ( .C1(n12715), .C2(n12749), .A(n12714), .B(n12713), .ZN(
        P3_U3178) );
  OAI211_X1 U15219 ( .C1(n12718), .C2(n12717), .A(n12716), .B(n12730), .ZN(
        n12726) );
  AOI21_X1 U15220 ( .B1(n12735), .B2(n12837), .A(n12719), .ZN(n12725) );
  AOI22_X1 U15221 ( .A1(n12741), .A2(n12977), .B1(n12721), .B2(n12720), .ZN(
        n12724) );
  NAND2_X1 U15222 ( .A1(n12747), .A2(n12722), .ZN(n12723) );
  NAND4_X1 U15223 ( .A1(n12726), .A2(n12725), .A3(n12724), .A4(n12723), .ZN(
        P3_U3179) );
  OAI21_X1 U15224 ( .B1(n12729), .B2(n12728), .A(n12727), .ZN(n12731) );
  NAND2_X1 U15225 ( .A1(n12731), .A2(n12730), .ZN(n12737) );
  AOI22_X1 U15226 ( .A1(n13201), .A2(n12747), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12732) );
  OAI21_X1 U15227 ( .B1(n13228), .B2(n12733), .A(n12732), .ZN(n12734) );
  AOI21_X1 U15228 ( .B1(n12961), .B2(n12735), .A(n12734), .ZN(n12736) );
  OAI211_X1 U15229 ( .C1(n13433), .C2(n12744), .A(n12737), .B(n12736), .ZN(
        P3_U3180) );
  XNOR2_X1 U15230 ( .A(n12738), .B(n13355), .ZN(n12739) );
  XNOR2_X1 U15231 ( .A(n12740), .B(n12739), .ZN(n12750) );
  NAND2_X1 U15232 ( .A1(n12741), .A2(n12970), .ZN(n12742) );
  NAND2_X1 U15233 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13037)
         );
  OAI211_X1 U15234 ( .C1(n13337), .C2(n12743), .A(n12742), .B(n13037), .ZN(
        n12746) );
  INV_X1 U15235 ( .A(n13410), .ZN(n13341) );
  NOR2_X1 U15236 ( .A1(n13341), .A2(n12744), .ZN(n12745) );
  AOI211_X1 U15237 ( .C1(n13338), .C2(n12747), .A(n12746), .B(n12745), .ZN(
        n12748) );
  OAI21_X1 U15238 ( .B1(n12750), .B2(n12749), .A(n12748), .ZN(P3_U3181) );
  XNOR2_X1 U15239 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12754) );
  XNOR2_X1 U15240 ( .A(n12755), .B(n12754), .ZN(n13501) );
  NAND2_X1 U15241 ( .A1(n13501), .A2(n12758), .ZN(n12757) );
  INV_X1 U15242 ( .A(SI_31_), .ZN(n13505) );
  OR2_X1 U15243 ( .A1(n12761), .A2(n13505), .ZN(n12756) );
  NAND2_X1 U15244 ( .A1(n12757), .A2(n12756), .ZN(n12786) );
  NAND2_X1 U15245 ( .A1(n12759), .A2(n12758), .ZN(n12763) );
  OR2_X1 U15246 ( .A1(n12761), .A2(n12760), .ZN(n12762) );
  NAND2_X1 U15247 ( .A1(n13158), .A2(n12764), .ZN(n12765) );
  INV_X1 U15248 ( .A(n12793), .ZN(n12951) );
  NAND2_X1 U15249 ( .A1(n12931), .A2(n12932), .ZN(n13199) );
  NAND2_X1 U15250 ( .A1(n12921), .A2(n12920), .ZN(n13224) );
  INV_X1 U15251 ( .A(n12914), .ZN(n12766) );
  INV_X1 U15252 ( .A(n13324), .ZN(n13322) );
  NAND2_X1 U15253 ( .A1(n12767), .A2(n12819), .ZN(n12770) );
  NOR4_X1 U15254 ( .A1(n12770), .A2(n11040), .A3(n12769), .A4(n12768), .ZN(
        n12772) );
  NAND4_X1 U15255 ( .A1(n12809), .A2(n12835), .A3(n12772), .A4(n12771), .ZN(
        n12774) );
  NOR3_X1 U15256 ( .A1(n12774), .A2(n12773), .A3(n12846), .ZN(n12776) );
  NAND4_X1 U15257 ( .A1(n12776), .A2(n12775), .A3(n12851), .A4(n12858), .ZN(
        n12777) );
  NOR4_X1 U15258 ( .A1(n13344), .A2(n13334), .A3(n12777), .A4(n12867), .ZN(
        n12778) );
  NAND4_X1 U15259 ( .A1(n13305), .A2(n12885), .A3(n13322), .A4(n12778), .ZN(
        n12779) );
  NAND3_X1 U15260 ( .A1(n12780), .A2(n13262), .A3(n13271), .ZN(n12781) );
  INV_X1 U15261 ( .A(n12789), .ZN(n12947) );
  NAND2_X1 U15262 ( .A1(n12786), .A2(n13153), .ZN(n12950) );
  NAND2_X1 U15263 ( .A1(n13158), .A2(n13153), .ZN(n12791) );
  NAND3_X1 U15264 ( .A1(n12791), .A2(n12943), .A3(n12939), .ZN(n12788) );
  OAI21_X1 U15265 ( .B1(n12789), .B2(n13153), .A(n12786), .ZN(n12795) );
  INV_X1 U15266 ( .A(n12948), .ZN(n12790) );
  NAND2_X1 U15267 ( .A1(n12791), .A2(n12790), .ZN(n12792) );
  INV_X1 U15268 ( .A(n13199), .ZN(n12929) );
  NAND2_X1 U15269 ( .A1(n12803), .A2(n12801), .ZN(n12802) );
  NAND2_X1 U15270 ( .A1(n12807), .A2(n12803), .ZN(n12804) );
  NAND2_X1 U15271 ( .A1(n12804), .A2(n12930), .ZN(n12805) );
  MUX2_X1 U15272 ( .A(n12807), .B(n12806), .S(n12930), .Z(n12808) );
  NAND3_X1 U15273 ( .A1(n12810), .A2(n12809), .A3(n12808), .ZN(n12814) );
  NAND2_X1 U15274 ( .A1(n12820), .A2(n12811), .ZN(n12812) );
  NAND2_X1 U15275 ( .A1(n12812), .A2(n12946), .ZN(n12813) );
  NAND2_X1 U15276 ( .A1(n10259), .A2(n12815), .ZN(n12816) );
  AOI21_X1 U15277 ( .B1(n12818), .B2(n12816), .A(n12946), .ZN(n12817) );
  OAI21_X1 U15278 ( .B1(n12946), .B2(n12820), .A(n12819), .ZN(n12825) );
  MUX2_X1 U15279 ( .A(n12822), .B(n12821), .S(n12946), .Z(n12823) );
  NAND2_X1 U15280 ( .A1(n12833), .A2(n12826), .ZN(n12829) );
  NAND2_X1 U15281 ( .A1(n12832), .A2(n12827), .ZN(n12828) );
  MUX2_X1 U15282 ( .A(n12829), .B(n12828), .S(n12930), .Z(n12830) );
  INV_X1 U15283 ( .A(n12830), .ZN(n12831) );
  MUX2_X1 U15284 ( .A(n12833), .B(n12832), .S(n12946), .Z(n12834) );
  NAND3_X1 U15285 ( .A1(n12836), .A2(n12835), .A3(n12834), .ZN(n12841) );
  NAND2_X1 U15286 ( .A1(n12838), .A2(n12837), .ZN(n12839) );
  MUX2_X1 U15287 ( .A(n12839), .B(n6498), .S(n12930), .Z(n12840) );
  NAND3_X1 U15288 ( .A1(n12841), .A2(n6437), .A3(n12840), .ZN(n12848) );
  NOR2_X1 U15289 ( .A1(n12843), .A2(n12842), .ZN(n12844) );
  MUX2_X1 U15290 ( .A(n6563), .B(n12844), .S(n12930), .Z(n12845) );
  NOR2_X1 U15291 ( .A1(n12846), .A2(n12845), .ZN(n12847) );
  NAND3_X1 U15292 ( .A1(n12848), .A2(n12851), .A3(n12847), .ZN(n12859) );
  MUX2_X1 U15293 ( .A(n6567), .B(n12849), .S(n12930), .Z(n12850) );
  NAND2_X1 U15294 ( .A1(n12851), .A2(n12850), .ZN(n12857) );
  NOR2_X1 U15295 ( .A1(n12852), .A2(n12974), .ZN(n12854) );
  MUX2_X1 U15296 ( .A(n12854), .B(n12853), .S(n12946), .Z(n12855) );
  INV_X1 U15297 ( .A(n12855), .ZN(n12856) );
  NAND2_X1 U15298 ( .A1(n12866), .A2(n12860), .ZN(n12861) );
  NAND2_X1 U15299 ( .A1(n12861), .A2(n12946), .ZN(n12862) );
  AOI21_X1 U15300 ( .B1(n12865), .B2(n12863), .A(n12946), .ZN(n12864) );
  NOR2_X1 U15301 ( .A1(n12866), .A2(n12946), .ZN(n12868) );
  MUX2_X1 U15302 ( .A(n12870), .B(n12869), .S(n12946), .Z(n12871) );
  INV_X1 U15303 ( .A(n12871), .ZN(n12872) );
  NAND3_X1 U15304 ( .A1(n12873), .A2(n13350), .A3(n12872), .ZN(n12877) );
  NOR2_X1 U15305 ( .A1(n13487), .A2(n13336), .ZN(n12875) );
  MUX2_X1 U15306 ( .A(n12875), .B(n12874), .S(n12930), .Z(n12876) );
  AOI21_X1 U15307 ( .B1(n12879), .B2(n12878), .A(n12930), .ZN(n12880) );
  NAND2_X1 U15308 ( .A1(n12882), .A2(n12881), .ZN(n12883) );
  NAND2_X1 U15309 ( .A1(n12883), .A2(n12930), .ZN(n12884) );
  NAND3_X1 U15310 ( .A1(n12886), .A2(n12885), .A3(n13305), .ZN(n12899) );
  INV_X1 U15311 ( .A(n12894), .ZN(n12887) );
  OR3_X1 U15312 ( .A1(n12888), .A2(n12930), .A3(n12887), .ZN(n12896) );
  AND2_X1 U15313 ( .A1(n13305), .A2(n12889), .ZN(n12892) );
  NAND2_X1 U15314 ( .A1(n12890), .A2(n12930), .ZN(n12891) );
  OAI21_X1 U15315 ( .B1(n12896), .B2(n12892), .A(n12891), .ZN(n12898) );
  INV_X1 U15316 ( .A(n12893), .ZN(n12895) );
  NAND3_X1 U15317 ( .A1(n12896), .A2(n12895), .A3(n12894), .ZN(n12897) );
  NAND3_X1 U15318 ( .A1(n12899), .A2(n12898), .A3(n12897), .ZN(n12903) );
  MUX2_X1 U15319 ( .A(n12901), .B(n12900), .S(n12930), .Z(n12902) );
  NAND3_X1 U15320 ( .A1(n13271), .A2(n12903), .A3(n12902), .ZN(n12907) );
  NAND2_X1 U15321 ( .A1(n13391), .A2(n12946), .ZN(n12905) );
  OR2_X1 U15322 ( .A1(n13391), .A2(n12946), .ZN(n12904) );
  MUX2_X1 U15323 ( .A(n12905), .B(n12904), .S(n13294), .Z(n12906) );
  INV_X1 U15324 ( .A(n13249), .ZN(n12908) );
  INV_X1 U15325 ( .A(n12909), .ZN(n12910) );
  MUX2_X1 U15326 ( .A(n12911), .B(n12910), .S(n12930), .Z(n12917) );
  INV_X1 U15327 ( .A(n13235), .ZN(n12916) );
  INV_X1 U15328 ( .A(n12912), .ZN(n12913) );
  NAND3_X1 U15329 ( .A1(n12918), .A2(n13227), .A3(n12930), .ZN(n12919) );
  INV_X1 U15330 ( .A(n12920), .ZN(n13207) );
  INV_X1 U15331 ( .A(n13218), .ZN(n13206) );
  NAND2_X1 U15332 ( .A1(n12920), .A2(n13206), .ZN(n12922) );
  NAND2_X1 U15333 ( .A1(n12922), .A2(n12921), .ZN(n12923) );
  MUX2_X1 U15334 ( .A(n13207), .B(n12923), .S(n12946), .Z(n12924) );
  OAI21_X1 U15335 ( .B1(n12925), .B2(n12924), .A(n13209), .ZN(n12928) );
  MUX2_X1 U15336 ( .A(n13196), .B(n12926), .S(n12946), .Z(n12927) );
  MUX2_X1 U15337 ( .A(n12932), .B(n12931), .S(n12930), .Z(n12933) );
  NAND2_X1 U15338 ( .A1(n12934), .A2(n12933), .ZN(n12935) );
  NAND2_X1 U15339 ( .A1(n12936), .A2(n12946), .ZN(n12938) );
  AND2_X1 U15340 ( .A1(n12938), .A2(n12937), .ZN(n12940) );
  OAI21_X1 U15341 ( .B1(n12941), .B2(n12940), .A(n12939), .ZN(n12942) );
  OAI211_X1 U15342 ( .C1(n12946), .C2(n12945), .A(n12944), .B(n12943), .ZN(
        n12949) );
  INV_X1 U15343 ( .A(n12953), .ZN(n12955) );
  NAND3_X1 U15344 ( .A1(n12955), .A2(n12954), .A3(n7029), .ZN(n12956) );
  OAI211_X1 U15345 ( .C1(n12957), .C2(n12959), .A(n12956), .B(P3_B_REG_SCAN_IN), .ZN(n12958) );
  MUX2_X1 U15346 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12960), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15347 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12961), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15348 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12962), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15349 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12963), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15350 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12964), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15351 ( .A(n13251), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12965), .Z(
        P3_U3514) );
  MUX2_X1 U15352 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12966), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15353 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13252), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15354 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13294), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15355 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12967), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15356 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12968), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15357 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12969), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15358 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12970), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15359 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12971), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15360 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12972), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15361 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12973), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15362 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12974), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15363 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12975), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15364 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12976), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15365 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12977), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15366 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12978), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15367 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12979), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15368 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n10259), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15369 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n9757), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15370 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15596), .S(P3_U3897), .Z(
        P3_U3491) );
  INV_X1 U15371 ( .A(n12983), .ZN(n12985) );
  AOI21_X1 U15372 ( .B1(n12985), .B2(n12984), .A(n13003), .ZN(n13002) );
  OAI21_X1 U15373 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n12987), .A(n13013), 
        .ZN(n13000) );
  MUX2_X1 U15374 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n7029), .Z(n13017) );
  XNOR2_X1 U15375 ( .A(n13017), .B(n13018), .ZN(n12991) );
  NAND2_X1 U15376 ( .A1(n12989), .A2(n12988), .ZN(n12992) );
  AND2_X1 U15377 ( .A1(n12991), .A2(n12992), .ZN(n12990) );
  INV_X1 U15378 ( .A(n13023), .ZN(n12995) );
  AOI21_X1 U15379 ( .B1(n12993), .B2(n12992), .A(n12991), .ZN(n12994) );
  OAI21_X1 U15380 ( .B1(n12995), .B2(n12994), .A(n13149), .ZN(n12998) );
  AOI21_X1 U15381 ( .B1(n15570), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12996), 
        .ZN(n12997) );
  OAI211_X1 U15382 ( .C1(n13147), .C2(n13004), .A(n12998), .B(n12997), .ZN(
        n12999) );
  AOI21_X1 U15383 ( .B1(n13000), .B2(n13112), .A(n12999), .ZN(n13001) );
  OAI21_X1 U15384 ( .B1(n13002), .B2(n13143), .A(n13001), .ZN(P3_U3195) );
  OR2_X1 U15385 ( .A1(n13028), .A2(n13006), .ZN(n13049) );
  NAND2_X1 U15386 ( .A1(n13028), .A2(n13006), .ZN(n13007) );
  AND2_X1 U15387 ( .A1(n13049), .A2(n13007), .ZN(n13048) );
  XNOR2_X1 U15388 ( .A(n13051), .B(n13048), .ZN(n13031) );
  INV_X1 U15389 ( .A(n13013), .ZN(n13009) );
  OR2_X1 U15390 ( .A1(n13028), .A2(n13359), .ZN(n13040) );
  NAND2_X1 U15391 ( .A1(n13028), .A2(n13359), .ZN(n13008) );
  NAND2_X1 U15392 ( .A1(n13040), .A2(n13008), .ZN(n13011) );
  INV_X1 U15393 ( .A(n13011), .ZN(n13020) );
  NOR3_X1 U15394 ( .A1(n13009), .A2(n13010), .A3(n13020), .ZN(n13014) );
  INV_X1 U15395 ( .A(n13010), .ZN(n13012) );
  OAI21_X1 U15396 ( .B1(n13014), .B2(n13033), .A(n13112), .ZN(n13030) );
  NAND2_X1 U15397 ( .A1(n15570), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n13016) );
  NAND2_X1 U15398 ( .A1(n13016), .A2(n13015), .ZN(n13027) );
  INV_X1 U15399 ( .A(n13017), .ZN(n13019) );
  NAND2_X1 U15400 ( .A1(n13019), .A2(n13018), .ZN(n13022) );
  MUX2_X1 U15401 ( .A(n13048), .B(n13020), .S(n13134), .Z(n13021) );
  INV_X1 U15402 ( .A(n13042), .ZN(n13025) );
  AOI21_X1 U15403 ( .B1(n13023), .B2(n13022), .A(n13021), .ZN(n13024) );
  NOR3_X1 U15404 ( .A1(n13025), .A2(n13024), .A3(n13125), .ZN(n13026) );
  AOI211_X1 U15405 ( .C1(n13100), .C2(n13028), .A(n13027), .B(n13026), .ZN(
        n13029) );
  OAI211_X1 U15406 ( .C1(n13031), .C2(n13143), .A(n13030), .B(n13029), .ZN(
        P3_U3196) );
  INV_X1 U15407 ( .A(n13040), .ZN(n13032) );
  AOI21_X1 U15408 ( .B1(n13036), .B2(n13035), .A(n13076), .ZN(n13056) );
  OAI21_X1 U15409 ( .B1(n13074), .B2(n13038), .A(n13037), .ZN(n13047) );
  MUX2_X1 U15410 ( .A(n13040), .B(n13049), .S(n7029), .Z(n13041) );
  MUX2_X1 U15411 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n7029), .Z(n13043) );
  AOI21_X1 U15412 ( .B1(n13044), .B2(n13043), .A(n13065), .ZN(n13045) );
  NOR2_X1 U15413 ( .A1(n13045), .A2(n13125), .ZN(n13046) );
  AOI211_X1 U15414 ( .C1(n13100), .C2(n13066), .A(n13047), .B(n13046), .ZN(
        n13055) );
  INV_X1 U15415 ( .A(n13048), .ZN(n13050) );
  OAI21_X1 U15416 ( .B1(n13052), .B2(P3_REG1_REG_15__SCAN_IN), .A(n13059), 
        .ZN(n13053) );
  NAND2_X1 U15417 ( .A1(n13053), .A2(n13122), .ZN(n13054) );
  OAI211_X1 U15418 ( .C1(n13056), .C2(n13151), .A(n13055), .B(n13054), .ZN(
        P3_U3197) );
  NAND2_X1 U15419 ( .A1(n13058), .A2(n13057), .ZN(n13060) );
  XNOR2_X1 U15420 ( .A(n13091), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13061) );
  OAI21_X1 U15421 ( .B1(n13062), .B2(n13061), .A(n13090), .ZN(n13063) );
  INV_X1 U15422 ( .A(n13063), .ZN(n13083) );
  INV_X1 U15423 ( .A(n13064), .ZN(n13067) );
  INV_X1 U15424 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13084) );
  INV_X1 U15425 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13407) );
  MUX2_X1 U15426 ( .A(n13084), .B(n13407), .S(n7029), .Z(n13068) );
  NOR2_X1 U15427 ( .A1(n13091), .A2(n13068), .ZN(n13095) );
  INV_X1 U15428 ( .A(n13095), .ZN(n13069) );
  NAND2_X1 U15429 ( .A1(n13091), .A2(n13068), .ZN(n13094) );
  NAND2_X1 U15430 ( .A1(n13069), .A2(n13094), .ZN(n13070) );
  XNOR2_X1 U15431 ( .A(n13096), .B(n13070), .ZN(n13081) );
  NAND2_X1 U15432 ( .A1(n13100), .A2(n13091), .ZN(n13072) );
  OAI211_X1 U15433 ( .C1(n13074), .C2(n13073), .A(n13072), .B(n13071), .ZN(
        n13080) );
  XNOR2_X1 U15434 ( .A(n13091), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13075) );
  OR3_X1 U15435 ( .A1(n13077), .A2(n13076), .A3(n13075), .ZN(n13078) );
  AOI21_X1 U15436 ( .B1(n13086), .B2(n13078), .A(n13151), .ZN(n13079) );
  AOI211_X1 U15437 ( .C1(n13149), .C2(n13081), .A(n13080), .B(n13079), .ZN(
        n13082) );
  OAI21_X1 U15438 ( .B1(n13083), .B2(n13143), .A(n13082), .ZN(P3_U3198) );
  INV_X1 U15439 ( .A(n13111), .ZN(n13087) );
  AOI21_X1 U15440 ( .B1(n13089), .B2(n13088), .A(n13087), .ZN(n13102) );
  INV_X1 U15441 ( .A(n13104), .ZN(n13116) );
  NAND2_X1 U15442 ( .A1(n15570), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n13092) );
  MUX2_X1 U15443 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n7029), .Z(n13105) );
  XNOR2_X1 U15444 ( .A(n13104), .B(n13105), .ZN(n13098) );
  AOI211_X1 U15445 ( .C1(n13098), .C2(n13097), .A(n13125), .B(n13103), .ZN(
        n13099) );
  OAI21_X1 U15446 ( .B1(n13102), .B2(n13151), .A(n13101), .ZN(P3_U3199) );
  MUX2_X1 U15447 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n7029), .Z(n13107) );
  AOI21_X1 U15448 ( .B1(n13107), .B2(n13106), .A(n13130), .ZN(n13126) );
  OR2_X1 U15449 ( .A1(n13131), .A2(n13309), .ZN(n13127) );
  NAND2_X1 U15450 ( .A1(n13131), .A2(n13309), .ZN(n13108) );
  NAND2_X1 U15451 ( .A1(n13127), .A2(n13108), .ZN(n13109) );
  AND3_X1 U15452 ( .A1(n13110), .A2(n13111), .A3(n13109), .ZN(n13113) );
  OAI21_X1 U15453 ( .B1(n13128), .B2(n13113), .A(n13112), .ZN(n13124) );
  INV_X1 U15454 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13403) );
  INV_X1 U15455 ( .A(n13114), .ZN(n13115) );
  OAI22_X1 U15456 ( .A1(n13117), .A2(n13403), .B1(n13116), .B2(n13115), .ZN(
        n13140) );
  XNOR2_X1 U15457 ( .A(n13131), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n13139) );
  XNOR2_X1 U15458 ( .A(n13140), .B(n13139), .ZN(n13121) );
  NAND2_X1 U15459 ( .A1(n15570), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13118) );
  OAI211_X1 U15460 ( .C1(n13147), .C2(n13138), .A(n13119), .B(n13118), .ZN(
        n13120) );
  AOI21_X1 U15461 ( .B1(n13122), .B2(n13121), .A(n13120), .ZN(n13123) );
  OAI211_X1 U15462 ( .C1(n13126), .C2(n13125), .A(n13124), .B(n13123), .ZN(
        P3_U3200) );
  XNOR2_X1 U15463 ( .A(n13146), .B(n13129), .ZN(n13133) );
  XNOR2_X1 U15464 ( .A(n13146), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13142) );
  INV_X1 U15465 ( .A(n13133), .ZN(n13135) );
  MUX2_X1 U15466 ( .A(n13142), .B(n13135), .S(n13134), .Z(n13136) );
  XNOR2_X1 U15467 ( .A(n13137), .B(n13136), .ZN(n13150) );
  AOI22_X1 U15468 ( .A1(n13140), .A2(n13139), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n13138), .ZN(n13141) );
  NAND2_X1 U15469 ( .A1(n15570), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13144) );
  OAI211_X1 U15470 ( .C1(n13147), .C2(n13146), .A(n13145), .B(n13144), .ZN(
        n13148) );
  NAND2_X1 U15471 ( .A1(n12786), .A2(n13347), .ZN(n13156) );
  NOR2_X1 U15472 ( .A1(n13153), .A2(n13152), .ZN(n13419) );
  NAND2_X1 U15473 ( .A1(n13154), .A2(n15604), .ZN(n13162) );
  INV_X1 U15474 ( .A(n13162), .ZN(n13155) );
  OAI21_X1 U15475 ( .B1(n13419), .B2(n13155), .A(n15608), .ZN(n13159) );
  OAI211_X1 U15476 ( .C1(n15608), .C2(n13157), .A(n13156), .B(n13159), .ZN(
        P3_U3202) );
  NAND2_X1 U15477 ( .A1(n13158), .A2(n13347), .ZN(n13160) );
  OAI211_X1 U15478 ( .C1(n15608), .C2(n13161), .A(n13160), .B(n13159), .ZN(
        P3_U3203) );
  OAI21_X1 U15479 ( .B1(n15608), .B2(n13163), .A(n13162), .ZN(n13164) );
  AOI21_X1 U15480 ( .B1(n13166), .B2(n13165), .A(n13164), .ZN(n13169) );
  NAND2_X1 U15481 ( .A1(n13167), .A2(n15608), .ZN(n13168) );
  OAI211_X1 U15482 ( .C1(n13170), .C2(n13363), .A(n13169), .B(n13168), .ZN(
        P3_U3204) );
  XOR2_X1 U15483 ( .A(n13171), .B(n13173), .Z(n13430) );
  INV_X1 U15484 ( .A(n13172), .ZN(n13175) );
  INV_X1 U15485 ( .A(n13173), .ZN(n13174) );
  AOI21_X1 U15486 ( .B1(n13175), .B2(n13174), .A(n15601), .ZN(n13179) );
  OAI22_X1 U15487 ( .A1(n13176), .A2(n15580), .B1(n13193), .B2(n15582), .ZN(
        n13177) );
  AOI21_X1 U15488 ( .B1(n13179), .B2(n13178), .A(n13177), .ZN(n13425) );
  MUX2_X1 U15489 ( .A(n13180), .B(n13425), .S(n15608), .Z(n13183) );
  AOI22_X1 U15490 ( .A1(n13427), .A2(n13347), .B1(n15604), .B2(n13181), .ZN(
        n13182) );
  OAI211_X1 U15491 ( .C1(n13363), .C2(n13430), .A(n13183), .B(n13182), .ZN(
        P3_U3205) );
  INV_X1 U15492 ( .A(n13184), .ZN(n13191) );
  AOI22_X1 U15493 ( .A1(n13185), .A2(n15604), .B1(n15610), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13186) );
  OAI21_X1 U15494 ( .B1(n13187), .B2(n13340), .A(n13186), .ZN(n13188) );
  AOI21_X1 U15495 ( .B1(n13189), .B2(n13245), .A(n13188), .ZN(n13190) );
  OAI21_X1 U15496 ( .B1(n13191), .B2(n15610), .A(n13190), .ZN(P3_U3206) );
  INV_X1 U15497 ( .A(n13371), .ZN(n13205) );
  AOI21_X1 U15498 ( .B1(n10311), .B2(n13195), .A(n13194), .ZN(n13198) );
  INV_X1 U15499 ( .A(n13196), .ZN(n13197) );
  NOR2_X1 U15500 ( .A1(n13198), .A2(n13197), .ZN(n13200) );
  XNOR2_X1 U15501 ( .A(n13200), .B(n13199), .ZN(n13373) );
  AOI22_X1 U15502 ( .A1(n13201), .A2(n15604), .B1(n15610), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13202) );
  OAI21_X1 U15503 ( .B1(n13433), .B2(n13340), .A(n13202), .ZN(n13203) );
  AOI21_X1 U15504 ( .B1(n13373), .B2(n13245), .A(n13203), .ZN(n13204) );
  OAI21_X1 U15505 ( .B1(n15610), .B2(n13205), .A(n13204), .ZN(P3_U3207) );
  INV_X1 U15506 ( .A(n10311), .ZN(n13234) );
  NOR3_X1 U15507 ( .A1(n13233), .A2(n13206), .A3(n13224), .ZN(n13220) );
  NOR2_X1 U15508 ( .A1(n13220), .A2(n13207), .ZN(n13208) );
  XNOR2_X1 U15509 ( .A(n13208), .B(n13209), .ZN(n13437) );
  XNOR2_X1 U15510 ( .A(n13210), .B(n13209), .ZN(n13211) );
  OAI222_X1 U15511 ( .A1(n15580), .A2(n13212), .B1(n15582), .B2(n13238), .C1(
        n13211), .C2(n15601), .ZN(n13375) );
  AOI22_X1 U15512 ( .A1(n13213), .A2(n15604), .B1(n15610), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13214) );
  OAI21_X1 U15513 ( .B1(n13215), .B2(n13340), .A(n13214), .ZN(n13216) );
  AOI21_X1 U15514 ( .B1(n13375), .B2(n15608), .A(n13216), .ZN(n13217) );
  OAI21_X1 U15515 ( .B1(n13437), .B2(n13363), .A(n13217), .ZN(P3_U3208) );
  INV_X1 U15516 ( .A(n13233), .ZN(n13219) );
  NAND2_X1 U15517 ( .A1(n13219), .A2(n13218), .ZN(n13221) );
  AOI22_X1 U15518 ( .A1(n13223), .A2(n13347), .B1(n15604), .B2(n13222), .ZN(
        n13232) );
  XOR2_X1 U15519 ( .A(n13225), .B(n13224), .Z(n13226) );
  OAI222_X1 U15520 ( .A1(n15580), .A2(n13228), .B1(n15582), .B2(n13227), .C1(
        n13226), .C2(n15601), .ZN(n13440) );
  INV_X1 U15521 ( .A(n13440), .ZN(n13229) );
  MUX2_X1 U15522 ( .A(n13230), .B(n13229), .S(n15608), .Z(n13231) );
  OAI211_X1 U15523 ( .C1(n13439), .C2(n13363), .A(n13232), .B(n13231), .ZN(
        P3_U3209) );
  AOI21_X1 U15524 ( .B1(n13234), .B2(n13235), .A(n13233), .ZN(n13381) );
  NOR2_X1 U15525 ( .A1(n6584), .A2(n13235), .ZN(n13237) );
  OR3_X1 U15526 ( .A1(n13237), .A2(n13236), .A3(n15601), .ZN(n13241) );
  OAI22_X1 U15527 ( .A1(n13238), .A2(n15580), .B1(n13264), .B2(n15582), .ZN(
        n13239) );
  INV_X1 U15528 ( .A(n13239), .ZN(n13240) );
  NAND2_X1 U15529 ( .A1(n13241), .A2(n13240), .ZN(n13446) );
  MUX2_X1 U15530 ( .A(n13446), .B(P3_REG2_REG_23__SCAN_IN), .S(n15610), .Z(
        n13244) );
  OAI22_X1 U15531 ( .A1(n13444), .A2(n13340), .B1(n13242), .B2(n15577), .ZN(
        n13243) );
  AOI211_X1 U15532 ( .C1(n13381), .C2(n13245), .A(n13244), .B(n13243), .ZN(
        n13246) );
  INV_X1 U15533 ( .A(n13246), .ZN(P3_U3210) );
  XNOR2_X1 U15534 ( .A(n13247), .B(n13249), .ZN(n13454) );
  AOI22_X1 U15535 ( .A1(n13451), .A2(n13347), .B1(n15604), .B2(n13248), .ZN(
        n13256) );
  XNOR2_X1 U15536 ( .A(n13250), .B(n13249), .ZN(n13253) );
  AOI222_X1 U15537 ( .A1(n10349), .A2(n13253), .B1(n13252), .B2(n15595), .C1(
        n13251), .C2(n15597), .ZN(n13449) );
  MUX2_X1 U15538 ( .A(n13254), .B(n13449), .S(n15608), .Z(n13255) );
  OAI211_X1 U15539 ( .C1(n13454), .C2(n13363), .A(n13256), .B(n13255), .ZN(
        P3_U3211) );
  XNOR2_X1 U15540 ( .A(n13257), .B(n13262), .ZN(n13459) );
  AOI22_X1 U15541 ( .A1(n13457), .A2(n13347), .B1(n15604), .B2(n13258), .ZN(
        n13269) );
  INV_X1 U15542 ( .A(n13259), .ZN(n13260) );
  AOI21_X1 U15543 ( .B1(n13262), .B2(n13261), .A(n13260), .ZN(n13263) );
  OAI222_X1 U15544 ( .A1(n15582), .A2(n13265), .B1(n15580), .B2(n13264), .C1(
        n15601), .C2(n13263), .ZN(n13455) );
  INV_X1 U15545 ( .A(n13455), .ZN(n13266) );
  MUX2_X1 U15546 ( .A(n13267), .B(n13266), .S(n15608), .Z(n13268) );
  OAI211_X1 U15547 ( .C1(n13459), .C2(n13363), .A(n13269), .B(n13268), .ZN(
        P3_U3212) );
  OAI21_X1 U15548 ( .B1(n13272), .B2(n13271), .A(n13270), .ZN(n13463) );
  INV_X1 U15549 ( .A(n13273), .ZN(n13275) );
  OAI22_X1 U15550 ( .A1(n13275), .A2(n15577), .B1(n15608), .B2(n13274), .ZN(
        n13276) );
  AOI21_X1 U15551 ( .B1(n13391), .B2(n13347), .A(n13276), .ZN(n13285) );
  NAND2_X1 U15552 ( .A1(n13291), .A2(n13279), .ZN(n13281) );
  XNOR2_X1 U15553 ( .A(n13281), .B(n13280), .ZN(n13282) );
  OAI222_X1 U15554 ( .A1(n15580), .A2(n13283), .B1(n15582), .B2(n13307), .C1(
        n15601), .C2(n13282), .ZN(n13390) );
  NAND2_X1 U15555 ( .A1(n13390), .A2(n15608), .ZN(n13284) );
  OAI211_X1 U15556 ( .C1(n13463), .C2(n13363), .A(n13285), .B(n13284), .ZN(
        P3_U3213) );
  NAND2_X1 U15557 ( .A1(n6925), .A2(n13287), .ZN(n13288) );
  XOR2_X1 U15558 ( .A(n13292), .B(n13288), .Z(n13467) );
  INV_X1 U15559 ( .A(n13289), .ZN(n13290) );
  NOR2_X1 U15560 ( .A1(n13304), .A2(n13290), .ZN(n13293) );
  OAI211_X1 U15561 ( .C1(n13293), .C2(n13292), .A(n13291), .B(n10349), .ZN(
        n13296) );
  NAND2_X1 U15562 ( .A1(n13294), .A2(n15597), .ZN(n13295) );
  OAI211_X1 U15563 ( .C1(n13316), .C2(n15582), .A(n13296), .B(n13295), .ZN(
        n13394) );
  AOI22_X1 U15564 ( .A1(n15610), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n13297), 
        .B2(n15604), .ZN(n13298) );
  OAI21_X1 U15565 ( .B1(n13299), .B2(n13340), .A(n13298), .ZN(n13300) );
  AOI21_X1 U15566 ( .B1(n13394), .B2(n15608), .A(n13300), .ZN(n13301) );
  OAI21_X1 U15567 ( .B1(n13467), .B2(n13363), .A(n13301), .ZN(P3_U3214) );
  OAI21_X1 U15568 ( .B1(n13302), .B2(n13305), .A(n6925), .ZN(n13472) );
  AOI22_X1 U15569 ( .A1(n13470), .A2(n13347), .B1(n15604), .B2(n13303), .ZN(
        n13311) );
  AOI21_X1 U15570 ( .B1(n13305), .B2(n13277), .A(n13304), .ZN(n13306) );
  OAI222_X1 U15571 ( .A1(n15580), .A2(n13307), .B1(n15582), .B2(n13326), .C1(
        n15601), .C2(n13306), .ZN(n13468) );
  INV_X1 U15572 ( .A(n13468), .ZN(n13308) );
  MUX2_X1 U15573 ( .A(n13309), .B(n13308), .S(n15608), .Z(n13310) );
  OAI211_X1 U15574 ( .C1(n13472), .C2(n13363), .A(n13311), .B(n13310), .ZN(
        P3_U3215) );
  XNOR2_X1 U15575 ( .A(n13312), .B(n13314), .ZN(n13476) );
  XNOR2_X1 U15576 ( .A(n13313), .B(n13314), .ZN(n13315) );
  OAI222_X1 U15577 ( .A1(n15580), .A2(n13316), .B1(n15582), .B2(n13337), .C1(
        n13315), .C2(n15601), .ZN(n13401) );
  AOI22_X1 U15578 ( .A1(n15610), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15604), 
        .B2(n13317), .ZN(n13318) );
  OAI21_X1 U15579 ( .B1(n13400), .B2(n13340), .A(n13318), .ZN(n13319) );
  AOI21_X1 U15580 ( .B1(n13401), .B2(n15608), .A(n13319), .ZN(n13320) );
  OAI21_X1 U15581 ( .B1(n13476), .B2(n13363), .A(n13320), .ZN(P3_U3216) );
  XNOR2_X1 U15582 ( .A(n13321), .B(n13322), .ZN(n13480) );
  XNOR2_X1 U15583 ( .A(n13323), .B(n13324), .ZN(n13325) );
  OAI222_X1 U15584 ( .A1(n15580), .A2(n13326), .B1(n15582), .B2(n13355), .C1(
        n13325), .C2(n15601), .ZN(n13405) );
  AOI22_X1 U15585 ( .A1(n15610), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15604), 
        .B2(n13327), .ZN(n13328) );
  OAI21_X1 U15586 ( .B1(n13329), .B2(n13340), .A(n13328), .ZN(n13330) );
  AOI21_X1 U15587 ( .B1(n13405), .B2(n15608), .A(n13330), .ZN(n13331) );
  OAI21_X1 U15588 ( .B1(n13480), .B2(n13363), .A(n13331), .ZN(P3_U3217) );
  AOI21_X1 U15589 ( .B1(n13332), .B2(n13334), .A(n6613), .ZN(n13484) );
  XNOR2_X1 U15590 ( .A(n13333), .B(n13334), .ZN(n13335) );
  OAI222_X1 U15591 ( .A1(n15580), .A2(n13337), .B1(n15582), .B2(n13336), .C1(
        n13335), .C2(n15601), .ZN(n13409) );
  AOI22_X1 U15592 ( .A1(n15610), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15604), 
        .B2(n13338), .ZN(n13339) );
  OAI21_X1 U15593 ( .B1(n13341), .B2(n13340), .A(n13339), .ZN(n13342) );
  AOI21_X1 U15594 ( .B1(n13409), .B2(n15608), .A(n13342), .ZN(n13343) );
  OAI21_X1 U15595 ( .B1(n13484), .B2(n13363), .A(n13343), .ZN(P3_U3218) );
  XNOR2_X1 U15596 ( .A(n13345), .B(n13344), .ZN(n13489) );
  AOI22_X1 U15597 ( .A1(n13487), .A2(n13347), .B1(n15604), .B2(n13346), .ZN(
        n13362) );
  NAND2_X1 U15598 ( .A1(n13349), .A2(n13348), .ZN(n13351) );
  NAND2_X1 U15599 ( .A1(n13351), .A2(n13350), .ZN(n13352) );
  NAND3_X1 U15600 ( .A1(n13353), .A2(n10349), .A3(n13352), .ZN(n13358) );
  OAI22_X1 U15601 ( .A1(n13355), .A2(n15580), .B1(n13354), .B2(n15582), .ZN(
        n13356) );
  INV_X1 U15602 ( .A(n13356), .ZN(n13357) );
  NAND2_X1 U15603 ( .A1(n13358), .A2(n13357), .ZN(n13485) );
  INV_X1 U15604 ( .A(n13485), .ZN(n13360) );
  MUX2_X1 U15605 ( .A(n13360), .B(n13359), .S(n15610), .Z(n13361) );
  OAI211_X1 U15606 ( .C1(n13489), .C2(n13363), .A(n13362), .B(n13361), .ZN(
        P3_U3219) );
  NAND2_X1 U15607 ( .A1(n12786), .A2(n13416), .ZN(n13364) );
  NAND2_X1 U15608 ( .A1(n13419), .A2(n15652), .ZN(n13366) );
  OAI211_X1 U15609 ( .C1(n15652), .C2(n13365), .A(n13364), .B(n13366), .ZN(
        P3_U3490) );
  NAND2_X1 U15610 ( .A1(n7202), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13367) );
  OAI211_X1 U15611 ( .C1(n13424), .C2(n13382), .A(n13367), .B(n13366), .ZN(
        P3_U3489) );
  INV_X1 U15612 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13368) );
  MUX2_X1 U15613 ( .A(n13368), .B(n13425), .S(n15652), .Z(n13370) );
  NAND2_X1 U15614 ( .A1(n13427), .A2(n13416), .ZN(n13369) );
  OAI211_X1 U15615 ( .C1(n13418), .C2(n13430), .A(n13370), .B(n13369), .ZN(
        P3_U3487) );
  INV_X1 U15616 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13374) );
  AOI21_X1 U15617 ( .B1(n13373), .B2(n13372), .A(n13371), .ZN(n13431) );
  INV_X1 U15618 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13377) );
  MUX2_X1 U15619 ( .A(n13377), .B(n13434), .S(n15652), .Z(n13378) );
  OAI22_X1 U15620 ( .A1(n13439), .A2(n13418), .B1(n13438), .B2(n13382), .ZN(
        n13380) );
  MUX2_X1 U15621 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13440), .S(n15652), .Z(
        n13379) );
  OR2_X1 U15622 ( .A1(n13380), .A2(n13379), .ZN(P3_U3483) );
  INV_X1 U15623 ( .A(n13381), .ZN(n13445) );
  OAI22_X1 U15624 ( .A1(n13445), .A2(n13418), .B1(n13444), .B2(n13382), .ZN(
        n13384) );
  MUX2_X1 U15625 ( .A(n13446), .B(P3_REG1_REG_23__SCAN_IN), .S(n7202), .Z(
        n13383) );
  OR2_X1 U15626 ( .A1(n13384), .A2(n13383), .ZN(P3_U3482) );
  INV_X1 U15627 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13385) );
  MUX2_X1 U15628 ( .A(n13385), .B(n13449), .S(n15652), .Z(n13387) );
  NAND2_X1 U15629 ( .A1(n13451), .A2(n13416), .ZN(n13386) );
  OAI211_X1 U15630 ( .C1(n13454), .C2(n13418), .A(n13387), .B(n13386), .ZN(
        P3_U3481) );
  MUX2_X1 U15631 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n13455), .S(n15652), .Z(
        n13388) );
  AOI21_X1 U15632 ( .B1(n13416), .B2(n13457), .A(n13388), .ZN(n13389) );
  OAI21_X1 U15633 ( .B1(n13459), .B2(n13418), .A(n13389), .ZN(P3_U3480) );
  INV_X1 U15634 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13392) );
  AOI21_X1 U15635 ( .B1(n15623), .B2(n13391), .A(n13390), .ZN(n13460) );
  MUX2_X1 U15636 ( .A(n13392), .B(n13460), .S(n15652), .Z(n13393) );
  OAI21_X1 U15637 ( .B1(n13463), .B2(n13418), .A(n13393), .ZN(P3_U3479) );
  INV_X1 U15638 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13396) );
  AOI21_X1 U15639 ( .B1(n13395), .B2(n15623), .A(n13394), .ZN(n13464) );
  MUX2_X1 U15640 ( .A(n13396), .B(n13464), .S(n15652), .Z(n13397) );
  OAI21_X1 U15641 ( .B1(n13467), .B2(n13418), .A(n13397), .ZN(P3_U3478) );
  MUX2_X1 U15642 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13468), .S(n15652), .Z(
        n13398) );
  AOI21_X1 U15643 ( .B1(n13416), .B2(n13470), .A(n13398), .ZN(n13399) );
  OAI21_X1 U15644 ( .B1(n13472), .B2(n13418), .A(n13399), .ZN(P3_U3477) );
  INV_X1 U15645 ( .A(n13400), .ZN(n13402) );
  AOI21_X1 U15646 ( .B1(n13402), .B2(n15623), .A(n13401), .ZN(n13473) );
  MUX2_X1 U15647 ( .A(n13403), .B(n13473), .S(n15652), .Z(n13404) );
  OAI21_X1 U15648 ( .B1(n13476), .B2(n13418), .A(n13404), .ZN(P3_U3476) );
  AOI21_X1 U15649 ( .B1(n15623), .B2(n13406), .A(n13405), .ZN(n13477) );
  MUX2_X1 U15650 ( .A(n13407), .B(n13477), .S(n15652), .Z(n13408) );
  OAI21_X1 U15651 ( .B1(n13480), .B2(n13418), .A(n13408), .ZN(P3_U3475) );
  INV_X1 U15652 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13411) );
  AOI21_X1 U15653 ( .B1(n15623), .B2(n13410), .A(n13409), .ZN(n13481) );
  MUX2_X1 U15654 ( .A(n13411), .B(n13481), .S(n15652), .Z(n13412) );
  OAI21_X1 U15655 ( .B1(n13484), .B2(n13418), .A(n13412), .ZN(P3_U3474) );
  MUX2_X1 U15656 ( .A(n13485), .B(P3_REG1_REG_14__SCAN_IN), .S(n7202), .Z(
        n13413) );
  AOI21_X1 U15657 ( .B1(n13416), .B2(n13487), .A(n13413), .ZN(n13414) );
  OAI21_X1 U15658 ( .B1(n13489), .B2(n13418), .A(n13414), .ZN(P3_U3473) );
  MUX2_X1 U15659 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n13490), .S(n15652), .Z(
        n13415) );
  AOI21_X1 U15660 ( .B1(n13416), .B2(n13492), .A(n13415), .ZN(n13417) );
  OAI21_X1 U15661 ( .B1(n13496), .B2(n13418), .A(n13417), .ZN(P3_U3472) );
  NAND2_X1 U15662 ( .A1(n12786), .A2(n13493), .ZN(n13420) );
  NAND2_X1 U15663 ( .A1(n13419), .A2(n15645), .ZN(n13422) );
  OAI211_X1 U15664 ( .C1(n15645), .C2(n13421), .A(n13420), .B(n13422), .ZN(
        P3_U3458) );
  NAND2_X1 U15665 ( .A1(n15643), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13423) );
  OAI211_X1 U15666 ( .C1(n13424), .C2(n13443), .A(n13423), .B(n13422), .ZN(
        P3_U3457) );
  INV_X1 U15667 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13426) );
  MUX2_X1 U15668 ( .A(n13426), .B(n13425), .S(n15645), .Z(n13429) );
  NAND2_X1 U15669 ( .A1(n13427), .A2(n13493), .ZN(n13428) );
  OAI211_X1 U15670 ( .C1(n13430), .C2(n13495), .A(n13429), .B(n13428), .ZN(
        P3_U3455) );
  INV_X1 U15671 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13432) );
  INV_X1 U15672 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13435) );
  MUX2_X1 U15673 ( .A(n13435), .B(n13434), .S(n15645), .Z(n13436) );
  OAI21_X1 U15674 ( .B1(n13437), .B2(n13495), .A(n13436), .ZN(P3_U3452) );
  OAI22_X1 U15675 ( .A1(n13439), .A2(n13495), .B1(n13438), .B2(n13443), .ZN(
        n13442) );
  MUX2_X1 U15676 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13440), .S(n15645), .Z(
        n13441) );
  OR2_X1 U15677 ( .A1(n13442), .A2(n13441), .ZN(P3_U3451) );
  OAI22_X1 U15678 ( .A1(n13445), .A2(n13495), .B1(n13444), .B2(n13443), .ZN(
        n13448) );
  MUX2_X1 U15679 ( .A(n13446), .B(P3_REG0_REG_23__SCAN_IN), .S(n15643), .Z(
        n13447) );
  OR2_X1 U15680 ( .A1(n13448), .A2(n13447), .ZN(P3_U3450) );
  INV_X1 U15681 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13450) );
  MUX2_X1 U15682 ( .A(n13450), .B(n13449), .S(n15645), .Z(n13453) );
  NAND2_X1 U15683 ( .A1(n13451), .A2(n13493), .ZN(n13452) );
  OAI211_X1 U15684 ( .C1(n13454), .C2(n13495), .A(n13453), .B(n13452), .ZN(
        P3_U3449) );
  MUX2_X1 U15685 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n13455), .S(n15645), .Z(
        n13456) );
  AOI21_X1 U15686 ( .B1(n13493), .B2(n13457), .A(n13456), .ZN(n13458) );
  OAI21_X1 U15687 ( .B1(n13459), .B2(n13495), .A(n13458), .ZN(P3_U3448) );
  INV_X1 U15688 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13461) );
  MUX2_X1 U15689 ( .A(n13461), .B(n13460), .S(n15645), .Z(n13462) );
  OAI21_X1 U15690 ( .B1(n13463), .B2(n13495), .A(n13462), .ZN(P3_U3447) );
  INV_X1 U15691 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13465) );
  MUX2_X1 U15692 ( .A(n13465), .B(n13464), .S(n15645), .Z(n13466) );
  OAI21_X1 U15693 ( .B1(n13467), .B2(n13495), .A(n13466), .ZN(P3_U3446) );
  MUX2_X1 U15694 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13468), .S(n15645), .Z(
        n13469) );
  AOI21_X1 U15695 ( .B1(n13493), .B2(n13470), .A(n13469), .ZN(n13471) );
  OAI21_X1 U15696 ( .B1(n13472), .B2(n13495), .A(n13471), .ZN(P3_U3444) );
  INV_X1 U15697 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13474) );
  MUX2_X1 U15698 ( .A(n13474), .B(n13473), .S(n15645), .Z(n13475) );
  OAI21_X1 U15699 ( .B1(n13476), .B2(n13495), .A(n13475), .ZN(P3_U3441) );
  INV_X1 U15700 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13478) );
  MUX2_X1 U15701 ( .A(n13478), .B(n13477), .S(n15645), .Z(n13479) );
  OAI21_X1 U15702 ( .B1(n13480), .B2(n13495), .A(n13479), .ZN(P3_U3438) );
  INV_X1 U15703 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13482) );
  MUX2_X1 U15704 ( .A(n13482), .B(n13481), .S(n15645), .Z(n13483) );
  OAI21_X1 U15705 ( .B1(n13484), .B2(n13495), .A(n13483), .ZN(P3_U3435) );
  MUX2_X1 U15706 ( .A(n13485), .B(P3_REG0_REG_14__SCAN_IN), .S(n15643), .Z(
        n13486) );
  AOI21_X1 U15707 ( .B1(n13493), .B2(n13487), .A(n13486), .ZN(n13488) );
  OAI21_X1 U15708 ( .B1(n13489), .B2(n13495), .A(n13488), .ZN(P3_U3432) );
  MUX2_X1 U15709 ( .A(P3_REG0_REG_13__SCAN_IN), .B(n13490), .S(n15645), .Z(
        n13491) );
  AOI21_X1 U15710 ( .B1(n13493), .B2(n13492), .A(n13491), .ZN(n13494) );
  OAI21_X1 U15711 ( .B1(n13496), .B2(n13495), .A(n13494), .ZN(P3_U3429) );
  MUX2_X1 U15712 ( .A(P3_D_REG_1__SCAN_IN), .B(n13497), .S(n13498), .Z(
        P3_U3377) );
  MUX2_X1 U15713 ( .A(P3_D_REG_0__SCAN_IN), .B(n13499), .S(n13498), .Z(
        P3_U3376) );
  NAND2_X1 U15714 ( .A1(n13501), .A2(n13500), .ZN(n13504) );
  OR4_X1 U15715 ( .A1(n7809), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), .A4(
        n13502), .ZN(n13503) );
  OAI211_X1 U15716 ( .C1(n13505), .C2(n13522), .A(n13504), .B(n13503), .ZN(
        P3_U3264) );
  INV_X1 U15717 ( .A(n13506), .ZN(n13508) );
  OAI222_X1 U15718 ( .A1(n13522), .A2(n13509), .B1(n13520), .B2(n13508), .C1(
        P3_U3151), .C2(n13507), .ZN(P3_U3266) );
  INV_X1 U15719 ( .A(n13510), .ZN(n13511) );
  OAI222_X1 U15720 ( .A1(P3_U3151), .A2(n13513), .B1(n13522), .B2(n13512), 
        .C1(n13520), .C2(n13511), .ZN(P3_U3267) );
  INV_X1 U15721 ( .A(n13514), .ZN(n13516) );
  OAI222_X1 U15722 ( .A1(n7029), .A2(P3_U3151), .B1(n13520), .B2(n13516), .C1(
        n13515), .C2(n13522), .ZN(P3_U3268) );
  INV_X1 U15723 ( .A(n13518), .ZN(n13519) );
  OAI222_X1 U15724 ( .A1(n13523), .A2(P3_U3151), .B1(n13522), .B2(n13521), 
        .C1(n13520), .C2(n13519), .ZN(P3_U3269) );
  MUX2_X1 U15725 ( .A(n13524), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  INV_X1 U15726 ( .A(n13525), .ZN(n13526) );
  AOI21_X1 U15727 ( .B1(n13528), .B2(n13527), .A(n13526), .ZN(n13534) );
  OAI21_X1 U15728 ( .B1(n13634), .B2(n13931), .A(n13529), .ZN(n13532) );
  OAI22_X1 U15729 ( .A1(n13645), .A2(n13976), .B1(n13530), .B2(n13623), .ZN(
        n13531) );
  AOI211_X1 U15730 ( .C1(n14084), .C2(n13647), .A(n13532), .B(n13531), .ZN(
        n13533) );
  OAI21_X1 U15731 ( .B1(n13534), .B2(n13649), .A(n13533), .ZN(P2_U3187) );
  NOR2_X1 U15732 ( .A1(n13535), .A2(n13609), .ZN(n13537) );
  XNOR2_X1 U15733 ( .A(n13537), .B(n13536), .ZN(n13540) );
  NAND2_X1 U15734 ( .A1(n13540), .A2(n13539), .ZN(n13538) );
  OAI211_X1 U15735 ( .C1(n13540), .C2(n13539), .A(n13538), .B(n13610), .ZN(
        n13545) );
  AOI22_X1 U15736 ( .A1(n13810), .A2(n13568), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13544) );
  AOI22_X1 U15737 ( .A1(n13654), .A2(n13630), .B1(n13815), .B2(n13631), .ZN(
        n13543) );
  NAND2_X1 U15738 ( .A1(n13541), .A2(n13647), .ZN(n13542) );
  NAND4_X1 U15739 ( .A1(n13545), .A2(n13544), .A3(n13543), .A4(n13542), .ZN(
        P2_U3188) );
  NOR2_X1 U15740 ( .A1(n6606), .A2(n13546), .ZN(n13547) );
  XNOR2_X1 U15741 ( .A(n13548), .B(n13547), .ZN(n13555) );
  INV_X1 U15742 ( .A(n13880), .ZN(n13552) );
  OAI22_X1 U15743 ( .A1(n13842), .A2(n13932), .B1(n13549), .B2(n13930), .ZN(
        n13876) );
  NOR2_X1 U15744 ( .A1(n13550), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13706) );
  AOI21_X1 U15745 ( .B1(n13876), .B2(n13643), .A(n13706), .ZN(n13551) );
  OAI21_X1 U15746 ( .B1(n13552), .B2(n13645), .A(n13551), .ZN(n13553) );
  AOI21_X1 U15747 ( .B1(n14059), .B2(n13647), .A(n13553), .ZN(n13554) );
  OAI21_X1 U15748 ( .B1(n13555), .B2(n13649), .A(n13554), .ZN(P2_U3191) );
  OAI211_X1 U15749 ( .C1(n13558), .C2(n13557), .A(n13556), .B(n13610), .ZN(
        n13562) );
  OAI22_X1 U15750 ( .A1(n13645), .A2(n13846), .B1(n13842), .B2(n13623), .ZN(
        n13560) );
  NOR2_X1 U15751 ( .A1(n13634), .A2(n13843), .ZN(n13559) );
  AOI211_X1 U15752 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(P2_U3088), .A(n13560), 
        .B(n13559), .ZN(n13561) );
  OAI211_X1 U15753 ( .C1(n14137), .C2(n13620), .A(n13562), .B(n13561), .ZN(
        P2_U3195) );
  INV_X1 U15754 ( .A(n13784), .ZN(n14126) );
  OAI211_X1 U15755 ( .C1(n13565), .C2(n13564), .A(n13563), .B(n13610), .ZN(
        n13570) );
  AOI22_X1 U15756 ( .A1(n13810), .A2(n13630), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13566) );
  OAI21_X1 U15757 ( .B1(n13782), .B2(n13645), .A(n13566), .ZN(n13567) );
  AOI21_X1 U15758 ( .B1(n13568), .B2(n13773), .A(n13567), .ZN(n13569) );
  OAI211_X1 U15759 ( .C1(n14126), .C2(n13620), .A(n13570), .B(n13569), .ZN(
        P2_U3197) );
  XNOR2_X1 U15760 ( .A(n13571), .B(n13572), .ZN(n13640) );
  AOI22_X1 U15761 ( .A1(n13640), .A2(n13639), .B1(n13571), .B2(n13573), .ZN(
        n13577) );
  NAND2_X1 U15762 ( .A1(n13575), .A2(n13574), .ZN(n13576) );
  XNOR2_X1 U15763 ( .A(n13577), .B(n13576), .ZN(n13581) );
  NAND2_X1 U15764 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n15505)
         );
  OAI21_X1 U15765 ( .B1(n13634), .B2(n13933), .A(n15505), .ZN(n13579) );
  OAI22_X1 U15766 ( .A1(n13645), .A2(n13937), .B1(n13931), .B2(n13623), .ZN(
        n13578) );
  AOI211_X1 U15767 ( .C1(n14074), .C2(n13647), .A(n13579), .B(n13578), .ZN(
        n13580) );
  OAI21_X1 U15768 ( .B1(n13581), .B2(n13649), .A(n13580), .ZN(P2_U3198) );
  OAI21_X1 U15769 ( .B1(n6993), .B2(n13583), .A(n13582), .ZN(n13585) );
  NAND2_X1 U15770 ( .A1(n13585), .A2(n13610), .ZN(n13589) );
  INV_X1 U15771 ( .A(n13586), .ZN(n13921) );
  AOI22_X1 U15772 ( .A1(n13657), .A2(n13968), .B1(n13966), .B2(n13658), .ZN(
        n13915) );
  NAND2_X1 U15773 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15520)
         );
  OAI21_X1 U15774 ( .B1(n13915), .B2(n13616), .A(n15520), .ZN(n13587) );
  AOI21_X1 U15775 ( .B1(n13921), .B2(n13631), .A(n13587), .ZN(n13588) );
  OAI211_X1 U15776 ( .C1(n14146), .C2(n13620), .A(n13589), .B(n13588), .ZN(
        P2_U3200) );
  OAI211_X1 U15777 ( .C1(n13592), .C2(n13591), .A(n13590), .B(n13610), .ZN(
        n13599) );
  OAI22_X1 U15778 ( .A1(n13594), .A2(n13634), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13593), .ZN(n13597) );
  OAI22_X1 U15779 ( .A1(n13595), .A2(n13623), .B1(n13798), .B2(n13645), .ZN(
        n13596) );
  AOI211_X1 U15780 ( .C1(n14036), .C2(n13647), .A(n13597), .B(n13596), .ZN(
        n13598) );
  NAND2_X1 U15781 ( .A1(n13599), .A2(n13598), .ZN(P2_U3201) );
  INV_X1 U15782 ( .A(n14140), .ZN(n13608) );
  OAI21_X1 U15783 ( .B1(n13602), .B2(n13601), .A(n13600), .ZN(n13603) );
  NAND2_X1 U15784 ( .A1(n13603), .A2(n13610), .ZN(n13607) );
  OAI22_X1 U15785 ( .A1(n13645), .A2(n13863), .B1(n13859), .B2(n13623), .ZN(
        n13605) );
  NOR2_X1 U15786 ( .A1(n13634), .A2(n13860), .ZN(n13604) );
  AOI211_X1 U15787 ( .C1(P2_REG3_REG_20__SCAN_IN), .C2(P2_U3088), .A(n13605), 
        .B(n13604), .ZN(n13606) );
  OAI211_X1 U15788 ( .C1(n13608), .C2(n13620), .A(n13607), .B(n13606), .ZN(
        P2_U3205) );
  INV_X1 U15789 ( .A(n13609), .ZN(n13611) );
  OAI211_X1 U15790 ( .C1(n13613), .C2(n13612), .A(n13611), .B(n13610), .ZN(
        n13619) );
  INV_X1 U15791 ( .A(n13614), .ZN(n13832) );
  AOI22_X1 U15792 ( .A1(n13794), .A2(n13968), .B1(n13966), .B2(n13655), .ZN(
        n13827) );
  OAI22_X1 U15793 ( .A1(n13827), .A2(n13616), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13615), .ZN(n13617) );
  AOI21_X1 U15794 ( .B1(n13832), .B2(n13631), .A(n13617), .ZN(n13618) );
  OAI211_X1 U15795 ( .C1(n14133), .C2(n13620), .A(n13619), .B(n13618), .ZN(
        P2_U3207) );
  XNOR2_X1 U15796 ( .A(n13622), .B(n13621), .ZN(n13627) );
  NAND2_X1 U15797 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13680)
         );
  OAI21_X1 U15798 ( .B1(n13634), .B2(n13859), .A(n13680), .ZN(n13625) );
  OAI22_X1 U15799 ( .A1(n13645), .A2(n13902), .B1(n13933), .B2(n13623), .ZN(
        n13624) );
  AOI211_X1 U15800 ( .C1(n14064), .C2(n13647), .A(n13625), .B(n13624), .ZN(
        n13626) );
  OAI21_X1 U15801 ( .B1(n13627), .B2(n13649), .A(n13626), .ZN(P2_U3210) );
  AOI21_X1 U15802 ( .B1(n13629), .B2(n13628), .A(n6524), .ZN(n13638) );
  AOI22_X1 U15803 ( .A1(n13795), .A2(n13630), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13633) );
  NAND2_X1 U15804 ( .A1(n13763), .A2(n13631), .ZN(n13632) );
  OAI211_X1 U15805 ( .C1(n13635), .C2(n13634), .A(n13633), .B(n13632), .ZN(
        n13636) );
  AOI21_X1 U15806 ( .B1(n14026), .B2(n13647), .A(n13636), .ZN(n13637) );
  OAI21_X1 U15807 ( .B1(n13638), .B2(n13649), .A(n13637), .ZN(P2_U3212) );
  XNOR2_X1 U15808 ( .A(n13640), .B(n13639), .ZN(n13650) );
  OAI22_X1 U15809 ( .A1(n13641), .A2(n13932), .B1(n13659), .B2(n13930), .ZN(
        n13949) );
  AOI21_X1 U15810 ( .B1(n13643), .B2(n13949), .A(n13642), .ZN(n13644) );
  OAI21_X1 U15811 ( .B1(n13645), .B2(n13957), .A(n13644), .ZN(n13646) );
  AOI21_X1 U15812 ( .B1(n13955), .B2(n13647), .A(n13646), .ZN(n13648) );
  OAI21_X1 U15813 ( .B1(n13650), .B2(n13649), .A(n13648), .ZN(P2_U3213) );
  MUX2_X1 U15814 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13651), .S(n13667), .Z(
        P2_U3562) );
  MUX2_X1 U15815 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13652), .S(n13667), .Z(
        P2_U3561) );
  CLKBUF_X2 U15816 ( .A(P2_U3947), .Z(n13667) );
  MUX2_X1 U15817 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13653), .S(n13667), .Z(
        P2_U3560) );
  MUX2_X1 U15818 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13742), .S(n13667), .Z(
        P2_U3559) );
  MUX2_X1 U15819 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13760), .S(n13667), .Z(
        P2_U3558) );
  MUX2_X1 U15820 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13773), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15821 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13795), .S(n13667), .Z(
        P2_U3556) );
  MUX2_X1 U15822 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13810), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15823 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13794), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15824 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13654), .S(n13667), .Z(
        P2_U3553) );
  MUX2_X1 U15825 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13655), .S(n13667), .Z(
        P2_U3552) );
  MUX2_X1 U15826 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13656), .S(n13667), .Z(
        P2_U3551) );
  MUX2_X1 U15827 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13894), .S(n13667), .Z(
        P2_U3550) );
  MUX2_X1 U15828 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13657), .S(n13667), .Z(
        P2_U3549) );
  MUX2_X1 U15829 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13893), .S(n13667), .Z(
        P2_U3548) );
  MUX2_X1 U15830 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13658), .S(n13667), .Z(
        P2_U3547) );
  MUX2_X1 U15831 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13969), .S(n13667), .Z(
        P2_U3546) );
  INV_X1 U15832 ( .A(n13659), .ZN(n13660) );
  MUX2_X1 U15833 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13660), .S(n13667), .Z(
        P2_U3545) );
  MUX2_X1 U15834 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13967), .S(n13667), .Z(
        P2_U3544) );
  MUX2_X1 U15835 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13661), .S(n13667), .Z(
        P2_U3543) );
  MUX2_X1 U15836 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13662), .S(P2_U3947), .Z(
        P2_U3542) );
  MUX2_X1 U15837 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13663), .S(P2_U3947), .Z(
        P2_U3541) );
  MUX2_X1 U15838 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13664), .S(P2_U3947), .Z(
        P2_U3540) );
  MUX2_X1 U15839 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13665), .S(P2_U3947), .Z(
        P2_U3539) );
  MUX2_X1 U15840 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13666), .S(P2_U3947), .Z(
        P2_U3538) );
  MUX2_X1 U15841 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13668), .S(n13667), .Z(
        P2_U3537) );
  MUX2_X1 U15842 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13669), .S(n13667), .Z(
        P2_U3536) );
  MUX2_X1 U15843 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13670), .S(n13667), .Z(
        P2_U3535) );
  MUX2_X1 U15844 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13671), .S(n13667), .Z(
        P2_U3534) );
  MUX2_X1 U15845 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8790), .S(n13667), .Z(
        P2_U3533) );
  MUX2_X1 U15846 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13672), .S(n13667), .Z(
        P2_U3532) );
  MUX2_X1 U15847 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13673), .S(n13667), .Z(
        P2_U3531) );
  NAND2_X1 U15848 ( .A1(n13674), .A2(n13685), .ZN(n13675) );
  NAND2_X1 U15849 ( .A1(n13676), .A2(n13675), .ZN(n15498) );
  INV_X1 U15850 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13940) );
  XNOR2_X1 U15851 ( .A(n15504), .B(n13940), .ZN(n15497) );
  NAND2_X1 U15852 ( .A1(n15498), .A2(n15497), .ZN(n15496) );
  NAND2_X1 U15853 ( .A1(n15504), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13677) );
  NAND2_X1 U15854 ( .A1(n15496), .A2(n13677), .ZN(n15511) );
  INV_X1 U15855 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13678) );
  MUX2_X1 U15856 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n13678), .S(n15518), .Z(
        n15510) );
  NAND2_X1 U15857 ( .A1(n15511), .A2(n15510), .ZN(n15509) );
  NAND2_X1 U15858 ( .A1(n15518), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13679) );
  NAND2_X1 U15859 ( .A1(n15509), .A2(n13679), .ZN(n13698) );
  XNOR2_X1 U15860 ( .A(n13698), .B(n13699), .ZN(n13700) );
  XNOR2_X1 U15861 ( .A(n13700), .B(n13903), .ZN(n13692) );
  INV_X1 U15862 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n13681) );
  OAI21_X1 U15863 ( .B1(n15522), .B2(n13681), .A(n13680), .ZN(n13690) );
  INV_X1 U15864 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13688) );
  INV_X1 U15865 ( .A(n13682), .ZN(n13684) );
  XNOR2_X1 U15866 ( .A(n15504), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15500) );
  XNOR2_X1 U15867 ( .A(n15518), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15514) );
  AOI211_X1 U15868 ( .C1(n13688), .C2(n13687), .A(n15513), .B(n13694), .ZN(
        n13689) );
  AOI211_X1 U15869 ( .C1(n15519), .C2(n13699), .A(n13690), .B(n13689), .ZN(
        n13691) );
  OAI21_X1 U15870 ( .B1(n15421), .B2(n13692), .A(n13691), .ZN(P2_U3232) );
  INV_X1 U15871 ( .A(n13693), .ZN(n13695) );
  OAI22_X1 U15872 ( .A1(n13700), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13699), 
        .B2(n13698), .ZN(n13701) );
  XNOR2_X1 U15873 ( .A(n13701), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13702) );
  NOR2_X1 U15874 ( .A1(n13702), .A2(n15421), .ZN(n13703) );
  AOI21_X1 U15875 ( .B1(n15441), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n13706), 
        .ZN(n13707) );
  NOR2_X1 U15876 ( .A1(n13909), .A2(n14000), .ZN(n13714) );
  NOR2_X1 U15877 ( .A1(n14116), .A2(n13979), .ZN(n13708) );
  AOI211_X1 U15878 ( .C1(n13909), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13714), 
        .B(n13708), .ZN(n13709) );
  OAI21_X1 U15879 ( .B1(n13868), .B2(n13710), .A(n13709), .ZN(P2_U3234) );
  AOI21_X1 U15880 ( .B1(n13727), .B2(n13999), .A(n13974), .ZN(n13712) );
  NAND2_X1 U15881 ( .A1(n13712), .A2(n13711), .ZN(n14001) );
  NOR2_X1 U15882 ( .A1(n13987), .A2(n13713), .ZN(n13715) );
  AOI211_X1 U15883 ( .C1(n13999), .C2(n13991), .A(n13715), .B(n13714), .ZN(
        n13716) );
  OAI21_X1 U15884 ( .B1(n14001), .B2(n13868), .A(n13716), .ZN(P2_U3235) );
  AND2_X1 U15885 ( .A1(n13720), .A2(n13742), .ZN(n14005) );
  INV_X1 U15886 ( .A(n14005), .ZN(n14010) );
  OAI21_X1 U15887 ( .B1(n14004), .B2(n14008), .A(n14010), .ZN(n13717) );
  INV_X1 U15888 ( .A(n14011), .ZN(n14006) );
  XNOR2_X1 U15889 ( .A(n13717), .B(n14006), .ZN(n13735) );
  OAI22_X1 U15890 ( .A1(n13723), .A2(n13930), .B1(n13722), .B2(n13721), .ZN(
        n13724) );
  INV_X1 U15891 ( .A(n13724), .ZN(n13725) );
  AND4_X2 U15892 ( .A1(n7828), .A2(n7827), .A3(n7826), .A4(n13725), .ZN(n14020) );
  INV_X1 U15893 ( .A(n14020), .ZN(n13733) );
  AOI21_X1 U15894 ( .B1(n13726), .B2(n14016), .A(n13974), .ZN(n13728) );
  NAND2_X1 U15895 ( .A1(n13728), .A2(n13727), .ZN(n14018) );
  AOI22_X1 U15896 ( .A1(n13729), .A2(n13990), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13909), .ZN(n13731) );
  NAND2_X1 U15897 ( .A1(n14016), .A2(n13991), .ZN(n13730) );
  OAI211_X1 U15898 ( .C1(n14018), .C2(n13868), .A(n13731), .B(n13730), .ZN(
        n13732) );
  AOI21_X1 U15899 ( .B1(n13733), .B2(n13987), .A(n13732), .ZN(n13734) );
  OAI21_X1 U15900 ( .B1(n13735), .B2(n13983), .A(n13734), .ZN(P2_U3236) );
  XNOR2_X1 U15901 ( .A(n13736), .B(n6696), .ZN(n14021) );
  INV_X1 U15902 ( .A(n14021), .ZN(n13756) );
  NAND3_X1 U15903 ( .A1(n13738), .A2(n6696), .A3(n13739), .ZN(n13740) );
  NAND2_X1 U15904 ( .A1(n13741), .A2(n13740), .ZN(n13746) );
  NAND2_X1 U15905 ( .A1(n13742), .A2(n13968), .ZN(n13743) );
  OAI21_X1 U15906 ( .B1(n13744), .B2(n13930), .A(n13743), .ZN(n13745) );
  INV_X1 U15907 ( .A(n14023), .ZN(n13754) );
  OAI211_X1 U15908 ( .C1(n13761), .C2(n14121), .A(n12569), .B(n13747), .ZN(
        n14022) );
  OAI22_X1 U15909 ( .A1(n13749), .A2(n13956), .B1(n13748), .B2(n13987), .ZN(
        n13750) );
  AOI21_X1 U15910 ( .B1(n13751), .B2(n13991), .A(n13750), .ZN(n13752) );
  OAI21_X1 U15911 ( .B1(n14022), .B2(n13868), .A(n13752), .ZN(n13753) );
  AOI21_X1 U15912 ( .B1(n13754), .B2(n13987), .A(n13753), .ZN(n13755) );
  OAI21_X1 U15913 ( .B1(n13756), .B2(n13983), .A(n13755), .ZN(P2_U3238) );
  XNOR2_X1 U15914 ( .A(n13757), .B(n13759), .ZN(n14029) );
  INV_X1 U15915 ( .A(n14028), .ZN(n13767) );
  OAI21_X1 U15916 ( .B1(n13779), .B2(n6692), .A(n12569), .ZN(n13762) );
  NOR2_X1 U15917 ( .A1(n13762), .A2(n13761), .ZN(n14025) );
  NAND2_X1 U15918 ( .A1(n14025), .A2(n13995), .ZN(n13765) );
  AOI22_X1 U15919 ( .A1(n13763), .A2(n13990), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13909), .ZN(n13764) );
  OAI211_X1 U15920 ( .C1(n6692), .C2(n13979), .A(n13765), .B(n13764), .ZN(
        n13766) );
  AOI21_X1 U15921 ( .B1(n13767), .B2(n13987), .A(n13766), .ZN(n13768) );
  OAI21_X1 U15922 ( .B1(n14029), .B2(n13983), .A(n13768), .ZN(P2_U3239) );
  XNOR2_X1 U15923 ( .A(n13769), .B(n7265), .ZN(n14032) );
  OAI21_X1 U15924 ( .B1(n13772), .B2(n13771), .A(n13770), .ZN(n13777) );
  NAND2_X1 U15925 ( .A1(n13773), .A2(n13968), .ZN(n13774) );
  OAI21_X1 U15926 ( .B1(n13775), .B2(n13930), .A(n13774), .ZN(n13776) );
  AOI21_X1 U15927 ( .B1(n13777), .B2(n13971), .A(n13776), .ZN(n14031) );
  INV_X1 U15928 ( .A(n14031), .ZN(n13787) );
  NAND2_X1 U15929 ( .A1(n13796), .A2(n13784), .ZN(n13778) );
  NAND2_X1 U15930 ( .A1(n13778), .A2(n12569), .ZN(n13780) );
  OR2_X1 U15931 ( .A1(n13780), .A2(n13779), .ZN(n14030) );
  OAI22_X1 U15932 ( .A1(n13782), .A2(n13956), .B1(n13781), .B2(n13987), .ZN(
        n13783) );
  AOI21_X1 U15933 ( .B1(n13784), .B2(n13991), .A(n13783), .ZN(n13785) );
  OAI21_X1 U15934 ( .B1(n14030), .B2(n13868), .A(n13785), .ZN(n13786) );
  AOI21_X1 U15935 ( .B1(n13787), .B2(n13987), .A(n13786), .ZN(n13788) );
  OAI21_X1 U15936 ( .B1(n13983), .B2(n14032), .A(n13788), .ZN(P2_U3240) );
  NAND3_X1 U15937 ( .A1(n13809), .A2(n13802), .A3(n13791), .ZN(n13793) );
  INV_X1 U15938 ( .A(n13796), .ZN(n13797) );
  AOI211_X1 U15939 ( .C1(n14036), .C2(n13814), .A(n13974), .B(n13797), .ZN(
        n14035) );
  INV_X1 U15940 ( .A(n13798), .ZN(n13799) );
  AOI22_X1 U15941 ( .A1(n13799), .A2(n13990), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13909), .ZN(n13800) );
  OAI21_X1 U15942 ( .B1(n7408), .B2(n13979), .A(n13800), .ZN(n13804) );
  OAI21_X1 U15943 ( .B1(n6589), .B2(n13802), .A(n13801), .ZN(n14039) );
  NOR2_X1 U15944 ( .A1(n14039), .A2(n13983), .ZN(n13803) );
  AOI211_X1 U15945 ( .C1(n14035), .C2(n13995), .A(n13804), .B(n13803), .ZN(
        n13805) );
  OAI21_X1 U15946 ( .B1(n14038), .B2(n13909), .A(n13805), .ZN(P2_U3241) );
  NAND2_X1 U15947 ( .A1(n13807), .A2(n9036), .ZN(n13808) );
  NAND2_X1 U15948 ( .A1(n13809), .A2(n13808), .ZN(n13813) );
  NAND2_X1 U15949 ( .A1(n13810), .A2(n13968), .ZN(n13811) );
  OAI21_X1 U15950 ( .B1(n13843), .B2(n13930), .A(n13811), .ZN(n13812) );
  OAI211_X1 U15951 ( .C1(n13829), .C2(n14129), .A(n12569), .B(n13814), .ZN(
        n14040) );
  INV_X1 U15952 ( .A(n14040), .ZN(n13820) );
  AOI22_X1 U15953 ( .A1(n13815), .A2(n13990), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n13909), .ZN(n13816) );
  OAI21_X1 U15954 ( .B1(n14129), .B2(n13979), .A(n13816), .ZN(n13819) );
  XNOR2_X1 U15955 ( .A(n13817), .B(n9036), .ZN(n14042) );
  NOR2_X1 U15956 ( .A1(n14042), .A2(n13983), .ZN(n13818) );
  AOI211_X1 U15957 ( .C1(n13820), .C2(n13995), .A(n13819), .B(n13818), .ZN(
        n13821) );
  OAI21_X1 U15958 ( .B1(n14041), .B2(n13909), .A(n13821), .ZN(P2_U3242) );
  NAND2_X1 U15959 ( .A1(n13822), .A2(n13826), .ZN(n13823) );
  AND2_X1 U15960 ( .A1(n13824), .A2(n13823), .ZN(n14045) );
  INV_X1 U15961 ( .A(n14045), .ZN(n13837) );
  OAI211_X1 U15962 ( .C1(n6523), .C2(n13826), .A(n13825), .B(n13971), .ZN(
        n13828) );
  NAND2_X1 U15963 ( .A1(n13828), .A2(n13827), .ZN(n14043) );
  NAND2_X1 U15964 ( .A1(n14043), .A2(n13987), .ZN(n13836) );
  INV_X1 U15965 ( .A(n13849), .ZN(n13830) );
  AOI211_X1 U15966 ( .C1(n13831), .C2(n13830), .A(n13974), .B(n13829), .ZN(
        n14044) );
  AOI22_X1 U15967 ( .A1(n13832), .A2(n13990), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n13909), .ZN(n13833) );
  OAI21_X1 U15968 ( .B1(n14133), .B2(n13979), .A(n13833), .ZN(n13834) );
  AOI21_X1 U15969 ( .B1(n14044), .B2(n13995), .A(n13834), .ZN(n13835) );
  OAI211_X1 U15970 ( .C1(n13837), .C2(n13983), .A(n13836), .B(n13835), .ZN(
        P2_U3243) );
  INV_X1 U15971 ( .A(n13838), .ZN(n13853) );
  NAND3_X1 U15972 ( .A1(n13858), .A2(n13853), .A3(n13839), .ZN(n13840) );
  NAND2_X1 U15973 ( .A1(n13841), .A2(n13840), .ZN(n13845) );
  OAI22_X1 U15974 ( .A1(n13843), .A2(n13932), .B1(n13842), .B2(n13930), .ZN(
        n13844) );
  AOI21_X1 U15975 ( .B1(n13845), .B2(n13971), .A(n13844), .ZN(n14049) );
  OAI22_X1 U15976 ( .A1(n13987), .A2(n13847), .B1(n13846), .B2(n13956), .ZN(
        n13851) );
  OAI21_X1 U15977 ( .B1(n13865), .B2(n14137), .A(n12569), .ZN(n13848) );
  OR2_X1 U15978 ( .A1(n13849), .A2(n13848), .ZN(n14048) );
  NOR2_X1 U15979 ( .A1(n14048), .A2(n13868), .ZN(n13850) );
  AOI211_X1 U15980 ( .C1(n13991), .C2(n7410), .A(n13851), .B(n13850), .ZN(
        n13855) );
  XNOR2_X1 U15981 ( .A(n13852), .B(n13853), .ZN(n14050) );
  OR2_X1 U15982 ( .A1(n14050), .A2(n13983), .ZN(n13854) );
  OAI211_X1 U15983 ( .C1(n14049), .C2(n13909), .A(n13855), .B(n13854), .ZN(
        P2_U3244) );
  NAND2_X1 U15984 ( .A1(n13856), .A2(n13871), .ZN(n13857) );
  NAND2_X1 U15985 ( .A1(n13858), .A2(n13857), .ZN(n13862) );
  OAI22_X1 U15986 ( .A1(n13860), .A2(n13932), .B1(n13859), .B2(n13930), .ZN(
        n13861) );
  AOI21_X1 U15987 ( .B1(n13862), .B2(n13971), .A(n13861), .ZN(n14054) );
  OAI22_X1 U15988 ( .A1(n13987), .A2(n13864), .B1(n13863), .B2(n13956), .ZN(
        n13870) );
  INV_X1 U15989 ( .A(n13865), .ZN(n13867) );
  AOI21_X1 U15990 ( .B1(n13878), .B2(n14140), .A(n13974), .ZN(n13866) );
  NAND2_X1 U15991 ( .A1(n13867), .A2(n13866), .ZN(n14053) );
  NOR2_X1 U15992 ( .A1(n14053), .A2(n13868), .ZN(n13869) );
  AOI211_X1 U15993 ( .C1(n13991), .C2(n14140), .A(n13870), .B(n13869), .ZN(
        n13874) );
  XNOR2_X1 U15994 ( .A(n13872), .B(n7787), .ZN(n14055) );
  OR2_X1 U15995 ( .A1(n14055), .A2(n13983), .ZN(n13873) );
  OAI211_X1 U15996 ( .C1(n14054), .C2(n13909), .A(n13874), .B(n13873), .ZN(
        P2_U3245) );
  XNOR2_X1 U15997 ( .A(n13875), .B(n13883), .ZN(n13877) );
  AOI21_X1 U15998 ( .B1(n13877), .B2(n13971), .A(n13876), .ZN(n14061) );
  INV_X1 U15999 ( .A(n13878), .ZN(n13879) );
  AOI211_X1 U16000 ( .C1(n14059), .C2(n13899), .A(n13974), .B(n13879), .ZN(
        n14058) );
  AOI22_X1 U16001 ( .A1(n13909), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13880), 
        .B2(n13990), .ZN(n13881) );
  OAI21_X1 U16002 ( .B1(n13882), .B2(n13979), .A(n13881), .ZN(n13886) );
  XNOR2_X1 U16003 ( .A(n13884), .B(n13883), .ZN(n14062) );
  NOR2_X1 U16004 ( .A1(n14062), .A2(n13983), .ZN(n13885) );
  AOI211_X1 U16005 ( .C1(n14058), .C2(n13995), .A(n13886), .B(n13885), .ZN(
        n13887) );
  OAI21_X1 U16006 ( .B1(n14061), .B2(n13909), .A(n13887), .ZN(P2_U3246) );
  XOR2_X1 U16007 ( .A(n13888), .B(n13892), .Z(n13898) );
  INV_X1 U16008 ( .A(n13889), .ZN(n13890) );
  AOI21_X1 U16009 ( .B1(n13892), .B2(n13891), .A(n13890), .ZN(n14067) );
  AOI22_X1 U16010 ( .A1(n13894), .A2(n13968), .B1(n13966), .B2(n13893), .ZN(
        n13895) );
  OAI21_X1 U16011 ( .B1(n14067), .B2(n13896), .A(n13895), .ZN(n13897) );
  AOI21_X1 U16012 ( .B1(n13898), .B2(n13971), .A(n13897), .ZN(n14066) );
  INV_X1 U16013 ( .A(n13899), .ZN(n13900) );
  AOI211_X1 U16014 ( .C1(n14064), .C2(n13917), .A(n13974), .B(n13900), .ZN(
        n14063) );
  NOR2_X1 U16015 ( .A1(n13901), .A2(n13979), .ZN(n13905) );
  OAI22_X1 U16016 ( .A1(n13987), .A2(n13903), .B1(n13902), .B2(n13956), .ZN(
        n13904) );
  AOI211_X1 U16017 ( .C1(n14063), .C2(n13995), .A(n13905), .B(n13904), .ZN(
        n13908) );
  INV_X1 U16018 ( .A(n14067), .ZN(n13906) );
  NAND2_X1 U16019 ( .A1(n13906), .A2(n13993), .ZN(n13907) );
  OAI211_X1 U16020 ( .C1(n14066), .C2(n13909), .A(n13908), .B(n13907), .ZN(
        P2_U3247) );
  AOI21_X1 U16021 ( .B1(n13927), .B2(n13928), .A(n13911), .ZN(n13912) );
  XOR2_X1 U16022 ( .A(n13913), .B(n13912), .Z(n14070) );
  INV_X1 U16023 ( .A(n14070), .ZN(n13926) );
  XNOR2_X1 U16024 ( .A(n13914), .B(n13913), .ZN(n13916) );
  OAI21_X1 U16025 ( .B1(n13916), .B2(n13951), .A(n13915), .ZN(n14068) );
  NAND2_X1 U16026 ( .A1(n14068), .A2(n13987), .ZN(n13925) );
  INV_X1 U16027 ( .A(n13939), .ZN(n13919) );
  INV_X1 U16028 ( .A(n13917), .ZN(n13918) );
  AOI211_X1 U16029 ( .C1(n13920), .C2(n13919), .A(n13974), .B(n13918), .ZN(
        n14069) );
  AOI22_X1 U16030 ( .A1(n13909), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13921), 
        .B2(n13990), .ZN(n13922) );
  OAI21_X1 U16031 ( .B1(n14146), .B2(n13979), .A(n13922), .ZN(n13923) );
  AOI21_X1 U16032 ( .B1(n14069), .B2(n13995), .A(n13923), .ZN(n13924) );
  OAI211_X1 U16033 ( .C1(n13926), .C2(n13983), .A(n13925), .B(n13924), .ZN(
        P2_U3248) );
  XNOR2_X1 U16034 ( .A(n13927), .B(n13928), .ZN(n14077) );
  AOI21_X1 U16035 ( .B1(n13929), .B2(n13928), .A(n13951), .ZN(n13936) );
  OAI22_X1 U16036 ( .A1(n13933), .A2(n13932), .B1(n13931), .B2(n13930), .ZN(
        n13934) );
  AOI21_X1 U16037 ( .B1(n13936), .B2(n13935), .A(n13934), .ZN(n14076) );
  OAI21_X1 U16038 ( .B1(n13937), .B2(n13956), .A(n14076), .ZN(n13938) );
  NAND2_X1 U16039 ( .A1(n13938), .A2(n13987), .ZN(n13944) );
  AOI211_X1 U16040 ( .C1(n14074), .C2(n13953), .A(n13974), .B(n13939), .ZN(
        n14073) );
  OAI22_X1 U16041 ( .A1(n13941), .A2(n13979), .B1(n13940), .B2(n13987), .ZN(
        n13942) );
  AOI21_X1 U16042 ( .B1(n14073), .B2(n13995), .A(n13942), .ZN(n13943) );
  OAI211_X1 U16043 ( .C1(n14077), .C2(n13983), .A(n13944), .B(n13943), .ZN(
        P2_U3249) );
  INV_X1 U16044 ( .A(n13947), .ZN(n13946) );
  OAI21_X1 U16045 ( .B1(n7812), .B2(n13946), .A(n13945), .ZN(n14080) );
  INV_X1 U16046 ( .A(n14080), .ZN(n13963) );
  XOR2_X1 U16047 ( .A(n13948), .B(n13947), .Z(n13952) );
  INV_X1 U16048 ( .A(n13949), .ZN(n13950) );
  OAI21_X1 U16049 ( .B1(n13952), .B2(n13951), .A(n13950), .ZN(n14078) );
  NAND2_X1 U16050 ( .A1(n14078), .A2(n13987), .ZN(n13962) );
  INV_X1 U16051 ( .A(n13953), .ZN(n13954) );
  AOI211_X1 U16052 ( .C1(n13955), .C2(n13973), .A(n13974), .B(n13954), .ZN(
        n14079) );
  NOR2_X1 U16053 ( .A1(n7172), .A2(n13979), .ZN(n13960) );
  OAI22_X1 U16054 ( .A1(n13987), .A2(n13958), .B1(n13957), .B2(n13956), .ZN(
        n13959) );
  AOI211_X1 U16055 ( .C1(n14079), .C2(n13995), .A(n13960), .B(n13959), .ZN(
        n13961) );
  OAI211_X1 U16056 ( .C1(n13963), .C2(n13983), .A(n13962), .B(n13961), .ZN(
        P2_U3250) );
  INV_X1 U16057 ( .A(n13982), .ZN(n13965) );
  OAI21_X1 U16058 ( .B1(n13965), .B2(n6616), .A(n13964), .ZN(n13970) );
  AOI222_X1 U16059 ( .A1(n13971), .A2(n13970), .B1(n13969), .B2(n13968), .C1(
        n13967), .C2(n13966), .ZN(n14086) );
  INV_X1 U16060 ( .A(n13972), .ZN(n13975) );
  AOI211_X1 U16061 ( .C1(n14084), .C2(n13975), .A(n13974), .B(n7401), .ZN(
        n14083) );
  INV_X1 U16062 ( .A(n13976), .ZN(n13977) );
  AOI22_X1 U16063 ( .A1(n13909), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n13977), 
        .B2(n13990), .ZN(n13978) );
  OAI21_X1 U16064 ( .B1(n13980), .B2(n13979), .A(n13978), .ZN(n13985) );
  XNOR2_X1 U16065 ( .A(n13981), .B(n13982), .ZN(n14087) );
  NOR2_X1 U16066 ( .A1(n14087), .A2(n13983), .ZN(n13984) );
  AOI211_X1 U16067 ( .C1(n14083), .C2(n13995), .A(n13985), .B(n13984), .ZN(
        n13986) );
  OAI21_X1 U16068 ( .B1(n14086), .B2(n13909), .A(n13986), .ZN(P2_U3251) );
  MUX2_X1 U16069 ( .A(n13989), .B(n13988), .S(n13987), .Z(n13998) );
  AOI22_X1 U16070 ( .A1(n13991), .A2(n6645), .B1(n13990), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n13997) );
  AOI22_X1 U16071 ( .A1(n13995), .A2(n13994), .B1(n13993), .B2(n13992), .ZN(
        n13996) );
  NAND3_X1 U16072 ( .A1(n13998), .A2(n13997), .A3(n13996), .ZN(P2_U3264) );
  MUX2_X1 U16073 ( .A(n14117), .B(n14002), .S(n15567), .Z(n14003) );
  OAI21_X1 U16074 ( .B1(n7406), .B2(n14104), .A(n14003), .ZN(P2_U3529) );
  NOR3_X2 U16075 ( .A1(n14004), .A2(n14008), .A3(n14011), .ZN(n14015) );
  NOR3_X1 U16076 ( .A1(n14007), .A2(n14006), .A3(n14005), .ZN(n14013) );
  NAND3_X1 U16077 ( .A1(n14011), .A2(n14008), .A3(n14010), .ZN(n14009) );
  OAI211_X1 U16078 ( .C1(n14011), .C2(n14010), .A(n14009), .B(n15541), .ZN(
        n14012) );
  NAND2_X1 U16079 ( .A1(n14016), .A2(n15553), .ZN(n14017) );
  NAND2_X1 U16080 ( .A1(n14021), .A2(n15541), .ZN(n14024) );
  AOI21_X1 U16081 ( .B1(n15553), .B2(n14026), .A(n14025), .ZN(n14027) );
  OAI211_X1 U16082 ( .C1(n15557), .C2(n14029), .A(n14028), .B(n14027), .ZN(
        n14122) );
  MUX2_X1 U16083 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14122), .S(n14101), .Z(
        P2_U3525) );
  OAI211_X1 U16084 ( .C1(n15557), .C2(n14032), .A(n14031), .B(n14030), .ZN(
        n14123) );
  MUX2_X1 U16085 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14123), .S(n14101), .Z(
        n14033) );
  INV_X1 U16086 ( .A(n14033), .ZN(n14034) );
  OAI21_X1 U16087 ( .B1(n14126), .B2(n14104), .A(n14034), .ZN(P2_U3524) );
  AOI21_X1 U16088 ( .B1(n15553), .B2(n14036), .A(n14035), .ZN(n14037) );
  MUX2_X1 U16089 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14127), .S(n14101), .Z(
        P2_U3523) );
  INV_X1 U16090 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14046) );
  AOI211_X1 U16091 ( .C1(n14045), .C2(n15541), .A(n14044), .B(n14043), .ZN(
        n14130) );
  MUX2_X1 U16092 ( .A(n14046), .B(n14130), .S(n14101), .Z(n14047) );
  OAI21_X1 U16093 ( .B1(n14133), .B2(n14104), .A(n14047), .ZN(P2_U3521) );
  OAI211_X1 U16094 ( .C1(n15557), .C2(n14050), .A(n14049), .B(n14048), .ZN(
        n14134) );
  MUX2_X1 U16095 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14134), .S(n14101), .Z(
        n14051) );
  AOI21_X1 U16096 ( .B1(n14096), .B2(n7410), .A(n14051), .ZN(n14052) );
  INV_X1 U16097 ( .A(n14052), .ZN(P2_U3520) );
  OAI211_X1 U16098 ( .C1(n15557), .C2(n14055), .A(n14054), .B(n14053), .ZN(
        n14138) );
  MUX2_X1 U16099 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14138), .S(n14101), .Z(
        n14056) );
  AOI21_X1 U16100 ( .B1(n14096), .B2(n14140), .A(n14056), .ZN(n14057) );
  INV_X1 U16101 ( .A(n14057), .ZN(P2_U3519) );
  AOI21_X1 U16102 ( .B1(n15553), .B2(n14059), .A(n14058), .ZN(n14060) );
  OAI211_X1 U16103 ( .C1(n15557), .C2(n14062), .A(n14061), .B(n14060), .ZN(
        n14142) );
  MUX2_X1 U16104 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14142), .S(n14101), .Z(
        P2_U3518) );
  AOI21_X1 U16105 ( .B1(n15553), .B2(n14064), .A(n14063), .ZN(n14065) );
  OAI211_X1 U16106 ( .C1(n14067), .C2(n15546), .A(n14066), .B(n14065), .ZN(
        n14143) );
  MUX2_X1 U16107 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14143), .S(n14101), .Z(
        P2_U3517) );
  INV_X1 U16108 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14071) );
  AOI211_X1 U16109 ( .C1(n15541), .C2(n14070), .A(n14069), .B(n14068), .ZN(
        n14144) );
  MUX2_X1 U16110 ( .A(n14071), .B(n14144), .S(n14101), .Z(n14072) );
  OAI21_X1 U16111 ( .B1(n14146), .B2(n14104), .A(n14072), .ZN(P2_U3516) );
  AOI21_X1 U16112 ( .B1(n15553), .B2(n14074), .A(n14073), .ZN(n14075) );
  OAI211_X1 U16113 ( .C1(n15557), .C2(n14077), .A(n14076), .B(n14075), .ZN(
        n14147) );
  MUX2_X1 U16114 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14147), .S(n14101), .Z(
        P2_U3515) );
  INV_X1 U16115 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14081) );
  AOI211_X1 U16116 ( .C1(n15541), .C2(n14080), .A(n14079), .B(n14078), .ZN(
        n14148) );
  MUX2_X1 U16117 ( .A(n14081), .B(n14148), .S(n14101), .Z(n14082) );
  OAI21_X1 U16118 ( .B1(n7172), .B2(n14104), .A(n14082), .ZN(P2_U3514) );
  AOI21_X1 U16119 ( .B1(n15553), .B2(n14084), .A(n14083), .ZN(n14085) );
  OAI211_X1 U16120 ( .C1(n15557), .C2(n14087), .A(n14086), .B(n14085), .ZN(
        n14151) );
  MUX2_X1 U16121 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14151), .S(n14101), .Z(
        P2_U3513) );
  AOI21_X1 U16122 ( .B1(n15553), .B2(n14089), .A(n14088), .ZN(n14090) );
  OAI211_X1 U16123 ( .C1(n15557), .C2(n14092), .A(n14091), .B(n14090), .ZN(
        n14152) );
  MUX2_X1 U16124 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14152), .S(n14101), .Z(
        P2_U3512) );
  AOI211_X1 U16125 ( .C1(n15541), .C2(n14095), .A(n14094), .B(n14093), .ZN(
        n14156) );
  AOI22_X1 U16126 ( .A1(n14154), .A2(n14096), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n15567), .ZN(n14097) );
  OAI21_X1 U16127 ( .B1(n14156), .B2(n15567), .A(n14097), .ZN(P2_U3511) );
  INV_X1 U16128 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n14102) );
  AOI211_X1 U16129 ( .C1(n15541), .C2(n14100), .A(n14099), .B(n14098), .ZN(
        n14157) );
  MUX2_X1 U16130 ( .A(n14102), .B(n14157), .S(n14101), .Z(n14103) );
  OAI21_X1 U16131 ( .B1(n14161), .B2(n14104), .A(n14103), .ZN(P2_U3510) );
  AOI21_X1 U16132 ( .B1(n15553), .B2(n14106), .A(n14105), .ZN(n14108) );
  OAI211_X1 U16133 ( .C1(n15557), .C2(n14109), .A(n14108), .B(n14107), .ZN(
        n14162) );
  MUX2_X1 U16134 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14162), .S(n15564), .Z(
        P2_U3508) );
  AOI21_X1 U16135 ( .B1(n15553), .B2(n14111), .A(n14110), .ZN(n14113) );
  OAI211_X1 U16136 ( .C1(n15557), .C2(n14114), .A(n14113), .B(n14112), .ZN(
        n14163) );
  MUX2_X1 U16137 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n14163), .S(n15564), .Z(
        P2_U3507) );
  MUX2_X1 U16138 ( .A(n14118), .B(n14117), .S(n15561), .Z(n14119) );
  OAI21_X1 U16139 ( .B1(n7406), .B2(n14160), .A(n14119), .ZN(P2_U3497) );
  INV_X2 U16140 ( .A(n15559), .ZN(n15561) );
  MUX2_X1 U16141 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14122), .S(n15561), .Z(
        P2_U3493) );
  MUX2_X1 U16142 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14123), .S(n15561), .Z(
        n14124) );
  INV_X1 U16143 ( .A(n14124), .ZN(n14125) );
  OAI21_X1 U16144 ( .B1(n14126), .B2(n14160), .A(n14125), .ZN(P2_U3492) );
  INV_X1 U16145 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14131) );
  MUX2_X1 U16146 ( .A(n14131), .B(n14130), .S(n15561), .Z(n14132) );
  OAI21_X1 U16147 ( .B1(n14133), .B2(n14160), .A(n14132), .ZN(P2_U3489) );
  MUX2_X1 U16148 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14134), .S(n15561), .Z(
        n14135) );
  INV_X1 U16149 ( .A(n14135), .ZN(n14136) );
  OAI21_X1 U16150 ( .B1(n14137), .B2(n14160), .A(n14136), .ZN(P2_U3488) );
  INV_X1 U16151 ( .A(n14160), .ZN(n14153) );
  MUX2_X1 U16152 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14138), .S(n15561), .Z(
        n14139) );
  AOI21_X1 U16153 ( .B1(n14153), .B2(n14140), .A(n14139), .ZN(n14141) );
  INV_X1 U16154 ( .A(n14141), .ZN(P2_U3487) );
  MUX2_X1 U16155 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14142), .S(n15561), .Z(
        P2_U3486) );
  MUX2_X1 U16156 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14143), .S(n15561), .Z(
        P2_U3484) );
  MUX2_X1 U16157 ( .A(n7769), .B(n14144), .S(n15561), .Z(n14145) );
  OAI21_X1 U16158 ( .B1(n14146), .B2(n14160), .A(n14145), .ZN(P2_U3481) );
  MUX2_X1 U16159 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14147), .S(n15561), .Z(
        P2_U3478) );
  MUX2_X1 U16160 ( .A(n14149), .B(n14148), .S(n15561), .Z(n14150) );
  OAI21_X1 U16161 ( .B1(n7172), .B2(n14160), .A(n14150), .ZN(P2_U3475) );
  MUX2_X1 U16162 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14151), .S(n15561), .Z(
        P2_U3472) );
  MUX2_X1 U16163 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n14152), .S(n15561), .Z(
        P2_U3469) );
  AOI22_X1 U16164 ( .A1(n14154), .A2(n14153), .B1(P2_REG0_REG_12__SCAN_IN), 
        .B2(n15559), .ZN(n14155) );
  OAI21_X1 U16165 ( .B1(n14156), .B2(n15559), .A(n14155), .ZN(P2_U3466) );
  MUX2_X1 U16166 ( .A(n14158), .B(n14157), .S(n15561), .Z(n14159) );
  OAI21_X1 U16167 ( .B1(n14161), .B2(n14160), .A(n14159), .ZN(P2_U3463) );
  MUX2_X1 U16168 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n14162), .S(n15561), .Z(
        P2_U3457) );
  MUX2_X1 U16169 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n14163), .S(n15561), .Z(
        P2_U3454) );
  INV_X1 U16170 ( .A(n14164), .ZN(n14171) );
  OR2_X1 U16171 ( .A1(n14165), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n14167) );
  NOR4_X1 U16172 ( .A1(n14167), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14166), .A4(
        P2_U3088), .ZN(n14168) );
  AOI21_X1 U16173 ( .B1(n14169), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14168), 
        .ZN(n14170) );
  OAI21_X1 U16174 ( .B1(n14171), .B2(n6438), .A(n14170), .ZN(P2_U3296) );
  INV_X1 U16175 ( .A(n14172), .ZN(n15180) );
  OAI222_X1 U16176 ( .A1(n14174), .A2(P2_U3088), .B1(n6438), .B2(n15180), .C1(
        n14173), .C2(n14184), .ZN(P2_U3298) );
  NAND2_X1 U16177 ( .A1(n14176), .A2(n14175), .ZN(n14178) );
  OAI211_X1 U16178 ( .C1(n14179), .C2(n14184), .A(n14178), .B(n14177), .ZN(
        P2_U3299) );
  INV_X1 U16179 ( .A(n14180), .ZN(n15183) );
  OAI222_X1 U16180 ( .A1(n14184), .A2(n14182), .B1(n6438), .B2(n15183), .C1(
        n14181), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U16181 ( .A(n14183), .ZN(n15187) );
  OAI222_X1 U16182 ( .A1(P2_U3088), .A2(n14186), .B1(n6438), .B2(n15187), .C1(
        n14185), .C2(n14184), .ZN(P2_U3301) );
  INV_X1 U16183 ( .A(n14187), .ZN(n14188) );
  MUX2_X1 U16184 ( .A(n14188), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U16185 ( .A(n14189), .ZN(n14190) );
  AOI21_X1 U16186 ( .B1(n14192), .B2(n14191), .A(n14190), .ZN(n14198) );
  NAND2_X1 U16187 ( .A1(n15221), .A2(n15223), .ZN(n14193) );
  OAI21_X1 U16188 ( .B1(n14975), .B2(n15052), .A(n14193), .ZN(n15004) );
  AOI21_X1 U16189 ( .B1(n15004), .B2(n14368), .A(n14194), .ZN(n14195) );
  OAI21_X1 U16190 ( .B1(n14353), .B2(n15007), .A(n14195), .ZN(n14196) );
  AOI21_X1 U16191 ( .B1(n15151), .B2(n14357), .A(n14196), .ZN(n14197) );
  OAI21_X1 U16192 ( .B1(n14198), .B2(n14359), .A(n14197), .ZN(P1_U3215) );
  INV_X1 U16193 ( .A(n15104), .ZN(n14211) );
  OR2_X1 U16194 ( .A1(n14240), .A2(n14199), .ZN(n14201) );
  NAND2_X1 U16195 ( .A1(n14201), .A2(n14200), .ZN(n14332) );
  INV_X1 U16196 ( .A(n14202), .ZN(n14204) );
  NOR3_X1 U16197 ( .A1(n14332), .A2(n14204), .A3(n14203), .ZN(n14205) );
  OAI21_X1 U16198 ( .B1(n14205), .B2(n6445), .A(n14370), .ZN(n14210) );
  OAI22_X1 U16199 ( .A1(n14266), .A2(n15052), .B1(n14241), .B2(n14976), .ZN(
        n14853) );
  INV_X1 U16200 ( .A(n14857), .ZN(n14207) );
  OAI22_X1 U16201 ( .A1(n14207), .A2(n14291), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14206), .ZN(n14208) );
  AOI21_X1 U16202 ( .B1(n14853), .B2(n14368), .A(n14208), .ZN(n14209) );
  OAI211_X1 U16203 ( .C1(n14211), .C2(n14380), .A(n14210), .B(n14209), .ZN(
        P1_U3216) );
  OAI211_X1 U16204 ( .C1(n14214), .C2(n14213), .A(n14212), .B(n14370), .ZN(
        n14218) );
  NAND2_X1 U16205 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(n6428), .ZN(n14734) );
  OAI21_X1 U16206 ( .B1(n14374), .B2(n15053), .A(n14734), .ZN(n14216) );
  NOR2_X1 U16207 ( .A1(n14291), .A2(n15056), .ZN(n14215) );
  AOI211_X1 U16208 ( .C1(n14377), .C2(n15048), .A(n14216), .B(n14215), .ZN(
        n14217) );
  OAI211_X1 U16209 ( .C1(n15058), .C2(n14380), .A(n14218), .B(n14217), .ZN(
        P1_U3217) );
  XNOR2_X1 U16210 ( .A(n14220), .B(n14219), .ZN(n14351) );
  NOR2_X1 U16211 ( .A1(n14352), .A2(n14351), .ZN(n14350) );
  NOR2_X1 U16212 ( .A1(n14350), .A2(n14221), .ZN(n14225) );
  XNOR2_X1 U16213 ( .A(n14223), .B(n14222), .ZN(n14224) );
  NAND2_X1 U16214 ( .A1(n14225), .A2(n14224), .ZN(n14310) );
  OAI211_X1 U16215 ( .C1(n14225), .C2(n14224), .A(n14310), .B(n14370), .ZN(
        n14229) );
  NOR2_X1 U16216 ( .A1(n14291), .A2(n14927), .ZN(n14227) );
  NAND2_X1 U16217 ( .A1(n6428), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14788) );
  OAI21_X1 U16218 ( .B1(n14923), .B2(n14374), .A(n14788), .ZN(n14226) );
  AOI211_X1 U16219 ( .C1(n14377), .C2(n14645), .A(n14227), .B(n14226), .ZN(
        n14228) );
  OAI211_X1 U16220 ( .C1(n14931), .C2(n14380), .A(n14229), .B(n14228), .ZN(
        P1_U3219) );
  OAI21_X1 U16221 ( .B1(n14232), .B2(n14231), .A(n14230), .ZN(n14233) );
  NAND2_X1 U16222 ( .A1(n14233), .A2(n14370), .ZN(n14238) );
  AOI22_X1 U16223 ( .A1(n14336), .A2(n11381), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14234), .ZN(n14237) );
  NAND2_X1 U16224 ( .A1(n14357), .A2(n11370), .ZN(n14236) );
  NAND2_X1 U16225 ( .A1(n14377), .A2(n11377), .ZN(n14235) );
  NAND4_X1 U16226 ( .A1(n14238), .A2(n14237), .A3(n14236), .A4(n14235), .ZN(
        P1_U3222) );
  AOI21_X1 U16227 ( .B1(n14240), .B2(n14239), .A(n7817), .ZN(n14249) );
  AND2_X1 U16228 ( .A1(n14889), .A2(n15400), .ZN(n15116) );
  INV_X1 U16229 ( .A(n14308), .ZN(n14247) );
  OAI22_X1 U16230 ( .A1(n14241), .A2(n15052), .B1(n14923), .B2(n14976), .ZN(
        n15115) );
  INV_X1 U16231 ( .A(n15115), .ZN(n14245) );
  AOI22_X1 U16232 ( .A1(n14893), .A2(n14242), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(n6428), .ZN(n14243) );
  OAI21_X1 U16233 ( .B1(n14245), .B2(n14244), .A(n14243), .ZN(n14246) );
  AOI21_X1 U16234 ( .B1(n15116), .B2(n14247), .A(n14246), .ZN(n14248) );
  OAI21_X1 U16235 ( .B1(n14249), .B2(n14359), .A(n14248), .ZN(P1_U3223) );
  INV_X1 U16236 ( .A(n15230), .ZN(n15239) );
  AOI21_X1 U16237 ( .B1(n14251), .B2(n14250), .A(n14359), .ZN(n14253) );
  NAND2_X1 U16238 ( .A1(n14253), .A2(n14252), .ZN(n14258) );
  OAI21_X1 U16239 ( .B1(n14374), .B2(n14443), .A(n14254), .ZN(n14256) );
  NOR2_X1 U16240 ( .A1(n14353), .A2(n15228), .ZN(n14255) );
  AOI211_X1 U16241 ( .C1(n14377), .C2(n15224), .A(n14256), .B(n14255), .ZN(
        n14257) );
  OAI211_X1 U16242 ( .C1(n15239), .C2(n14380), .A(n14258), .B(n14257), .ZN(
        P1_U3224) );
  INV_X1 U16243 ( .A(n14259), .ZN(n14300) );
  INV_X1 U16244 ( .A(n14260), .ZN(n14262) );
  NOR3_X1 U16245 ( .A1(n14300), .A2(n14262), .A3(n14261), .ZN(n14265) );
  INV_X1 U16246 ( .A(n14263), .ZN(n14264) );
  OAI21_X1 U16247 ( .B1(n14265), .B2(n14264), .A(n14370), .ZN(n14273) );
  NOR2_X1 U16248 ( .A1(n14266), .A2(n14976), .ZN(n14267) );
  AOI21_X1 U16249 ( .B1(n14639), .B2(n15222), .A(n14267), .ZN(n14820) );
  INV_X1 U16250 ( .A(n14820), .ZN(n14271) );
  INV_X1 U16251 ( .A(n14268), .ZN(n14823) );
  OAI22_X1 U16252 ( .A1(n14823), .A2(n14353), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14269), .ZN(n14270) );
  AOI21_X1 U16253 ( .B1(n14271), .B2(n14368), .A(n14270), .ZN(n14272) );
  OAI211_X1 U16254 ( .C1(n15093), .C2(n14308), .A(n14273), .B(n14272), .ZN(
        P1_U3225) );
  XOR2_X1 U16255 ( .A(n14275), .B(n14276), .Z(n14373) );
  INV_X1 U16256 ( .A(n14274), .ZN(n14372) );
  NAND2_X1 U16257 ( .A1(n14373), .A2(n14372), .ZN(n14371) );
  OAI21_X1 U16258 ( .B1(n14276), .B2(n14275), .A(n14371), .ZN(n14280) );
  XOR2_X1 U16259 ( .A(n14278), .B(n14277), .Z(n14279) );
  XNOR2_X1 U16260 ( .A(n14280), .B(n14279), .ZN(n14286) );
  OAI21_X1 U16261 ( .B1(n14374), .B2(n14974), .A(n14281), .ZN(n14282) );
  AOI21_X1 U16262 ( .B1(n14377), .B2(n14647), .A(n14282), .ZN(n14283) );
  OAI21_X1 U16263 ( .B1(n14291), .B2(n14979), .A(n14283), .ZN(n14284) );
  AOI21_X1 U16264 ( .B1(n15142), .B2(n14357), .A(n14284), .ZN(n14285) );
  OAI21_X1 U16265 ( .B1(n14286), .B2(n14359), .A(n14285), .ZN(P1_U3226) );
  XNOR2_X1 U16266 ( .A(n14288), .B(n14287), .ZN(n14289) );
  XNOR2_X1 U16267 ( .A(n14290), .B(n14289), .ZN(n14296) );
  NOR2_X1 U16268 ( .A1(n14291), .A2(n14959), .ZN(n14294) );
  NAND2_X1 U16269 ( .A1(n14377), .A2(n14987), .ZN(n14292) );
  NAND2_X1 U16270 ( .A1(n6428), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14746) );
  OAI211_X1 U16271 ( .C1(n14957), .C2(n14374), .A(n14292), .B(n14746), .ZN(
        n14293) );
  AOI211_X1 U16272 ( .C1(n15137), .C2(n14357), .A(n14294), .B(n14293), .ZN(
        n14295) );
  OAI21_X1 U16273 ( .B1(n14296), .B2(n14359), .A(n14295), .ZN(P1_U3228) );
  NAND2_X1 U16274 ( .A1(n14838), .A2(n15400), .ZN(n15098) );
  INV_X1 U16275 ( .A(n14297), .ZN(n14299) );
  NOR3_X1 U16276 ( .A1(n6445), .A2(n14299), .A3(n14298), .ZN(n14301) );
  OAI21_X1 U16277 ( .B1(n14301), .B2(n14300), .A(n14370), .ZN(n14307) );
  AND2_X1 U16278 ( .A1(n14871), .A2(n15223), .ZN(n14302) );
  AOI21_X1 U16279 ( .B1(n14640), .B2(n15222), .A(n14302), .ZN(n15100) );
  INV_X1 U16280 ( .A(n15100), .ZN(n14305) );
  OAI22_X1 U16281 ( .A1(n14841), .A2(n14291), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14303), .ZN(n14304) );
  AOI21_X1 U16282 ( .B1(n14305), .B2(n14368), .A(n14304), .ZN(n14306) );
  OAI211_X1 U16283 ( .C1(n15098), .C2(n14308), .A(n14307), .B(n14306), .ZN(
        P1_U3229) );
  NAND2_X1 U16284 ( .A1(n14310), .A2(n14309), .ZN(n14312) );
  XNOR2_X1 U16285 ( .A(n14312), .B(n14311), .ZN(n14319) );
  OAI22_X1 U16286 ( .A1(n14901), .A2(n14374), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14313), .ZN(n14314) );
  AOI21_X1 U16287 ( .B1(n14377), .B2(n14644), .A(n14314), .ZN(n14315) );
  OAI21_X1 U16288 ( .B1(n14353), .B2(n14316), .A(n14315), .ZN(n14317) );
  AOI21_X1 U16289 ( .B1(n15122), .B2(n14357), .A(n14317), .ZN(n14318) );
  OAI21_X1 U16290 ( .B1(n14319), .B2(n14359), .A(n14318), .ZN(P1_U3233) );
  OAI211_X1 U16291 ( .C1(n14322), .C2(n14321), .A(n14320), .B(n14370), .ZN(
        n14328) );
  OAI21_X1 U16292 ( .B1(n14374), .B2(n14324), .A(n14323), .ZN(n14326) );
  NOR2_X1 U16293 ( .A1(n14291), .A2(n15033), .ZN(n14325) );
  AOI211_X1 U16294 ( .C1(n14377), .C2(n15027), .A(n14326), .B(n14325), .ZN(
        n14327) );
  OAI211_X1 U16295 ( .C1(n15252), .C2(n14380), .A(n14328), .B(n14327), .ZN(
        P1_U3234) );
  INV_X1 U16296 ( .A(n14329), .ZN(n14331) );
  NOR3_X1 U16297 ( .A1(n7817), .A2(n14331), .A3(n14330), .ZN(n14333) );
  OAI21_X1 U16298 ( .B1(n14333), .B2(n14332), .A(n14370), .ZN(n14338) );
  AOI22_X1 U16299 ( .A1(n14870), .A2(n14377), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14334) );
  OAI21_X1 U16300 ( .B1(n14353), .B2(n14875), .A(n14334), .ZN(n14335) );
  AOI21_X1 U16301 ( .B1(n14336), .B2(n14871), .A(n14335), .ZN(n14337) );
  OAI211_X1 U16302 ( .C1(n14380), .C2(n14878), .A(n14338), .B(n14337), .ZN(
        P1_U3235) );
  INV_X1 U16303 ( .A(n14339), .ZN(n14340) );
  AOI21_X1 U16304 ( .B1(n14342), .B2(n14341), .A(n14340), .ZN(n14349) );
  NOR2_X1 U16305 ( .A1(n14353), .A2(n14343), .ZN(n14347) );
  NAND2_X1 U16306 ( .A1(n14377), .A2(n14437), .ZN(n14345) );
  OAI211_X1 U16307 ( .C1(n14445), .C2(n14374), .A(n14345), .B(n14344), .ZN(
        n14346) );
  AOI211_X1 U16308 ( .C1(n14438), .C2(n14357), .A(n14347), .B(n14346), .ZN(
        n14348) );
  OAI21_X1 U16309 ( .B1(n14349), .B2(n14359), .A(n14348), .ZN(P1_U3236) );
  AOI21_X1 U16310 ( .B1(n14352), .B2(n14351), .A(n14350), .ZN(n14360) );
  NOR2_X1 U16311 ( .A1(n14353), .A2(n14938), .ZN(n14356) );
  NAND2_X1 U16312 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14758)
         );
  NAND2_X1 U16313 ( .A1(n14377), .A2(n14646), .ZN(n14354) );
  OAI211_X1 U16314 ( .C1(n14944), .C2(n14374), .A(n14758), .B(n14354), .ZN(
        n14355) );
  AOI211_X1 U16315 ( .C1(n15131), .C2(n14357), .A(n14356), .B(n14355), .ZN(
        n14358) );
  OAI21_X1 U16316 ( .B1(n14360), .B2(n14359), .A(n14358), .ZN(P1_U3238) );
  OAI21_X1 U16317 ( .B1(n14363), .B2(n14362), .A(n14361), .ZN(n14364) );
  OAI22_X1 U16318 ( .A1(n14365), .A2(n15052), .B1(n14802), .B2(n14976), .ZN(
        n14804) );
  OAI22_X1 U16319 ( .A1(n14808), .A2(n14291), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14366), .ZN(n14367) );
  AOI21_X1 U16320 ( .B1(n14804), .B2(n14368), .A(n14367), .ZN(n14369) );
  OAI211_X1 U16321 ( .C1(n14373), .C2(n14372), .A(n14371), .B(n14370), .ZN(
        n14379) );
  NAND2_X1 U16322 ( .A1(n6428), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15317) );
  OAI21_X1 U16323 ( .B1(n14374), .B2(n14956), .A(n15317), .ZN(n14376) );
  NOR2_X1 U16324 ( .A1(n14291), .A2(n14992), .ZN(n14375) );
  AOI211_X1 U16325 ( .C1(n14377), .C2(n15026), .A(n14376), .B(n14375), .ZN(
        n14378) );
  OAI211_X1 U16326 ( .C1(n14995), .C2(n14380), .A(n14379), .B(n14378), .ZN(
        P1_U3241) );
  NAND2_X1 U16327 ( .A1(n14381), .A2(n14575), .ZN(n14382) );
  MUX2_X1 U16328 ( .A(n14638), .B(n15082), .S(n14549), .Z(n14529) );
  XNOR2_X1 U16329 ( .A(n14385), .B(n14467), .ZN(n14386) );
  OAI211_X1 U16330 ( .C1(n14388), .C2(n14387), .A(n14583), .B(n14386), .ZN(
        n14393) );
  INV_X1 U16331 ( .A(n14389), .ZN(n14390) );
  MUX2_X1 U16332 ( .A(n14391), .B(n14390), .S(n14467), .Z(n14392) );
  NAND2_X1 U16333 ( .A1(n14393), .A2(n14392), .ZN(n14394) );
  NAND2_X1 U16334 ( .A1(n14541), .A2(n15330), .ZN(n14396) );
  NAND2_X1 U16335 ( .A1(n14467), .A2(n15348), .ZN(n14395) );
  MUX2_X1 U16336 ( .A(n14396), .B(n14395), .S(n11381), .Z(n14397) );
  NAND2_X1 U16337 ( .A1(n14398), .A2(n14467), .ZN(n14401) );
  NAND2_X1 U16338 ( .A1(n14652), .A2(n14446), .ZN(n14400) );
  MUX2_X1 U16339 ( .A(n14401), .B(n14400), .S(n14399), .Z(n14402) );
  MUX2_X1 U16340 ( .A(n14404), .B(n14651), .S(n14530), .Z(n14403) );
  INV_X1 U16341 ( .A(n14403), .ZN(n14406) );
  MUX2_X1 U16342 ( .A(n14651), .B(n14404), .S(n14530), .Z(n14405) );
  NAND2_X1 U16343 ( .A1(n14407), .A2(n14406), .ZN(n14408) );
  MUX2_X1 U16344 ( .A(n14650), .B(n15355), .S(n14530), .Z(n14411) );
  MUX2_X1 U16345 ( .A(n15355), .B(n14650), .S(n14530), .Z(n14410) );
  INV_X1 U16346 ( .A(n14411), .ZN(n14412) );
  MUX2_X1 U16347 ( .A(n14413), .B(n14649), .S(n14530), .Z(n14416) );
  MUX2_X1 U16348 ( .A(n14649), .B(n14413), .S(n14530), .Z(n14414) );
  INV_X1 U16349 ( .A(n14416), .ZN(n14417) );
  MUX2_X1 U16350 ( .A(n14419), .B(n14418), .S(n14549), .Z(n14422) );
  MUX2_X1 U16351 ( .A(n14419), .B(n14418), .S(n14530), .Z(n14420) );
  MUX2_X1 U16352 ( .A(n14648), .B(n14424), .S(n14549), .Z(n14426) );
  MUX2_X1 U16353 ( .A(n14648), .B(n14424), .S(n14530), .Z(n14425) );
  INV_X1 U16354 ( .A(n14426), .ZN(n14427) );
  MUX2_X1 U16355 ( .A(n15048), .B(n14428), .S(n14530), .Z(n14432) );
  MUX2_X1 U16356 ( .A(n15048), .B(n14428), .S(n14549), .Z(n14429) );
  NAND2_X1 U16357 ( .A1(n14430), .A2(n14429), .ZN(n14436) );
  INV_X1 U16358 ( .A(n14431), .ZN(n14434) );
  INV_X1 U16359 ( .A(n14432), .ZN(n14433) );
  NAND2_X1 U16360 ( .A1(n14434), .A2(n14433), .ZN(n14435) );
  MUX2_X1 U16361 ( .A(n14437), .B(n15399), .S(n14446), .Z(n14441) );
  MUX2_X1 U16362 ( .A(n15053), .B(n15259), .S(n14530), .Z(n14448) );
  MUX2_X1 U16363 ( .A(n15224), .B(n14438), .S(n14446), .Z(n14447) );
  MUX2_X1 U16364 ( .A(n14439), .B(n15058), .S(n14530), .Z(n14440) );
  AND2_X1 U16365 ( .A1(n14471), .A2(n14442), .ZN(n14456) );
  MUX2_X1 U16366 ( .A(n14443), .B(n15252), .S(n14530), .Z(n14459) );
  OR2_X1 U16367 ( .A1(n15036), .A2(n14530), .ZN(n14460) );
  NAND2_X1 U16368 ( .A1(n14443), .A2(n14530), .ZN(n14454) );
  NAND3_X1 U16369 ( .A1(n14459), .A2(n14460), .A3(n14454), .ZN(n14444) );
  AND2_X1 U16370 ( .A1(n14456), .A2(n14444), .ZN(n14458) );
  MUX2_X1 U16371 ( .A(n14445), .B(n15239), .S(n14530), .Z(n14451) );
  MUX2_X1 U16372 ( .A(n15027), .B(n15230), .S(n14446), .Z(n14450) );
  AOI22_X1 U16373 ( .A1(n14451), .A2(n14450), .B1(n14448), .B2(n14447), .ZN(
        n14449) );
  INV_X1 U16374 ( .A(n14450), .ZN(n14453) );
  INV_X1 U16375 ( .A(n14451), .ZN(n14452) );
  AND2_X1 U16376 ( .A1(n14453), .A2(n14452), .ZN(n14457) );
  OAI21_X1 U16377 ( .B1(n14459), .B2(n14454), .A(n15011), .ZN(n14455) );
  INV_X1 U16378 ( .A(n14459), .ZN(n14462) );
  INV_X1 U16379 ( .A(n14460), .ZN(n14461) );
  NAND2_X1 U16380 ( .A1(n14462), .A2(n14461), .ZN(n14463) );
  OAI211_X1 U16381 ( .C1(n15011), .C2(n14467), .A(n14466), .B(n14463), .ZN(
        n14464) );
  INV_X1 U16382 ( .A(n14464), .ZN(n14465) );
  OAI21_X1 U16383 ( .B1(n15010), .B2(n15026), .A(n14466), .ZN(n14468) );
  INV_X1 U16384 ( .A(n14467), .ZN(n14549) );
  NAND2_X1 U16385 ( .A1(n14468), .A2(n14549), .ZN(n14469) );
  INV_X1 U16386 ( .A(n15142), .ZN(n14470) );
  MUX2_X1 U16387 ( .A(n14956), .B(n14470), .S(n14549), .Z(n14483) );
  MUX2_X1 U16388 ( .A(n14987), .B(n15142), .S(n14467), .Z(n14482) );
  INV_X1 U16389 ( .A(n14471), .ZN(n14472) );
  AOI22_X1 U16390 ( .A1(n14483), .A2(n14482), .B1(n14472), .B2(n14549), .ZN(
        n14473) );
  MUX2_X1 U16391 ( .A(n14475), .B(n14474), .S(n14467), .Z(n14478) );
  OAI21_X1 U16392 ( .B1(n14643), .B2(n15122), .A(n14476), .ZN(n14477) );
  AND2_X1 U16393 ( .A1(n14478), .A2(n14477), .ZN(n14500) );
  NAND2_X1 U16394 ( .A1(n14974), .A2(n14530), .ZN(n14489) );
  NAND2_X1 U16395 ( .A1(n14596), .A2(n14489), .ZN(n14479) );
  NAND3_X1 U16396 ( .A1(n14492), .A2(n14496), .A3(n14479), .ZN(n14481) );
  NOR2_X1 U16397 ( .A1(n15137), .A2(n14467), .ZN(n14494) );
  NAND2_X1 U16398 ( .A1(n14496), .A2(n14494), .ZN(n14480) );
  NAND2_X1 U16399 ( .A1(n14481), .A2(n14480), .ZN(n14487) );
  INV_X1 U16400 ( .A(n14482), .ZN(n14485) );
  INV_X1 U16401 ( .A(n14483), .ZN(n14484) );
  NAND2_X1 U16402 ( .A1(n14485), .A2(n14484), .ZN(n14486) );
  NAND4_X1 U16403 ( .A1(n14488), .A2(n14500), .A3(n14487), .A4(n14486), .ZN(
        n14505) );
  NOR2_X1 U16404 ( .A1(n14598), .A2(n14489), .ZN(n14490) );
  NAND2_X1 U16405 ( .A1(n14492), .A2(n14490), .ZN(n14491) );
  OAI21_X1 U16406 ( .B1(n14492), .B2(n14467), .A(n14491), .ZN(n14498) );
  INV_X1 U16407 ( .A(n14598), .ZN(n14493) );
  NAND3_X1 U16408 ( .A1(n14496), .A2(n14494), .A3(n14493), .ZN(n14495) );
  OAI21_X1 U16409 ( .B1(n14541), .B2(n14496), .A(n14495), .ZN(n14497) );
  NAND2_X1 U16410 ( .A1(n14500), .A2(n14499), .ZN(n14504) );
  NOR2_X1 U16411 ( .A1(n14923), .A2(n14467), .ZN(n14502) );
  OAI21_X1 U16412 ( .B1(n14549), .B2(n14643), .A(n15122), .ZN(n14501) );
  OAI21_X1 U16413 ( .B1(n14502), .B2(n15122), .A(n14501), .ZN(n14503) );
  NAND3_X1 U16414 ( .A1(n14505), .A2(n14504), .A3(n14503), .ZN(n14508) );
  INV_X1 U16415 ( .A(n14889), .ZN(n14895) );
  MUX2_X1 U16416 ( .A(n14901), .B(n14895), .S(n14549), .Z(n14507) );
  MUX2_X1 U16417 ( .A(n14870), .B(n14889), .S(n14467), .Z(n14506) );
  OAI21_X1 U16418 ( .B1(n14508), .B2(n14507), .A(n14506), .ZN(n14510) );
  NAND2_X1 U16419 ( .A1(n14508), .A2(n14507), .ZN(n14509) );
  MUX2_X1 U16420 ( .A(n15111), .B(n14642), .S(n14549), .Z(n14512) );
  MUX2_X1 U16421 ( .A(n15111), .B(n14642), .S(n14467), .Z(n14511) );
  INV_X1 U16422 ( .A(n14512), .ZN(n14513) );
  MUX2_X1 U16423 ( .A(n14871), .B(n15104), .S(n14549), .Z(n14515) );
  MUX2_X1 U16424 ( .A(n14871), .B(n15104), .S(n14467), .Z(n14514) );
  INV_X1 U16425 ( .A(n14515), .ZN(n14516) );
  MUX2_X1 U16426 ( .A(n14641), .B(n14838), .S(n14467), .Z(n14518) );
  MUX2_X1 U16427 ( .A(n14641), .B(n14838), .S(n14549), .Z(n14517) );
  MUX2_X1 U16428 ( .A(n14640), .B(n14829), .S(n14549), .Z(n14520) );
  MUX2_X1 U16429 ( .A(n14640), .B(n14829), .S(n14467), .Z(n14519) );
  INV_X1 U16430 ( .A(n14520), .ZN(n14521) );
  MUX2_X1 U16431 ( .A(n14639), .B(n15087), .S(n14467), .Z(n14524) );
  MUX2_X1 U16432 ( .A(n14522), .B(n14811), .S(n14549), .Z(n14523) );
  MUX2_X1 U16433 ( .A(n14638), .B(n15082), .S(n14467), .Z(n14526) );
  MUX2_X1 U16434 ( .A(n14637), .B(n15077), .S(n14530), .Z(n14532) );
  MUX2_X1 U16435 ( .A(n14637), .B(n15077), .S(n14549), .Z(n14531) );
  INV_X1 U16436 ( .A(n14532), .ZN(n14533) );
  XNOR2_X1 U16437 ( .A(n14534), .B(n14634), .ZN(n14609) );
  INV_X1 U16438 ( .A(n14535), .ZN(n14536) );
  NAND2_X1 U16439 ( .A1(n14537), .A2(n14536), .ZN(n14539) );
  AND2_X1 U16440 ( .A1(n14539), .A2(n14538), .ZN(n14554) );
  NAND2_X1 U16441 ( .A1(n14609), .A2(n14554), .ZN(n14573) );
  OAI21_X1 U16442 ( .B1(n14634), .B2(n14540), .A(n14635), .ZN(n14542) );
  MUX2_X1 U16443 ( .A(n14542), .B(n15066), .S(n14541), .Z(n14553) );
  INV_X1 U16444 ( .A(n14635), .ZN(n14547) );
  AOI22_X1 U16445 ( .A1(n14634), .A2(n14549), .B1(n14544), .B2(n14543), .ZN(
        n14546) );
  INV_X1 U16446 ( .A(n15066), .ZN(n14800) );
  NAND2_X1 U16447 ( .A1(n14800), .A2(n14467), .ZN(n14545) );
  OAI21_X1 U16448 ( .B1(n14547), .B2(n14546), .A(n14545), .ZN(n14552) );
  NOR2_X1 U16449 ( .A1(n14553), .A2(n14552), .ZN(n14569) );
  NOR2_X1 U16450 ( .A1(n14573), .A2(n14569), .ZN(n14564) );
  MUX2_X1 U16451 ( .A(n14548), .B(n15070), .S(n14467), .Z(n14557) );
  MUX2_X1 U16452 ( .A(n14636), .B(n14550), .S(n14549), .Z(n14556) );
  AND2_X1 U16453 ( .A1(n14557), .A2(n14556), .ZN(n14561) );
  NOR3_X1 U16454 ( .A1(n14551), .A2(n14564), .A3(n14561), .ZN(n14633) );
  AND2_X1 U16455 ( .A1(n14553), .A2(n14552), .ZN(n14568) );
  NAND2_X1 U16456 ( .A1(n14634), .A2(n14467), .ZN(n14619) );
  INV_X1 U16457 ( .A(n14554), .ZN(n14622) );
  AND2_X1 U16458 ( .A1(n14622), .A2(n14614), .ZN(n14620) );
  NOR2_X1 U16459 ( .A1(n14634), .A2(n14467), .ZN(n14618) );
  NAND2_X1 U16460 ( .A1(n14534), .A2(n14618), .ZN(n14555) );
  OAI211_X1 U16461 ( .C1(n14534), .C2(n14619), .A(n14620), .B(n14555), .ZN(
        n14571) );
  INV_X1 U16462 ( .A(n14556), .ZN(n14559) );
  INV_X1 U16463 ( .A(n14557), .ZN(n14558) );
  NAND2_X1 U16464 ( .A1(n14559), .A2(n14558), .ZN(n14563) );
  AOI21_X1 U16465 ( .B1(n14562), .B2(n14561), .A(n14560), .ZN(n14566) );
  INV_X1 U16466 ( .A(n14568), .ZN(n14572) );
  INV_X1 U16467 ( .A(n14569), .ZN(n14570) );
  OAI22_X1 U16468 ( .A1(n14573), .A2(n14572), .B1(n14571), .B2(n14570), .ZN(
        n14580) );
  AOI21_X1 U16469 ( .B1(n14627), .B2(n14575), .A(n14574), .ZN(n14579) );
  NAND3_X1 U16470 ( .A1(n14577), .A2(n14576), .A3(n15223), .ZN(n14578) );
  AOI22_X1 U16471 ( .A1(n14580), .A2(n14627), .B1(n14579), .B2(n14578), .ZN(
        n14631) );
  XOR2_X1 U16472 ( .A(n14635), .B(n15066), .Z(n14608) );
  INV_X1 U16473 ( .A(n14999), .ZN(n14986) );
  NAND4_X1 U16474 ( .A1(n14585), .A2(n14584), .A3(n14583), .A4(n14582), .ZN(
        n14587) );
  NOR2_X1 U16475 ( .A1(n14587), .A2(n14586), .ZN(n14591) );
  NAND4_X1 U16476 ( .A1(n14591), .A2(n14590), .A3(n14589), .A4(n14588), .ZN(
        n14594) );
  OR4_X1 U16477 ( .A1(n14594), .A2(n14593), .A3(n14592), .A4(n15046), .ZN(
        n14595) );
  NOR4_X1 U16478 ( .A1(n14986), .A2(n15218), .A3(n15022), .A4(n14595), .ZN(
        n14599) );
  INV_X1 U16479 ( .A(n14596), .ZN(n14597) );
  NAND4_X1 U16480 ( .A1(n14599), .A2(n7743), .A3(n15011), .A4(n14962), .ZN(
        n14600) );
  NOR4_X1 U16481 ( .A1(n14601), .A2(n14921), .A3(n14942), .A4(n14600), .ZN(
        n14602) );
  NAND4_X1 U16482 ( .A1(n14602), .A2(n14863), .A3(n14886), .A4(n14909), .ZN(
        n14604) );
  NOR4_X1 U16484 ( .A1(n14814), .A2(n14604), .A3(n14830), .A4(n7632), .ZN(
        n14606) );
  NAND4_X1 U16485 ( .A1(n14608), .A2(n14607), .A3(n14606), .A4(n14605), .ZN(
        n14612) );
  INV_X1 U16486 ( .A(n14609), .ZN(n14611) );
  XNOR2_X1 U16487 ( .A(n14613), .B(n14381), .ZN(n14615) );
  NOR2_X1 U16488 ( .A1(n14615), .A2(n14614), .ZN(n14629) );
  INV_X1 U16489 ( .A(n14634), .ZN(n14616) );
  AOI21_X1 U16490 ( .B1(n14616), .B2(n14620), .A(n14618), .ZN(n14617) );
  AOI21_X1 U16491 ( .B1(n14618), .B2(n14622), .A(n14617), .ZN(n14626) );
  INV_X1 U16492 ( .A(n14619), .ZN(n14623) );
  AOI21_X1 U16493 ( .B1(n14620), .B2(n14634), .A(n14623), .ZN(n14621) );
  AOI21_X1 U16494 ( .B1(n14623), .B2(n14622), .A(n14621), .ZN(n14625) );
  MUX2_X1 U16495 ( .A(n14626), .B(n14625), .S(n14624), .Z(n14628) );
  OAI211_X1 U16496 ( .C1(n14633), .C2(n14632), .A(n14631), .B(n14630), .ZN(
        P1_U3242) );
  MUX2_X1 U16497 ( .A(n14634), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14653), .Z(
        P1_U3591) );
  MUX2_X1 U16498 ( .A(n14635), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14653), .Z(
        P1_U3590) );
  MUX2_X1 U16499 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14636), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16500 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14637), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16501 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14638), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16502 ( .A(n14639), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14653), .Z(
        P1_U3586) );
  MUX2_X1 U16503 ( .A(n14640), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14653), .Z(
        P1_U3585) );
  MUX2_X1 U16504 ( .A(n14641), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14653), .Z(
        P1_U3584) );
  MUX2_X1 U16505 ( .A(n14871), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14653), .Z(
        P1_U3583) );
  MUX2_X1 U16506 ( .A(n14642), .B(P1_DATAO_REG_22__SCAN_IN), .S(n14653), .Z(
        P1_U3582) );
  MUX2_X1 U16507 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14870), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16508 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14643), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16509 ( .A(n14644), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14653), .Z(
        P1_U3579) );
  MUX2_X1 U16510 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14645), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16511 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14646), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16512 ( .A(n14987), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14653), .Z(
        P1_U3576) );
  MUX2_X1 U16513 ( .A(n14647), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14653), .Z(
        P1_U3575) );
  MUX2_X1 U16514 ( .A(n15026), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14653), .Z(
        P1_U3574) );
  MUX2_X1 U16515 ( .A(n15221), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14653), .Z(
        P1_U3573) );
  MUX2_X1 U16516 ( .A(n15027), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14653), .Z(
        P1_U3572) );
  MUX2_X1 U16517 ( .A(n14648), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14653), .Z(
        P1_U3568) );
  MUX2_X1 U16518 ( .A(n14649), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14653), .Z(
        P1_U3566) );
  MUX2_X1 U16519 ( .A(n14650), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14653), .Z(
        P1_U3565) );
  MUX2_X1 U16520 ( .A(n14651), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14653), .Z(
        P1_U3564) );
  MUX2_X1 U16521 ( .A(n14652), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14653), .Z(
        P1_U3563) );
  MUX2_X1 U16522 ( .A(n11381), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14653), .Z(
        P1_U3562) );
  MUX2_X1 U16523 ( .A(n11380), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14653), .Z(
        P1_U3561) );
  MUX2_X1 U16524 ( .A(n11377), .B(P1_DATAO_REG_0__SCAN_IN), .S(n14653), .Z(
        P1_U3560) );
  NAND2_X1 U16525 ( .A1(n15193), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14669) );
  INV_X1 U16526 ( .A(n14669), .ZN(n14659) );
  MUX2_X1 U16527 ( .A(n14655), .B(P1_REG2_REG_1__SCAN_IN), .S(n14654), .Z(
        n14658) );
  INV_X1 U16528 ( .A(n14656), .ZN(n14657) );
  OAI211_X1 U16529 ( .C1(n14659), .C2(n14658), .A(n14785), .B(n14657), .ZN(
        n14667) );
  AOI22_X1 U16530 ( .A1(n15299), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14666) );
  NAND2_X1 U16531 ( .A1(n14783), .A2(n14660), .ZN(n14665) );
  OAI211_X1 U16532 ( .C1(n14663), .C2(n14662), .A(n15310), .B(n14661), .ZN(
        n14664) );
  NAND4_X1 U16533 ( .A1(n14667), .A2(n14666), .A3(n14665), .A4(n14664), .ZN(
        P1_U3244) );
  MUX2_X1 U16534 ( .A(n14669), .B(n14668), .S(n15291), .Z(n14672) );
  NOR2_X1 U16535 ( .A1(n15291), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14670) );
  OR2_X1 U16536 ( .A1(n14670), .A2(n14671), .ZN(n15289) );
  NAND2_X1 U16537 ( .A1(n15289), .A2(n15293), .ZN(n15296) );
  OAI211_X1 U16538 ( .C1(n14672), .C2(n14671), .A(P1_U4016), .B(n15296), .ZN(
        n14714) );
  OAI22_X1 U16539 ( .A1(n15319), .A2(n9098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9257), .ZN(n14673) );
  AOI21_X1 U16540 ( .B1(n14674), .B2(n14783), .A(n14673), .ZN(n14685) );
  MUX2_X1 U16541 ( .A(n14676), .B(P1_REG2_REG_2__SCAN_IN), .S(n14675), .Z(
        n14679) );
  INV_X1 U16542 ( .A(n14677), .ZN(n14678) );
  OAI211_X1 U16543 ( .C1(n14679), .C2(n14678), .A(n14785), .B(n14688), .ZN(
        n14684) );
  OAI211_X1 U16544 ( .C1(n14682), .C2(n14681), .A(n15310), .B(n14680), .ZN(
        n14683) );
  NAND4_X1 U16545 ( .A1(n14714), .A2(n14685), .A3(n14684), .A4(n14683), .ZN(
        P1_U3245) );
  INV_X1 U16546 ( .A(n14708), .ZN(n14690) );
  NAND3_X1 U16547 ( .A1(n14688), .A2(n14687), .A3(n14686), .ZN(n14689) );
  NAND3_X1 U16548 ( .A1(n14785), .A2(n14690), .A3(n14689), .ZN(n14698) );
  AOI22_X1 U16549 ( .A1(n15299), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(n6428), .ZN(n14697) );
  NAND2_X1 U16550 ( .A1(n14783), .A2(n14691), .ZN(n14696) );
  OAI211_X1 U16551 ( .C1(n14694), .C2(n14693), .A(n15310), .B(n14692), .ZN(
        n14695) );
  NAND4_X1 U16552 ( .A1(n14698), .A2(n14697), .A3(n14696), .A4(n14695), .ZN(
        P1_U3246) );
  NAND2_X1 U16553 ( .A1(n15299), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n14700) );
  NAND2_X1 U16554 ( .A1(n14700), .A2(n14699), .ZN(n14701) );
  AOI21_X1 U16555 ( .B1(n14702), .B2(n14783), .A(n14701), .ZN(n14713) );
  OAI211_X1 U16556 ( .C1(n14705), .C2(n14704), .A(n15310), .B(n14703), .ZN(
        n14712) );
  OR3_X1 U16557 ( .A1(n14708), .A2(n14707), .A3(n14706), .ZN(n14709) );
  NAND3_X1 U16558 ( .A1(n14785), .A2(n14710), .A3(n14709), .ZN(n14711) );
  NAND4_X1 U16559 ( .A1(n14714), .A2(n14713), .A3(n14712), .A4(n14711), .ZN(
        P1_U3247) );
  OR3_X1 U16560 ( .A1(n14717), .A2(n14716), .A3(n14715), .ZN(n14718) );
  NAND3_X1 U16561 ( .A1(n14719), .A2(n14785), .A3(n14718), .ZN(n14728) );
  NOR2_X1 U16562 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9311), .ZN(n14720) );
  AOI21_X1 U16563 ( .B1(n15299), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n14720), .ZN(
        n14727) );
  OAI211_X1 U16564 ( .C1(n14723), .C2(n14722), .A(n15310), .B(n14721), .ZN(
        n14726) );
  NAND2_X1 U16565 ( .A1(n14783), .A2(n14724), .ZN(n14725) );
  NAND4_X1 U16566 ( .A1(n14728), .A2(n14727), .A3(n14726), .A4(n14725), .ZN(
        P1_U3249) );
  OR3_X1 U16567 ( .A1(n14731), .A2(n14730), .A3(n14729), .ZN(n14732) );
  NAND3_X1 U16568 ( .A1(n14733), .A2(n14785), .A3(n14732), .ZN(n14743) );
  INV_X1 U16569 ( .A(n14734), .ZN(n14735) );
  AOI21_X1 U16570 ( .B1(n15299), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n14735), 
        .ZN(n14742) );
  OAI211_X1 U16571 ( .C1(n14738), .C2(n14737), .A(n14736), .B(n15310), .ZN(
        n14741) );
  NAND2_X1 U16572 ( .A1(n14783), .A2(n14739), .ZN(n14740) );
  NAND4_X1 U16573 ( .A1(n14743), .A2(n14742), .A3(n14741), .A4(n14740), .ZN(
        P1_U3253) );
  AOI22_X1 U16574 ( .A1(n14745), .A2(n14744), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n14749), .ZN(n14761) );
  XNOR2_X1 U16575 ( .A(n14762), .B(n14960), .ZN(n14760) );
  XNOR2_X1 U16576 ( .A(n14761), .B(n14760), .ZN(n14757) );
  INV_X1 U16577 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14747) );
  OAI21_X1 U16578 ( .B1(n15319), .B2(n14747), .A(n14746), .ZN(n14748) );
  AOI21_X1 U16579 ( .B1(n14765), .B2(n14783), .A(n14748), .ZN(n14756) );
  XNOR2_X1 U16580 ( .A(n14762), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14754) );
  NAND2_X1 U16581 ( .A1(n14749), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n14750) );
  INV_X1 U16582 ( .A(n14764), .ZN(n14752) );
  OAI211_X1 U16583 ( .C1(n14754), .C2(n14753), .A(n14752), .B(n15310), .ZN(
        n14755) );
  OAI211_X1 U16584 ( .C1(n14757), .C2(n15305), .A(n14756), .B(n14755), .ZN(
        P1_U3260) );
  OAI21_X1 U16585 ( .B1(n15319), .B2(n9185), .A(n14758), .ZN(n14759) );
  AOI21_X1 U16586 ( .B1(n14779), .B2(n14783), .A(n14759), .ZN(n14772) );
  OAI211_X1 U16587 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14763), .A(n14785), 
        .B(n14781), .ZN(n14771) );
  INV_X1 U16588 ( .A(n14766), .ZN(n14769) );
  INV_X1 U16589 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14767) );
  INV_X1 U16590 ( .A(n14776), .ZN(n14768) );
  OAI211_X1 U16591 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14769), .A(n15310), 
        .B(n14768), .ZN(n14770) );
  NAND3_X1 U16592 ( .A1(n14772), .A2(n14771), .A3(n14770), .ZN(P1_U3261) );
  NOR2_X1 U16593 ( .A1(n14774), .A2(n14773), .ZN(n14775) );
  NAND2_X1 U16594 ( .A1(n14779), .A2(n14778), .ZN(n14780) );
  NAND2_X1 U16595 ( .A1(n14781), .A2(n14780), .ZN(n14782) );
  AOI22_X1 U16596 ( .A1(n14786), .A2(n15310), .B1(n14785), .B2(n14784), .ZN(
        n14787) );
  NOR2_X1 U16597 ( .A1(n15049), .A2(n14791), .ZN(n14792) );
  NOR2_X1 U16598 ( .A1(n15340), .A2(n15064), .ZN(n14798) );
  AOI211_X1 U16599 ( .C1(n14534), .C2(n15329), .A(n14792), .B(n14798), .ZN(
        n14793) );
  OAI21_X1 U16600 ( .B1(n14794), .B2(n14860), .A(n14793), .ZN(P1_U3263) );
  OAI211_X1 U16601 ( .C1(n14796), .C2(n15066), .A(n15333), .B(n14795), .ZN(
        n15065) );
  NOR2_X1 U16602 ( .A1(n15049), .A2(n14797), .ZN(n14799) );
  AOI211_X1 U16603 ( .C1(n14800), .C2(n15329), .A(n14799), .B(n14798), .ZN(
        n14801) );
  OAI21_X1 U16604 ( .B1(n15065), .B2(n14860), .A(n14801), .ZN(P1_U3264) );
  AOI21_X1 U16605 ( .B1(n14802), .B2(n14829), .A(n14819), .ZN(n14803) );
  XNOR2_X1 U16606 ( .A(n14803), .B(n14814), .ZN(n14805) );
  AOI21_X2 U16607 ( .B1(n14805), .B2(n15024), .A(n14804), .ZN(n15089) );
  INV_X1 U16608 ( .A(n14825), .ZN(n14807) );
  INV_X1 U16609 ( .A(n12435), .ZN(n14806) );
  INV_X1 U16610 ( .A(n14808), .ZN(n14809) );
  AOI22_X1 U16611 ( .A1(n14809), .A2(n15331), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15340), .ZN(n14810) );
  OAI21_X1 U16612 ( .B1(n14811), .B2(n15057), .A(n14810), .ZN(n14816) );
  INV_X1 U16613 ( .A(n14832), .ZN(n14812) );
  NAND2_X1 U16614 ( .A1(n15092), .A2(n14813), .ZN(n14815) );
  AND2_X1 U16615 ( .A1(n14817), .A2(n14830), .ZN(n14818) );
  OAI21_X1 U16616 ( .B1(n14819), .B2(n14818), .A(n15024), .ZN(n14821) );
  NAND2_X1 U16617 ( .A1(n14821), .A2(n14820), .ZN(n15097) );
  INV_X1 U16618 ( .A(n15097), .ZN(n14835) );
  OAI22_X1 U16619 ( .A1(n14823), .A2(n15055), .B1(n14822), .B2(n15049), .ZN(
        n14828) );
  NAND2_X1 U16620 ( .A1(n14839), .A2(n14829), .ZN(n14824) );
  NAND2_X1 U16621 ( .A1(n14824), .A2(n15333), .ZN(n14826) );
  NOR2_X1 U16622 ( .A1(n15094), .A2(n14860), .ZN(n14827) );
  AOI211_X1 U16623 ( .C1(n15329), .C2(n14829), .A(n14828), .B(n14827), .ZN(
        n14834) );
  INV_X1 U16624 ( .A(n14830), .ZN(n14831) );
  NAND2_X1 U16625 ( .A1(n14832), .A2(n14831), .ZN(n15091) );
  NAND3_X1 U16626 ( .A1(n15092), .A2(n14865), .A3(n15091), .ZN(n14833) );
  OAI211_X1 U16627 ( .C1(n14835), .C2(n15340), .A(n14834), .B(n14833), .ZN(
        P1_U3268) );
  XNOR2_X1 U16628 ( .A(n14836), .B(n7632), .ZN(n15103) );
  AOI21_X1 U16629 ( .B1(n7814), .B2(n14838), .A(n15365), .ZN(n14840) );
  NAND2_X1 U16630 ( .A1(n14840), .A2(n14839), .ZN(n15099) );
  INV_X1 U16631 ( .A(n15099), .ZN(n14850) );
  INV_X1 U16632 ( .A(n14841), .ZN(n14842) );
  AOI22_X1 U16633 ( .A1(n14842), .A2(n15331), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15340), .ZN(n14843) );
  OAI21_X1 U16634 ( .B1(n14844), .B2(n15057), .A(n14843), .ZN(n14849) );
  OAI211_X1 U16635 ( .C1(n14847), .C2(n14846), .A(n15024), .B(n14845), .ZN(
        n15101) );
  AOI21_X1 U16636 ( .B1(n15101), .B2(n15100), .A(n15340), .ZN(n14848) );
  AOI211_X1 U16637 ( .C1(n14850), .C2(n15235), .A(n14849), .B(n14848), .ZN(
        n14851) );
  OAI21_X1 U16638 ( .B1(n15103), .B2(n14952), .A(n14851), .ZN(P1_U3269) );
  XNOR2_X1 U16639 ( .A(n14852), .B(n14863), .ZN(n14854) );
  AOI21_X1 U16640 ( .B1(n14854), .B2(n15024), .A(n14853), .ZN(n15109) );
  AOI21_X1 U16641 ( .B1(n14855), .B2(n15104), .A(n15365), .ZN(n14856) );
  NAND2_X1 U16642 ( .A1(n14856), .A2(n7814), .ZN(n15106) );
  AOI22_X1 U16643 ( .A1(n14857), .A2(n15331), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15340), .ZN(n14859) );
  NAND2_X1 U16644 ( .A1(n15104), .A2(n15329), .ZN(n14858) );
  OAI211_X1 U16645 ( .C1(n15106), .C2(n14860), .A(n14859), .B(n14858), .ZN(
        n14861) );
  INV_X1 U16646 ( .A(n14861), .ZN(n14867) );
  NAND2_X1 U16647 ( .A1(n14864), .A2(n14863), .ZN(n15105) );
  NAND3_X1 U16648 ( .A1(n14862), .A2(n15105), .A3(n14865), .ZN(n14866) );
  OAI211_X1 U16649 ( .C1(n15109), .C2(n15340), .A(n14867), .B(n14866), .ZN(
        P1_U3270) );
  OAI21_X1 U16650 ( .B1(n14880), .B2(n14869), .A(n14868), .ZN(n14872) );
  AOI222_X1 U16651 ( .A1(n14872), .A2(n15024), .B1(n14871), .B2(n15222), .C1(
        n14870), .C2(n15223), .ZN(n15113) );
  INV_X1 U16652 ( .A(n14892), .ZN(n14874) );
  INV_X1 U16653 ( .A(n14855), .ZN(n14873) );
  AOI211_X1 U16654 ( .C1(n15111), .C2(n14874), .A(n15365), .B(n14873), .ZN(
        n15110) );
  INV_X1 U16655 ( .A(n14875), .ZN(n14876) );
  AOI22_X1 U16656 ( .A1(n14876), .A2(n15331), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15340), .ZN(n14877) );
  OAI21_X1 U16657 ( .B1(n14878), .B2(n15057), .A(n14877), .ZN(n14882) );
  XNOR2_X1 U16658 ( .A(n14879), .B(n14880), .ZN(n15114) );
  NOR2_X1 U16659 ( .A1(n15114), .A2(n15062), .ZN(n14881) );
  AOI211_X1 U16660 ( .C1(n15110), .C2(n15235), .A(n14882), .B(n14881), .ZN(
        n14883) );
  OAI21_X1 U16661 ( .B1(n15113), .B2(n15340), .A(n14883), .ZN(P1_U3271) );
  XOR2_X1 U16662 ( .A(n14884), .B(n14886), .Z(n15120) );
  OAI211_X1 U16663 ( .C1(n14887), .C2(n14886), .A(n15024), .B(n14885), .ZN(
        n14888) );
  INV_X1 U16664 ( .A(n14888), .ZN(n15118) );
  OAI21_X1 U16665 ( .B1(n15118), .B2(n15115), .A(n15049), .ZN(n14898) );
  NAND2_X1 U16666 ( .A1(n14906), .A2(n14889), .ZN(n14890) );
  NAND2_X1 U16667 ( .A1(n14890), .A2(n15333), .ZN(n14891) );
  NOR2_X1 U16668 ( .A1(n14892), .A2(n14891), .ZN(n15117) );
  AOI22_X1 U16669 ( .A1(n14893), .A2(n15331), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15340), .ZN(n14894) );
  OAI21_X1 U16670 ( .B1(n14895), .B2(n15057), .A(n14894), .ZN(n14896) );
  AOI21_X1 U16671 ( .B1(n15117), .B2(n15235), .A(n14896), .ZN(n14897) );
  OAI211_X1 U16672 ( .C1(n15120), .C2(n15062), .A(n14898), .B(n14897), .ZN(
        P1_U3272) );
  AOI21_X1 U16673 ( .B1(n14900), .B2(n14899), .A(n15325), .ZN(n14903) );
  OAI22_X1 U16674 ( .A1(n14901), .A2(n15052), .B1(n14944), .B2(n14976), .ZN(
        n14902) );
  AOI21_X1 U16675 ( .B1(n14904), .B2(n14903), .A(n14902), .ZN(n15124) );
  AOI211_X1 U16676 ( .C1(n15122), .C2(n14926), .A(n15365), .B(n7030), .ZN(
        n15121) );
  NAND2_X1 U16677 ( .A1(n15121), .A2(n14958), .ZN(n14907) );
  AOI21_X1 U16678 ( .B1(n15124), .B2(n14907), .A(n15340), .ZN(n14916) );
  NAND2_X1 U16679 ( .A1(n14908), .A2(n14909), .ZN(n14910) );
  NAND2_X1 U16680 ( .A1(n14911), .A2(n14910), .ZN(n15125) );
  AOI22_X1 U16681 ( .A1(n14912), .A2(n15331), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n15340), .ZN(n14914) );
  NAND2_X1 U16682 ( .A1(n15122), .A2(n15329), .ZN(n14913) );
  OAI211_X1 U16683 ( .C1(n15125), .C2(n15062), .A(n14914), .B(n14913), .ZN(
        n14915) );
  OR2_X1 U16684 ( .A1(n14916), .A2(n14915), .ZN(P1_U3273) );
  XOR2_X1 U16685 ( .A(n14917), .B(n14921), .Z(n15130) );
  INV_X1 U16686 ( .A(n14918), .ZN(n14919) );
  AOI21_X1 U16687 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(n14922) );
  OAI222_X1 U16688 ( .A1(n15052), .A2(n14923), .B1(n14976), .B2(n14957), .C1(
        n14922), .C2(n15325), .ZN(n15126) );
  OR2_X1 U16689 ( .A1(n14937), .A2(n14931), .ZN(n14925) );
  AND3_X1 U16690 ( .A1(n14926), .A2(n14925), .A3(n15333), .ZN(n15127) );
  NAND2_X1 U16691 ( .A1(n15127), .A2(n15235), .ZN(n14930) );
  INV_X1 U16692 ( .A(n14927), .ZN(n14928) );
  AOI22_X1 U16693 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(n15340), .B1(n14928), 
        .B2(n15331), .ZN(n14929) );
  OAI211_X1 U16694 ( .C1(n14931), .C2(n15057), .A(n14930), .B(n14929), .ZN(
        n14932) );
  AOI21_X1 U16695 ( .B1(n15126), .B2(n15049), .A(n14932), .ZN(n14933) );
  OAI21_X1 U16696 ( .B1(n15130), .B2(n15062), .A(n14933), .ZN(P1_U3274) );
  XNOR2_X1 U16697 ( .A(n14934), .B(n14942), .ZN(n15134) );
  NOR2_X1 U16698 ( .A1(n14935), .A2(n14941), .ZN(n14936) );
  INV_X1 U16699 ( .A(n14938), .ZN(n14939) );
  AOI22_X1 U16700 ( .A1(n15340), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14939), 
        .B2(n15331), .ZN(n14940) );
  OAI21_X1 U16701 ( .B1(n14941), .B2(n15057), .A(n14940), .ZN(n14949) );
  AOI21_X1 U16702 ( .B1(n14943), .B2(n14942), .A(n15325), .ZN(n14947) );
  OAI22_X1 U16703 ( .A1(n14944), .A2(n15052), .B1(n14974), .B2(n14976), .ZN(
        n14945) );
  AOI21_X1 U16704 ( .B1(n14947), .B2(n14946), .A(n14945), .ZN(n15133) );
  NOR2_X1 U16705 ( .A1(n15133), .A2(n15340), .ZN(n14948) );
  AOI211_X1 U16706 ( .C1(n7815), .C2(n14950), .A(n14949), .B(n14948), .ZN(
        n14951) );
  OAI21_X1 U16707 ( .B1(n14952), .B2(n15134), .A(n14951), .ZN(P1_U3275) );
  XNOR2_X1 U16708 ( .A(n7811), .B(n15137), .ZN(n14953) );
  NOR2_X1 U16709 ( .A1(n14953), .A2(n15365), .ZN(n15136) );
  XOR2_X1 U16710 ( .A(n14954), .B(n14962), .Z(n14955) );
  OAI222_X1 U16711 ( .A1(n15052), .A2(n14957), .B1(n14976), .B2(n14956), .C1(
        n14955), .C2(n15325), .ZN(n15135) );
  AOI21_X1 U16712 ( .B1(n15136), .B2(n14958), .A(n15135), .ZN(n14967) );
  OAI22_X1 U16713 ( .A1(n15049), .A2(n14960), .B1(n14959), .B2(n15055), .ZN(
        n14965) );
  XNOR2_X1 U16714 ( .A(n14963), .B(n14962), .ZN(n15139) );
  NOR2_X1 U16715 ( .A1(n15139), .A2(n15062), .ZN(n14964) );
  AOI211_X1 U16716 ( .C1(n15329), .C2(n15137), .A(n14965), .B(n14964), .ZN(
        n14966) );
  OAI21_X1 U16717 ( .B1(n14967), .B2(n15340), .A(n14966), .ZN(P1_U3276) );
  XNOR2_X1 U16718 ( .A(n14968), .B(n7743), .ZN(n15144) );
  INV_X1 U16719 ( .A(n14969), .ZN(n14970) );
  AOI21_X1 U16720 ( .B1(n14972), .B2(n14971), .A(n14970), .ZN(n14973) );
  OAI222_X1 U16721 ( .A1(n14976), .A2(n14975), .B1(n15052), .B2(n14974), .C1(
        n14973), .C2(n15325), .ZN(n15140) );
  AOI21_X1 U16722 ( .B1(n14989), .B2(n15142), .A(n15365), .ZN(n14977) );
  AND2_X1 U16723 ( .A1(n14977), .A2(n7811), .ZN(n15141) );
  NAND2_X1 U16724 ( .A1(n15141), .A2(n15235), .ZN(n14982) );
  NAND2_X1 U16725 ( .A1(n15340), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14978) );
  OAI21_X1 U16726 ( .B1(n15055), .B2(n14979), .A(n14978), .ZN(n14980) );
  AOI21_X1 U16727 ( .B1(n15142), .B2(n15329), .A(n14980), .ZN(n14981) );
  NAND2_X1 U16728 ( .A1(n14982), .A2(n14981), .ZN(n14983) );
  AOI21_X1 U16729 ( .B1(n15140), .B2(n15049), .A(n14983), .ZN(n14984) );
  OAI21_X1 U16730 ( .B1(n15062), .B2(n15144), .A(n14984), .ZN(P1_U3277) );
  XNOR2_X1 U16731 ( .A(n14985), .B(n14986), .ZN(n14988) );
  AOI222_X1 U16732 ( .A1(n14988), .A2(n15024), .B1(n14987), .B2(n15222), .C1(
        n15026), .C2(n15223), .ZN(n15148) );
  INV_X1 U16733 ( .A(n15006), .ZN(n14991) );
  INV_X1 U16734 ( .A(n14989), .ZN(n14990) );
  AOI211_X1 U16735 ( .C1(n15146), .C2(n14991), .A(n15365), .B(n14990), .ZN(
        n15145) );
  INV_X1 U16736 ( .A(n14992), .ZN(n14993) );
  AOI22_X1 U16737 ( .A1(n15340), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14993), 
        .B2(n15331), .ZN(n14994) );
  OAI21_X1 U16738 ( .B1(n14995), .B2(n15057), .A(n14994), .ZN(n15001) );
  INV_X1 U16739 ( .A(n14997), .ZN(n14998) );
  AOI21_X1 U16740 ( .B1(n14999), .B2(n14996), .A(n14998), .ZN(n15149) );
  NOR2_X1 U16741 ( .A1(n15149), .A2(n15062), .ZN(n15000) );
  AOI211_X1 U16742 ( .C1(n15145), .C2(n15235), .A(n15001), .B(n15000), .ZN(
        n15002) );
  OAI21_X1 U16743 ( .B1(n15340), .B2(n15148), .A(n15002), .ZN(P1_U3278) );
  XOR2_X1 U16744 ( .A(n15003), .B(n15011), .Z(n15005) );
  AOI21_X1 U16745 ( .B1(n15005), .B2(n15024), .A(n15004), .ZN(n15153) );
  AOI211_X1 U16746 ( .C1(n15151), .C2(n15030), .A(n15365), .B(n15006), .ZN(
        n15150) );
  INV_X1 U16747 ( .A(n15007), .ZN(n15008) );
  AOI22_X1 U16748 ( .A1(n15340), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n15008), 
        .B2(n15331), .ZN(n15009) );
  OAI21_X1 U16749 ( .B1(n15010), .B2(n15057), .A(n15009), .ZN(n15016) );
  NAND2_X1 U16750 ( .A1(n15012), .A2(n15011), .ZN(n15013) );
  NAND2_X1 U16751 ( .A1(n15014), .A2(n15013), .ZN(n15154) );
  NOR2_X1 U16752 ( .A1(n15154), .A2(n15062), .ZN(n15015) );
  AOI211_X1 U16753 ( .C1(n15150), .C2(n15235), .A(n15016), .B(n15015), .ZN(
        n15017) );
  OAI21_X1 U16754 ( .B1(n15340), .B2(n15153), .A(n15017), .ZN(P1_U3279) );
  XNOR2_X1 U16755 ( .A(n15018), .B(n15019), .ZN(n15250) );
  NAND2_X1 U16756 ( .A1(n15021), .A2(n15020), .ZN(n15023) );
  XNOR2_X1 U16757 ( .A(n15023), .B(n15022), .ZN(n15025) );
  NAND2_X1 U16758 ( .A1(n15025), .A2(n15024), .ZN(n15029) );
  AOI22_X1 U16759 ( .A1(n15223), .A2(n15027), .B1(n15026), .B2(n15222), .ZN(
        n15028) );
  NAND2_X1 U16760 ( .A1(n15029), .A2(n15028), .ZN(n15255) );
  AOI21_X1 U16761 ( .B1(n15232), .B2(n15036), .A(n15365), .ZN(n15031) );
  NAND2_X1 U16762 ( .A1(n15031), .A2(n15030), .ZN(n15251) );
  NOR2_X1 U16763 ( .A1(n15251), .A2(n14381), .ZN(n15032) );
  OAI21_X1 U16764 ( .B1(n15255), .B2(n15032), .A(n15049), .ZN(n15038) );
  OAI22_X1 U16765 ( .A1(n15049), .A2(n15034), .B1(n15033), .B2(n15055), .ZN(
        n15035) );
  AOI21_X1 U16766 ( .B1(n15036), .B2(n15329), .A(n15035), .ZN(n15037) );
  OAI211_X1 U16767 ( .C1(n15250), .C2(n15062), .A(n15038), .B(n15037), .ZN(
        P1_U3280) );
  XOR2_X1 U16768 ( .A(n15039), .B(n15046), .Z(n15403) );
  INV_X1 U16769 ( .A(n15043), .ZN(n15040) );
  NAND2_X1 U16770 ( .A1(n15040), .A2(n15041), .ZN(n15045) );
  INV_X1 U16771 ( .A(n15041), .ZN(n15042) );
  NOR3_X1 U16772 ( .A1(n15043), .A2(n15042), .A3(n15046), .ZN(n15044) );
  AOI211_X1 U16773 ( .C1(n15046), .C2(n15045), .A(n15325), .B(n15044), .ZN(
        n15047) );
  AOI21_X1 U16774 ( .B1(n15223), .B2(n15048), .A(n15047), .ZN(n15402) );
  MUX2_X1 U16775 ( .A(n15050), .B(n15402), .S(n15049), .Z(n15061) );
  OAI21_X1 U16776 ( .B1(n15051), .B2(n15058), .A(n15333), .ZN(n15054) );
  OAI22_X1 U16777 ( .A1(n15054), .A2(n11937), .B1(n15053), .B2(n15052), .ZN(
        n15398) );
  OAI22_X1 U16778 ( .A1(n15058), .A2(n15057), .B1(n15056), .B2(n15055), .ZN(
        n15059) );
  AOI21_X1 U16779 ( .B1(n15398), .B2(n15235), .A(n15059), .ZN(n15060) );
  OAI211_X1 U16780 ( .C1(n15403), .C2(n15062), .A(n15061), .B(n15060), .ZN(
        P1_U3283) );
  MUX2_X1 U16781 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15063), .S(n15420), .Z(
        P1_U3559) );
  OAI211_X1 U16782 ( .C1(n15066), .C2(n15363), .A(n15065), .B(n15064), .ZN(
        n15155) );
  MUX2_X1 U16783 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15155), .S(n15420), .Z(
        P1_U3558) );
  OAI211_X1 U16784 ( .C1(n15070), .C2(n15363), .A(n15069), .B(n15068), .ZN(
        n15071) );
  NAND3_X1 U16785 ( .A1(n15075), .A2(n15074), .A3(n15395), .ZN(n15080) );
  AOI21_X1 U16786 ( .B1(n15400), .B2(n15077), .A(n15076), .ZN(n15078) );
  NAND3_X1 U16787 ( .A1(n15080), .A2(n15079), .A3(n15078), .ZN(n15157) );
  MUX2_X1 U16788 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15157), .S(n15420), .Z(
        P1_U3556) );
  AOI21_X1 U16789 ( .B1(n15400), .B2(n15082), .A(n15081), .ZN(n15083) );
  OAI211_X1 U16790 ( .C1(n15404), .C2(n15085), .A(n15084), .B(n15083), .ZN(
        n15158) );
  MUX2_X1 U16791 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15158), .S(n15420), .Z(
        P1_U3555) );
  AOI21_X1 U16792 ( .B1(n15400), .B2(n15087), .A(n15086), .ZN(n15088) );
  OAI211_X1 U16793 ( .C1(n15404), .C2(n15090), .A(n15089), .B(n15088), .ZN(
        n15159) );
  MUX2_X1 U16794 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15159), .S(n15420), .Z(
        P1_U3554) );
  NAND2_X1 U16795 ( .A1(n15094), .A2(n15093), .ZN(n15095) );
  OR3_X2 U16796 ( .A1(n15097), .A2(n15096), .A3(n15095), .ZN(n15160) );
  MUX2_X1 U16797 ( .A(n15160), .B(P1_REG1_REG_25__SCAN_IN), .S(n15418), .Z(
        P1_U3553) );
  OAI21_X1 U16798 ( .B1(n15404), .B2(n15103), .A(n15102), .ZN(n15161) );
  MUX2_X1 U16799 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15161), .S(n15420), .Z(
        P1_U3552) );
  NAND2_X1 U16800 ( .A1(n15104), .A2(n15400), .ZN(n15108) );
  NAND3_X1 U16801 ( .A1(n14862), .A2(n15395), .A3(n15105), .ZN(n15107) );
  NAND4_X1 U16802 ( .A1(n15109), .A2(n15108), .A3(n15107), .A4(n15106), .ZN(
        n15162) );
  MUX2_X1 U16803 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15162), .S(n15420), .Z(
        P1_U3551) );
  AOI21_X1 U16804 ( .B1(n15400), .B2(n15111), .A(n15110), .ZN(n15112) );
  OAI211_X1 U16805 ( .C1(n15404), .C2(n15114), .A(n15113), .B(n15112), .ZN(
        n15163) );
  MUX2_X1 U16806 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15163), .S(n15420), .Z(
        P1_U3550) );
  NOR4_X1 U16807 ( .A1(n15118), .A2(n15117), .A3(n15116), .A4(n15115), .ZN(
        n15119) );
  OAI21_X1 U16808 ( .B1(n15404), .B2(n15120), .A(n15119), .ZN(n15164) );
  MUX2_X1 U16809 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15164), .S(n15420), .Z(
        P1_U3549) );
  AOI21_X1 U16810 ( .B1(n15400), .B2(n15122), .A(n15121), .ZN(n15123) );
  OAI211_X1 U16811 ( .C1(n15404), .C2(n15125), .A(n15124), .B(n15123), .ZN(
        n15165) );
  MUX2_X1 U16812 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15165), .S(n15420), .Z(
        P1_U3548) );
  AOI211_X1 U16813 ( .C1(n15400), .C2(n15128), .A(n15127), .B(n15126), .ZN(
        n15129) );
  OAI21_X1 U16814 ( .B1(n15404), .B2(n15130), .A(n15129), .ZN(n15166) );
  MUX2_X1 U16815 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15166), .S(n15420), .Z(
        P1_U3547) );
  AOI22_X1 U16816 ( .A1(n7815), .A2(n15333), .B1(n15400), .B2(n15131), .ZN(
        n15132) );
  OAI211_X1 U16817 ( .C1(n15404), .C2(n15134), .A(n15133), .B(n15132), .ZN(
        n15167) );
  MUX2_X1 U16818 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15167), .S(n15420), .Z(
        P1_U3546) );
  AOI211_X1 U16819 ( .C1(n15400), .C2(n15137), .A(n15136), .B(n15135), .ZN(
        n15138) );
  OAI21_X1 U16820 ( .B1(n15404), .B2(n15139), .A(n15138), .ZN(n15168) );
  MUX2_X1 U16821 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15168), .S(n15420), .Z(
        P1_U3545) );
  AOI211_X1 U16822 ( .C1(n15400), .C2(n15142), .A(n15141), .B(n15140), .ZN(
        n15143) );
  OAI21_X1 U16823 ( .B1(n15404), .B2(n15144), .A(n15143), .ZN(n15169) );
  MUX2_X1 U16824 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15169), .S(n15420), .Z(
        P1_U3544) );
  AOI21_X1 U16825 ( .B1(n15400), .B2(n15146), .A(n15145), .ZN(n15147) );
  OAI211_X1 U16826 ( .C1(n15404), .C2(n15149), .A(n15148), .B(n15147), .ZN(
        n15170) );
  MUX2_X1 U16827 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15170), .S(n15420), .Z(
        P1_U3543) );
  AOI21_X1 U16828 ( .B1(n15400), .B2(n15151), .A(n15150), .ZN(n15152) );
  OAI211_X1 U16829 ( .C1(n15404), .C2(n15154), .A(n15153), .B(n15152), .ZN(
        n15171) );
  MUX2_X1 U16830 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15171), .S(n15420), .Z(
        P1_U3542) );
  MUX2_X1 U16831 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15155), .S(n15408), .Z(
        P1_U3526) );
  MUX2_X1 U16832 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15157), .S(n15408), .Z(
        P1_U3524) );
  MUX2_X1 U16833 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15158), .S(n15408), .Z(
        P1_U3523) );
  MUX2_X1 U16834 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15159), .S(n15408), .Z(
        P1_U3522) );
  MUX2_X1 U16835 ( .A(n15160), .B(P1_REG0_REG_25__SCAN_IN), .S(n15406), .Z(
        P1_U3521) );
  MUX2_X1 U16836 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15161), .S(n15408), .Z(
        P1_U3520) );
  MUX2_X1 U16837 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15162), .S(n15408), .Z(
        P1_U3519) );
  MUX2_X1 U16838 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15163), .S(n15408), .Z(
        P1_U3518) );
  MUX2_X1 U16839 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15164), .S(n15408), .Z(
        P1_U3517) );
  MUX2_X1 U16840 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15165), .S(n15408), .Z(
        P1_U3516) );
  MUX2_X1 U16841 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15166), .S(n15408), .Z(
        P1_U3515) );
  MUX2_X1 U16842 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15167), .S(n15408), .Z(
        P1_U3513) );
  MUX2_X1 U16843 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15168), .S(n15408), .Z(
        P1_U3510) );
  MUX2_X1 U16844 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15169), .S(n15408), .Z(
        P1_U3507) );
  MUX2_X1 U16845 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15170), .S(n15408), .Z(
        P1_U3504) );
  MUX2_X1 U16846 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15171), .S(n15408), .Z(
        P1_U3501) );
  NAND3_X1 U16847 ( .A1(n15173), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n15176) );
  OAI22_X1 U16848 ( .A1(n15172), .A2(n15176), .B1(n15175), .B2(n15174), .ZN(
        n15177) );
  AOI21_X1 U16849 ( .B1(n14164), .B2(n15178), .A(n15177), .ZN(n15179) );
  INV_X1 U16850 ( .A(n15179), .ZN(P1_U3324) );
  OAI222_X1 U16851 ( .A1(n15185), .A2(n15182), .B1(n6428), .B2(n15181), .C1(
        n15188), .C2(n15180), .ZN(P1_U3326) );
  OAI222_X1 U16852 ( .A1(n15185), .A2(n15184), .B1(P1_U3086), .B2(n15291), 
        .C1(n15188), .C2(n15183), .ZN(P1_U3328) );
  OAI222_X1 U16853 ( .A1(n6428), .A2(n15189), .B1(n15188), .B2(n15187), .C1(
        n15186), .C2(n15185), .ZN(P1_U3329) );
  MUX2_X1 U16854 ( .A(n15191), .B(n15190), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16855 ( .A(n15192), .ZN(n15194) );
  MUX2_X1 U16856 ( .A(n15194), .B(n15193), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  XNOR2_X1 U16857 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n15195), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16858 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15196) );
  OAI21_X1 U16859 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n15196), 
        .ZN(U28) );
  AOI21_X1 U16860 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15197) );
  OAI21_X1 U16861 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15197), 
        .ZN(U29) );
  INV_X1 U16862 ( .A(n15198), .ZN(n15200) );
  AOI222_X1 U16863 ( .A1(n15201), .A2(n15200), .B1(n15201), .B2(n15199), .C1(
        n15661), .C2(n15198), .ZN(SUB_1596_U61) );
  XOR2_X1 U16864 ( .A(n15202), .B(n15203), .Z(SUB_1596_U57) );
  OAI21_X1 U16865 ( .B1(n15206), .B2(n15205), .A(n15204), .ZN(n15207) );
  XNOR2_X1 U16866 ( .A(n15207), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  OAI21_X1 U16867 ( .B1(n15210), .B2(n15209), .A(n15208), .ZN(n15211) );
  XNOR2_X1 U16868 ( .A(n15211), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  AOI21_X1 U16869 ( .B1(n15214), .B2(n15213), .A(n15212), .ZN(n15216) );
  XNOR2_X1 U16870 ( .A(n15216), .B(n15215), .ZN(SUB_1596_U70) );
  XNOR2_X1 U16871 ( .A(n15217), .B(n15218), .ZN(n15243) );
  XNOR2_X1 U16872 ( .A(n15220), .B(n15219), .ZN(n15226) );
  AOI22_X1 U16873 ( .A1(n15224), .A2(n15223), .B1(n15222), .B2(n15221), .ZN(
        n15225) );
  OAI21_X1 U16874 ( .B1(n15226), .B2(n15325), .A(n15225), .ZN(n15227) );
  AOI21_X1 U16875 ( .B1(n15361), .B2(n15243), .A(n15227), .ZN(n15240) );
  INV_X1 U16876 ( .A(n15228), .ZN(n15229) );
  AOI222_X1 U16877 ( .A1(n15230), .A2(n15329), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n15340), .C1(n15229), .C2(n15331), .ZN(n15237) );
  INV_X1 U16878 ( .A(n15231), .ZN(n15337) );
  INV_X1 U16879 ( .A(n11938), .ZN(n15233) );
  OAI211_X1 U16880 ( .C1(n15233), .C2(n15239), .A(n15333), .B(n15232), .ZN(
        n15238) );
  INV_X1 U16881 ( .A(n15238), .ZN(n15234) );
  AOI22_X1 U16882 ( .A1(n15243), .A2(n15337), .B1(n15235), .B2(n15234), .ZN(
        n15236) );
  OAI211_X1 U16883 ( .C1(n15340), .C2(n15240), .A(n15237), .B(n15236), .ZN(
        P1_U3281) );
  INV_X1 U16884 ( .A(n15374), .ZN(n15353) );
  OAI21_X1 U16885 ( .B1(n15239), .B2(n15363), .A(n15238), .ZN(n15242) );
  INV_X1 U16886 ( .A(n15240), .ZN(n15241) );
  AOI211_X1 U16887 ( .C1(n15353), .C2(n15243), .A(n15242), .B(n15241), .ZN(
        n15245) );
  INV_X1 U16888 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n15244) );
  AOI22_X1 U16889 ( .A1(n15408), .A2(n15245), .B1(n15244), .B2(n15406), .ZN(
        P1_U3495) );
  AOI22_X1 U16890 ( .A1(n15420), .A2(n15245), .B1(n11288), .B2(n15418), .ZN(
        P1_U3540) );
  AOI21_X1 U16891 ( .B1(n15248), .B2(n15247), .A(n15246), .ZN(n15249) );
  XNOR2_X1 U16892 ( .A(n15249), .B(n15523), .ZN(SUB_1596_U63) );
  NOR2_X1 U16893 ( .A1(n15250), .A2(n15404), .ZN(n15254) );
  OAI21_X1 U16894 ( .B1(n15252), .B2(n15363), .A(n15251), .ZN(n15253) );
  NOR3_X1 U16895 ( .A1(n15255), .A2(n15254), .A3(n15253), .ZN(n15263) );
  AOI22_X1 U16896 ( .A1(n15420), .A2(n15263), .B1(n15256), .B2(n15418), .ZN(
        P1_U3541) );
  AND2_X1 U16897 ( .A1(n15257), .A2(n15395), .ZN(n15261) );
  OAI21_X1 U16898 ( .B1(n15259), .B2(n15363), .A(n15258), .ZN(n15260) );
  NOR3_X1 U16899 ( .A1(n15262), .A2(n15261), .A3(n15260), .ZN(n15265) );
  AOI22_X1 U16900 ( .A1(n15420), .A2(n15265), .B1(n9357), .B2(n15418), .ZN(
        P1_U3539) );
  AOI22_X1 U16901 ( .A1(n15408), .A2(n15263), .B1(n9384), .B2(n15406), .ZN(
        P1_U3498) );
  INV_X1 U16902 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15264) );
  AOI22_X1 U16903 ( .A1(n15408), .A2(n15265), .B1(n15264), .B2(n15406), .ZN(
        P1_U3492) );
  AOI21_X1 U16904 ( .B1(n15268), .B2(n15267), .A(n15266), .ZN(n15270) );
  XNOR2_X1 U16905 ( .A(n15270), .B(n15269), .ZN(SUB_1596_U69) );
  XNOR2_X1 U16906 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n15271), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16907 ( .B1(n15274), .B2(n15273), .A(n15272), .ZN(n15276) );
  XNOR2_X1 U16908 ( .A(n15276), .B(n15275), .ZN(SUB_1596_U67) );
  AOI21_X1 U16909 ( .B1(n15279), .B2(n15278), .A(n15277), .ZN(n15281) );
  XNOR2_X1 U16910 ( .A(n15281), .B(n15280), .ZN(SUB_1596_U66) );
  NOR2_X1 U16911 ( .A1(n15283), .A2(n15282), .ZN(n15284) );
  XOR2_X1 U16912 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15284), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16913 ( .B1(n15287), .B2(n15286), .A(n15285), .ZN(n15288) );
  XNOR2_X1 U16914 ( .A(n15288), .B(n15507), .ZN(SUB_1596_U64) );
  INV_X1 U16915 ( .A(n15289), .ZN(n15292) );
  NAND2_X1 U16916 ( .A1(n15291), .A2(n15290), .ZN(n15294) );
  NAND2_X1 U16917 ( .A1(n15292), .A2(n15294), .ZN(n15295) );
  MUX2_X1 U16918 ( .A(n15295), .B(n15294), .S(n15293), .Z(n15297) );
  NAND2_X1 U16919 ( .A1(n15297), .A2(n15296), .ZN(n15301) );
  AOI22_X1 U16920 ( .A1(n15299), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n6428), .ZN(n15300) );
  OAI21_X1 U16921 ( .B1(n15302), .B2(n15301), .A(n15300), .ZN(P1_U3243) );
  AOI21_X1 U16922 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n15304), .A(n15303), 
        .ZN(n15306) );
  OR2_X1 U16923 ( .A1(n15306), .A2(n15305), .ZN(n15313) );
  OAI21_X1 U16924 ( .B1(n15309), .B2(n15308), .A(n15307), .ZN(n15311) );
  NAND2_X1 U16925 ( .A1(n15311), .A2(n15310), .ZN(n15312) );
  OAI211_X1 U16926 ( .C1(n15315), .C2(n15314), .A(n15313), .B(n15312), .ZN(
        n15316) );
  INV_X1 U16927 ( .A(n15316), .ZN(n15318) );
  OAI211_X1 U16928 ( .C1(n15320), .C2(n15319), .A(n15318), .B(n15317), .ZN(
        P1_U3258) );
  OAI21_X1 U16929 ( .B1(n15322), .B2(n15323), .A(n15321), .ZN(n15352) );
  XNOR2_X1 U16930 ( .A(n15324), .B(n15323), .ZN(n15326) );
  NOR2_X1 U16931 ( .A1(n15326), .A2(n15325), .ZN(n15327) );
  AOI211_X1 U16932 ( .C1(n15361), .C2(n15352), .A(n15328), .B(n15327), .ZN(
        n15349) );
  AOI222_X1 U16933 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n15340), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n15331), .C1(n15330), .C2(n15329), .ZN(
        n15339) );
  INV_X1 U16934 ( .A(n15332), .ZN(n15335) );
  OAI211_X1 U16935 ( .C1(n15348), .C2(n15335), .A(n15334), .B(n15333), .ZN(
        n15347) );
  INV_X1 U16936 ( .A(n15347), .ZN(n15336) );
  AOI22_X1 U16937 ( .A1(n15352), .A2(n15337), .B1(n15235), .B2(n15336), .ZN(
        n15338) );
  OAI211_X1 U16938 ( .C1(n15340), .C2(n15349), .A(n15339), .B(n15338), .ZN(
        P1_U3291) );
  AND2_X1 U16939 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15341), .ZN(P1_U3294) );
  AND2_X1 U16940 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15341), .ZN(P1_U3295) );
  AND2_X1 U16941 ( .A1(n15341), .A2(P1_D_REG_29__SCAN_IN), .ZN(P1_U3296) );
  AND2_X1 U16942 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15341), .ZN(P1_U3297) );
  AND2_X1 U16943 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15341), .ZN(P1_U3298) );
  AND2_X1 U16944 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15341), .ZN(P1_U3299) );
  AND2_X1 U16945 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15341), .ZN(P1_U3300) );
  AND2_X1 U16946 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15341), .ZN(P1_U3301) );
  AND2_X1 U16947 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15341), .ZN(P1_U3302) );
  AND2_X1 U16948 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15341), .ZN(P1_U3303) );
  AND2_X1 U16949 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15341), .ZN(P1_U3304) );
  AND2_X1 U16950 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15341), .ZN(P1_U3305) );
  AND2_X1 U16951 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15341), .ZN(P1_U3306) );
  AND2_X1 U16952 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15341), .ZN(P1_U3307) );
  AND2_X1 U16953 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15341), .ZN(P1_U3308) );
  AND2_X1 U16954 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15341), .ZN(P1_U3309) );
  AND2_X1 U16955 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15341), .ZN(P1_U3310) );
  AND2_X1 U16956 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15341), .ZN(P1_U3311) );
  AND2_X1 U16957 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15341), .ZN(P1_U3312) );
  AND2_X1 U16958 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15341), .ZN(P1_U3313) );
  AND2_X1 U16959 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15341), .ZN(P1_U3314) );
  AND2_X1 U16960 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15341), .ZN(P1_U3315) );
  AND2_X1 U16961 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15341), .ZN(P1_U3316) );
  AND2_X1 U16962 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15341), .ZN(P1_U3317) );
  AND2_X1 U16963 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15341), .ZN(P1_U3318) );
  AND2_X1 U16964 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15341), .ZN(P1_U3319) );
  AND2_X1 U16965 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15341), .ZN(P1_U3320) );
  AND2_X1 U16966 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15341), .ZN(P1_U3321) );
  AND2_X1 U16967 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15341), .ZN(P1_U3322) );
  AND2_X1 U16968 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15341), .ZN(P1_U3323) );
  OAI21_X1 U16969 ( .B1(n15343), .B2(n15363), .A(n15342), .ZN(n15345) );
  AOI211_X1 U16970 ( .C1(n15353), .C2(n15346), .A(n15345), .B(n15344), .ZN(
        n15410) );
  AOI22_X1 U16971 ( .A1(n15408), .A2(n15410), .B1(n9238), .B2(n15406), .ZN(
        P1_U3462) );
  OAI21_X1 U16972 ( .B1(n15348), .B2(n15363), .A(n15347), .ZN(n15351) );
  INV_X1 U16973 ( .A(n15349), .ZN(n15350) );
  AOI211_X1 U16974 ( .C1(n15353), .C2(n15352), .A(n15351), .B(n15350), .ZN(
        n15412) );
  AOI22_X1 U16975 ( .A1(n15408), .A2(n15412), .B1(n9258), .B2(n15406), .ZN(
        P1_U3465) );
  INV_X1 U16976 ( .A(n15358), .ZN(n15360) );
  AOI21_X1 U16977 ( .B1(n15400), .B2(n15355), .A(n15354), .ZN(n15356) );
  OAI211_X1 U16978 ( .C1(n15358), .C2(n15374), .A(n15357), .B(n15356), .ZN(
        n15359) );
  AOI21_X1 U16979 ( .B1(n15361), .B2(n15360), .A(n15359), .ZN(n15413) );
  INV_X1 U16980 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15362) );
  AOI22_X1 U16981 ( .A1(n15408), .A2(n15413), .B1(n15362), .B2(n15406), .ZN(
        P1_U3474) );
  NOR2_X1 U16982 ( .A1(n15369), .A2(n15375), .ZN(n15371) );
  OAI22_X1 U16983 ( .A1(n15366), .A2(n15365), .B1(n15364), .B2(n15363), .ZN(
        n15367) );
  INV_X1 U16984 ( .A(n15367), .ZN(n15368) );
  OAI21_X1 U16985 ( .B1(n15369), .B2(n15374), .A(n15368), .ZN(n15370) );
  NOR3_X1 U16986 ( .A1(n15372), .A2(n15371), .A3(n15370), .ZN(n15414) );
  AOI22_X1 U16987 ( .A1(n15408), .A2(n15414), .B1(n9310), .B2(n15406), .ZN(
        P1_U3477) );
  OAI21_X1 U16988 ( .B1(n15374), .B2(n15376), .A(n15373), .ZN(n15380) );
  NOR2_X1 U16989 ( .A1(n15376), .A2(n15375), .ZN(n15377) );
  NOR4_X1 U16990 ( .A1(n15380), .A2(n15379), .A3(n15378), .A4(n15377), .ZN(
        n15415) );
  INV_X1 U16991 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15381) );
  AOI22_X1 U16992 ( .A1(n15408), .A2(n15415), .B1(n15381), .B2(n15406), .ZN(
        P1_U3480) );
  NAND4_X1 U16993 ( .A1(n15385), .A2(n15384), .A3(n15383), .A4(n15382), .ZN(
        n15386) );
  AOI21_X1 U16994 ( .B1(n15387), .B2(n15395), .A(n15386), .ZN(n15416) );
  INV_X1 U16995 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15388) );
  AOI22_X1 U16996 ( .A1(n15408), .A2(n15416), .B1(n15388), .B2(n15406), .ZN(
        P1_U3483) );
  INV_X1 U16997 ( .A(n15389), .ZN(n15396) );
  AOI21_X1 U16998 ( .B1(n15396), .B2(n15395), .A(n15394), .ZN(n15417) );
  INV_X1 U16999 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15397) );
  AOI22_X1 U17000 ( .A1(n15408), .A2(n15417), .B1(n15397), .B2(n15406), .ZN(
        P1_U3486) );
  AOI21_X1 U17001 ( .B1(n15400), .B2(n15399), .A(n15398), .ZN(n15401) );
  OAI211_X1 U17002 ( .C1(n15404), .C2(n15403), .A(n15402), .B(n15401), .ZN(
        n15405) );
  INV_X1 U17003 ( .A(n15405), .ZN(n15419) );
  INV_X1 U17004 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U17005 ( .A1(n15408), .A2(n15419), .B1(n15407), .B2(n15406), .ZN(
        P1_U3489) );
  AOI22_X1 U17006 ( .A1(n15420), .A2(n15410), .B1(n15409), .B2(n15418), .ZN(
        P1_U3529) );
  AOI22_X1 U17007 ( .A1(n15420), .A2(n15412), .B1(n15411), .B2(n15418), .ZN(
        P1_U3530) );
  AOI22_X1 U17008 ( .A1(n15420), .A2(n15413), .B1(n10684), .B2(n15418), .ZN(
        P1_U3533) );
  AOI22_X1 U17009 ( .A1(n15420), .A2(n15414), .B1(n10687), .B2(n15418), .ZN(
        P1_U3534) );
  AOI22_X1 U17010 ( .A1(n15420), .A2(n15415), .B1(n9229), .B2(n15418), .ZN(
        P1_U3535) );
  AOI22_X1 U17011 ( .A1(n15420), .A2(n15416), .B1(n9328), .B2(n15418), .ZN(
        P1_U3536) );
  AOI22_X1 U17012 ( .A1(n15420), .A2(n15417), .B1(n10873), .B2(n15418), .ZN(
        P1_U3537) );
  AOI22_X1 U17013 ( .A1(n15420), .A2(n15419), .B1(n9341), .B2(n15418), .ZN(
        P1_U3538) );
  NOR2_X1 U17014 ( .A1(n15441), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U17015 ( .A1(n15508), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n15471), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15425) );
  OAI22_X1 U17016 ( .A1(n15513), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n15421), .ZN(n15422) );
  NOR2_X1 U17017 ( .A1(n15519), .A2(n15422), .ZN(n15424) );
  AOI22_X1 U17018 ( .A1(n15441), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15423) );
  OAI221_X1 U17019 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n15425), .C1(n6686), .C2(
        n15424), .A(n15423), .ZN(P2_U3214) );
  OAI21_X1 U17020 ( .B1(n15428), .B2(n15427), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15429) );
  OAI21_X1 U17021 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15429), .ZN(n15443) );
  OAI211_X1 U17022 ( .C1(n15432), .C2(n15431), .A(n15508), .B(n15430), .ZN(
        n15433) );
  INV_X1 U17023 ( .A(n15433), .ZN(n15440) );
  INV_X1 U17024 ( .A(n15434), .ZN(n15437) );
  INV_X1 U17025 ( .A(n15435), .ZN(n15436) );
  AOI211_X1 U17026 ( .C1(n15438), .C2(n15437), .A(n15436), .B(n15513), .ZN(
        n15439) );
  AOI211_X1 U17027 ( .C1(n15441), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n15440), .B(
        n15439), .ZN(n15442) );
  NAND2_X1 U17028 ( .A1(n15443), .A2(n15442), .ZN(P2_U3215) );
  OAI211_X1 U17029 ( .C1(n15446), .C2(n15445), .A(n15508), .B(n15444), .ZN(
        n15451) );
  OAI211_X1 U17030 ( .C1(n15449), .C2(n15448), .A(n15471), .B(n15447), .ZN(
        n15450) );
  NAND2_X1 U17031 ( .A1(n15451), .A2(n15450), .ZN(n15452) );
  AOI21_X1 U17032 ( .B1(n15453), .B2(n15519), .A(n15452), .ZN(n15455) );
  NAND2_X1 U17033 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n15454) );
  OAI211_X1 U17034 ( .C1(n15522), .C2(n15456), .A(n15455), .B(n15454), .ZN(
        P2_U3217) );
  OAI211_X1 U17035 ( .C1(n15459), .C2(n15458), .A(n15508), .B(n15457), .ZN(
        n15464) );
  OAI211_X1 U17036 ( .C1(n15462), .C2(n15461), .A(n15471), .B(n15460), .ZN(
        n15463) );
  NAND2_X1 U17037 ( .A1(n15464), .A2(n15463), .ZN(n15465) );
  AOI21_X1 U17038 ( .B1(n15466), .B2(n15519), .A(n15465), .ZN(n15468) );
  OAI211_X1 U17039 ( .C1(n15522), .C2(n15469), .A(n15468), .B(n15467), .ZN(
        P2_U3219) );
  OAI211_X1 U17040 ( .C1(n15473), .C2(n15472), .A(n15471), .B(n15470), .ZN(
        n15478) );
  OAI211_X1 U17041 ( .C1(n15476), .C2(n15475), .A(n15508), .B(n15474), .ZN(
        n15477) );
  OAI211_X1 U17042 ( .C1(n15490), .C2(n15479), .A(n15478), .B(n15477), .ZN(
        n15480) );
  INV_X1 U17043 ( .A(n15480), .ZN(n15482) );
  NAND2_X1 U17044 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n15481) );
  OAI211_X1 U17045 ( .C1(n15522), .C2(n9149), .A(n15482), .B(n15481), .ZN(
        P2_U3220) );
  AOI211_X1 U17046 ( .C1(n15484), .C2(n15483), .A(n15513), .B(n6502), .ZN(
        n15492) );
  OAI211_X1 U17047 ( .C1(n15487), .C2(n15486), .A(n15508), .B(n15485), .ZN(
        n15488) );
  OAI21_X1 U17048 ( .B1(n15490), .B2(n15489), .A(n15488), .ZN(n15491) );
  NOR2_X1 U17049 ( .A1(n15492), .A2(n15491), .ZN(n15494) );
  NAND2_X1 U17050 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n15493) );
  OAI211_X1 U17051 ( .C1(n15495), .C2(n15522), .A(n15494), .B(n15493), .ZN(
        P2_U3222) );
  OAI211_X1 U17052 ( .C1(n15498), .C2(n15497), .A(n15496), .B(n15508), .ZN(
        n15499) );
  INV_X1 U17053 ( .A(n15499), .ZN(n15503) );
  AOI211_X1 U17054 ( .C1(n15501), .C2(n15500), .A(n15513), .B(n6514), .ZN(
        n15502) );
  AOI211_X1 U17055 ( .C1(n15519), .C2(n15504), .A(n15503), .B(n15502), .ZN(
        n15506) );
  OAI211_X1 U17056 ( .C1(n15507), .C2(n15522), .A(n15506), .B(n15505), .ZN(
        P2_U3230) );
  OAI211_X1 U17057 ( .C1(n15511), .C2(n15510), .A(n15509), .B(n15508), .ZN(
        n15512) );
  INV_X1 U17058 ( .A(n15512), .ZN(n15517) );
  AOI211_X1 U17059 ( .C1(n15515), .C2(n15514), .A(n15513), .B(n6494), .ZN(
        n15516) );
  AOI211_X1 U17060 ( .C1(n15519), .C2(n15518), .A(n15517), .B(n15516), .ZN(
        n15521) );
  OAI211_X1 U17061 ( .C1(n15523), .C2(n15522), .A(n15521), .B(n15520), .ZN(
        P2_U3231) );
  INV_X1 U17062 ( .A(n15533), .ZN(n15530) );
  NOR2_X1 U17063 ( .A1(n15530), .A2(n15524), .ZN(n15526) );
  AND2_X1 U17064 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15527), .ZN(P2_U3266) );
  AND2_X1 U17065 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15527), .ZN(P2_U3267) );
  AND2_X1 U17066 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15527), .ZN(P2_U3268) );
  AND2_X1 U17067 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15527), .ZN(P2_U3269) );
  AND2_X1 U17068 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15527), .ZN(P2_U3270) );
  AND2_X1 U17069 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15527), .ZN(P2_U3271) );
  AND2_X1 U17070 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15527), .ZN(P2_U3272) );
  AND2_X1 U17071 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15527), .ZN(P2_U3273) );
  AND2_X1 U17072 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15527), .ZN(P2_U3274) );
  AND2_X1 U17073 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15527), .ZN(P2_U3275) );
  AND2_X1 U17074 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15527), .ZN(P2_U3276) );
  AND2_X1 U17075 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15527), .ZN(P2_U3277) );
  AND2_X1 U17076 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15527), .ZN(P2_U3278) );
  AND2_X1 U17077 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15527), .ZN(P2_U3279) );
  AND2_X1 U17078 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15527), .ZN(P2_U3280) );
  AND2_X1 U17079 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15527), .ZN(P2_U3281) );
  AND2_X1 U17080 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15527), .ZN(P2_U3282) );
  AND2_X1 U17081 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15527), .ZN(P2_U3283) );
  AND2_X1 U17082 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15527), .ZN(P2_U3284) );
  AND2_X1 U17083 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15527), .ZN(P2_U3285) );
  AND2_X1 U17084 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15527), .ZN(P2_U3286) );
  AND2_X1 U17085 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15527), .ZN(P2_U3287) );
  AND2_X1 U17086 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15527), .ZN(P2_U3288) );
  AND2_X1 U17087 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15527), .ZN(P2_U3289) );
  AND2_X1 U17088 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15527), .ZN(P2_U3290) );
  NOR2_X1 U17089 ( .A1(n15526), .A2(n15525), .ZN(P2_U3291) );
  AND2_X1 U17090 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15527), .ZN(P2_U3292) );
  AND2_X1 U17091 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15527), .ZN(P2_U3293) );
  AND2_X1 U17092 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15527), .ZN(P2_U3294) );
  AND2_X1 U17093 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15527), .ZN(P2_U3295) );
  AOI22_X1 U17094 ( .A1(n15533), .A2(n15529), .B1(n15528), .B2(n15530), .ZN(
        P2_U3416) );
  AOI22_X1 U17095 ( .A1(n15533), .A2(n15532), .B1(n15531), .B2(n15530), .ZN(
        P2_U3417) );
  AOI22_X1 U17096 ( .A1(n15561), .A2(n15534), .B1(n7621), .B2(n15559), .ZN(
        P2_U3430) );
  OAI21_X1 U17097 ( .B1(n15537), .B2(n15536), .A(n15535), .ZN(n15539) );
  AOI211_X1 U17098 ( .C1(n15541), .C2(n15540), .A(n15539), .B(n15538), .ZN(
        n15563) );
  AOI22_X1 U17099 ( .A1(n15561), .A2(n15563), .B1(n7900), .B2(n15559), .ZN(
        P2_U3436) );
  INV_X1 U17100 ( .A(n15547), .ZN(n15549) );
  AOI21_X1 U17101 ( .B1(n15553), .B2(n15543), .A(n15542), .ZN(n15544) );
  OAI211_X1 U17102 ( .C1(n15547), .C2(n15546), .A(n15545), .B(n15544), .ZN(
        n15548) );
  AOI21_X1 U17103 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(n15566) );
  AOI22_X1 U17104 ( .A1(n15561), .A2(n15566), .B1(n8005), .B2(n15559), .ZN(
        P2_U3448) );
  AOI21_X1 U17105 ( .B1(n15553), .B2(n15552), .A(n15551), .ZN(n15555) );
  OAI211_X1 U17106 ( .C1(n15557), .C2(n15556), .A(n15555), .B(n15554), .ZN(
        n15558) );
  INV_X1 U17107 ( .A(n15558), .ZN(n15568) );
  INV_X1 U17108 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15560) );
  AOI22_X1 U17109 ( .A1(n15561), .A2(n15568), .B1(n15560), .B2(n15559), .ZN(
        P2_U3451) );
  AOI22_X1 U17110 ( .A1(n15564), .A2(n15563), .B1(n15562), .B2(n15567), .ZN(
        P2_U3501) );
  AOI22_X1 U17111 ( .A1(n15569), .A2(n15566), .B1(n15565), .B2(n15567), .ZN(
        P2_U3505) );
  AOI22_X1 U17112 ( .A1(n15569), .A2(n15568), .B1(n8019), .B2(n15567), .ZN(
        P2_U3506) );
  NOR2_X1 U17113 ( .A1(P3_U3897), .A2(n15570), .ZN(P3_U3150) );
  INV_X1 U17114 ( .A(n15571), .ZN(n15590) );
  XNOR2_X1 U17115 ( .A(n15572), .B(n15578), .ZN(n15587) );
  INV_X1 U17116 ( .A(n15587), .ZN(n15616) );
  AND2_X1 U17117 ( .A1(n15573), .A2(n15623), .ZN(n15615) );
  INV_X1 U17118 ( .A(n15615), .ZN(n15574) );
  OAI22_X1 U17119 ( .A1(n15577), .A2(n15576), .B1(n15575), .B2(n15574), .ZN(
        n15589) );
  XNOR2_X1 U17120 ( .A(n15579), .B(n15578), .ZN(n15585) );
  OAI22_X1 U17121 ( .A1(n15583), .A2(n15582), .B1(n15581), .B2(n15580), .ZN(
        n15584) );
  AOI21_X1 U17122 ( .B1(n15585), .B2(n10349), .A(n15584), .ZN(n15586) );
  OAI21_X1 U17123 ( .B1(n15588), .B2(n15587), .A(n15586), .ZN(n15614) );
  AOI211_X1 U17124 ( .C1(n15590), .C2(n15616), .A(n15589), .B(n15614), .ZN(
        n15591) );
  AOI22_X1 U17125 ( .A1(n15610), .A2(n15592), .B1(n15591), .B2(n15608), .ZN(
        P3_U3231) );
  NOR2_X1 U17126 ( .A1(n15593), .A2(n15638), .ZN(n15612) );
  XOR2_X1 U17127 ( .A(n15594), .B(n11040), .Z(n15602) );
  AOI22_X1 U17128 ( .A1(n15597), .A2(n10259), .B1(n15596), .B2(n15595), .ZN(
        n15600) );
  XNOR2_X1 U17129 ( .A(n15598), .B(n11040), .ZN(n15613) );
  NAND2_X1 U17130 ( .A1(n15613), .A2(n15642), .ZN(n15599) );
  OAI211_X1 U17131 ( .C1(n15602), .C2(n15601), .A(n15600), .B(n15599), .ZN(
        n15611) );
  AOI21_X1 U17132 ( .B1(n15612), .B2(n15603), .A(n15611), .ZN(n15609) );
  AOI22_X1 U17133 ( .A1(n15605), .A2(n15613), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15604), .ZN(n15606) );
  OAI221_X1 U17134 ( .B1(n15610), .B2(n15609), .C1(n15608), .C2(n15607), .A(
        n15606), .ZN(P3_U3232) );
  AOI211_X1 U17135 ( .C1(n15635), .C2(n15613), .A(n15612), .B(n15611), .ZN(
        n15646) );
  AOI22_X1 U17136 ( .A1(n15645), .A2(n15646), .B1(n9724), .B2(n15643), .ZN(
        P3_U3393) );
  AOI211_X1 U17137 ( .C1(n15616), .C2(n15635), .A(n15615), .B(n15614), .ZN(
        n15647) );
  INV_X1 U17138 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U17139 ( .A1(n15645), .A2(n15647), .B1(n15617), .B2(n15643), .ZN(
        P3_U3396) );
  INV_X1 U17140 ( .A(n15618), .ZN(n15619) );
  AOI211_X1 U17141 ( .C1(n15635), .C2(n15621), .A(n15620), .B(n15619), .ZN(
        n15648) );
  AOI22_X1 U17142 ( .A1(n15645), .A2(n15648), .B1(n9780), .B2(n15643), .ZN(
        P3_U3399) );
  AOI21_X1 U17143 ( .B1(n15624), .B2(n15623), .A(n15622), .ZN(n15625) );
  OAI21_X1 U17144 ( .B1(n15627), .B2(n15626), .A(n15625), .ZN(n15628) );
  AOI21_X1 U17145 ( .B1(n15642), .B2(n15629), .A(n15628), .ZN(n15649) );
  AOI22_X1 U17146 ( .A1(n15645), .A2(n15649), .B1(n9801), .B2(n15643), .ZN(
        P3_U3402) );
  INV_X1 U17147 ( .A(n15630), .ZN(n15632) );
  AOI211_X1 U17148 ( .C1(n15633), .C2(n15635), .A(n15632), .B(n15631), .ZN(
        n15650) );
  INV_X1 U17149 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15634) );
  AOI22_X1 U17150 ( .A1(n15645), .A2(n15650), .B1(n15634), .B2(n15643), .ZN(
        P3_U3405) );
  NAND2_X1 U17151 ( .A1(n15641), .A2(n15635), .ZN(n15636) );
  OAI211_X1 U17152 ( .C1(n15639), .C2(n15638), .A(n15637), .B(n15636), .ZN(
        n15640) );
  AOI21_X1 U17153 ( .B1(n15642), .B2(n15641), .A(n15640), .ZN(n15651) );
  INV_X1 U17154 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15644) );
  AOI22_X1 U17155 ( .A1(n15645), .A2(n15651), .B1(n15644), .B2(n15643), .ZN(
        P3_U3408) );
  AOI22_X1 U17156 ( .A1(n15652), .A2(n15646), .B1(n10968), .B2(n7202), .ZN(
        P3_U3460) );
  AOI22_X1 U17157 ( .A1(n15652), .A2(n15647), .B1(n10919), .B2(n7202), .ZN(
        P3_U3461) );
  AOI22_X1 U17158 ( .A1(n15652), .A2(n15648), .B1(n11003), .B2(n7202), .ZN(
        P3_U3462) );
  AOI22_X1 U17159 ( .A1(n15652), .A2(n15649), .B1(n10901), .B2(n7202), .ZN(
        P3_U3463) );
  AOI22_X1 U17160 ( .A1(n15652), .A2(n15650), .B1(n9827), .B2(n7202), .ZN(
        P3_U3464) );
  AOI22_X1 U17161 ( .A1(n15652), .A2(n15651), .B1(n10906), .B2(n7202), .ZN(
        P3_U3465) );
  XNOR2_X1 U17162 ( .A(n15653), .B(n15654), .ZN(SUB_1596_U59) );
  XNOR2_X1 U17163 ( .A(n15655), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17164 ( .B1(n15657), .B2(n15656), .A(n15665), .ZN(SUB_1596_U53) );
  XNOR2_X1 U17165 ( .A(n15659), .B(n15658), .ZN(SUB_1596_U56) );
  OAI21_X1 U17166 ( .B1(n15662), .B2(n15661), .A(n15660), .ZN(n15663) );
  XNOR2_X1 U17167 ( .A(n15663), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U17168 ( .A(n15665), .B(n15664), .Z(SUB_1596_U5) );
  CLKBUF_X3 U7193 ( .A(n8579), .Z(n8726) );
  INV_X2 U9125 ( .A(n9284), .ZN(n9649) );
  CLKBUF_X2 U9275 ( .A(n8856), .Z(n8948) );
endmodule

