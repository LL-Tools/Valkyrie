

module b15_C_SARLock_k_128_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954;

  OR2_X1 U3581 ( .A1(n5381), .A2(n4299), .ZN(n5545) );
  NAND2_X1 U3582 ( .A1(n5070), .A2(n5069), .ZN(n5068) );
  NAND2_X1 U3583 ( .A1(n3921), .A2(n4336), .ZN(n3934) );
  NAND2_X2 U3584 ( .A1(n3976), .A2(n4672), .ZN(n4069) );
  AND2_X1 U3585 ( .A1(n3891), .A2(n4688), .ZN(n3921) );
  CLKBUF_X2 U3586 ( .A(n3722), .Z(n4250) );
  CLKBUF_X2 U3588 ( .A(n3335), .Z(n4246) );
  CLKBUF_X2 U3589 ( .A(n3406), .Z(n3135) );
  CLKBUF_X2 U3590 ( .A(n3336), .Z(n4247) );
  CLKBUF_X2 U3591 ( .A(n3372), .Z(n3358) );
  NOR2_X2 U3592 ( .A1(n3300), .A2(n3301), .ZN(n5247) );
  CLKBUF_X1 U3593 ( .A(n3304), .Z(n4688) );
  CLKBUF_X1 U3594 ( .A(n3292), .Z(n3301) );
  NAND4_X2 U3595 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3160), .ZN(n3300)
         );
  AND4_X1 U3596 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3250)
         );
  AND2_X1 U3597 ( .A1(n3170), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3178)
         );
  AOI22_X1 U3598 ( .A1(n6904), .A2(keyinput36), .B1(ADDRESS_REG_18__SCAN_IN), 
        .B2(n6903), .ZN(n6902) );
  AND2_X1 U3599 ( .A1(n3170), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3141)
         );
  OAI221_X1 U3600 ( .B1(n6904), .B2(keyinput36), .C1(n6903), .C2(
        ADDRESS_REG_18__SCAN_IN), .A(n6902), .ZN(n6913) );
  CLKBUF_X2 U3601 ( .A(n3270), .Z(n4249) );
  AOI22_X1 U3602 ( .A1(n6842), .A2(keyinput43), .B1(n6841), .B2(keyinput72), 
        .ZN(n6840) );
  AND4_X1 U3603 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3231)
         );
  INV_X1 U3604 ( .A(n3301), .ZN(n4362) );
  OAI221_X1 U3605 ( .B1(n6842), .B2(keyinput43), .C1(n6841), .C2(keyinput72), 
        .A(n6840), .ZN(n6937) );
  NAND3_X1 U3606 ( .A1(n5990), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5965) );
  NAND4_X1 U3607 ( .A1(n3253), .A2(n3252), .A3(n3251), .A4(n3250), .ZN(n3292)
         );
  INV_X1 U3608 ( .A(n4238), .ZN(n4217) );
  OR2_X2 U3609 ( .A1(n4621), .A2(n4620), .ZN(n5034) );
  AND2_X1 U3610 ( .A1(n5800), .A2(n3974), .ZN(n5773) );
  OR2_X1 U3611 ( .A1(n3214), .A2(n3213), .ZN(n4648) );
  CLKBUF_X3 U3612 ( .A(n3292), .Z(n4672) );
  INV_X1 U3613 ( .A(n5588), .ZN(n6283) );
  NAND2_X1 U3614 ( .A1(n4290), .A2(n4289), .ZN(n5569) );
  INV_X1 U3615 ( .A(n6070), .ZN(n6081) );
  INV_X1 U3616 ( .A(n6120), .ZN(n6108) );
  OR2_X2 U3617 ( .A1(n5068), .A2(n5059), .ZN(n3132) );
  AND2_X2 U3618 ( .A1(n3143), .A2(n3144), .ZN(n4159) );
  NAND2_X2 U3620 ( .A1(n4186), .A2(n3161), .ZN(n4290) );
  BUF_X4 U3621 ( .A(n3285), .Z(n3303) );
  OAI21_X2 U3622 ( .B1(n3325), .B2(n4346), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3329) );
  NOR2_X2 U3623 ( .A1(n6561), .A2(n5965), .ZN(n5845) );
  XNOR2_X2 U3624 ( .A(n3423), .B(n3422), .ZN(n4511) );
  NAND2_X2 U3625 ( .A1(n3396), .A2(n3395), .ZN(n3423) );
  NOR2_X1 U3626 ( .A1(n5515), .A2(n4199), .ZN(n4313) );
  CLKBUF_X2 U3627 ( .A(n6184), .Z(n6202) );
  OR2_X2 U3628 ( .A1(n6611), .A2(n3949), .ZN(n5262) );
  CLKBUF_X1 U3629 ( .A(n3397), .Z(n3398) );
  NAND2_X2 U3630 ( .A1(n4149), .A2(n3429), .ZN(n3930) );
  INV_X4 U3631 ( .A(n4535), .ZN(n5455) );
  OR2_X2 U3632 ( .A1(n3287), .A2(n3976), .ZN(n3310) );
  NAND2_X1 U3633 ( .A1(n3195), .A2(n3194), .ZN(n3285) );
  CLKBUF_X2 U3635 ( .A(n3369), .Z(n4251) );
  CLKBUF_X2 U3636 ( .A(n3370), .Z(n4259) );
  CLKBUF_X2 U3637 ( .A(n3407), .Z(n3357) );
  CLKBUF_X2 U3638 ( .A(n3337), .Z(n4258) );
  NOR2_X1 U3639 ( .A1(n5556), .A2(n4396), .ZN(n4325) );
  CLKBUF_X1 U3640 ( .A(n4290), .Z(n5653) );
  CLKBUF_X1 U3641 ( .A(n4291), .Z(n4292) );
  NAND2_X1 U3642 ( .A1(n4306), .A2(n4304), .ZN(n5681) );
  CLKBUF_X1 U3643 ( .A(n5571), .Z(n5787) );
  CLKBUF_X1 U3644 ( .A(n5353), .Z(n5598) );
  OR2_X1 U3645 ( .A1(n5383), .A2(n5382), .ZN(n5470) );
  INV_X1 U3646 ( .A(n4315), .ZN(n5497) );
  NOR2_X2 U3647 ( .A1(n5515), .A2(n5517), .ZN(n5516) );
  NAND2_X1 U3648 ( .A1(n5518), .A2(n5520), .ZN(n5515) );
  CLKBUF_X1 U3649 ( .A(n5518), .Z(n5532) );
  NAND2_X1 U3650 ( .A1(n5278), .A2(n5277), .ZN(n6206) );
  NOR2_X1 U3651 ( .A1(n5336), .A2(n5335), .ZN(n5334) );
  CLKBUF_X1 U3652 ( .A(n5295), .Z(n5304) );
  NAND2_X1 U3653 ( .A1(n5295), .A2(n5303), .ZN(n5336) );
  NAND2_X1 U3654 ( .A1(n5232), .A2(n5236), .ZN(n5297) );
  CLKBUF_X1 U3655 ( .A(n5232), .Z(n5237) );
  NOR2_X2 U3656 ( .A1(n5343), .A2(n5342), .ZN(n5348) );
  OAI21_X1 U3657 ( .B1(n4110), .B2(n4139), .A(n4109), .ZN(n4111) );
  NAND2_X2 U3658 ( .A1(n3150), .A2(n3528), .ZN(n4110) );
  XNOR2_X1 U3659 ( .A(n3151), .B(n3489), .ZN(n4626) );
  OAI21_X2 U3660 ( .B1(n4090), .B2(n4139), .A(n4089), .ZN(n4465) );
  XNOR2_X1 U3661 ( .A(n3491), .B(n3494), .ZN(n4082) );
  NAND2_X1 U3662 ( .A1(n4532), .A2(n4425), .ZN(n6611) );
  CLKBUF_X1 U3663 ( .A(n4471), .Z(n6368) );
  NAND2_X1 U3664 ( .A1(n3501), .A2(n3502), .ZN(n3505) );
  INV_X2 U3665 ( .A(n6134), .ZN(n3133) );
  OR2_X2 U3666 ( .A1(n4489), .A2(n6510), .ZN(n4566) );
  CLKBUF_X1 U3667 ( .A(n4600), .Z(n5447) );
  NOR2_X1 U3668 ( .A1(n4580), .A2(n4614), .ZN(n4002) );
  NAND2_X1 U3669 ( .A1(n3405), .A2(n3404), .ZN(n3422) );
  NAND2_X1 U3670 ( .A1(n3993), .A2(n3992), .ZN(n4607) );
  CLKBUF_X1 U3671 ( .A(n4346), .Z(n5929) );
  CLKBUF_X1 U3672 ( .A(n4329), .Z(n4537) );
  NAND2_X1 U3673 ( .A1(n3324), .A2(n3323), .ZN(n3939) );
  OAI21_X1 U3674 ( .B1(n4333), .B2(n5540), .A(n4534), .ZN(n3266) );
  OR2_X1 U3675 ( .A1(n4572), .A2(n3320), .ZN(n4357) );
  NAND2_X1 U3676 ( .A1(n3305), .A2(n4431), .ZN(n4509) );
  AND4_X1 U3677 ( .A1(n4335), .A2(n4362), .A3(n4648), .A4(n4688), .ZN(n3305)
         );
  AND3_X1 U3678 ( .A1(n3269), .A2(n4648), .A3(n3284), .ZN(n4370) );
  MUX2_X1 U3679 ( .A(n3288), .B(n3286), .S(n3303), .Z(n3291) );
  NAND2_X1 U3680 ( .A1(n4570), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4149) );
  INV_X1 U3681 ( .A(n3303), .ZN(n4335) );
  INV_X1 U3682 ( .A(n4648), .ZN(n5540) );
  AND4_X1 U3683 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(n3233)
         );
  AND4_X1 U3684 ( .A1(n3237), .A2(n3236), .A3(n3235), .A4(n3234), .ZN(n3253)
         );
  CLKBUF_X2 U3685 ( .A(n3276), .Z(n4257) );
  AND4_X1 U3686 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), .ZN(n3194)
         );
  AND4_X1 U3687 ( .A1(n3189), .A2(n3187), .A3(n3188), .A4(n3186), .ZN(n3195)
         );
  AND4_X1 U3688 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(n3281)
         );
  AND4_X1 U3689 ( .A1(n3222), .A2(n3221), .A3(n3220), .A4(n3219), .ZN(n3232)
         );
  AND4_X1 U3690 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3251)
         );
  AOI22_X1 U3691 ( .A1(n3406), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3186) );
  BUF_X2 U3692 ( .A(n3805), .Z(n4256) );
  INV_X2 U3693 ( .A(n6581), .ZN(n3134) );
  AND2_X2 U3694 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4483) );
  INV_X1 U3695 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3177) );
  OR2_X2 U3696 ( .A1(n5472), .A2(n5473), .ZN(n5469) );
  CLKBUF_X1 U3697 ( .A(n6252), .Z(n3136) );
  CLKBUF_X1 U3698 ( .A(n6244), .Z(n3137) );
  NOR2_X1 U3699 ( .A1(n5556), .A2(n4396), .ZN(n3138) );
  INV_X1 U3700 ( .A(n5889), .ZN(n3139) );
  NAND2_X1 U3701 ( .A1(n3351), .A2(n3350), .ZN(n3140) );
  INV_X1 U3702 ( .A(n4845), .ZN(n3142) );
  NAND2_X1 U3703 ( .A1(n3505), .A2(n3504), .ZN(n4090) );
  NOR2_X4 U3704 ( .A1(n5034), .A2(n5035), .ZN(n5070) );
  OR2_X2 U3705 ( .A1(n5307), .A2(n5306), .ZN(n5343) );
  NOR2_X2 U3706 ( .A1(n3132), .A2(n5230), .ZN(n5229) );
  NAND2_X1 U3708 ( .A1(n6222), .A2(n3146), .ZN(n3143) );
  OR2_X1 U3709 ( .A1(n3145), .A2(n4158), .ZN(n3144) );
  INV_X1 U3710 ( .A(n6215), .ZN(n3145) );
  AND2_X1 U3711 ( .A1(n6224), .A2(n6215), .ZN(n3146) );
  NAND2_X1 U3712 ( .A1(n4159), .A2(n6216), .ZN(n3147) );
  OAI21_X1 U3713 ( .B1(n6206), .B2(n4163), .A(n4162), .ZN(n3148) );
  AOI21_X1 U3714 ( .B1(n5681), .B2(n5683), .A(n5682), .ZN(n3149) );
  OR2_X2 U3715 ( .A1(n3527), .A2(n4627), .ZN(n3150) );
  XNOR2_X1 U3716 ( .A(n3152), .B(n3420), .ZN(n3151) );
  OAI22_X1 U3717 ( .A1(n4511), .A2(STATE2_REG_0__SCAN_IN), .B1(n4105), .B2(
        n4149), .ZN(n3152) );
  OAI21_X1 U3718 ( .B1(n5353), .B2(n4170), .A(n5599), .ZN(n4174) );
  AOI21_X1 U3719 ( .B1(n5681), .B2(n5683), .A(n5682), .ZN(n5592) );
  OAI21_X1 U3720 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5423), .A(n5422), 
        .ZN(n5424) );
  AND2_X1 U3721 ( .A1(n3141), .A2(n5450), .ZN(n3153) );
  AND2_X1 U3722 ( .A1(n3178), .A2(n5450), .ZN(n3154) );
  AND2_X2 U3723 ( .A1(n3141), .A2(n5450), .ZN(n3407) );
  AND2_X1 U3724 ( .A1(n5450), .A2(n3179), .ZN(n3155) );
  AND2_X1 U3725 ( .A1(n5450), .A2(n3179), .ZN(n3156) );
  AND2_X4 U3726 ( .A1(n5443), .A2(n4484), .ZN(n3369) );
  AND2_X1 U3727 ( .A1(n5443), .A2(n4483), .ZN(n3157) );
  AND2_X1 U3728 ( .A1(n4589), .A2(n4483), .ZN(n3158) );
  AND2_X1 U3729 ( .A1(n4589), .A2(n4483), .ZN(n3159) );
  NAND2_X1 U3730 ( .A1(n3284), .A2(n3268), .ZN(n3288) );
  OR2_X1 U3731 ( .A1(n3925), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3945)
         );
  AND2_X1 U3732 ( .A1(n5392), .A2(n5393), .ZN(n3885) );
  INV_X1 U3733 ( .A(n3304), .ZN(n3268) );
  AND2_X1 U3734 ( .A1(n4370), .A2(n4195), .ZN(n4347) );
  NAND2_X1 U3735 ( .A1(n3929), .A2(n3928), .ZN(n3944) );
  OR2_X1 U3736 ( .A1(n4377), .A2(n4482), .ZN(n5317) );
  OR2_X1 U3737 ( .A1(n4149), .A2(n3388), .ZN(n3344) );
  OR2_X1 U3738 ( .A1(n3927), .A2(n3926), .ZN(n3925) );
  AND2_X1 U3739 ( .A1(n4375), .A2(n4374), .ZN(n4429) );
  AND2_X1 U3740 ( .A1(n3884), .A2(n3885), .ZN(n4222) );
  NAND2_X1 U3741 ( .A1(n4535), .A2(n5460), .ZN(n4354) );
  NAND2_X1 U3742 ( .A1(n3204), .A2(n3166), .ZN(n3304) );
  AND2_X1 U3743 ( .A1(n4415), .A2(n3947), .ZN(n4411) );
  INV_X1 U3744 ( .A(n3938), .ZN(n4495) );
  OR2_X1 U3745 ( .A1(n6502), .A2(n3948), .ZN(n3949) );
  NAND2_X1 U3746 ( .A1(n4568), .A2(n6194), .ZN(n5373) );
  AND2_X1 U3747 ( .A1(n3883), .A2(n3882), .ZN(n5393) );
  AND2_X2 U3748 ( .A1(n5516), .A2(n5507), .ZN(n5496) );
  NAND2_X1 U3749 ( .A1(n3704), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3731)
         );
  NOR2_X1 U3750 ( .A1(n4896), .A2(n4897), .ZN(n5058) );
  NOR2_X1 U3751 ( .A1(n3557), .A2(n3556), .ZN(n3558) );
  NOR2_X1 U3752 ( .A1(n4618), .A2(n4619), .ZN(n4965) );
  NAND2_X1 U3753 ( .A1(n4613), .A2(n4611), .ZN(n4619) );
  AND2_X1 U3754 ( .A1(n4345), .A2(n4344), .ZN(n4377) );
  OR2_X1 U3755 ( .A1(n5730), .A2(n4794), .ZN(n5073) );
  OR2_X1 U3757 ( .A1(n3934), .A2(n3933), .ZN(n3935) );
  OAI21_X1 U3758 ( .B1(n5497), .B2(n4316), .A(n5490), .ZN(n5807) );
  AND2_X1 U3759 ( .A1(n5539), .A2(n5374), .ZN(n6948) );
  INV_X1 U3760 ( .A(n5539), .ZN(n6947) );
  XNOR2_X1 U3761 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .B(n3951), .ZN(n4285)
         );
  OR2_X1 U3762 ( .A1(n6779), .A2(n4245), .ZN(n3951) );
  AND2_X1 U3763 ( .A1(n5588), .A2(n4282), .ZN(n6257) );
  NOR2_X2 U3764 ( .A1(n4566), .A2(n6489), .ZN(n6272) );
  NAND2_X1 U3765 ( .A1(n4192), .A2(n4191), .ZN(n4193) );
  MUX2_X1 U3766 ( .A(n5457), .B(n3987), .S(n5469), .Z(n4356) );
  XNOR2_X1 U3767 ( .A(n4328), .B(n5609), .ZN(n4407) );
  NAND2_X1 U3768 ( .A1(n4327), .A2(n4326), .ZN(n4328) );
  XNOR2_X1 U3769 ( .A(n4311), .B(n4310), .ZN(n5435) );
  NAND2_X1 U3770 ( .A1(n5423), .A2(n4309), .ZN(n4311) );
  OR2_X1 U3771 ( .A1(n4306), .A2(n4308), .ZN(n4309) );
  NAND2_X1 U3772 ( .A1(n3386), .A2(n3503), .ZN(n3504) );
  NAND2_X1 U3773 ( .A1(n3140), .A2(n3503), .ZN(n3501) );
  INV_X1 U3774 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6485) );
  INV_X1 U3775 ( .A(n6368), .ZN(n5077) );
  OR2_X1 U3776 ( .A1(n3321), .A2(n4684), .ZN(n3282) );
  CLKBUF_X2 U3777 ( .A(n3371), .Z(n4248) );
  NAND2_X1 U3778 ( .A1(n3746), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3226)
         );
  INV_X1 U3779 ( .A(n3545), .ZN(n3468) );
  OR2_X1 U3780 ( .A1(n3478), .A2(n3477), .ZN(n4142) );
  OR2_X1 U3781 ( .A1(n3465), .A2(n3464), .ZN(n4132) );
  AND2_X1 U3782 ( .A1(n4509), .A2(n3306), .ZN(n3314) );
  AND2_X1 U3783 ( .A1(n4672), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3891) );
  NAND2_X1 U3784 ( .A1(n3284), .A2(n3319), .ZN(n3286) );
  AOI22_X1 U3785 ( .A1(n3412), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3203) );
  AOI22_X1 U3786 ( .A1(n3407), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3182) );
  AND2_X1 U3787 ( .A1(n3319), .A2(n4676), .ZN(n4365) );
  INV_X1 U3788 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3926) );
  AND2_X1 U3789 ( .A1(n4222), .A2(n4297), .ZN(n4296) );
  NOR2_X2 U3790 ( .A1(n5297), .A2(n5296), .ZN(n5295) );
  AND2_X1 U3791 ( .A1(n4164), .A2(n6679), .ZN(n4173) );
  OR2_X1 U3792 ( .A1(n3418), .A2(n3417), .ZN(n4097) );
  AND2_X1 U3793 ( .A1(n4684), .A2(n4361), .ZN(n4336) );
  INV_X1 U3794 ( .A(n4154), .ZN(n3382) );
  XNOR2_X1 U3795 ( .A(n3493), .B(n3492), .ZN(n3494) );
  OR2_X1 U3796 ( .A1(n3439), .A2(n3438), .ZN(n4114) );
  INV_X1 U3797 ( .A(n5730), .ZN(n5131) );
  XNOR2_X1 U3798 ( .A(n4591), .B(n4967), .ZN(n4471) );
  AOI22_X1 U3799 ( .A1(n3412), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3262) );
  AND2_X2 U3800 ( .A1(n5443), .A2(n3179), .ZN(n3371) );
  AOI21_X1 U3801 ( .B1(n4597), .B2(n4633), .A(n6592), .ZN(n4647) );
  INV_X1 U3802 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4790) );
  INV_X1 U3803 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5075) );
  OR2_X1 U3804 ( .A1(n6600), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4278) );
  AND2_X1 U3805 ( .A1(n3946), .A2(n3945), .ZN(n4414) );
  INV_X1 U3806 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5847) );
  INV_X1 U3807 ( .A(n6063), .ZN(n6004) );
  NOR2_X1 U3808 ( .A1(n6096), .A2(n3970), .ZN(n6044) );
  AND3_X1 U3809 ( .A1(n4028), .A2(n4059), .A3(n4027), .ZN(n5342) );
  OR2_X1 U3810 ( .A1(n5489), .A2(n5479), .ZN(n5480) );
  NOR2_X1 U3811 ( .A1(n4566), .A2(n4439), .ZN(n6135) );
  NAND2_X1 U3812 ( .A1(n4539), .A2(n4495), .ZN(n4532) );
  AND2_X1 U3813 ( .A1(n3950), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4200)
         );
  OR2_X1 U3814 ( .A1(n3833), .A2(n5788), .ZN(n3875) );
  OR2_X1 U3815 ( .A1(n3847), .A2(n5577), .ZN(n3833) );
  AND2_X1 U3816 ( .A1(n3845), .A2(n3844), .ZN(n5491) );
  OR2_X1 U3817 ( .A1(n4315), .A2(n4314), .ZN(n5490) );
  NOR2_X1 U3818 ( .A1(n3731), .A2(n5847), .ZN(n3732) );
  NAND2_X1 U3819 ( .A1(n3732), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3856)
         );
  CLKBUF_X1 U3820 ( .A(n5515), .Z(n5519) );
  OAI21_X1 U3821 ( .B1(n4273), .B2(n5958), .A(n3717), .ZN(n5534) );
  NAND2_X1 U3822 ( .A1(n3690), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3691)
         );
  NOR2_X1 U3823 ( .A1(n6904), .A2(n3691), .ZN(n3704) );
  NAND2_X1 U3824 ( .A1(n5367), .A2(n5368), .ZN(n5533) );
  NOR2_X1 U3825 ( .A1(n3685), .A2(n5988), .ZN(n3690) );
  NOR2_X2 U3826 ( .A1(n5361), .A2(n5362), .ZN(n5367) );
  CLKBUF_X1 U3827 ( .A(n5334), .Z(n5339) );
  OR2_X1 U3828 ( .A1(n3630), .A2(n6025), .ZN(n3631) );
  NOR2_X1 U3829 ( .A1(n6842), .A2(n3631), .ZN(n3657) );
  INV_X1 U3830 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6842) );
  INV_X1 U3831 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6025) );
  AND2_X1 U3832 ( .A1(n3602), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3605)
         );
  INV_X1 U3833 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6684) );
  NOR2_X1 U3834 ( .A1(n6684), .A2(n3575), .ZN(n3602) );
  NAND2_X1 U3835 ( .A1(n3562), .A2(n3561), .ZN(n4964) );
  AND2_X1 U3836 ( .A1(n3560), .A2(n3559), .ZN(n3561) );
  INV_X1 U3837 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3556) );
  AOI21_X1 U3838 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n4197), .A(n3486), 
        .ZN(n4618) );
  NAND2_X1 U3839 ( .A1(n3547), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3557)
         );
  INV_X1 U3840 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3539) );
  NOR2_X1 U3841 ( .A1(n3540), .A2(n3539), .ZN(n3547) );
  INV_X1 U3842 ( .A(n3516), .ZN(n3529) );
  NAND2_X1 U3843 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3529), .ZN(n3540)
         );
  NAND2_X1 U3844 ( .A1(n3526), .A2(n3525), .ZN(n4605) );
  NAND2_X1 U3845 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3516) );
  NAND2_X1 U3846 ( .A1(n4069), .A2(n5460), .ZN(n5456) );
  NAND2_X1 U3847 ( .A1(n4074), .A2(n4075), .ZN(n5472) );
  AND2_X1 U3848 ( .A1(n4066), .A2(n4065), .ZN(n5483) );
  NOR2_X2 U3849 ( .A1(n5484), .A2(n5483), .ZN(n5482) );
  AND2_X1 U3850 ( .A1(n5508), .A2(n4057), .ZN(n5502) );
  NAND2_X1 U3851 ( .A1(n5502), .A2(n5432), .ZN(n5434) );
  INV_X1 U3852 ( .A(n3987), .ZN(n5511) );
  AND2_X1 U3853 ( .A1(n4040), .A2(n4039), .ZN(n5524) );
  OR2_X1 U3854 ( .A1(n5402), .A2(n4173), .ZN(n5597) );
  AND2_X1 U3855 ( .A1(n4032), .A2(n4031), .ZN(n5347) );
  XNOR2_X1 U3856 ( .A(n4164), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5893)
         );
  NAND2_X1 U3857 ( .A1(n5300), .A2(n5299), .ZN(n5307) );
  AND2_X1 U3858 ( .A1(n6207), .A2(n4161), .ZN(n4162) );
  OR2_X1 U3859 ( .A1(n4164), .A2(n6293), .ZN(n4161) );
  INV_X1 U3860 ( .A(n5690), .ZN(n5321) );
  AND3_X1 U3861 ( .A1(n4015), .A2(n4059), .A3(n4014), .ZN(n5230) );
  AND2_X1 U3862 ( .A1(n4006), .A2(n4005), .ZN(n4620) );
  INV_X1 U3863 ( .A(n4557), .ZN(n3992) );
  INV_X1 U3864 ( .A(n4558), .ZN(n3993) );
  AND2_X1 U3865 ( .A1(n4378), .A2(n5724), .ZN(n5688) );
  AND2_X1 U3866 ( .A1(n5910), .A2(n4376), .ZN(n5690) );
  CLKBUF_X1 U3867 ( .A(n4082), .Z(n4795) );
  OR2_X1 U3868 ( .A1(n4110), .A2(n5730), .ZN(n5039) );
  AND2_X1 U3869 ( .A1(n3678), .A2(n3680), .ZN(n6473) );
  NOR2_X1 U3870 ( .A1(n3939), .A2(n4361), .ZN(n4346) );
  AOI211_X1 U3871 ( .C1(n4503), .C2(n4502), .A(n4501), .B(n4500), .ZN(n6479)
         );
  OR2_X1 U3872 ( .A1(n4641), .A2(n5073), .ZN(n4646) );
  NOR2_X1 U3873 ( .A1(n5039), .A2(n4795), .ZN(n4846) );
  AND2_X1 U3874 ( .A1(n5076), .A2(n6368), .ZN(n5040) );
  NOR2_X1 U3875 ( .A1(n5073), .A2(n4110), .ZN(n4927) );
  INV_X1 U3876 ( .A(n4649), .ZN(n4899) );
  INV_X1 U3877 ( .A(n4698), .ZN(n4762) );
  INV_X1 U3878 ( .A(n4090), .ZN(n4845) );
  INV_X1 U3879 ( .A(n4766), .ZN(n4830) );
  NOR2_X1 U3880 ( .A1(n6590), .A2(n4647), .ZN(n4829) );
  NOR2_X1 U3881 ( .A1(n4666), .A2(n4845), .ZN(n4763) );
  INV_X2 U3882 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6497) );
  AND2_X1 U3883 ( .A1(n6501), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3937) );
  NAND2_X1 U3884 ( .A1(n5773), .A2(n3975), .ZN(n4079) );
  INV_X1 U3885 ( .A(n5781), .ZN(n5800) );
  NOR2_X1 U3886 ( .A1(n5843), .A2(n3966), .ZN(n5842) );
  INV_X1 U3887 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6904) );
  INV_X1 U3888 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5988) );
  AND2_X1 U3889 ( .A1(n4535), .A2(n4078), .ZN(n6087) );
  AND2_X1 U3890 ( .A1(n6044), .A2(REIP_REG_9__SCAN_IN), .ZN(n6032) );
  AND2_X1 U3891 ( .A1(n5262), .A2(n3952), .ZN(n6070) );
  AND2_X1 U3892 ( .A1(n4285), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3952) );
  INV_X1 U3893 ( .A(n5262), .ZN(n6109) );
  INV_X1 U3894 ( .A(n6087), .ZN(n6123) );
  INV_X1 U3895 ( .A(n6099), .ZN(n6110) );
  AND2_X1 U3896 ( .A1(n5262), .A2(n3959), .ZN(n6120) );
  NAND2_X1 U3897 ( .A1(n4434), .A2(n4569), .ZN(n5492) );
  NAND2_X1 U3898 ( .A1(n4491), .A2(n4433), .ZN(n4434) );
  AND2_X1 U3899 ( .A1(n5373), .A2(n5372), .ZN(n6946) );
  NOR2_X1 U3900 ( .A1(n4576), .A2(n4575), .ZN(n5340) );
  OR2_X1 U3901 ( .A1(n5373), .A2(n4573), .ZN(n5539) );
  INV_X1 U3902 ( .A(n5340), .ZN(n5246) );
  INV_X1 U3904 ( .A(n6194), .ZN(n6203) );
  NAND2_X1 U3905 ( .A1(n5395), .A2(n3886), .ZN(n3887) );
  NAND2_X1 U3906 ( .A1(n5396), .A2(n5395), .ZN(n5571) );
  OR2_X1 U3907 ( .A1(n5394), .A2(n5393), .ZN(n5396) );
  AND2_X1 U3908 ( .A1(n5439), .A2(n4393), .ZN(n5656) );
  AND2_X1 U3909 ( .A1(n5436), .A2(n4387), .ZN(n5655) );
  CLKBUF_X1 U3910 ( .A(n5884), .Z(n5889) );
  NOR2_X1 U3911 ( .A1(n5912), .A2(n5322), .ZN(n6288) );
  INV_X1 U3912 ( .A(n5317), .ZN(n6353) );
  OR2_X1 U3913 ( .A1(n4377), .A2(n5445), .ZN(n5910) );
  CLKBUF_X1 U3914 ( .A(n3506), .Z(n3507) );
  CLKBUF_X1 U3915 ( .A(n4626), .Z(n5730) );
  CLKBUF_X1 U3916 ( .A(n4511), .Z(n4512) );
  NOR2_X1 U3917 ( .A1(n4794), .A2(n5939), .ZN(n5731) );
  INV_X1 U3918 ( .A(n6371), .ZN(n5733) );
  OAI221_X1 U3919 ( .B1(n5082), .B2(n3296), .C1(n5082), .C2(n5081), .A(n5080), 
        .ZN(n5122) );
  INV_X1 U3920 ( .A(n6370), .ZN(n6413) );
  OR3_X1 U3921 ( .A1(n6378), .A2(n6377), .A3(n6376), .ZN(n6415) );
  NAND2_X1 U3922 ( .A1(n4971), .A2(n4845), .ZN(n6419) );
  NAND2_X1 U3923 ( .A1(n4846), .A2(n4845), .ZN(n4958) );
  NOR2_X1 U3924 ( .A1(n6177), .A2(n4830), .ZN(n6440) );
  INV_X1 U3925 ( .A(n5096), .ZN(n6384) );
  NOR2_X1 U3926 ( .A1(n6179), .A2(n4830), .ZN(n6383) );
  INV_X1 U3927 ( .A(n5091), .ZN(n6445) );
  NOR2_X1 U3928 ( .A1(n6181), .A2(n4830), .ZN(n6446) );
  INV_X1 U3929 ( .A(n5113), .ZN(n6451) );
  NOR2_X1 U3930 ( .A1(n6183), .A2(n4830), .ZN(n6452) );
  INV_X1 U3931 ( .A(n5118), .ZN(n6457) );
  NOR2_X1 U3932 ( .A1(n6186), .A2(n4830), .ZN(n6458) );
  NOR2_X1 U3933 ( .A1(n6188), .A2(n4830), .ZN(n6467) );
  INV_X1 U3934 ( .A(n5101), .ZN(n6406) );
  NOR2_X1 U3935 ( .A1(n6815), .A2(n4830), .ZN(n6405) );
  INV_X1 U3936 ( .A(n5108), .ZN(n6428) );
  NOR2_X1 U3937 ( .A1(n6191), .A2(n4830), .ZN(n6432) );
  INV_X1 U3938 ( .A(n6383), .ZN(n5095) );
  INV_X1 U3939 ( .A(n6446), .ZN(n5090) );
  INV_X1 U3940 ( .A(n6452), .ZN(n5112) );
  INV_X1 U3941 ( .A(n6458), .ZN(n5117) );
  INV_X1 U3942 ( .A(n6467), .ZN(n5123) );
  INV_X1 U3943 ( .A(n6405), .ZN(n5100) );
  INV_X1 U3944 ( .A(n6432), .ZN(n5107) );
  NOR2_X1 U3945 ( .A1(n4666), .A2(n3142), .ZN(n5029) );
  NAND2_X1 U3946 ( .A1(n3937), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6510) );
  AND2_X1 U3947 ( .A1(n4287), .A2(n4286), .ZN(n4288) );
  OR2_X1 U3948 ( .A1(n5748), .A2(n6286), .ZN(n4409) );
  AND2_X1 U3949 ( .A1(n4320), .A2(n4319), .ZN(n4321) );
  INV_X1 U3950 ( .A(n4401), .ZN(n4402) );
  NAND2_X1 U3951 ( .A1(n4407), .A2(n6356), .ZN(n4403) );
  OAI21_X1 U3952 ( .B1(n5749), .B2(n6351), .A(n4400), .ZN(n4401) );
  NAND2_X4 U3953 ( .A1(n4152), .A2(n4151), .ZN(n4164) );
  AND4_X1 U3954 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3160)
         );
  XNOR2_X1 U3955 ( .A(n5382), .B(n4408), .ZN(n5748) );
  INV_X1 U3956 ( .A(n3508), .ZN(n4238) );
  OAI21_X1 U3957 ( .B1(n6206), .B2(n4163), .A(n4162), .ZN(n5312) );
  XOR2_X1 U3958 ( .A(n4164), .B(n5645), .Z(n3161) );
  INV_X1 U3959 ( .A(n3939), .ZN(n4415) );
  AND2_X1 U3960 ( .A1(n6497), .A2(n5939), .ZN(n4243) );
  INV_X1 U3961 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5993) );
  AND2_X1 U3962 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3162) );
  AND3_X1 U3963 ( .A1(n4177), .A2(n4176), .A3(n4175), .ZN(n3163) );
  AND4_X1 U3964 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3164)
         );
  OR2_X1 U3965 ( .A1(n5635), .A2(n6123), .ZN(n3165) );
  AND4_X1 U3966 ( .A1(n3203), .A2(n3202), .A3(n3201), .A4(n3200), .ZN(n3166)
         );
  OR2_X1 U3967 ( .A1(n4173), .A2(n4172), .ZN(n5599) );
  AND4_X1 U3968 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3167)
         );
  OR2_X1 U3969 ( .A1(n3327), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3168)
         );
  NAND2_X1 U3970 ( .A1(n4277), .A2(n6371), .ZN(n6286) );
  AND4_X1 U3971 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3169)
         );
  INV_X1 U3972 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4310) );
  AND2_X2 U3973 ( .A1(n4589), .A2(n3179), .ZN(n3258) );
  INV_X1 U3974 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n3296) );
  AND2_X1 U3975 ( .A1(n4092), .A2(n4093), .ZN(n4525) );
  INV_X1 U3976 ( .A(n3502), .ZN(n3386) );
  INV_X1 U3977 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n3350) );
  INV_X1 U3978 ( .A(n4164), .ZN(n4187) );
  OR2_X1 U3979 ( .A1(n3678), .A2(n4570), .ZN(n3307) );
  AND2_X1 U3980 ( .A1(n5179), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3902)
         );
  OR2_X1 U3981 ( .A1(n5597), .A2(n4169), .ZN(n4170) );
  OR2_X1 U3982 ( .A1(n3451), .A2(n3450), .ZN(n4122) );
  INV_X1 U3983 ( .A(n4096), .ZN(n3388) );
  INV_X1 U3984 ( .A(n4097), .ZN(n4105) );
  AND2_X1 U3985 ( .A1(n3270), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U3986 ( .A1(n3412), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3193) );
  OR2_X1 U3987 ( .A1(n3364), .A2(n3363), .ZN(n4154) );
  NAND2_X1 U3988 ( .A1(n4362), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3429) );
  AOI21_X1 U3989 ( .B1(n3258), .B2(INSTQUEUE_REG_4__2__SCAN_IN), .A(n3271), 
        .ZN(n3275) );
  BUF_X1 U3990 ( .A(n3288), .Z(n4333) );
  NAND2_X1 U3991 ( .A1(n3454), .A2(n3535), .ZN(n3546) );
  OR2_X1 U3992 ( .A1(n4164), .A2(n4183), .ZN(n4184) );
  NOR2_X1 U3993 ( .A1(n3546), .A2(n3468), .ZN(n3553) );
  OR2_X1 U3994 ( .A1(n3378), .A2(n3377), .ZN(n4095) );
  AND4_X1 U3995 ( .A1(n3199), .A2(n3198), .A3(n3197), .A4(n3196), .ZN(n3204)
         );
  NAND2_X1 U3996 ( .A1(n5511), .A2(n3984), .ZN(n3986) );
  NOR2_X1 U3997 ( .A1(n3316), .A2(n4333), .ZN(n3317) );
  NOR2_X1 U3998 ( .A1(n4648), .A2(n6497), .ZN(n3508) );
  NAND2_X1 U3999 ( .A1(n3553), .A2(n3552), .ZN(n4152) );
  OR2_X1 U4000 ( .A1(n3343), .A2(n3342), .ZN(n4096) );
  INV_X1 U4001 ( .A(n3348), .ZN(n3394) );
  AND2_X2 U4002 ( .A1(n4483), .A2(n4478), .ZN(n3372) );
  OR2_X1 U4003 ( .A1(n3986), .A2(EBX_REG_1__SCAN_IN), .ZN(n3981) );
  AND2_X1 U4004 ( .A1(n4019), .A2(n4018), .ZN(n5238) );
  NOR2_X1 U4006 ( .A1(n3856), .A2(n3760), .ZN(n3858) );
  AND2_X1 U4007 ( .A1(n6473), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4240) );
  OR2_X1 U4008 ( .A1(n4140), .A2(n3555), .ZN(n3562) );
  NOR2_X1 U4009 ( .A1(n5565), .A2(n4189), .ZN(n4323) );
  CLKBUF_X2 U4010 ( .A(n3268), .Z(n4570) );
  NAND2_X1 U4011 ( .A1(n4127), .A2(n4126), .ZN(n4128) );
  NOR2_X1 U4012 ( .A1(n4473), .A2(n4480), .ZN(n4375) );
  AND2_X2 U4013 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4478) );
  AND2_X1 U4014 ( .A1(n4850), .A2(n6371), .ZN(n4852) );
  AND2_X1 U4015 ( .A1(n3441), .A2(n3440), .ZN(n4627) );
  NAND2_X1 U4016 ( .A1(n3428), .A2(n3427), .ZN(n4967) );
  INV_X1 U4017 ( .A(n3267), .ZN(n4684) );
  AND2_X1 U4018 ( .A1(n4200), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4223)
         );
  NAND2_X1 U4019 ( .A1(n3858), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3847)
         );
  OR2_X1 U4020 ( .A1(n3660), .A2(n5993), .ZN(n3685) );
  NAND2_X1 U4021 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n3657), .ZN(n3660)
         );
  BUF_X2 U4022 ( .A(n3984), .Z(n4535) );
  INV_X1 U4023 ( .A(n6112), .ZN(n6073) );
  CLKBUF_X1 U4024 ( .A(n5229), .Z(n5239) );
  INV_X1 U4025 ( .A(n6510), .ZN(n4569) );
  AND2_X1 U4026 ( .A1(n5496), .A2(n4222), .ZN(n4298) );
  NOR2_X1 U4027 ( .A1(n3678), .A2(n5540), .ZN(n4574) );
  NOR2_X1 U4028 ( .A1(n3875), .A2(n5570), .ZN(n3950) );
  AND2_X1 U4029 ( .A1(n5497), .A2(n5478), .ZN(n5489) );
  NOR2_X2 U4030 ( .A1(n5533), .A2(n5534), .ZN(n5518) );
  NAND2_X1 U4031 ( .A1(n3605), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3630)
         );
  OR2_X1 U4032 ( .A1(n6272), .A2(n4279), .ZN(n5588) );
  INV_X1 U4033 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U4034 ( .A1(n5590), .A2(n5582), .ZN(n5423) );
  AND2_X1 U4035 ( .A1(n4164), .A2(n5419), .ZN(n5420) );
  OR2_X1 U4036 ( .A1(n5598), .A2(n5402), .ZN(n5404) );
  AOI21_X1 U4037 ( .B1(n4626), .B2(n4336), .A(n4100), .ZN(n6271) );
  CLKBUF_X1 U4038 ( .A(n4478), .Z(n4508) );
  AND2_X1 U4039 ( .A1(n5077), .A2(n5076), .ZN(n5135) );
  OR2_X1 U4040 ( .A1(n5188), .A2(n3142), .ZN(n6370) );
  INV_X1 U4041 ( .A(n4795), .ZN(n4794) );
  AOI21_X1 U4042 ( .B1(n5179), .B2(STATE2_REG_3__SCAN_IN), .A(n4830), .ZN(
        n4973) );
  INV_X1 U4043 ( .A(n4243), .ZN(n4273) );
  NAND2_X1 U4044 ( .A1(n4411), .A2(n4569), .ZN(n4425) );
  NAND2_X1 U4045 ( .A1(n4223), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4245)
         );
  OR2_X1 U4046 ( .A1(n5998), .A2(n3963), .ZN(n5843) );
  AND2_X1 U4047 ( .A1(n6032), .A2(n3971), .ZN(n6018) );
  INV_X1 U4048 ( .A(n6066), .ZN(n6083) );
  NAND2_X1 U4049 ( .A1(n5737), .A2(n3958), .ZN(n6112) );
  NAND2_X1 U4050 ( .A1(n5262), .A2(n6096), .ZN(n6063) );
  NAND2_X1 U4051 ( .A1(n5364), .A2(n5363), .ZN(n5369) );
  AND2_X1 U4052 ( .A1(n5496), .A2(n4296), .ZN(n5381) );
  OAI21_X1 U4053 ( .B1(n4534), .B2(n6613), .A(n4533), .ZN(n6184) );
  INV_X1 U4054 ( .A(n4566), .ZN(n4539) );
  INV_X1 U4055 ( .A(n6166), .ZN(n6201) );
  OR2_X1 U4056 ( .A1(n5807), .A2(n6286), .ZN(n4320) );
  NAND2_X1 U4057 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n3558), .ZN(n3575)
         );
  AND3_X1 U4058 ( .A1(n4605), .A2(n4604), .A3(n4577), .ZN(n4613) );
  AND2_X1 U4059 ( .A1(n5656), .A2(n4395), .ZN(n5631) );
  NOR2_X1 U4060 ( .A1(n5664), .A2(n5675), .ZN(n5439) );
  NOR2_X1 U4061 ( .A1(n6288), .A2(n5407), .ZN(n5905) );
  NOR2_X1 U4062 ( .A1(n6319), .A2(n5320), .ZN(n5322) );
  INV_X1 U4063 ( .A(n6351), .ZN(n6323) );
  INV_X1 U4064 ( .A(n5913), .ZN(n6356) );
  NOR2_X1 U4065 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4647), .ZN(n4766) );
  NOR2_X1 U4066 ( .A1(n3296), .A2(n4489), .ZN(n6592) );
  INV_X1 U4067 ( .A(n4895), .ZN(n5009) );
  INV_X1 U4068 ( .A(n5106), .ZN(n5128) );
  INV_X1 U4069 ( .A(n4646), .ZN(n5169) );
  INV_X1 U4070 ( .A(n4973), .ZN(n5183) );
  AND2_X1 U4071 ( .A1(n4642), .A2(n6371), .ZN(n5184) );
  NOR3_X1 U4072 ( .A1(n5131), .A2(n4794), .A3(n4793), .ZN(n4971) );
  INV_X1 U4073 ( .A(n4889), .ZN(n4835) );
  INV_X1 U4074 ( .A(n4958), .ZN(n4886) );
  INV_X1 U4075 ( .A(n6471), .ZN(n4960) );
  INV_X1 U4076 ( .A(n5046), .ZN(n6463) );
  OR2_X1 U4077 ( .A1(n4703), .A2(n4702), .ZN(n5016) );
  INV_X1 U4078 ( .A(n5086), .ZN(n6439) );
  INV_X1 U4079 ( .A(n5126), .ZN(n6465) );
  INV_X1 U4080 ( .A(n4926), .ZN(n4990) );
  OAI211_X1 U4081 ( .C1(n3296), .C2(n4770), .A(n4769), .B(n4768), .ZN(n4986)
         );
  INV_X1 U4082 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6501) );
  INV_X1 U4083 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6529) );
  INV_X1 U4084 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5939) );
  NAND2_X1 U4085 ( .A1(n4079), .A2(n3165), .ZN(n4080) );
  NAND2_X1 U4086 ( .A1(n5262), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U4087 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6018), .ZN(n6014) );
  NAND2_X1 U4088 ( .A1(n3888), .A2(n3887), .ZN(n5558) );
  OR2_X1 U4089 ( .A1(n6135), .A2(n6614), .ZN(n6134) );
  INV_X1 U4090 ( .A(n6135), .ZN(n6164) );
  NAND2_X1 U4091 ( .A1(n4539), .A2(n4538), .ZN(n6194) );
  OR2_X1 U4092 ( .A1(n4532), .A2(n4361), .ZN(n6166) );
  AOI211_X1 U4093 ( .C1(n6257), .C2(n5778), .A(n5573), .B(n5572), .ZN(n5574)
         );
  INV_X1 U4094 ( .A(n6272), .ZN(n6278) );
  INV_X1 U4095 ( .A(n6257), .ZN(n6280) );
  OR2_X1 U4096 ( .A1(n4377), .A2(n4360), .ZN(n6351) );
  INV_X1 U4097 ( .A(n4283), .ZN(n6349) );
  OR2_X1 U4098 ( .A1(n4377), .A2(n4350), .ZN(n5913) );
  INV_X1 U4099 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5179) );
  INV_X1 U4100 ( .A(n5029), .ZN(n5012) );
  NAND2_X1 U4101 ( .A1(n4734), .A2(n3142), .ZN(n4895) );
  OR2_X1 U4102 ( .A1(n4856), .A2(n4090), .ZN(n5106) );
  OR2_X1 U4103 ( .A1(n5074), .A2(n5073), .ZN(n5172) );
  NAND2_X1 U4104 ( .A1(n4639), .A2(n3142), .ZN(n5222) );
  NAND2_X1 U4105 ( .A1(n4971), .A2(n3142), .ZN(n6436) );
  NOR2_X1 U4106 ( .A1(n4799), .A2(n4798), .ZN(n4837) );
  NAND2_X1 U4107 ( .A1(n4846), .A2(n3142), .ZN(n4889) );
  INV_X1 U4108 ( .A(n6440), .ZN(n5085) );
  AOI21_X1 U4109 ( .B1(n4932), .B2(n5040), .A(n4929), .ZN(n4963) );
  NAND2_X1 U4110 ( .A1(n4927), .A2(n3142), .ZN(n6471) );
  NAND2_X1 U4111 ( .A1(n4927), .A2(n4845), .ZN(n5046) );
  NAND2_X1 U4112 ( .A1(n4762), .A2(n4845), .ZN(n4926) );
  INV_X1 U4113 ( .A(n4763), .ZN(n5033) );
  INV_X1 U4114 ( .A(n6588), .ZN(n6518) );
  INV_X1 U4115 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6525) );
  INV_X1 U4116 ( .A(n6579), .ZN(n6577) );
  OR2_X1 U4117 ( .A1(n4081), .A2(n4080), .ZN(U2800) );
  NOR2_X2 U4118 ( .A1(n5939), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4197) );
  INV_X1 U4119 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3170) );
  NOR2_X4 U4120 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4589) );
  AND2_X2 U4121 ( .A1(n3141), .A2(n4589), .ZN(n3335) );
  INV_X1 U4122 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3171) );
  AND2_X4 U4123 ( .A1(n3171), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5443)
         );
  INV_X1 U4124 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3172) );
  AND2_X2 U4125 ( .A1(n3172), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3179)
         );
  AOI22_X1 U4126 ( .A1(n3335), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3176) );
  AND2_X4 U4127 ( .A1(n3179), .A2(n4478), .ZN(n3805) );
  AOI22_X1 U4128 ( .A1(n3805), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3175) );
  NOR2_X4 U4129 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4484) );
  AND2_X2 U4130 ( .A1(n4589), .A2(n4484), .ZN(n3336) );
  AND2_X2 U4131 ( .A1(n4484), .A2(n4478), .ZN(n3270) );
  AOI22_X1 U4132 ( .A1(n3336), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3174) );
  AND2_X4 U4133 ( .A1(n3178), .A2(n4478), .ZN(n3746) );
  AOI22_X1 U4134 ( .A1(n3746), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3173) );
  AND2_X4 U4135 ( .A1(n3177), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5450)
         );
  AND2_X2 U4136 ( .A1(n5450), .A2(n4484), .ZN(n3406) );
  AND2_X4 U4137 ( .A1(n5443), .A2(n4483), .ZN(n3722) );
  AOI22_X1 U4138 ( .A1(n3406), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3183) );
  AND2_X2 U4139 ( .A1(n3178), .A2(n5443), .ZN(n3276) );
  AND2_X4 U4140 ( .A1(n5450), .A2(n4483), .ZN(n3412) );
  AOI22_X1 U4141 ( .A1(n3412), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3181) );
  AND2_X4 U4142 ( .A1(n5450), .A2(n3179), .ZN(n3370) );
  AND2_X2 U4143 ( .A1(n4589), .A2(n4483), .ZN(n3337) );
  AOI22_X1 U4144 ( .A1(n3370), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3337), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3180) );
  NAND4_X1 U4145 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3184)
         );
  INV_X1 U4146 ( .A(n3184), .ZN(n3185) );
  AND2_X2 U4147 ( .A1(n3167), .A2(n3185), .ZN(n3267) );
  AOI22_X1 U4148 ( .A1(n3746), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3189) );
  AOI22_X1 U4149 ( .A1(n3153), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4150 ( .A1(n3805), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4151 ( .A1(n3335), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U4152 ( .A1(n3371), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U4153 ( .A1(n3258), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3190) );
  NAND2_X2 U4154 ( .A1(n3267), .A2(n3285), .ZN(n3284) );
  AOI22_X1 U4155 ( .A1(n3407), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4156 ( .A1(n3805), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U4157 ( .A1(n3406), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4158 ( .A1(n3276), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3746), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4159 ( .A1(n3335), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3337), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3202) );
  AOI22_X1 U4160 ( .A1(n3371), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4161 ( .A1(n3258), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4162 ( .A1(n3406), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3208) );
  AOI22_X1 U4163 ( .A1(n3276), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3746), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3207) );
  AOI22_X1 U4164 ( .A1(n3154), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4165 ( .A1(n3805), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3205) );
  NAND4_X1 U4166 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n3214)
         );
  AOI22_X1 U4167 ( .A1(n3412), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4168 ( .A1(n3335), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4169 ( .A1(n3371), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4170 ( .A1(n3258), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3209) );
  NAND4_X1 U4171 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3213)
         );
  NAND2_X1 U4172 ( .A1(n3335), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4173 ( .A1(n3412), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3217)
         );
  NAND2_X1 U4174 ( .A1(n3370), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3216) );
  NAND2_X1 U4175 ( .A1(n3337), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3215)
         );
  NAND2_X1 U4176 ( .A1(n3406), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4177 ( .A1(n3407), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4178 ( .A1(n3722), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3220)
         );
  NAND2_X1 U4179 ( .A1(n3369), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4180 ( .A1(n3276), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3225)
         );
  NAND2_X1 U4181 ( .A1(n3805), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4182 ( .A1(n3372), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3223)
         );
  NAND2_X1 U4183 ( .A1(n3270), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U4184 ( .A1(n3336), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4185 ( .A1(n3371), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U4186 ( .A1(n3258), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3227) );
  INV_X2 U4187 ( .A(n3300), .ZN(n3892) );
  NAND2_X1 U4188 ( .A1(n3412), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3237)
         );
  NAND2_X1 U4189 ( .A1(n3370), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3236) );
  NAND2_X1 U4190 ( .A1(n3258), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U4191 ( .A1(n3336), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4192 ( .A1(n3746), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3241)
         );
  NAND2_X1 U4193 ( .A1(n3406), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4194 ( .A1(n3276), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3239)
         );
  NAND2_X1 U4195 ( .A1(n3805), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U4197 ( .A1(n3407), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3245) );
  NAND2_X1 U4198 ( .A1(n3369), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3244) );
  NAND2_X1 U4199 ( .A1(n3157), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3243)
         );
  NAND2_X1 U4200 ( .A1(n3372), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3242)
         );
  NAND2_X1 U4201 ( .A1(n3335), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3249) );
  NAND2_X1 U4202 ( .A1(n3371), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3248) );
  NAND2_X1 U4203 ( .A1(n3337), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3247)
         );
  NAND2_X1 U4204 ( .A1(n3270), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U4206 ( .A1(n4570), .A2(n4684), .ZN(n3322) );
  AOI22_X1 U4207 ( .A1(n3276), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3746), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4208 ( .A1(n3406), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4209 ( .A1(n3154), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4210 ( .A1(n3805), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3254) );
  NAND4_X1 U4211 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3264)
         );
  AOI22_X1 U4212 ( .A1(n3335), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4213 ( .A1(n3371), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4214 ( .A1(n3258), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3259) );
  NAND4_X1 U4215 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), .ZN(n3263)
         );
  OR2_X2 U4216 ( .A1(n3264), .A2(n3263), .ZN(n4676) );
  NAND2_X2 U4217 ( .A1(n4676), .A2(n3300), .ZN(n3987) );
  OR2_X2 U4218 ( .A1(n3322), .A2(n3987), .ZN(n3265) );
  NAND2_X1 U4219 ( .A1(n3266), .A2(n3265), .ZN(n3309) );
  NOR2_X2 U4220 ( .A1(n3267), .A2(n3285), .ZN(n3287) );
  NAND2_X1 U4221 ( .A1(n3287), .A2(n3268), .ZN(n3269) );
  BUF_X2 U4222 ( .A(n3287), .Z(n3678) );
  AOI22_X1 U4223 ( .A1(n3412), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4224 ( .A1(n3407), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4225 ( .A1(n3746), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4226 ( .A1(n3276), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4227 ( .A1(n3722), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4228 ( .A1(n3370), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4229 ( .A1(n3335), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3337), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3277) );
  AND2_X2 U4230 ( .A1(n3281), .A2(n3169), .ZN(n3319) );
  XNOR2_X1 U4231 ( .A(n6525), .B(STATE_REG_2__SCAN_IN), .ZN(n3953) );
  NOR2_X1 U4232 ( .A1(n3300), .A2(n3953), .ZN(n3321) );
  NAND4_X1 U4233 ( .A1(n4370), .A2(n3307), .A3(n4365), .A4(n3282), .ZN(n3283)
         );
  OAI21_X1 U4234 ( .B1(n3309), .B2(n3283), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3295) );
  INV_X2 U4236 ( .A(n3319), .ZN(n4680) );
  NAND2_X1 U4237 ( .A1(n3288), .A2(n4680), .ZN(n3289) );
  AND2_X2 U4238 ( .A1(n3291), .A2(n3290), .ZN(n3324) );
  NAND2_X1 U4239 ( .A1(n3324), .A2(n3892), .ZN(n3293) );
  INV_X1 U4240 ( .A(n3429), .ZN(n3419) );
  NAND2_X1 U4241 ( .A1(n3293), .A2(n3419), .ZN(n3294) );
  NAND2_X1 U4242 ( .A1(n3295), .A2(n3294), .ZN(n3397) );
  NAND2_X1 U4243 ( .A1(n3397), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3299) );
  INV_X1 U4244 ( .A(n3937), .ZN(n3402) );
  NAND2_X1 U4245 ( .A1(n6501), .A2(n3296), .ZN(n6600) );
  INV_X1 U4246 ( .A(n4278), .ZN(n3403) );
  MUX2_X1 U4247 ( .A(n3402), .B(n3403), .S(n5179), .Z(n3297) );
  INV_X1 U4248 ( .A(n3297), .ZN(n3298) );
  NAND2_X1 U4249 ( .A1(n3299), .A2(n3298), .ZN(n3347) );
  INV_X1 U4250 ( .A(n5247), .ZN(n3302) );
  INV_X1 U4251 ( .A(n3322), .ZN(n4196) );
  NAND2_X1 U4252 ( .A1(n4362), .A2(n4361), .ZN(n5251) );
  OAI22_X1 U4253 ( .A1(n3324), .A2(n3302), .B1(n4196), .B2(n5251), .ZN(n4372)
         );
  INV_X1 U4254 ( .A(n4372), .ZN(n3315) );
  NOR2_X1 U4255 ( .A1(n4676), .A2(n4680), .ZN(n4431) );
  OR2_X1 U4256 ( .A1(n6600), .A2(n3350), .ZN(n6511) );
  AOI21_X1 U4257 ( .B1(n4680), .B2(n4672), .A(n6511), .ZN(n3306) );
  NAND3_X1 U4258 ( .A1(n4370), .A2(n4676), .A3(n3307), .ZN(n3308) );
  NAND2_X1 U4259 ( .A1(n3308), .A2(n4361), .ZN(n3313) );
  INV_X1 U4260 ( .A(n3309), .ZN(n3312) );
  NAND2_X1 U4261 ( .A1(n3310), .A2(n4534), .ZN(n3311) );
  NAND2_X1 U4262 ( .A1(n3315), .A2(n3164), .ZN(n3346) );
  NAND2_X1 U4263 ( .A1(n3347), .A2(n3346), .ZN(n3348) );
  NAND2_X1 U4264 ( .A1(n4365), .A2(n4335), .ZN(n3316) );
  NAND2_X1 U4265 ( .A1(n3317), .A2(n4574), .ZN(n4329) );
  INV_X1 U4266 ( .A(n4329), .ZN(n3318) );
  NAND2_X1 U4267 ( .A1(n3318), .A2(n3301), .ZN(n3938) );
  INV_X1 U4268 ( .A(n4684), .ZN(n5372) );
  NAND4_X1 U4269 ( .A1(n3319), .A2(n5372), .A3(n5247), .A4(n3976), .ZN(n4572)
         );
  AND2_X1 U4270 ( .A1(n4648), .A2(n3303), .ZN(n5374) );
  INV_X1 U4271 ( .A(n5374), .ZN(n3320) );
  OAI21_X1 U4272 ( .B1(n3938), .B2(n3321), .A(n4357), .ZN(n3325) );
  NOR2_X1 U4273 ( .A1(n3322), .A2(n4672), .ZN(n3323) );
  INV_X2 U4274 ( .A(n3892), .ZN(n4361) );
  INV_X1 U4275 ( .A(n3329), .ZN(n3326) );
  XNOR2_X1 U4276 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5083) );
  OAI22_X1 U4277 ( .A1(n4278), .A2(n5083), .B1(n3937), .B2(n4790), .ZN(n3327)
         );
  NAND2_X1 U4278 ( .A1(n3326), .A2(n3168), .ZN(n3395) );
  AOI21_X1 U4279 ( .B1(n3397), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3327), 
        .ZN(n3328) );
  NAND2_X1 U4280 ( .A1(n3329), .A2(n3328), .ZN(n3393) );
  NAND2_X1 U4281 ( .A1(n3395), .A2(n3393), .ZN(n3330) );
  XNOR2_X1 U4282 ( .A(n3394), .B(n3330), .ZN(n4600) );
  NAND2_X1 U4283 ( .A1(n4600), .A2(n3350), .ZN(n3345) );
  AOI22_X1 U4284 ( .A1(n3352), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4285 ( .A1(n4257), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4287 ( .A1(n4202), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4288 ( .A1(n3154), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3331) );
  NAND4_X1 U4289 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3343)
         );
  AOI22_X1 U4290 ( .A1(n4246), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4291 ( .A1(n3135), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4292 ( .A1(n4248), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4293 ( .A1(n3337), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3338) );
  NAND4_X1 U4294 ( .A1(n3341), .A2(n3340), .A3(n3339), .A4(n3338), .ZN(n3342)
         );
  NAND2_X1 U4295 ( .A1(n3345), .A2(n3344), .ZN(n3491) );
  OR2_X1 U4296 ( .A1(n3347), .A2(n3346), .ZN(n3349) );
  NAND2_X1 U4297 ( .A1(n3349), .A2(n3348), .ZN(n3506) );
  INV_X1 U4298 ( .A(n3506), .ZN(n3351) );
  NAND2_X1 U4299 ( .A1(n3351), .A2(n3350), .ZN(n3500) );
  INV_X1 U4300 ( .A(n4149), .ZN(n3380) );
  AOI22_X1 U4301 ( .A1(n4246), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4302 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n3864), .B1(n3135), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4303 ( .A1(n4248), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4304 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n4202), .B1(n4249), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3353) );
  NAND4_X1 U4305 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3364)
         );
  AOI22_X1 U4306 ( .A1(n3153), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4307 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n3369), .B1(n3157), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4308 ( .A1(n3370), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3337), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4309 ( .A1(n4256), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3359) );
  NAND4_X1 U4310 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3363)
         );
  AOI22_X1 U4311 ( .A1(n4246), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4312 ( .A1(n3407), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4313 ( .A1(n3135), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4314 ( .A1(n4202), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3365) );
  NAND4_X1 U4315 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3378)
         );
  AOI22_X1 U4316 ( .A1(n4257), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4317 ( .A1(n3370), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4318 ( .A1(n4248), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4319 ( .A1(n4256), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3373) );
  NAND4_X1 U4320 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3377)
         );
  XNOR2_X1 U4321 ( .A(n3382), .B(n4095), .ZN(n3379) );
  NAND2_X1 U4322 ( .A1(n3380), .A2(n3379), .ZN(n3503) );
  AND2_X1 U4323 ( .A1(n3503), .A2(n4149), .ZN(n3387) );
  NAND2_X1 U4324 ( .A1(n3921), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3385) );
  NAND2_X1 U4325 ( .A1(n4362), .A2(n4095), .ZN(n3381) );
  OAI211_X1 U4326 ( .C1(n3382), .C2(n4688), .A(STATE2_REG_0__SCAN_IN), .B(
        n3381), .ZN(n3383) );
  INV_X1 U4327 ( .A(n3383), .ZN(n3384) );
  NAND2_X1 U4328 ( .A1(n3385), .A2(n3384), .ZN(n3502) );
  AOI21_X2 U4329 ( .B1(n3500), .B2(n3387), .A(n3386), .ZN(n3493) );
  NAND2_X1 U4330 ( .A1(n3921), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3390) );
  OR2_X1 U4331 ( .A1(n3429), .A2(n3388), .ZN(n3389) );
  OAI211_X1 U4332 ( .C1(n4149), .C2(n4154), .A(n3390), .B(n3389), .ZN(n3492)
         );
  OAI21_X1 U4333 ( .B1(n3491), .B2(n3493), .A(n3492), .ZN(n3392) );
  NAND2_X1 U4334 ( .A1(n3491), .A2(n3493), .ZN(n3391) );
  NAND2_X1 U4335 ( .A1(n3392), .A2(n3391), .ZN(n3488) );
  NAND2_X1 U4336 ( .A1(n3394), .A2(n3393), .ZN(n3396) );
  NAND2_X1 U4337 ( .A1(n3398), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3405) );
  AND2_X1 U4338 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3399) );
  NAND2_X1 U4339 ( .A1(n3399), .A2(n5075), .ZN(n5134) );
  INV_X1 U4340 ( .A(n3399), .ZN(n3400) );
  NAND2_X1 U4341 ( .A1(n3400), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3401) );
  NAND2_X1 U4342 ( .A1(n5134), .A2(n3401), .ZN(n4650) );
  AOI22_X1 U4343 ( .A1(n3403), .A2(n4650), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3402), .ZN(n3404) );
  AOI22_X1 U4344 ( .A1(n3135), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3411) );
  INV_X1 U4345 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6800) );
  AOI22_X1 U4346 ( .A1(n4257), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3746), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4347 ( .A1(n3407), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4348 ( .A1(n3805), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3408) );
  NAND4_X1 U4349 ( .A1(n3411), .A2(n3410), .A3(n3409), .A4(n3408), .ZN(n3418)
         );
  AOI22_X1 U4350 ( .A1(n3352), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4351 ( .A1(n4246), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4352 ( .A1(n4248), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4353 ( .A1(n4202), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3413) );
  NAND4_X1 U4354 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3417)
         );
  OAI22_X1 U4355 ( .A1(n4511), .A2(STATE2_REG_0__SCAN_IN), .B1(n4105), .B2(
        n4149), .ZN(n3421) );
  AOI22_X1 U4356 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n3921), .B1(n3419), 
        .B2(n4097), .ZN(n3420) );
  XNOR2_X1 U4357 ( .A(n3421), .B(n3420), .ZN(n3487) );
  NAND2_X1 U4358 ( .A1(n3488), .A2(n3487), .ZN(n3527) );
  NAND2_X1 U4359 ( .A1(n3423), .A2(n3422), .ZN(n4591) );
  NAND2_X1 U4360 ( .A1(n3398), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3428) );
  NAND3_X1 U4361 ( .A1(n6485), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6363) );
  INV_X1 U4362 ( .A(n6363), .ZN(n3424) );
  NAND2_X1 U4363 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3424), .ZN(n6420) );
  NAND2_X1 U4364 ( .A1(n6485), .A2(n6420), .ZN(n3425) );
  NOR3_X1 U4365 ( .A1(n6485), .A2(n5075), .A3(n4790), .ZN(n4760) );
  NAND2_X1 U4366 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4760), .ZN(n5027) );
  NAND2_X1 U4367 ( .A1(n3425), .A2(n5027), .ZN(n4640) );
  OAI22_X1 U4368 ( .A1(n4278), .A2(n4640), .B1(n3937), .B2(n6485), .ZN(n3426)
         );
  INV_X1 U4369 ( .A(n3426), .ZN(n3427) );
  NAND2_X1 U4370 ( .A1(n4471), .A2(n3350), .ZN(n3441) );
  INV_X1 U4371 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6746) );
  AOI22_X1 U4372 ( .A1(n3864), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4373 ( .A1(n3153), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4202), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4374 ( .A1(n4257), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4375 ( .A1(n3370), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3430) );
  NAND4_X1 U4376 ( .A1(n3433), .A2(n3432), .A3(n3431), .A4(n3430), .ZN(n3439)
         );
  AOI22_X1 U4377 ( .A1(n3352), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4248), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3437) );
  AOI22_X1 U4378 ( .A1(n3135), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4379 ( .A1(n4246), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4380 ( .A1(n4250), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3434) );
  NAND4_X1 U4381 ( .A1(n3437), .A2(n3436), .A3(n3435), .A4(n3434), .ZN(n3438)
         );
  AOI22_X1 U4382 ( .A1(n3930), .A2(n4114), .B1(n3921), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3440) );
  INV_X1 U4383 ( .A(n3150), .ZN(n3454) );
  AOI22_X1 U4384 ( .A1(n3135), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4385 ( .A1(n4257), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4386 ( .A1(n3407), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4387 ( .A1(n4256), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3442) );
  NAND4_X1 U4388 ( .A1(n3445), .A2(n3444), .A3(n3443), .A4(n3442), .ZN(n3451)
         );
  AOI22_X1 U4389 ( .A1(n3352), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4390 ( .A1(n4246), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4391 ( .A1(n4248), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4392 ( .A1(n4202), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3446) );
  NAND4_X1 U4393 ( .A1(n3449), .A2(n3448), .A3(n3447), .A4(n3446), .ZN(n3450)
         );
  NAND2_X1 U4394 ( .A1(n3930), .A2(n4122), .ZN(n3453) );
  NAND2_X1 U4395 ( .A1(n3921), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3452) );
  NAND2_X1 U4396 ( .A1(n3453), .A2(n3452), .ZN(n3535) );
  AOI22_X1 U4397 ( .A1(n3352), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U4398 ( .A1(n3357), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4399 ( .A1(n4257), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3457) );
  INV_X1 U4400 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4401 ( .A1(n4251), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3456) );
  NAND4_X1 U4402 ( .A1(n3459), .A2(n3458), .A3(n3457), .A4(n3456), .ZN(n3465)
         );
  AOI22_X1 U4403 ( .A1(n4246), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4248), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4404 ( .A1(n3135), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4202), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4405 ( .A1(n4249), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4406 ( .A1(n3156), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3460) );
  NAND4_X1 U4407 ( .A1(n3463), .A2(n3462), .A3(n3461), .A4(n3460), .ZN(n3464)
         );
  NAND2_X1 U4408 ( .A1(n3930), .A2(n4132), .ZN(n3467) );
  NAND2_X1 U4409 ( .A1(n3921), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3466) );
  NAND2_X1 U4410 ( .A1(n3467), .A2(n3466), .ZN(n3545) );
  INV_X1 U4411 ( .A(n3553), .ZN(n3482) );
  AOI22_X1 U4412 ( .A1(n3135), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4413 ( .A1(n4257), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4414 ( .A1(n3357), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4415 ( .A1(n4256), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3469) );
  NAND4_X1 U4416 ( .A1(n3472), .A2(n3471), .A3(n3470), .A4(n3469), .ZN(n3478)
         );
  AOI22_X1 U4417 ( .A1(n3352), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4418 ( .A1(n4246), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4419 ( .A1(n4248), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4420 ( .A1(n4202), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3473) );
  NAND4_X1 U4421 ( .A1(n3476), .A2(n3475), .A3(n3474), .A4(n3473), .ZN(n3477)
         );
  NAND2_X1 U4422 ( .A1(n3930), .A2(n4142), .ZN(n3480) );
  NAND2_X1 U4423 ( .A1(n3921), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3479) );
  NAND2_X1 U4424 ( .A1(n3480), .A2(n3479), .ZN(n3552) );
  INV_X1 U4425 ( .A(n3552), .ZN(n3481) );
  NAND2_X1 U4426 ( .A1(n3482), .A2(n3481), .ZN(n4130) );
  INV_X1 U4427 ( .A(n4130), .ZN(n3485) );
  NOR2_X2 U4428 ( .A1(n3303), .A2(n6497), .ZN(n3669) );
  INV_X1 U4429 ( .A(n3669), .ZN(n3555) );
  XOR2_X1 U4430 ( .A(n3556), .B(n3557), .Z(n6239) );
  INV_X1 U4431 ( .A(n6239), .ZN(n3483) );
  AOI22_X1 U4432 ( .A1(n3483), .A2(n4243), .B1(n4217), .B2(EAX_REG_6__SCAN_IN), 
        .ZN(n3484) );
  OAI21_X1 U4433 ( .B1(n3485), .B2(n3555), .A(n3484), .ZN(n3486) );
  INV_X1 U4434 ( .A(n3488), .ZN(n3489) );
  NAND2_X1 U4435 ( .A1(n4626), .A2(n3669), .ZN(n3490) );
  INV_X1 U4436 ( .A(n4197), .ZN(n3839) );
  NAND2_X1 U4437 ( .A1(n3490), .A2(n3839), .ZN(n4556) );
  NAND2_X1 U4438 ( .A1(n4082), .A2(n3669), .ZN(n3499) );
  NAND2_X1 U4439 ( .A1(n5374), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3538) );
  INV_X1 U4440 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U4441 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6497), .ZN(n3496)
         );
  NAND2_X1 U4442 ( .A1(n4217), .A2(EAX_REG_1__SCAN_IN), .ZN(n3495) );
  OAI211_X1 U4443 ( .C1(n3538), .C2(n5454), .A(n3496), .B(n3495), .ZN(n3497)
         );
  INV_X1 U4444 ( .A(n3497), .ZN(n3498) );
  NAND2_X1 U4445 ( .A1(n3499), .A2(n3498), .ZN(n4460) );
  AOI21_X1 U4446 ( .B1(n4090), .B2(n4335), .A(n6497), .ZN(n4437) );
  OR2_X1 U4447 ( .A1(n3507), .A2(n3555), .ZN(n3512) );
  INV_X1 U4448 ( .A(n3538), .ZN(n3515) );
  NAND2_X1 U4449 ( .A1(n3515), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4450 ( .A1(n3508), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6497), .ZN(n3509) );
  AND2_X1 U4451 ( .A1(n3510), .A2(n3509), .ZN(n3511) );
  NAND2_X1 U4452 ( .A1(n3512), .A2(n3511), .ZN(n4436) );
  NAND2_X1 U4453 ( .A1(n4437), .A2(n4436), .ZN(n4435) );
  INV_X1 U4454 ( .A(n4436), .ZN(n3513) );
  NAND2_X1 U4455 ( .A1(n3513), .A2(n4243), .ZN(n3514) );
  NAND2_X1 U4456 ( .A1(n4435), .A2(n3514), .ZN(n4459) );
  NAND2_X1 U4457 ( .A1(n4460), .A2(n4459), .ZN(n4462) );
  NAND2_X1 U4458 ( .A1(n3515), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3521) );
  OAI21_X1 U4459 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3516), .ZN(n6277) );
  NAND2_X1 U4460 ( .A1(n6277), .A2(n4243), .ZN(n3518) );
  NAND2_X1 U4461 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n4197), .ZN(n3517)
         );
  NAND2_X1 U4462 ( .A1(n3518), .A2(n3517), .ZN(n3519) );
  AOI21_X1 U4463 ( .B1(n4217), .B2(EAX_REG_2__SCAN_IN), .A(n3519), .ZN(n3520)
         );
  AND2_X1 U4464 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  NAND2_X1 U4465 ( .A1(n4462), .A2(n3522), .ZN(n4555) );
  NAND2_X1 U4466 ( .A1(n4556), .A2(n4555), .ZN(n3526) );
  INV_X1 U4467 ( .A(n4462), .ZN(n3524) );
  INV_X1 U4468 ( .A(n3522), .ZN(n3523) );
  NAND2_X1 U4469 ( .A1(n3524), .A2(n3523), .ZN(n3525) );
  NAND2_X1 U4470 ( .A1(n3527), .A2(n4627), .ZN(n3528) );
  OR2_X1 U4471 ( .A1(n4110), .A2(n3555), .ZN(n3534) );
  INV_X1 U4472 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4506) );
  OAI21_X1 U4473 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3529), .A(n3540), 
        .ZN(n6268) );
  AOI22_X1 U4474 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n4197), .B1(n4243), 
        .B2(n6268), .ZN(n3531) );
  NAND2_X1 U4475 ( .A1(n4217), .A2(EAX_REG_3__SCAN_IN), .ZN(n3530) );
  OAI211_X1 U4476 ( .C1(n3538), .C2(n4506), .A(n3531), .B(n3530), .ZN(n3532)
         );
  INV_X1 U4477 ( .A(n3532), .ZN(n3533) );
  NAND2_X1 U4478 ( .A1(n3534), .A2(n3533), .ZN(n4604) );
  XNOR2_X1 U4479 ( .A(n3150), .B(n3535), .ZN(n4113) );
  NAND2_X1 U4480 ( .A1(n4113), .A2(n3669), .ZN(n3544) );
  INV_X1 U4481 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4592) );
  OAI21_X1 U4482 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n5939), .A(n6497), 
        .ZN(n3537) );
  NAND2_X1 U4483 ( .A1(n4217), .A2(EAX_REG_4__SCAN_IN), .ZN(n3536) );
  OAI211_X1 U4484 ( .C1(n3538), .C2(n4592), .A(n3537), .B(n3536), .ZN(n3542)
         );
  AOI21_X1 U4485 ( .B1(n3540), .B2(n3539), .A(n3547), .ZN(n6256) );
  NAND2_X1 U4486 ( .A1(n6256), .A2(n4243), .ZN(n3541) );
  NAND2_X1 U4487 ( .A1(n3542), .A2(n3541), .ZN(n3543) );
  NAND2_X1 U4488 ( .A1(n3544), .A2(n3543), .ZN(n4577) );
  XNOR2_X1 U4489 ( .A(n3546), .B(n3545), .ZN(n4121) );
  NAND2_X1 U4490 ( .A1(n4121), .A2(n3669), .ZN(n3551) );
  NAND2_X1 U4491 ( .A1(n4217), .A2(EAX_REG_5__SCAN_IN), .ZN(n3549) );
  OAI21_X1 U4492 ( .B1(n3547), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3557), 
        .ZN(n6251) );
  AOI22_X1 U4493 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4197), .B1(n4243), 
        .B2(n6251), .ZN(n3548) );
  AND2_X1 U4494 ( .A1(n3549), .A2(n3548), .ZN(n3550) );
  NAND2_X1 U4495 ( .A1(n3551), .A2(n3550), .ZN(n4611) );
  AOI22_X1 U4496 ( .A1(n3930), .A2(n4154), .B1(n3921), .B2(
        INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3554) );
  XNOR2_X1 U4497 ( .A(n4152), .B(n3554), .ZN(n4140) );
  OAI21_X1 U4498 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3558), .A(n3575), 
        .ZN(n6237) );
  AOI22_X1 U4499 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n4197), .B1(n4243), 
        .B2(n6237), .ZN(n3560) );
  NAND2_X1 U4500 ( .A1(n4217), .A2(EAX_REG_7__SCAN_IN), .ZN(n3559) );
  NAND2_X1 U4501 ( .A1(n4965), .A2(n4964), .ZN(n4896) );
  AOI22_X1 U4502 ( .A1(n3135), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4503 ( .A1(n4256), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4504 ( .A1(n3352), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4505 ( .A1(n4248), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4506 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3572)
         );
  AOI22_X1 U4507 ( .A1(n4246), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4508 ( .A1(n3357), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4509 ( .A1(n4202), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4510 ( .A1(n4257), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4511 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3571)
         );
  OAI21_X1 U4512 ( .B1(n3572), .B2(n3571), .A(n3669), .ZN(n3574) );
  NAND2_X1 U4513 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n4197), .ZN(n3573)
         );
  NAND2_X1 U4514 ( .A1(n3574), .A2(n3573), .ZN(n3577) );
  AOI21_X1 U4515 ( .B1(n6684), .B2(n3575), .A(n3602), .ZN(n6226) );
  NOR2_X1 U4516 ( .A1(n6226), .A2(n4273), .ZN(n3576) );
  AOI211_X1 U4517 ( .C1(n4217), .C2(EAX_REG_8__SCAN_IN), .A(n3577), .B(n3576), 
        .ZN(n4897) );
  XOR2_X1 U4518 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3602), .Z(n6218) );
  AOI22_X1 U4519 ( .A1(n3508), .A2(EAX_REG_9__SCAN_IN), .B1(n4197), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4520 ( .A1(n4257), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4521 ( .A1(n3135), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4522 ( .A1(n3352), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4523 ( .A1(n4256), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3578) );
  NAND4_X1 U4524 ( .A1(n3581), .A2(n3580), .A3(n3579), .A4(n3578), .ZN(n3587)
         );
  AOI22_X1 U4525 ( .A1(n4259), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4526 ( .A1(n3357), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4527 ( .A1(n4202), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4528 ( .A1(n4248), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3582) );
  NAND4_X1 U4529 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3586)
         );
  OAI21_X1 U4530 ( .B1(n3587), .B2(n3586), .A(n3669), .ZN(n3588) );
  OAI211_X1 U4531 ( .C1(n6218), .C2(n4273), .A(n3589), .B(n3588), .ZN(n5057)
         );
  NAND2_X1 U4532 ( .A1(n5058), .A2(n5057), .ZN(n5234) );
  INV_X1 U4533 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4534 ( .A1(n3352), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4248), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4535 ( .A1(n4257), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4202), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4536 ( .A1(n4246), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4537 ( .A1(n4256), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3590) );
  NAND4_X1 U4538 ( .A1(n3593), .A2(n3592), .A3(n3591), .A4(n3590), .ZN(n3599)
         );
  AOI22_X1 U4539 ( .A1(n3357), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4540 ( .A1(n4250), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4541 ( .A1(n4259), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4542 ( .A1(n3135), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3594) );
  NAND4_X1 U4543 ( .A1(n3597), .A2(n3596), .A3(n3595), .A4(n3594), .ZN(n3598)
         );
  OAI21_X1 U4544 ( .B1(n3599), .B2(n3598), .A(n3669), .ZN(n3600) );
  OAI21_X1 U4545 ( .B1(n3601), .B2(n3839), .A(n3600), .ZN(n3604) );
  XOR2_X1 U4546 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3605), .Z(n6038) );
  NOR2_X1 U4547 ( .A1(n6038), .A2(n4273), .ZN(n3603) );
  AOI211_X1 U4548 ( .C1(n3508), .C2(EAX_REG_10__SCAN_IN), .A(n3604), .B(n3603), 
        .ZN(n5233) );
  NOR2_X2 U4549 ( .A1(n5234), .A2(n5233), .ZN(n5232) );
  XOR2_X1 U4550 ( .A(n6025), .B(n3630), .Z(n6210) );
  AOI22_X1 U4551 ( .A1(n3508), .A2(EAX_REG_11__SCAN_IN), .B1(n4197), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4552 ( .A1(n3357), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4553 ( .A1(n4259), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4554 ( .A1(n3352), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4555 ( .A1(n4202), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3606) );
  NAND4_X1 U4556 ( .A1(n3609), .A2(n3608), .A3(n3607), .A4(n3606), .ZN(n3615)
         );
  AOI22_X1 U4557 ( .A1(n4246), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4248), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4558 ( .A1(n3135), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4559 ( .A1(n3864), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4560 ( .A1(n4257), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3610) );
  NAND4_X1 U4561 ( .A1(n3613), .A2(n3612), .A3(n3611), .A4(n3610), .ZN(n3614)
         );
  OAI21_X1 U4562 ( .B1(n3615), .B2(n3614), .A(n3669), .ZN(n3616) );
  OAI211_X1 U4563 ( .C1(n6210), .C2(n4273), .A(n3617), .B(n3616), .ZN(n5236)
         );
  AOI22_X1 U4564 ( .A1(n3352), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4248), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4565 ( .A1(n3135), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4566 ( .A1(n4259), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4567 ( .A1(n3357), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3618) );
  NAND4_X1 U4568 ( .A1(n3621), .A2(n3620), .A3(n3619), .A4(n3618), .ZN(n3627)
         );
  AOI22_X1 U4569 ( .A1(n4257), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4570 ( .A1(n3864), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4571 ( .A1(n4246), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4572 ( .A1(n4202), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3622) );
  NAND4_X1 U4573 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n3626)
         );
  OAI21_X1 U4574 ( .B1(n3627), .B2(n3626), .A(n3669), .ZN(n3629) );
  NAND2_X1 U4575 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n4197), .ZN(n3628)
         );
  NAND2_X1 U4576 ( .A1(n3629), .A2(n3628), .ZN(n3633) );
  AOI21_X1 U4577 ( .B1(n6842), .B2(n3631), .A(n3657), .ZN(n6020) );
  NOR2_X1 U4578 ( .A1(n6020), .A2(n4273), .ZN(n3632) );
  AOI211_X1 U4579 ( .C1(n3508), .C2(EAX_REG_12__SCAN_IN), .A(n3633), .B(n3632), 
        .ZN(n5296) );
  XOR2_X1 U4580 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3657), .Z(n6012) );
  AOI22_X1 U4581 ( .A1(n3508), .A2(EAX_REG_13__SCAN_IN), .B1(n4197), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4582 ( .A1(n3352), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4248), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4583 ( .A1(n3357), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4584 ( .A1(n4250), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4585 ( .A1(n3864), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3634) );
  NAND4_X1 U4586 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3643)
         );
  AOI22_X1 U4587 ( .A1(n3135), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4202), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4588 ( .A1(n4257), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4589 ( .A1(n4246), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4590 ( .A1(n4259), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4591 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3642)
         );
  OAI21_X1 U4592 ( .B1(n3643), .B2(n3642), .A(n3669), .ZN(n3644) );
  OAI211_X1 U4593 ( .C1(n6012), .C2(n4273), .A(n3645), .B(n3644), .ZN(n5303)
         );
  AOI22_X1 U4594 ( .A1(n3135), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4248), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4595 ( .A1(n3357), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4596 ( .A1(n4250), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4597 ( .A1(n4257), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3646) );
  NAND4_X1 U4598 ( .A1(n3649), .A2(n3648), .A3(n3647), .A4(n3646), .ZN(n3655)
         );
  AOI22_X1 U4599 ( .A1(n4259), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4600 ( .A1(n4202), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4601 ( .A1(n4246), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4602 ( .A1(n4247), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3650) );
  NAND4_X1 U4603 ( .A1(n3653), .A2(n3652), .A3(n3651), .A4(n3650), .ZN(n3654)
         );
  OAI21_X1 U4604 ( .B1(n3655), .B2(n3654), .A(n3669), .ZN(n3656) );
  OAI21_X1 U4605 ( .B1(n5993), .B2(n3839), .A(n3656), .ZN(n3659) );
  XOR2_X1 U4606 ( .A(n5993), .B(n3660), .Z(n5999) );
  NOR2_X1 U4607 ( .A1(n5999), .A2(n4273), .ZN(n3658) );
  AOI211_X1 U4608 ( .C1(n3508), .C2(EAX_REG_14__SCAN_IN), .A(n3659), .B(n3658), 
        .ZN(n5335) );
  XOR2_X1 U4609 ( .A(n5988), .B(n3685), .Z(n5984) );
  AOI22_X1 U4610 ( .A1(n3508), .A2(EAX_REG_15__SCAN_IN), .B1(n4197), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4611 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n4202), .B1(n4250), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4612 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n4257), .B1(n4256), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4613 ( .A1(n3357), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4614 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n4248), .B1(n4258), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3661) );
  NAND4_X1 U4615 ( .A1(n3664), .A2(n3663), .A3(n3662), .A4(n3661), .ZN(n3671)
         );
  AOI22_X1 U4616 ( .A1(n4259), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4617 ( .A1(n3352), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4618 ( .A1(n3135), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4619 ( .A1(n3864), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3665) );
  NAND4_X1 U4620 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(n3670)
         );
  OAI21_X1 U4621 ( .B1(n3671), .B2(n3670), .A(n3669), .ZN(n3672) );
  OAI211_X1 U4622 ( .C1(n5984), .C2(n4273), .A(n3673), .B(n3672), .ZN(n5338)
         );
  NAND2_X1 U4623 ( .A1(n5334), .A2(n5338), .ZN(n5361) );
  AOI22_X1 U4624 ( .A1(n4257), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3746), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4625 ( .A1(n4250), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4626 ( .A1(n4259), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4627 ( .A1(n4202), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3674) );
  NAND4_X1 U4628 ( .A1(n3677), .A2(n3676), .A3(n3675), .A4(n3674), .ZN(n3689)
         );
  NAND2_X1 U4629 ( .A1(n4648), .A2(n4688), .ZN(n3679) );
  NOR2_X1 U4630 ( .A1(n3679), .A2(n4680), .ZN(n3680) );
  AOI22_X1 U4631 ( .A1(n3357), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4632 ( .A1(n3352), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4248), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4633 ( .A1(n4246), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4634 ( .A1(n3805), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3681) );
  NAND4_X1 U4635 ( .A1(n3684), .A2(n3683), .A3(n3682), .A4(n3681), .ZN(n3688)
         );
  XOR2_X1 U4636 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3690), .Z(n5973) );
  AOI22_X1 U4637 ( .A1(n3508), .A2(EAX_REG_16__SCAN_IN), .B1(n4197), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3686) );
  OAI21_X1 U4638 ( .B1(n5973), .B2(n4273), .A(n3686), .ZN(n3687) );
  AOI221_X1 U4639 ( .B1(n3689), .B2(n4240), .C1(n3688), .C2(n4240), .A(n3687), 
        .ZN(n5362) );
  AOI21_X1 U4640 ( .B1(n6904), .B2(n3691), .A(n3704), .ZN(n5966) );
  AOI22_X1 U4641 ( .A1(n3508), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6497), .ZN(n3703) );
  AOI22_X1 U4642 ( .A1(n3135), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4643 ( .A1(n4248), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4644 ( .A1(n4246), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4645 ( .A1(n3357), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3692) );
  NAND4_X1 U4646 ( .A1(n3695), .A2(n3694), .A3(n3693), .A4(n3692), .ZN(n3701)
         );
  AOI22_X1 U4647 ( .A1(n4259), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4648 ( .A1(n4257), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4649 ( .A1(n3864), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4650 ( .A1(n4202), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3696) );
  NAND4_X1 U4651 ( .A1(n3699), .A2(n3698), .A3(n3697), .A4(n3696), .ZN(n3700)
         );
  AOI221_X1 U4652 ( .B1(n3701), .B2(n4240), .C1(n3700), .C2(n4240), .A(n4243), 
        .ZN(n3702) );
  AOI22_X1 U4653 ( .A1(n4243), .A2(n5966), .B1(n3703), .B2(n3702), .ZN(n5368)
         );
  OAI21_X1 U4654 ( .B1(n3704), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n3731), 
        .ZN(n5958) );
  AOI22_X1 U4655 ( .A1(n4217), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6497), .ZN(n3716) );
  AOI22_X1 U4656 ( .A1(n4246), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4657 ( .A1(n4257), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4658 ( .A1(n4248), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4659 ( .A1(n4202), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3705) );
  NAND4_X1 U4660 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .ZN(n3714)
         );
  AOI22_X1 U4661 ( .A1(n3357), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3746), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4662 ( .A1(n3135), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4663 ( .A1(n4259), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4664 ( .A1(n3805), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3709) );
  NAND4_X1 U4665 ( .A1(n3712), .A2(n3711), .A3(n3710), .A4(n3709), .ZN(n3713)
         );
  OAI21_X1 U4666 ( .B1(n3714), .B2(n3713), .A(n4240), .ZN(n3715) );
  NAND3_X1 U4667 ( .A1(n4273), .A2(n3716), .A3(n3715), .ZN(n3717) );
  XOR2_X1 U4668 ( .A(n5847), .B(n3731), .Z(n5874) );
  AOI22_X1 U4669 ( .A1(n4217), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6497), .ZN(n3730) );
  AOI22_X1 U4670 ( .A1(n3357), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4671 ( .A1(n3135), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4672 ( .A1(n4202), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4673 ( .A1(n4259), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3718) );
  NAND4_X1 U4674 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(n3728)
         );
  AOI22_X1 U4675 ( .A1(n4246), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4676 ( .A1(n3864), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4677 ( .A1(n4248), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4678 ( .A1(n4257), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3723) );
  NAND4_X1 U4679 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3727)
         );
  AOI221_X1 U4680 ( .B1(n3728), .B2(n4240), .C1(n3727), .C2(n4240), .A(n4243), 
        .ZN(n3729) );
  AOI22_X1 U4681 ( .A1(n4243), .A2(n5874), .B1(n3730), .B2(n3729), .ZN(n5520)
         );
  OAI21_X1 U4682 ( .B1(n3732), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n3856), 
        .ZN(n5873) );
  AOI22_X1 U4683 ( .A1(n4217), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6497), .ZN(n3744) );
  AOI22_X1 U4684 ( .A1(n4259), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4685 ( .A1(n3357), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4202), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4686 ( .A1(n4248), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4687 ( .A1(n3805), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3733) );
  NAND4_X1 U4688 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3742)
         );
  AOI22_X1 U4689 ( .A1(n4257), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3746), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4690 ( .A1(n4250), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4691 ( .A1(n3135), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4692 ( .A1(n3412), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3737) );
  NAND4_X1 U4693 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .ZN(n3741)
         );
  OAI21_X1 U4694 ( .B1(n3742), .B2(n3741), .A(n4240), .ZN(n3743) );
  NAND3_X1 U4695 ( .A1(n4273), .A2(n3744), .A3(n3743), .ZN(n3745) );
  OAI21_X1 U4696 ( .B1(n4273), .B2(n5873), .A(n3745), .ZN(n5517) );
  XNOR2_X1 U4697 ( .A(n3856), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5824)
         );
  INV_X1 U4698 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5826) );
  AOI22_X1 U4699 ( .A1(n4246), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4700 ( .A1(n3412), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4248), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4701 ( .A1(n4250), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4702 ( .A1(n3357), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3746), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3747) );
  NAND4_X1 U4703 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n3756)
         );
  AOI22_X1 U4704 ( .A1(n4259), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4705 ( .A1(n4202), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4706 ( .A1(n4251), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4707 ( .A1(n3358), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3751) );
  NAND4_X1 U4708 ( .A1(n3754), .A2(n3753), .A3(n3752), .A4(n3751), .ZN(n3755)
         );
  AOI221_X1 U4709 ( .B1(n3756), .B2(n4240), .C1(n3755), .C2(n4240), .A(n4243), 
        .ZN(n3757) );
  OAI21_X1 U4710 ( .B1(n5826), .B2(STATE2_REG_2__SCAN_IN), .A(n3757), .ZN(
        n3758) );
  AOI21_X1 U4711 ( .B1(n4217), .B2(EAX_REG_21__SCAN_IN), .A(n3758), .ZN(n3759)
         );
  AOI21_X1 U4712 ( .B1(n5824), .B2(n4243), .A(n3759), .ZN(n5507) );
  NAND2_X1 U4713 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3760) );
  INV_X1 U4714 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5577) );
  INV_X1 U4715 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5788) );
  INV_X1 U4716 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5570) );
  INV_X1 U4717 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5561) );
  XNOR2_X1 U4718 ( .A(n3950), .B(n5561), .ZN(n5559) );
  NAND2_X1 U4719 ( .A1(n5559), .A2(n4243), .ZN(n3827) );
  AOI22_X1 U4720 ( .A1(n4259), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4721 ( .A1(n4246), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4722 ( .A1(n4248), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4723 ( .A1(n4202), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3761) );
  NAND4_X1 U4724 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3770)
         );
  AOI22_X1 U4725 ( .A1(n3135), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4726 ( .A1(n4257), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4727 ( .A1(n3357), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4728 ( .A1(n4256), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4729 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3769)
         );
  NOR2_X1 U4730 ( .A1(n3770), .A2(n3769), .ZN(n3828) );
  AOI22_X1 U4731 ( .A1(n4259), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4732 ( .A1(n3357), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4733 ( .A1(n4202), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4734 ( .A1(n3864), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3771) );
  NAND4_X1 U4735 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3780)
         );
  AOI22_X1 U4736 ( .A1(n4257), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4737 ( .A1(n3135), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4738 ( .A1(n4248), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4739 ( .A1(n3352), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4740 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3779)
         );
  NOR2_X1 U4741 ( .A1(n3780), .A2(n3779), .ZN(n3848) );
  AOI22_X1 U4742 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n4259), .B1(n4246), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4743 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4257), .B1(n4256), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4744 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n3135), .B1(n4250), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4745 ( .A1(n4202), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3781) );
  NAND4_X1 U4746 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3790)
         );
  AOI22_X1 U4747 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n3357), .B1(n4251), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4748 ( .A1(n3352), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4749 ( .A1(n4248), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4750 ( .A1(n3864), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4751 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3789)
         );
  NOR2_X1 U4752 ( .A1(n3790), .A2(n3789), .ZN(n3849) );
  NOR2_X1 U4753 ( .A1(n3848), .A2(n3849), .ZN(n3837) );
  AOI22_X1 U4754 ( .A1(n3135), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4755 ( .A1(n4257), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4756 ( .A1(n3357), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4757 ( .A1(n3805), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4758 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3800)
         );
  AOI22_X1 U4759 ( .A1(n3352), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4760 ( .A1(n4246), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4761 ( .A1(n4248), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4762 ( .A1(n4202), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3795) );
  NAND4_X1 U4763 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3799)
         );
  OR2_X1 U4764 ( .A1(n3800), .A2(n3799), .ZN(n3836) );
  NAND2_X1 U4765 ( .A1(n3837), .A2(n3836), .ZN(n3842) );
  NOR2_X1 U4766 ( .A1(n3828), .A2(n3842), .ZN(n3877) );
  AOI22_X1 U4767 ( .A1(n4259), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4768 ( .A1(n4246), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4769 ( .A1(n4248), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4770 ( .A1(n4202), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3801) );
  NAND4_X1 U4771 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3811)
         );
  AOI22_X1 U4772 ( .A1(n3135), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4773 ( .A1(n4257), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4774 ( .A1(n3357), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4775 ( .A1(n3805), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3806) );
  NAND4_X1 U4776 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3810)
         );
  OR2_X1 U4777 ( .A1(n3811), .A2(n3810), .ZN(n3878) );
  NAND2_X1 U4778 ( .A1(n3877), .A2(n3878), .ZN(n4213) );
  AOI22_X1 U4779 ( .A1(n3357), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4780 ( .A1(n4246), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4781 ( .A1(n4247), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4782 ( .A1(n4256), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3812) );
  NAND4_X1 U4783 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3821)
         );
  AOI22_X1 U4784 ( .A1(n4259), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4785 ( .A1(n4257), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4786 ( .A1(n4248), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4202), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4787 ( .A1(n3135), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3816) );
  NAND4_X1 U4788 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3820)
         );
  NOR2_X1 U4789 ( .A1(n3821), .A2(n3820), .ZN(n4214) );
  XOR2_X1 U4790 ( .A(n4213), .B(n4214), .Z(n3822) );
  NAND2_X1 U4791 ( .A1(n3822), .A2(n4240), .ZN(n3825) );
  OAI21_X1 U4792 ( .B1(n5561), .B2(STATE2_REG_2__SCAN_IN), .A(n4273), .ZN(
        n3823) );
  AOI21_X1 U4793 ( .B1(n4217), .B2(EAX_REG_27__SCAN_IN), .A(n3823), .ZN(n3824)
         );
  NAND2_X1 U4794 ( .A1(n3825), .A2(n3824), .ZN(n3826) );
  NAND2_X1 U4795 ( .A1(n3827), .A2(n3826), .ZN(n3886) );
  INV_X1 U4796 ( .A(n3886), .ZN(n3884) );
  XOR2_X1 U4797 ( .A(n3828), .B(n3842), .Z(n3829) );
  AOI21_X1 U4798 ( .B1(n3829), .B2(n4240), .A(n4243), .ZN(n3832) );
  NAND2_X1 U4799 ( .A1(n6497), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3831)
         );
  NAND2_X1 U4800 ( .A1(n4217), .A2(EAX_REG_25__SCAN_IN), .ZN(n3830) );
  NAND3_X1 U4801 ( .A1(n3832), .A2(n3831), .A3(n3830), .ZN(n3835) );
  XOR2_X1 U4802 ( .A(n5788), .B(n3833), .Z(n5864) );
  NAND2_X1 U4803 ( .A1(n4243), .A2(n5864), .ZN(n3834) );
  AND2_X1 U4804 ( .A1(n3835), .A2(n3834), .ZN(n5479) );
  XNOR2_X1 U4805 ( .A(n3847), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5799)
         );
  OR2_X1 U4806 ( .A1(n5799), .A2(n4273), .ZN(n3845) );
  OR2_X1 U4807 ( .A1(n3837), .A2(n3836), .ZN(n3838) );
  AND2_X1 U4808 ( .A1(n4240), .A2(n3838), .ZN(n3843) );
  INV_X1 U4809 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3840) );
  OAI22_X1 U4810 ( .A1(n4238), .A2(n3840), .B1(n3839), .B2(n5577), .ZN(n3841)
         );
  AOI21_X1 U4811 ( .B1(n3843), .B2(n3842), .A(n3841), .ZN(n3844) );
  OR2_X1 U4812 ( .A1(n3858), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3846)
         );
  NAND2_X1 U4813 ( .A1(n3847), .A2(n3846), .ZN(n5805) );
  XOR2_X1 U4814 ( .A(n3849), .B(n3848), .Z(n3850) );
  NAND2_X1 U4815 ( .A1(n3850), .A2(n4240), .ZN(n3853) );
  INV_X1 U4816 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6785) );
  OAI21_X1 U4817 ( .B1(n6785), .B2(STATE2_REG_2__SCAN_IN), .A(n4273), .ZN(
        n3851) );
  AOI21_X1 U4818 ( .B1(n4217), .B2(EAX_REG_23__SCAN_IN), .A(n3851), .ZN(n3852)
         );
  NAND2_X1 U4819 ( .A1(n3853), .A2(n3852), .ZN(n3854) );
  OAI21_X1 U4820 ( .B1(n5805), .B2(n4273), .A(n3854), .ZN(n4314) );
  NOR2_X1 U4821 ( .A1(n5491), .A2(n4314), .ZN(n5478) );
  AND2_X1 U4822 ( .A1(n5479), .A2(n5478), .ZN(n3874) );
  INV_X1 U4823 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3855) );
  OAI21_X1 U4824 ( .B1(n3856), .B2(n5826), .A(n3855), .ZN(n3857) );
  INV_X1 U4825 ( .A(n3857), .ZN(n3859) );
  OR2_X1 U4826 ( .A1(n3859), .A2(n3858), .ZN(n5816) );
  INV_X1 U4827 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4455) );
  AOI22_X1 U4828 ( .A1(n4202), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4829 ( .A1(n4257), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4830 ( .A1(n4259), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4831 ( .A1(n4248), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3860) );
  NAND4_X1 U4832 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3870)
         );
  AOI22_X1 U4833 ( .A1(n4246), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4834 ( .A1(n3357), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4835 ( .A1(n3135), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4836 ( .A1(n4256), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3865) );
  NAND4_X1 U4837 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3869)
         );
  OAI21_X1 U4838 ( .B1(n3870), .B2(n3869), .A(n4240), .ZN(n3872) );
  OAI21_X1 U4839 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5939), .A(n6497), 
        .ZN(n3871) );
  OAI211_X1 U4840 ( .C1(n4455), .C2(n4238), .A(n3872), .B(n3871), .ZN(n3873)
         );
  OAI21_X1 U4841 ( .B1(n5816), .B2(n4273), .A(n3873), .ZN(n5499) );
  INV_X1 U4842 ( .A(n5499), .ZN(n4312) );
  AND2_X1 U4843 ( .A1(n3874), .A2(n4312), .ZN(n5392) );
  AND2_X1 U4844 ( .A1(n3875), .A2(n5570), .ZN(n3876) );
  NOR2_X1 U4845 ( .A1(n3950), .A2(n3876), .ZN(n5778) );
  NAND2_X1 U4846 ( .A1(n5778), .A2(n4243), .ZN(n3883) );
  XNOR2_X1 U4847 ( .A(n3878), .B(n3877), .ZN(n3881) );
  INV_X1 U4848 ( .A(n4240), .ZN(n4271) );
  OAI21_X1 U4849 ( .B1(n5570), .B2(STATE2_REG_2__SCAN_IN), .A(n4273), .ZN(
        n3879) );
  AOI21_X1 U4850 ( .B1(n4217), .B2(EAX_REG_26__SCAN_IN), .A(n3879), .ZN(n3880)
         );
  OAI21_X1 U4851 ( .B1(n3881), .B2(n4271), .A(n3880), .ZN(n3882) );
  INV_X1 U4852 ( .A(n4298), .ZN(n3888) );
  NAND2_X1 U4853 ( .A1(n5496), .A2(n3885), .ZN(n5395) );
  XNOR2_X1 U4854 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3901) );
  XOR2_X1 U4855 ( .A(n3901), .B(n3902), .Z(n3941) );
  INV_X1 U4856 ( .A(n3930), .ZN(n3889) );
  OAI21_X1 U4857 ( .B1(n3889), .B2(n3892), .A(n4684), .ZN(n3898) );
  INV_X1 U4858 ( .A(n3902), .ZN(n3890) );
  OAI21_X1 U4859 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5179), .A(n3890), 
        .ZN(n3893) );
  OAI21_X1 U4860 ( .B1(n4196), .B2(n3893), .A(n3891), .ZN(n3896) );
  OAI21_X1 U4861 ( .B1(n4362), .B2(n4684), .A(n3892), .ZN(n3912) );
  INV_X1 U4862 ( .A(n3893), .ZN(n3894) );
  NAND2_X1 U4863 ( .A1(n3930), .A2(n3894), .ZN(n3895) );
  AOI22_X1 U4864 ( .A1(n3896), .A2(n3912), .B1(n3934), .B2(n3895), .ZN(n3897)
         );
  OAI21_X1 U4865 ( .B1(n3898), .B2(n3941), .A(n3897), .ZN(n3900) );
  NAND3_X1 U4866 ( .A1(n3898), .A2(STATE2_REG_0__SCAN_IN), .A3(n3941), .ZN(
        n3899) );
  OAI211_X1 U4867 ( .C1(n3941), .C2(n3934), .A(n3900), .B(n3899), .ZN(n3916)
         );
  INV_X1 U4868 ( .A(n3921), .ZN(n3906) );
  NAND2_X1 U4869 ( .A1(n3902), .A2(n3901), .ZN(n3904) );
  NAND2_X1 U4870 ( .A1(n4790), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3903) );
  NAND2_X1 U4871 ( .A1(n3904), .A2(n3903), .ZN(n3908) );
  XNOR2_X1 U4872 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3907) );
  INV_X1 U4873 ( .A(n3907), .ZN(n3905) );
  XNOR2_X1 U4874 ( .A(n3908), .B(n3905), .ZN(n3942) );
  NAND2_X1 U4875 ( .A1(n3930), .A2(n3942), .ZN(n3913) );
  OAI211_X1 U4876 ( .C1(n3906), .C2(n3942), .A(n3913), .B(n3912), .ZN(n3915)
         );
  NAND2_X1 U4877 ( .A1(n3908), .A2(n3907), .ZN(n3910) );
  NAND2_X1 U4878 ( .A1(n5075), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3909) );
  NAND2_X1 U4879 ( .A1(n3910), .A2(n3909), .ZN(n3918) );
  XNOR2_X1 U4880 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3917) );
  INV_X1 U4881 ( .A(n3917), .ZN(n3911) );
  XNOR2_X1 U4882 ( .A(n3918), .B(n3911), .ZN(n3940) );
  INV_X1 U4883 ( .A(n4336), .ZN(n4139) );
  OAI22_X1 U4884 ( .A1(n3913), .A2(n3912), .B1(n3940), .B2(n4139), .ZN(n3914)
         );
  AOI21_X1 U4885 ( .B1(n3916), .B2(n3915), .A(n3914), .ZN(n3923) );
  NAND2_X1 U4886 ( .A1(n3918), .A2(n3917), .ZN(n3920) );
  NAND2_X1 U4887 ( .A1(n6485), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3919) );
  NAND2_X1 U4888 ( .A1(n3920), .A2(n3919), .ZN(n3927) );
  AOI21_X1 U4889 ( .B1(n3940), .B2(n3945), .A(n3921), .ZN(n3922) );
  OAI22_X1 U4890 ( .A1(n3923), .A2(n3922), .B1(n3934), .B2(n3945), .ZN(n3924)
         );
  AOI21_X1 U4891 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n3350), .A(n3924), 
        .ZN(n3932) );
  NAND2_X1 U4892 ( .A1(n3925), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3929) );
  NAND2_X1 U4893 ( .A1(n3927), .A2(n3926), .ZN(n3928) );
  NAND2_X1 U4894 ( .A1(n3930), .A2(n3944), .ZN(n3931) );
  NAND2_X1 U4895 ( .A1(n3932), .A2(n3931), .ZN(n3936) );
  INV_X1 U4896 ( .A(n3944), .ZN(n3933) );
  AND3_X1 U4897 ( .A1(n3942), .A2(n3941), .A3(n3940), .ZN(n3943) );
  OR2_X1 U4898 ( .A1(n3944), .A2(n3943), .ZN(n3946) );
  INV_X1 U4899 ( .A(n4414), .ZN(n3947) );
  NOR2_X1 U4900 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6617) );
  INV_X1 U4901 ( .A(n6617), .ZN(n4597) );
  NOR3_X1 U4902 ( .A1(n3350), .A2(n3296), .A3(n4597), .ZN(n6502) );
  NOR2_X1 U4903 ( .A1(n4278), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4283) );
  NOR3_X1 U4904 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6501), .A3(n4273), .ZN(
        n6512) );
  OR2_X1 U4905 ( .A1(n4283), .A2(n6512), .ZN(n3948) );
  INV_X1 U4906 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U4907 ( .A1(n3953), .A2(n6529), .ZN(n6524) );
  NOR2_X1 U4908 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3960) );
  INV_X1 U4909 ( .A(n3960), .ZN(n3954) );
  NOR2_X4 U4910 ( .A1(n6497), .A2(n6109), .ZN(n5249) );
  OAI21_X1 U4911 ( .B1(n6524), .B2(n3954), .A(n5249), .ZN(n3955) );
  INV_X1 U4912 ( .A(n3955), .ZN(n3956) );
  NAND2_X1 U4913 ( .A1(n4534), .A2(n3956), .ZN(n5737) );
  OAI21_X1 U4914 ( .B1(READY_N), .B2(STATEBS16_REG_SCAN_IN), .A(n5249), .ZN(
        n4077) );
  NOR2_X1 U4915 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4077), .ZN(n3957) );
  NAND2_X1 U4916 ( .A1(n4672), .A2(n3957), .ZN(n3958) );
  AOI22_X1 U4917 ( .A1(n6112), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6110), .ZN(n3969) );
  NOR2_X1 U4918 ( .A1(n4285), .A2(n6501), .ZN(n3959) );
  INV_X1 U4919 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6703) );
  INV_X1 U4920 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6857) );
  NOR3_X1 U4921 ( .A1(n6703), .A2(n6857), .A3(n5658), .ZN(n3974) );
  INV_X1 U4922 ( .A(n6524), .ZN(n4494) );
  NOR2_X1 U4923 ( .A1(n4361), .A2(n4494), .ZN(n4330) );
  NAND3_X1 U4924 ( .A1(n4672), .A2(n5249), .A3(n3960), .ZN(n3961) );
  OR2_X2 U4925 ( .A1(n4330), .A2(n3961), .ZN(n6096) );
  NAND3_X1 U4926 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n3967) );
  INV_X1 U4927 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6920) );
  INV_X1 U4928 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6819) );
  NOR2_X1 U4929 ( .A1(n6920), .A2(n6819), .ZN(n3972) );
  INV_X1 U4930 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6694) );
  INV_X1 U4931 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6542) );
  NAND3_X1 U4932 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6094) );
  NOR2_X1 U4933 ( .A1(n6542), .A2(n6094), .ZN(n6082) );
  NAND2_X1 U4934 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6082), .ZN(n6064) );
  NAND2_X1 U4935 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n6058) );
  NOR2_X1 U4936 ( .A1(n6064), .A2(n6058), .ZN(n6051) );
  NAND2_X1 U4937 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6051), .ZN(n3970) );
  INV_X1 U4938 ( .A(n3970), .ZN(n6033) );
  INV_X1 U4939 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6553) );
  INV_X1 U4940 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6551) );
  NOR2_X1 U4941 ( .A1(n6553), .A2(n6551), .ZN(n3971) );
  NAND4_X1 U4942 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6033), .A3(n3971), .A4(n5262), .ZN(n6015) );
  NOR2_X1 U4943 ( .A1(n6694), .A2(n6015), .ZN(n6003) );
  AOI21_X1 U4944 ( .B1(n3972), .B2(n6003), .A(n6004), .ZN(n5998) );
  NAND2_X1 U4945 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5979) );
  INV_X1 U4946 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6561) );
  OAI21_X1 U4947 ( .B1(n5979), .B2(n6561), .A(n6063), .ZN(n3962) );
  INV_X1 U4948 ( .A(n3962), .ZN(n3963) );
  INV_X1 U4949 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5854) );
  INV_X1 U4950 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6563) );
  NOR2_X1 U4951 ( .A1(n5854), .A2(n6563), .ZN(n3964) );
  AND2_X1 U4952 ( .A1(n3964), .A2(REIP_REG_20__SCAN_IN), .ZN(n3965) );
  NOR2_X1 U4953 ( .A1(n6096), .A2(n3965), .ZN(n3966) );
  INV_X1 U4954 ( .A(n5842), .ZN(n5828) );
  AOI21_X1 U4955 ( .B1(n3967), .B2(n6063), .A(n5828), .ZN(n5811) );
  OAI21_X1 U4956 ( .B1(n3974), .B2(n6004), .A(n5811), .ZN(n5783) );
  AOI22_X1 U4957 ( .A1(n5559), .A2(n6120), .B1(REIP_REG_27__SCAN_IN), .B2(
        n5783), .ZN(n3968) );
  OAI211_X1 U4958 ( .C1(n5558), .C2(n6081), .A(n3969), .B(n3968), .ZN(n4081)
         );
  INV_X1 U4959 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6566) );
  INV_X1 U4960 ( .A(n3972), .ZN(n3973) );
  NOR2_X2 U4961 ( .A1(n6014), .A2(n3973), .ZN(n5990) );
  NAND3_X1 U4962 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5845), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5841) );
  NOR2_X2 U4963 ( .A1(n6566), .A2(n5841), .ZN(n5829) );
  NAND4_X1 U4964 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5829), .ZN(n5781) );
  INV_X1 U4965 ( .A(REIP_REG_27__SCAN_IN), .ZN(n3975) );
  INV_X1 U4967 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U4968 ( .A1(n4069), .A2(n4657), .ZN(n3979) );
  CLKBUF_X3 U4969 ( .A(n3987), .Z(n5460) );
  INV_X1 U4970 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3977) );
  NAND2_X1 U4971 ( .A1(n3984), .A2(n3977), .ZN(n3978) );
  NAND3_X1 U4972 ( .A1(n3979), .A2(n5460), .A3(n3978), .ZN(n3980) );
  NAND2_X2 U4973 ( .A1(n3981), .A2(n3980), .ZN(n3985) );
  NAND2_X1 U4974 ( .A1(n4069), .A2(EBX_REG_0__SCAN_IN), .ZN(n3983) );
  INV_X1 U4975 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U4976 ( .A1(n4023), .A2(n5271), .ZN(n3982) );
  AND2_X1 U4977 ( .A1(n3983), .A2(n3982), .ZN(n4428) );
  XNOR2_X2 U4978 ( .A(n3985), .B(n4428), .ZN(n4463) );
  OAI21_X1 U4979 ( .B1(n4463), .B2(n5455), .A(n3985), .ZN(n4558) );
  OR2_X1 U4980 ( .A1(n5458), .A2(EBX_REG_2__SCAN_IN), .ZN(n3991) );
  INV_X1 U4981 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U4982 ( .A1(n4069), .A2(n6360), .ZN(n3989) );
  INV_X1 U4983 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4560) );
  NAND2_X1 U4984 ( .A1(n4535), .A2(n4560), .ZN(n3988) );
  NAND3_X1 U4985 ( .A1(n3989), .A2(n4023), .A3(n3988), .ZN(n3990) );
  AND2_X1 U4986 ( .A1(n3991), .A2(n3990), .ZN(n4557) );
  INV_X1 U4987 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U4988 ( .A1(n4535), .A2(n6695), .ZN(n3995) );
  NAND2_X1 U4989 ( .A1(n5460), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3994)
         );
  NAND3_X1 U4990 ( .A1(n3995), .A2(n4069), .A3(n3994), .ZN(n3996) );
  OAI21_X1 U4991 ( .B1(n4354), .B2(EBX_REG_3__SCAN_IN), .A(n3996), .ZN(n4606)
         );
  NOR2_X2 U4992 ( .A1(n4607), .A2(n4606), .ZN(n4582) );
  MUX2_X1 U4993 ( .A(n5458), .B(n4069), .S(EBX_REG_4__SCAN_IN), .Z(n4000) );
  INV_X1 U4994 ( .A(n4069), .ZN(n3997) );
  NAND2_X1 U4995 ( .A1(n3997), .A2(n5455), .ZN(n4059) );
  NAND2_X1 U4996 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n5455), .ZN(n3998)
         );
  AND2_X1 U4997 ( .A1(n4059), .A2(n3998), .ZN(n3999) );
  NAND2_X1 U4998 ( .A1(n4000), .A2(n3999), .ZN(n4581) );
  NAND2_X1 U4999 ( .A1(n4582), .A2(n4581), .ZN(n4580) );
  MUX2_X1 U5000 ( .A(n4354), .B(n5460), .S(EBX_REG_5__SCAN_IN), .Z(n4001) );
  OAI21_X1 U5001 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5456), .A(n4001), 
        .ZN(n4614) );
  INV_X1 U5002 ( .A(n4002), .ZN(n4621) );
  OR2_X1 U5003 ( .A1(n5458), .A2(EBX_REG_6__SCAN_IN), .ZN(n4006) );
  INV_X1 U5004 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4660) );
  NAND2_X1 U5005 ( .A1(n4069), .A2(n4660), .ZN(n4004) );
  INV_X1 U5006 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U5007 ( .A1(n4535), .A2(n6074), .ZN(n4003) );
  NAND3_X1 U5008 ( .A1(n4004), .A2(n4023), .A3(n4003), .ZN(n4005) );
  MUX2_X1 U5009 ( .A(n4354), .B(n5460), .S(EBX_REG_7__SCAN_IN), .Z(n4007) );
  OAI21_X1 U5010 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5456), .A(n4007), 
        .ZN(n5035) );
  OR2_X1 U5011 ( .A1(n5458), .A2(EBX_REG_8__SCAN_IN), .ZN(n4012) );
  INV_X1 U5012 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U5013 ( .A1(n4069), .A2(n6310), .ZN(n4010) );
  INV_X1 U5014 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4008) );
  NAND2_X1 U5015 ( .A1(n4535), .A2(n4008), .ZN(n4009) );
  NAND3_X1 U5016 ( .A1(n4010), .A2(n4023), .A3(n4009), .ZN(n4011) );
  NAND2_X1 U5017 ( .A1(n4012), .A2(n4011), .ZN(n5069) );
  MUX2_X1 U5018 ( .A(n4354), .B(n5460), .S(EBX_REG_9__SCAN_IN), .Z(n4013) );
  OAI21_X1 U5019 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5456), .A(n4013), 
        .ZN(n5059) );
  MUX2_X1 U5020 ( .A(n5458), .B(n4069), .S(EBX_REG_10__SCAN_IN), .Z(n4015) );
  NAND2_X1 U5021 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5455), .ZN(n4014) );
  INV_X1 U5022 ( .A(n4354), .ZN(n4052) );
  INV_X1 U5023 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U5024 ( .A1(n4052), .A2(n6877), .ZN(n4019) );
  NAND2_X1 U5025 ( .A1(n4535), .A2(n6877), .ZN(n4017) );
  NAND2_X1 U5026 ( .A1(n5460), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4016) );
  NAND3_X1 U5027 ( .A1(n4017), .A2(n4069), .A3(n4016), .ZN(n4018) );
  AND2_X2 U5028 ( .A1(n5229), .A2(n5238), .ZN(n5300) );
  MUX2_X1 U5029 ( .A(n5458), .B(n4069), .S(EBX_REG_12__SCAN_IN), .Z(n4022) );
  NAND2_X1 U5030 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5455), .ZN(n4020) );
  AND2_X1 U5031 ( .A1(n4059), .A2(n4020), .ZN(n4021) );
  NAND2_X1 U5032 ( .A1(n4022), .A2(n4021), .ZN(n5299) );
  INV_X1 U5033 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U5034 ( .A1(n4535), .A2(n5309), .ZN(n4025) );
  NAND2_X1 U5035 ( .A1(n4023), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4024) );
  NAND3_X1 U5036 ( .A1(n4025), .A2(n4069), .A3(n4024), .ZN(n4026) );
  OAI21_X1 U5037 ( .B1(n4354), .B2(EBX_REG_13__SCAN_IN), .A(n4026), .ZN(n5306)
         );
  MUX2_X1 U5038 ( .A(n5458), .B(n4069), .S(EBX_REG_14__SCAN_IN), .Z(n4028) );
  NAND2_X1 U5039 ( .A1(n5455), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4027) );
  INV_X1 U5040 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U5041 ( .A1(n4052), .A2(n5350), .ZN(n4032) );
  NAND2_X1 U5042 ( .A1(n4535), .A2(n5350), .ZN(n4030) );
  NAND2_X1 U5043 ( .A1(n5460), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4029) );
  NAND3_X1 U5044 ( .A1(n4030), .A2(n4069), .A3(n4029), .ZN(n4031) );
  AND2_X2 U5045 ( .A1(n5348), .A2(n5347), .ZN(n5364) );
  MUX2_X1 U5046 ( .A(n5458), .B(n4069), .S(EBX_REG_16__SCAN_IN), .Z(n4035) );
  NAND2_X1 U5047 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5455), .ZN(n4033) );
  AND2_X1 U5048 ( .A1(n4059), .A2(n4033), .ZN(n4034) );
  NAND2_X1 U5049 ( .A1(n4035), .A2(n4034), .ZN(n5363) );
  MUX2_X1 U5050 ( .A(n4354), .B(n4023), .S(EBX_REG_17__SCAN_IN), .Z(n4036) );
  OAI21_X1 U5051 ( .B1(n5456), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n4036), 
        .ZN(n5370) );
  OR2_X2 U5052 ( .A1(n5369), .A2(n5370), .ZN(n5523) );
  OR2_X1 U5053 ( .A1(n5458), .A2(EBX_REG_19__SCAN_IN), .ZN(n4040) );
  INV_X1 U5054 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4303) );
  NAND2_X1 U5055 ( .A1(n4069), .A2(n4303), .ZN(n4038) );
  INV_X1 U5056 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U5057 ( .A1(n4535), .A2(n5525), .ZN(n4037) );
  NAND3_X1 U5058 ( .A1(n4038), .A2(n5460), .A3(n4037), .ZN(n4039) );
  OR2_X2 U5059 ( .A1(n5523), .A2(n5524), .ZN(n5510) );
  NAND2_X1 U5060 ( .A1(n5456), .A2(EBX_REG_18__SCAN_IN), .ZN(n4042) );
  NAND2_X1 U5061 ( .A1(n5455), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U5062 ( .A1(n4042), .A2(n4041), .ZN(n5512) );
  OR2_X1 U5063 ( .A1(n5512), .A2(n4023), .ZN(n5522) );
  OR2_X1 U5064 ( .A1(n5456), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4044)
         );
  INV_X1 U5065 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U5066 ( .A1(n4535), .A2(n5834), .ZN(n4043) );
  NAND2_X1 U5067 ( .A1(n4044), .A2(n4043), .ZN(n4045) );
  NAND2_X1 U5068 ( .A1(n5522), .A2(n4045), .ZN(n4047) );
  NAND2_X1 U5069 ( .A1(n5512), .A2(n5460), .ZN(n5521) );
  INV_X1 U5070 ( .A(n4045), .ZN(n5513) );
  NAND2_X1 U5071 ( .A1(n5521), .A2(n5513), .ZN(n4046) );
  NAND2_X1 U5072 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  NOR2_X4 U5073 ( .A1(n5510), .A2(n4048), .ZN(n5508) );
  MUX2_X1 U5074 ( .A(n5458), .B(n4069), .S(EBX_REG_21__SCAN_IN), .Z(n4051) );
  NAND2_X1 U5075 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n5455), .ZN(n4049) );
  AND2_X1 U5076 ( .A1(n4059), .A2(n4049), .ZN(n4050) );
  NAND2_X1 U5077 ( .A1(n4051), .A2(n4050), .ZN(n5509) );
  INV_X1 U5078 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U5079 ( .A1(n4052), .A2(n5503), .ZN(n4056) );
  NAND2_X1 U5080 ( .A1(n4535), .A2(n5503), .ZN(n4054) );
  NAND2_X1 U5081 ( .A1(n3987), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4053) );
  NAND3_X1 U5082 ( .A1(n4054), .A2(n4069), .A3(n4053), .ZN(n4055) );
  AND2_X1 U5083 ( .A1(n4056), .A2(n4055), .ZN(n5500) );
  AND2_X1 U5084 ( .A1(n5509), .A2(n5500), .ZN(n4057) );
  MUX2_X1 U5085 ( .A(n5458), .B(n4069), .S(EBX_REG_23__SCAN_IN), .Z(n4061) );
  NAND2_X1 U5086 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n5455), .ZN(n4058) );
  AND2_X1 U5087 ( .A1(n4059), .A2(n4058), .ZN(n4060) );
  NAND2_X1 U5088 ( .A1(n4061), .A2(n4060), .ZN(n5432) );
  MUX2_X1 U5089 ( .A(n4354), .B(n5460), .S(EBX_REG_24__SCAN_IN), .Z(n4062) );
  OAI21_X1 U5090 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n5456), .A(n4062), 
        .ZN(n5426) );
  OR2_X2 U5091 ( .A1(n5434), .A2(n5426), .ZN(n5484) );
  OR2_X1 U5092 ( .A1(n5458), .A2(EBX_REG_25__SCAN_IN), .ZN(n4066) );
  INV_X1 U5093 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U5094 ( .A1(n4069), .A2(n5645), .ZN(n4064) );
  INV_X1 U5095 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U5096 ( .A1(n4535), .A2(n6795), .ZN(n4063) );
  NAND3_X1 U5097 ( .A1(n4064), .A2(n3987), .A3(n4063), .ZN(n4065) );
  MUX2_X1 U5098 ( .A(n4354), .B(n3987), .S(EBX_REG_26__SCAN_IN), .Z(n4067) );
  OAI21_X1 U5099 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5456), .A(n4067), 
        .ZN(n4068) );
  INV_X1 U5100 ( .A(n4068), .ZN(n5399) );
  AND2_X2 U5101 ( .A1(n5482), .A2(n5399), .ZN(n4074) );
  OR2_X1 U5102 ( .A1(n5458), .A2(EBX_REG_27__SCAN_IN), .ZN(n4073) );
  INV_X1 U5103 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U5104 ( .A1(n4069), .A2(n5638), .ZN(n4071) );
  INV_X1 U5105 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U5106 ( .A1(n4535), .A2(n5475), .ZN(n4070) );
  NAND3_X1 U5107 ( .A1(n4071), .A2(n5460), .A3(n4070), .ZN(n4072) );
  NAND2_X1 U5108 ( .A1(n4073), .A2(n4072), .ZN(n4075) );
  OR2_X1 U5109 ( .A1(n4074), .A2(n4075), .ZN(n4076) );
  NAND2_X1 U5110 ( .A1(n5472), .A2(n4076), .ZN(n5635) );
  INV_X1 U5111 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6716) );
  NOR2_X1 U5112 ( .A1(n4077), .A2(n6716), .ZN(n4078) );
  NAND2_X1 U5113 ( .A1(n4082), .A2(n4336), .ZN(n4087) );
  INV_X1 U5114 ( .A(n4095), .ZN(n4083) );
  XNOR2_X1 U5115 ( .A(n4083), .B(n4096), .ZN(n4085) );
  NAND2_X1 U5116 ( .A1(n3319), .A2(n4684), .ZN(n4084) );
  AOI21_X1 U5117 ( .B1(n4085), .B2(n4534), .A(n4084), .ZN(n4086) );
  NAND2_X1 U5118 ( .A1(n4087), .A2(n4086), .ZN(n4526) );
  INV_X1 U5119 ( .A(n4534), .ZN(n6616) );
  NAND2_X1 U5120 ( .A1(n4362), .A2(n4676), .ZN(n4098) );
  OAI21_X1 U5121 ( .B1(n6616), .B2(n4095), .A(n4098), .ZN(n4088) );
  INV_X1 U5122 ( .A(n4088), .ZN(n4089) );
  NAND2_X1 U5123 ( .A1(n4465), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4091)
         );
  NAND2_X1 U5124 ( .A1(n4091), .A2(n4657), .ZN(n4092) );
  AND2_X1 U5125 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U5126 ( .A1(n4465), .A2(n6348), .ZN(n4093) );
  NAND2_X1 U5127 ( .A1(n4526), .A2(n4525), .ZN(n4094) );
  NAND2_X1 U5128 ( .A1(n4094), .A2(n4093), .ZN(n6269) );
  NAND2_X1 U5129 ( .A1(n6269), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4101)
         );
  NAND2_X1 U5130 ( .A1(n4096), .A2(n4095), .ZN(n4106) );
  XNOR2_X1 U5131 ( .A(n4106), .B(n4097), .ZN(n4099) );
  OAI21_X1 U5132 ( .B1(n4099), .B2(n6616), .A(n4098), .ZN(n4100) );
  NAND2_X1 U5133 ( .A1(n4101), .A2(n6271), .ZN(n4104) );
  INV_X1 U5134 ( .A(n6269), .ZN(n4102) );
  NAND2_X1 U5135 ( .A1(n4102), .A2(n6360), .ZN(n4103) );
  AND2_X1 U5136 ( .A1(n4104), .A2(n4103), .ZN(n6262) );
  NAND2_X1 U5137 ( .A1(n4106), .A2(n4105), .ZN(n4115) );
  INV_X1 U5138 ( .A(n4114), .ZN(n4107) );
  XNOR2_X1 U5139 ( .A(n4115), .B(n4107), .ZN(n4108) );
  NAND2_X1 U5140 ( .A1(n4108), .A2(n4534), .ZN(n4109) );
  INV_X1 U5141 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6344) );
  XNOR2_X1 U5142 ( .A(n4111), .B(n6344), .ZN(n6263) );
  NAND2_X1 U5143 ( .A1(n6262), .A2(n6263), .ZN(n6261) );
  NAND2_X1 U5144 ( .A1(n4111), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4112)
         );
  NAND2_X1 U5145 ( .A1(n6261), .A2(n4112), .ZN(n6254) );
  NAND2_X1 U5146 ( .A1(n4113), .A2(n4336), .ZN(n4118) );
  NAND2_X1 U5147 ( .A1(n4115), .A2(n4114), .ZN(n4124) );
  XNOR2_X1 U5148 ( .A(n4124), .B(n4122), .ZN(n4116) );
  NAND2_X1 U5149 ( .A1(n4116), .A2(n4534), .ZN(n4117) );
  NAND2_X1 U5150 ( .A1(n4118), .A2(n4117), .ZN(n4119) );
  INV_X1 U5151 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6337) );
  XNOR2_X1 U5152 ( .A(n4119), .B(n6337), .ZN(n6253) );
  NAND2_X1 U5153 ( .A1(n6254), .A2(n6253), .ZN(n6252) );
  NAND2_X1 U5154 ( .A1(n4119), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4120)
         );
  NAND2_X1 U5155 ( .A1(n6252), .A2(n4120), .ZN(n6246) );
  NAND2_X1 U5156 ( .A1(n4121), .A2(n4336), .ZN(n4127) );
  INV_X1 U5157 ( .A(n4122), .ZN(n4123) );
  OR2_X1 U5158 ( .A1(n4124), .A2(n4123), .ZN(n4131) );
  XNOR2_X1 U5159 ( .A(n4131), .B(n4132), .ZN(n4125) );
  NAND2_X1 U5160 ( .A1(n4125), .A2(n4534), .ZN(n4126) );
  INV_X1 U5161 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6317) );
  XNOR2_X1 U5162 ( .A(n4128), .B(n6317), .ZN(n6245) );
  NAND2_X1 U5163 ( .A1(n6246), .A2(n6245), .ZN(n6244) );
  NAND2_X1 U5164 ( .A1(n4128), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4129)
         );
  NAND2_X1 U5165 ( .A1(n6244), .A2(n4129), .ZN(n4656) );
  NAND3_X1 U5166 ( .A1(n4152), .A2(n4130), .A3(n4336), .ZN(n4136) );
  INV_X1 U5167 ( .A(n4131), .ZN(n4133) );
  NAND2_X1 U5168 ( .A1(n4133), .A2(n4132), .ZN(n4141) );
  XNOR2_X1 U5169 ( .A(n4141), .B(n4142), .ZN(n4134) );
  NAND2_X1 U5170 ( .A1(n4134), .A2(n4534), .ZN(n4135) );
  NAND2_X1 U5171 ( .A1(n4136), .A2(n4135), .ZN(n4137) );
  XNOR2_X1 U5172 ( .A(n4137), .B(n4660), .ZN(n4655) );
  NAND2_X1 U5173 ( .A1(n4656), .A2(n4655), .ZN(n4654) );
  NAND2_X1 U5174 ( .A1(n4137), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4138)
         );
  NAND2_X1 U5175 ( .A1(n4654), .A2(n4138), .ZN(n6231) );
  OR2_X1 U5176 ( .A1(n4140), .A2(n4139), .ZN(n4146) );
  INV_X1 U5177 ( .A(n4141), .ZN(n4143) );
  NAND2_X1 U5178 ( .A1(n4143), .A2(n4142), .ZN(n4153) );
  XNOR2_X1 U5179 ( .A(n4153), .B(n4154), .ZN(n4144) );
  NAND2_X1 U5180 ( .A1(n4144), .A2(n4534), .ZN(n4145) );
  NAND2_X1 U5181 ( .A1(n4146), .A2(n4145), .ZN(n4147) );
  INV_X1 U5182 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6315) );
  XNOR2_X1 U5183 ( .A(n4147), .B(n6315), .ZN(n6230) );
  NAND2_X1 U5184 ( .A1(n6231), .A2(n6230), .ZN(n6233) );
  NAND2_X1 U5185 ( .A1(n4147), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4148)
         );
  NAND2_X1 U5186 ( .A1(n6233), .A2(n4148), .ZN(n6222) );
  NAND2_X1 U5187 ( .A1(n4336), .A2(n4154), .ZN(n4150) );
  NOR2_X1 U5188 ( .A1(n4150), .A2(n4149), .ZN(n4151) );
  INV_X1 U5189 ( .A(n4153), .ZN(n4155) );
  NAND3_X1 U5190 ( .A1(n4155), .A2(n4534), .A3(n4154), .ZN(n4156) );
  NAND2_X1 U5191 ( .A1(n4164), .A2(n4156), .ZN(n4157) );
  XNOR2_X1 U5192 ( .A(n4157), .B(n6310), .ZN(n6224) );
  NAND2_X1 U5193 ( .A1(n6222), .A2(n6224), .ZN(n6223) );
  NAND2_X1 U5194 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4158)
         );
  NAND2_X1 U5195 ( .A1(n6223), .A2(n4158), .ZN(n6214) );
  INV_X1 U5196 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U5197 ( .A1(n4164), .A2(n6302), .ZN(n6215) );
  OR2_X1 U5198 ( .A1(n4164), .A2(n6302), .ZN(n6216) );
  NAND2_X1 U5199 ( .A1(n4159), .A2(n6216), .ZN(n5278) );
  INV_X1 U5200 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4160) );
  NAND2_X1 U5201 ( .A1(n4164), .A2(n4160), .ZN(n5277) );
  INV_X1 U5202 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6293) );
  AND2_X1 U5203 ( .A1(n4164), .A2(n6293), .ZN(n4163) );
  OR2_X1 U5204 ( .A1(n4164), .A2(n4160), .ZN(n6207) );
  INV_X1 U5205 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6782) );
  NOR2_X1 U5206 ( .A1(n4164), .A2(n6782), .ZN(n5315) );
  OR2_X1 U5207 ( .A1(n5312), .A2(n5315), .ZN(n4165) );
  NAND2_X1 U5208 ( .A1(n4164), .A2(n6782), .ZN(n5313) );
  NAND2_X1 U5209 ( .A1(n4165), .A2(n5313), .ZN(n5892) );
  NAND2_X1 U5210 ( .A1(n5892), .A2(n5893), .ZN(n4168) );
  INV_X1 U5211 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4166) );
  NAND2_X1 U5212 ( .A1(n4164), .A2(n4166), .ZN(n4167) );
  NAND2_X1 U5213 ( .A1(n4168), .A2(n4167), .ZN(n5353) );
  INV_X1 U5214 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5354) );
  AND2_X1 U5215 ( .A1(n4164), .A2(n5354), .ZN(n5402) );
  INV_X1 U5216 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6679) );
  INV_X1 U5217 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4176) );
  AND2_X1 U5218 ( .A1(n4164), .A2(n4176), .ZN(n4169) );
  OR2_X1 U5219 ( .A1(n4164), .A2(n5354), .ZN(n5403) );
  XNOR2_X1 U5220 ( .A(n4164), .B(n6679), .ZN(n5406) );
  INV_X1 U5221 ( .A(n5406), .ZN(n4171) );
  AND2_X1 U5222 ( .A1(n5403), .A2(n4171), .ZN(n4172) );
  INV_X1 U5223 ( .A(n4174), .ZN(n5712) );
  INV_X1 U5224 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4177) );
  INV_X1 U5225 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4175) );
  NAND2_X1 U5226 ( .A1(n5712), .A2(n3163), .ZN(n4178) );
  NAND2_X1 U5227 ( .A1(n4178), .A2(n4187), .ZN(n4180) );
  INV_X1 U5228 ( .A(n5712), .ZN(n5884) );
  AND2_X1 U5229 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U5230 ( .A1(n5884), .A2(n5701), .ZN(n4179) );
  NAND2_X1 U5231 ( .A1(n4180), .A2(n4179), .ZN(n5703) );
  NAND2_X1 U5232 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U5233 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5694) );
  NOR2_X1 U5234 ( .A1(n5664), .A2(n5694), .ZN(n4307) );
  AND2_X1 U5235 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4393) );
  NAND2_X1 U5236 ( .A1(n4307), .A2(n4393), .ZN(n4181) );
  NAND2_X1 U5237 ( .A1(n4164), .A2(n4181), .ZN(n4182) );
  NAND2_X1 U5238 ( .A1(n5703), .A2(n4182), .ZN(n4185) );
  NOR2_X1 U5239 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5666) );
  NOR2_X1 U5240 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5427) );
  NOR2_X1 U5241 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5692) );
  AND3_X1 U5242 ( .A1(n5666), .A2(n5427), .A3(n5692), .ZN(n4183) );
  NAND2_X1 U5243 ( .A1(n4185), .A2(n4184), .ZN(n4291) );
  INV_X1 U5244 ( .A(n4291), .ZN(n4186) );
  INV_X1 U5245 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5649) );
  NOR2_X1 U5246 ( .A1(n4187), .A2(n5649), .ZN(n5567) );
  NAND2_X1 U5247 ( .A1(n4164), .A2(n5645), .ZN(n4289) );
  AND2_X1 U5248 ( .A1(n5567), .A2(n4289), .ZN(n4188) );
  NAND2_X1 U5249 ( .A1(n4290), .A2(n4188), .ZN(n5556) );
  NAND2_X1 U5250 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U5251 ( .A1(n3138), .A2(n3162), .ZN(n4192) );
  INV_X1 U5252 ( .A(n5653), .ZN(n4190) );
  OR2_X1 U5253 ( .A1(n4164), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5565)
         );
  INV_X1 U5254 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U5255 ( .A1(n5627), .A2(n5638), .ZN(n4189) );
  INV_X1 U5256 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6714) );
  NAND4_X1 U5257 ( .A1(n4190), .A2(n4323), .A3(n6714), .A4(n5609), .ZN(n4191)
         );
  XNOR2_X1 U5258 ( .A(n4193), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5617)
         );
  OAI21_X1 U5259 ( .B1(n3678), .B2(n4672), .A(n4365), .ZN(n4194) );
  INV_X1 U5260 ( .A(n4194), .ZN(n4195) );
  NAND2_X1 U5261 ( .A1(n4347), .A2(n4196), .ZN(n6489) );
  AOI22_X1 U5262 ( .A1(n4217), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4197), .ZN(n4276) );
  INV_X1 U5263 ( .A(n5517), .ZN(n4198) );
  NAND2_X1 U5264 ( .A1(n4198), .A2(n5507), .ZN(n4199) );
  NOR2_X1 U5265 ( .A1(n4200), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4201)
         );
  OR2_X1 U5266 ( .A1(n4223), .A2(n4201), .ZN(n5769) );
  AOI22_X1 U5267 ( .A1(n4259), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U5268 ( .A1(n4246), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5269 ( .A1(n4248), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U5270 ( .A1(n4202), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4203) );
  NAND4_X1 U5271 ( .A1(n4206), .A2(n4205), .A3(n4204), .A4(n4203), .ZN(n4212)
         );
  AOI22_X1 U5272 ( .A1(n3135), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U5273 ( .A1(n4257), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U5274 ( .A1(n3357), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U5275 ( .A1(n4256), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4207) );
  NAND4_X1 U5276 ( .A1(n4210), .A2(n4209), .A3(n4208), .A4(n4207), .ZN(n4211)
         );
  OR2_X1 U5277 ( .A1(n4212), .A2(n4211), .ZN(n4224) );
  NOR2_X1 U5278 ( .A1(n4214), .A2(n4213), .ZN(n4225) );
  XNOR2_X1 U5279 ( .A(n4224), .B(n4225), .ZN(n4219) );
  INV_X1 U5280 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4215) );
  OAI21_X1 U5281 ( .B1(n4215), .B2(STATE2_REG_2__SCAN_IN), .A(n4273), .ZN(
        n4216) );
  AOI21_X1 U5282 ( .B1(n4217), .B2(EAX_REG_28__SCAN_IN), .A(n4216), .ZN(n4218)
         );
  OAI21_X1 U5283 ( .B1(n4219), .B2(n4271), .A(n4218), .ZN(n4220) );
  OAI21_X1 U5284 ( .B1(n5769), .B2(n4273), .A(n4220), .ZN(n4221) );
  INV_X1 U5285 ( .A(n4221), .ZN(n4297) );
  INV_X1 U5286 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5385) );
  XNOR2_X1 U5287 ( .A(n4223), .B(n5385), .ZN(n5759) );
  NAND2_X1 U5288 ( .A1(n4225), .A2(n4224), .ZN(n4266) );
  AOI22_X1 U5289 ( .A1(n3135), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4202), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4229) );
  AOI22_X1 U5290 ( .A1(n4257), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U5291 ( .A1(n3357), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4227) );
  AOI22_X1 U5292 ( .A1(n4259), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4226) );
  NAND4_X1 U5293 ( .A1(n4229), .A2(n4228), .A3(n4227), .A4(n4226), .ZN(n4235)
         );
  AOI22_X1 U5294 ( .A1(n4246), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U5295 ( .A1(n4248), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4232) );
  AOI22_X1 U5296 ( .A1(n4250), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4231) );
  AOI22_X1 U5297 ( .A1(n4256), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4230) );
  NAND4_X1 U5298 ( .A1(n4233), .A2(n4232), .A3(n4231), .A4(n4230), .ZN(n4234)
         );
  NOR2_X1 U5299 ( .A1(n4235), .A2(n4234), .ZN(n4267) );
  XOR2_X1 U5300 ( .A(n4266), .B(n4267), .Z(n4241) );
  INV_X1 U5301 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4237) );
  AOI21_X1 U5302 ( .B1(n6497), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4243), 
        .ZN(n4236) );
  OAI21_X1 U5303 ( .B1(n4238), .B2(n4237), .A(n4236), .ZN(n4239) );
  AOI21_X1 U5304 ( .B1(n4241), .B2(n4240), .A(n4239), .ZN(n4242) );
  AOI21_X1 U5305 ( .B1(n5759), .B2(n4243), .A(n4242), .ZN(n5380) );
  AND2_X1 U5306 ( .A1(n4296), .A2(n5380), .ZN(n4244) );
  AND2_X2 U5307 ( .A1(n4313), .A2(n4244), .ZN(n5382) );
  XOR2_X1 U5308 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .B(n4245), .Z(n5758) );
  AOI22_X1 U5309 ( .A1(n4246), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U5310 ( .A1(n4248), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U5311 ( .A1(n4250), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U5312 ( .A1(n4251), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4252) );
  NAND4_X1 U5313 ( .A1(n4255), .A2(n4254), .A3(n4253), .A4(n4252), .ZN(n4265)
         );
  AOI22_X1 U5314 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n3135), .B1(n4202), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U5315 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n3357), .B1(n3864), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4262) );
  AOI22_X1 U5316 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n4257), .B1(n4256), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4261) );
  AOI22_X1 U5317 ( .A1(n4259), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4260) );
  NAND4_X1 U5318 ( .A1(n4263), .A2(n4262), .A3(n4261), .A4(n4260), .ZN(n4264)
         );
  NOR2_X1 U5319 ( .A1(n4265), .A2(n4264), .ZN(n4269) );
  NOR2_X1 U5320 ( .A1(n4267), .A2(n4266), .ZN(n4268) );
  XOR2_X1 U5321 ( .A(n4269), .B(n4268), .Z(n4272) );
  AOI22_X1 U5322 ( .A1(n4217), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6497), .ZN(n4270) );
  OAI21_X1 U5323 ( .B1(n4272), .B2(n4271), .A(n4270), .ZN(n4274) );
  MUX2_X1 U5324 ( .A(n5758), .B(n4274), .S(n4273), .Z(n4408) );
  NAND2_X1 U5325 ( .A1(n5382), .A2(n4408), .ZN(n4275) );
  XOR2_X1 U5326 ( .A(n4276), .B(n4275), .Z(n5739) );
  NAND3_X1 U5327 ( .A1(n3350), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6516) );
  INV_X1 U5328 ( .A(n6516), .ZN(n4277) );
  NOR2_X2 U5329 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6371) );
  INV_X2 U5330 ( .A(n6286), .ZN(n6273) );
  NAND2_X1 U5331 ( .A1(n5739), .A2(n6273), .ZN(n4287) );
  NAND2_X1 U5332 ( .A1(n5733), .A2(n4278), .ZN(n6612) );
  AND2_X1 U5333 ( .A1(n6612), .A2(n3350), .ZN(n4279) );
  NAND2_X1 U5334 ( .A1(n3350), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4281) );
  NAND2_X1 U5335 ( .A1(n5939), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4280) );
  AND2_X1 U5336 ( .A1(n4281), .A2(n4280), .ZN(n4466) );
  INV_X1 U5337 ( .A(n4466), .ZN(n4282) );
  INV_X1 U5338 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5736) );
  INV_X2 U5339 ( .A(n6349), .ZN(n6325) );
  NAND2_X1 U5340 ( .A1(n6325), .A2(REIP_REG_31__SCAN_IN), .ZN(n5612) );
  OAI21_X1 U5341 ( .B1(n5588), .B2(n5736), .A(n5612), .ZN(n4284) );
  AOI21_X1 U5342 ( .B1(n6257), .B2(n4285), .A(n4284), .ZN(n4286) );
  OAI21_X1 U5343 ( .B1(n5617), .B2(n6278), .A(n4288), .ZN(U2955) );
  NOR3_X1 U5344 ( .A1(n5569), .A2(n4187), .A3(n5638), .ZN(n4294) );
  OR2_X1 U5345 ( .A1(n5565), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4293)
         );
  NOR2_X1 U5346 ( .A1(n4292), .A2(n4293), .ZN(n5554) );
  OAI22_X1 U5347 ( .A1(n4294), .A2(n5554), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5638), .ZN(n4295) );
  XNOR2_X1 U5348 ( .A(n4295), .B(n5627), .ZN(n5634) );
  NOR2_X1 U5349 ( .A1(n4298), .A2(n4297), .ZN(n4299) );
  INV_X1 U5350 ( .A(n5545), .ZN(n5772) );
  INV_X1 U5351 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6862) );
  NOR2_X1 U5352 ( .A1(n6349), .A2(n6862), .ZN(n5629) );
  AOI21_X1 U5353 ( .B1(n6283), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5629), 
        .ZN(n4300) );
  OAI21_X1 U5354 ( .B1(n5769), .B2(n6280), .A(n4300), .ZN(n4301) );
  AOI21_X1 U5355 ( .B1(n5772), .B2(n6273), .A(n4301), .ZN(n4302) );
  OAI21_X1 U5356 ( .B1(n5634), .B2(n6278), .A(n4302), .ZN(U2958) );
  XNOR2_X1 U5357 ( .A(n4164), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5704)
         );
  NAND2_X1 U5358 ( .A1(n5703), .A2(n5704), .ZN(n4306) );
  OR2_X1 U5359 ( .A1(n4164), .A2(n4303), .ZN(n4304) );
  INV_X1 U5360 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4305) );
  NAND2_X1 U5361 ( .A1(n4164), .A2(n4305), .ZN(n5683) );
  NOR2_X1 U5362 ( .A1(n4164), .A2(n4305), .ZN(n5682) );
  XNOR2_X1 U5363 ( .A(n4164), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5593)
         );
  AND2_X2 U5364 ( .A1(n5592), .A2(n5593), .ZN(n5590) );
  NOR2_X1 U5365 ( .A1(n4164), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5582)
         );
  INV_X1 U5366 ( .A(n4307), .ZN(n4308) );
  NAND2_X1 U5367 ( .A1(n5435), .A2(n6272), .ZN(n4322) );
  NAND2_X1 U5368 ( .A1(n4313), .A2(n4312), .ZN(n4315) );
  INV_X1 U5369 ( .A(n4314), .ZN(n4316) );
  INV_X1 U5370 ( .A(REIP_REG_23__SCAN_IN), .ZN(n4317) );
  NOR2_X1 U5371 ( .A1(n6349), .A2(n4317), .ZN(n5438) );
  NOR2_X1 U5372 ( .A1(n6280), .A2(n5805), .ZN(n4318) );
  AOI211_X1 U5373 ( .C1(n6283), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5438), 
        .B(n4318), .ZN(n4319) );
  NAND2_X1 U5374 ( .A1(n4322), .A2(n4321), .ZN(U2963) );
  NAND2_X1 U5375 ( .A1(n5569), .A2(n4323), .ZN(n5377) );
  INV_X1 U5376 ( .A(n5377), .ZN(n4324) );
  NAND2_X1 U5377 ( .A1(n4324), .A2(n6714), .ZN(n4327) );
  NAND2_X1 U5378 ( .A1(n4325), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4326) );
  OR3_X1 U5379 ( .A1(n4537), .A2(n4330), .A3(READY_N), .ZN(n4492) );
  NOR2_X1 U5380 ( .A1(n5374), .A2(n4362), .ZN(n4331) );
  AOI21_X1 U5381 ( .B1(n4492), .B2(n4331), .A(n4680), .ZN(n4332) );
  NAND2_X1 U5382 ( .A1(n4539), .A2(n4332), .ZN(n4345) );
  NAND3_X1 U5383 ( .A1(n4489), .A2(n6473), .A3(n4361), .ZN(n4342) );
  INV_X1 U5384 ( .A(n4333), .ZN(n4334) );
  NAND2_X1 U5385 ( .A1(n4574), .A2(n4334), .ZN(n4338) );
  NAND2_X1 U5386 ( .A1(n4336), .A2(n4335), .ZN(n4373) );
  AND2_X1 U5387 ( .A1(n4373), .A2(n4672), .ZN(n4337) );
  NAND2_X1 U5388 ( .A1(n4338), .A2(n4337), .ZN(n4369) );
  NAND2_X1 U5389 ( .A1(n4347), .A2(n4369), .ZN(n4339) );
  NAND2_X1 U5390 ( .A1(n3939), .A2(n4339), .ZN(n4497) );
  NAND2_X1 U5391 ( .A1(n4361), .A2(n6524), .ZN(n4340) );
  NOR2_X1 U5392 ( .A1(READY_N), .A2(n4414), .ZN(n4563) );
  NAND3_X1 U5393 ( .A1(n4340), .A2(n4563), .A3(n4680), .ZN(n4341) );
  NAND3_X1 U5394 ( .A1(n4342), .A2(n4497), .A3(n4341), .ZN(n4343) );
  NAND2_X1 U5395 ( .A1(n4343), .A2(n4569), .ZN(n4344) );
  NAND2_X1 U5396 ( .A1(n4347), .A2(n5247), .ZN(n4565) );
  NAND2_X1 U5397 ( .A1(n4565), .A2(n6489), .ZN(n4413) );
  OAI22_X1 U5398 ( .A1(n4537), .A2(n5455), .B1(n4570), .B2(n4357), .ZN(n4348)
         );
  OR2_X1 U5399 ( .A1(n4413), .A2(n4348), .ZN(n4349) );
  NOR2_X1 U5400 ( .A1(n5929), .A2(n4349), .ZN(n4350) );
  OR2_X1 U5401 ( .A1(n5456), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4353)
         );
  INV_X1 U5402 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4351) );
  NAND2_X1 U5403 ( .A1(n4535), .A2(n4351), .ZN(n4352) );
  NAND2_X1 U5404 ( .A1(n4353), .A2(n4352), .ZN(n5457) );
  MUX2_X1 U5405 ( .A(n4354), .B(n5460), .S(EBX_REG_28__SCAN_IN), .Z(n4355) );
  OAI21_X1 U5406 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5456), .A(n4355), 
        .ZN(n5473) );
  AOI22_X1 U5407 ( .A1(n5456), .A2(EBX_REG_30__SCAN_IN), .B1(n5455), .B2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5462) );
  XNOR2_X2 U5408 ( .A(n4356), .B(n5462), .ZN(n5749) );
  OR2_X1 U5409 ( .A1(n4537), .A2(n6616), .ZN(n6496) );
  INV_X1 U5410 ( .A(n4357), .ZN(n4358) );
  NAND2_X1 U5411 ( .A1(n4358), .A2(n4570), .ZN(n4359) );
  AND2_X1 U5412 ( .A1(n6496), .A2(n4359), .ZN(n4360) );
  NAND2_X1 U5413 ( .A1(n4415), .A2(n4361), .ZN(n5445) );
  INV_X1 U5414 ( .A(n5456), .ZN(n4366) );
  NAND2_X1 U5415 ( .A1(n5374), .A2(n4362), .ZN(n4363) );
  NAND2_X1 U5416 ( .A1(n4363), .A2(n4680), .ZN(n4364) );
  OR2_X1 U5417 ( .A1(n5251), .A2(n4680), .ZN(n4498) );
  OAI211_X1 U5418 ( .C1(n4366), .C2(n4365), .A(n4364), .B(n4498), .ZN(n4367)
         );
  INV_X1 U5419 ( .A(n4367), .ZN(n4368) );
  OAI211_X1 U5420 ( .C1(n4370), .C2(n4023), .A(n4369), .B(n4368), .ZN(n4371)
         );
  OR2_X1 U5421 ( .A1(n4372), .A2(n4371), .ZN(n4473) );
  INV_X1 U5422 ( .A(n4509), .ZN(n4480) );
  OR2_X1 U5423 ( .A1(n4377), .A2(n4375), .ZN(n4376) );
  INV_X1 U5424 ( .A(n4373), .ZN(n4374) );
  INV_X1 U5425 ( .A(n4429), .ZN(n4482) );
  NAND2_X1 U5426 ( .A1(n5690), .A2(n5317), .ZN(n5608) );
  INV_X1 U5427 ( .A(n5608), .ZN(n5691) );
  INV_X1 U5428 ( .A(n4376), .ZN(n5911) );
  INV_X1 U5429 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U5430 ( .A1(n5911), .A2(n6594), .ZN(n4378) );
  NAND2_X1 U5431 ( .A1(n6349), .A2(n4377), .ZN(n5724) );
  NAND4_X1 U5432 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A3(INSTADDRPOINTER_REG_17__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4390) );
  NOR2_X1 U5433 ( .A1(n6315), .A2(n6310), .ZN(n6304) );
  INV_X1 U5434 ( .A(n6304), .ZN(n5285) );
  NAND2_X1 U5435 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5286) );
  NOR2_X1 U5436 ( .A1(n5285), .A2(n5286), .ZN(n4381) );
  NAND4_X1 U5437 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6318) );
  NOR3_X1 U5438 ( .A1(n6317), .A2(n4660), .A3(n6318), .ZN(n5287) );
  NAND2_X1 U5439 ( .A1(n4381), .A2(n5287), .ZN(n5320) );
  NAND2_X1 U5440 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5908) );
  NOR2_X1 U5441 ( .A1(n4166), .A2(n5908), .ZN(n5918) );
  NAND2_X1 U5442 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5918), .ZN(n5407) );
  NAND2_X1 U5443 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5904) );
  NOR2_X1 U5444 ( .A1(n5407), .A2(n5904), .ZN(n4382) );
  INV_X1 U5445 ( .A(n4382), .ZN(n4379) );
  NOR2_X1 U5446 ( .A1(n5320), .A2(n4379), .ZN(n5689) );
  INV_X1 U5447 ( .A(n5689), .ZN(n4380) );
  OAI21_X1 U5448 ( .B1(n4390), .B2(n4380), .A(n5321), .ZN(n4384) );
  AOI21_X1 U5449 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6352) );
  NAND2_X1 U5450 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6334) );
  NOR2_X1 U5451 ( .A1(n6352), .A2(n6334), .ZN(n6321) );
  NAND2_X1 U5452 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6321), .ZN(n4659)
         );
  NOR2_X1 U5453 ( .A1(n4660), .A2(n4659), .ZN(n5288) );
  NAND2_X1 U5454 ( .A1(n5288), .A2(n4381), .ZN(n4391) );
  INV_X1 U5455 ( .A(n4391), .ZN(n5318) );
  NAND2_X1 U5456 ( .A1(n5318), .A2(n4382), .ZN(n5686) );
  OAI21_X1 U5457 ( .B1(n4390), .B2(n5686), .A(n6353), .ZN(n4383) );
  NAND3_X1 U5458 ( .A1(n5688), .A2(n4384), .A3(n4383), .ZN(n5677) );
  AND2_X1 U5459 ( .A1(n5608), .A2(n5664), .ZN(n4385) );
  NOR2_X1 U5460 ( .A1(n5677), .A2(n4385), .ZN(n5436) );
  NAND2_X1 U5461 ( .A1(n6594), .A2(n5910), .ZN(n4527) );
  NAND2_X1 U5462 ( .A1(n5321), .A2(n4527), .ZN(n6319) );
  INV_X1 U5463 ( .A(n6319), .ZN(n6346) );
  NOR2_X1 U5464 ( .A1(n6353), .A2(n6346), .ZN(n4386) );
  OR2_X1 U5465 ( .A1(n4386), .A2(n4393), .ZN(n4387) );
  NAND2_X1 U5466 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U5467 ( .A1(n5608), .A2(n4394), .ZN(n4388) );
  NAND2_X1 U5468 ( .A1(n5655), .A2(n4388), .ZN(n5626) );
  AND2_X1 U5469 ( .A1(n5608), .A2(n4396), .ZN(n4389) );
  NOR2_X1 U5470 ( .A1(n5626), .A2(n4389), .ZN(n5621) );
  OAI21_X1 U5471 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5691), .A(n5621), 
        .ZN(n5607) );
  NAND2_X1 U5472 ( .A1(n6325), .A2(REIP_REG_30__SCAN_IN), .ZN(n4405) );
  INV_X1 U5473 ( .A(n4405), .ZN(n4399) );
  INV_X1 U5474 ( .A(n4390), .ZN(n4392) );
  NOR2_X1 U5475 ( .A1(n5317), .A2(n4391), .ZN(n5912) );
  NAND3_X1 U5476 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5905), .ZN(n5900) );
  INV_X1 U5477 ( .A(n5900), .ZN(n5693) );
  NAND2_X1 U5478 ( .A1(n4392), .A2(n5693), .ZN(n5675) );
  INV_X1 U5479 ( .A(n4394), .ZN(n4395) );
  INV_X1 U5480 ( .A(n4396), .ZN(n4397) );
  NAND2_X1 U5481 ( .A1(n5631), .A2(n4397), .ZN(n5610) );
  NOR3_X1 U5482 ( .A1(n5610), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6714), 
        .ZN(n4398) );
  AOI211_X1 U5483 ( .C1(n5607), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4399), .B(n4398), .ZN(n4400) );
  NAND2_X1 U5484 ( .A1(n4403), .A2(n4402), .ZN(U2988) );
  NAND2_X1 U5485 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4404)
         );
  OAI211_X1 U5486 ( .C1(n5758), .C2(n6280), .A(n4405), .B(n4404), .ZN(n4406)
         );
  AOI21_X1 U5487 ( .B1(n4407), .B2(n6272), .A(n4406), .ZN(n4410) );
  NAND2_X1 U5488 ( .A1(n4410), .A2(n4409), .ZN(U2956) );
  INV_X1 U5489 ( .A(n4489), .ZN(n4502) );
  OAI22_X1 U5490 ( .A1(n4502), .A2(n5247), .B1(n4495), .B2(n4411), .ZN(n5934)
         );
  INV_X1 U5491 ( .A(n5251), .ZN(n4412) );
  OR2_X1 U5492 ( .A1(n4534), .A2(n4412), .ZN(n4423) );
  AOI21_X1 U5493 ( .B1(n4423), .B2(n6524), .A(READY_N), .ZN(n6615) );
  NOR2_X1 U5494 ( .A1(n5934), .A2(n6615), .ZN(n6488) );
  NOR2_X1 U5495 ( .A1(n6488), .A2(n6510), .ZN(n5941) );
  INV_X1 U5496 ( .A(MORE_REG_SCAN_IN), .ZN(n4421) );
  OR2_X1 U5497 ( .A1(n4489), .A2(n4482), .ZN(n4418) );
  OAI21_X1 U5498 ( .B1(n4495), .B2(n4413), .A(n4489), .ZN(n4417) );
  NAND2_X1 U5499 ( .A1(n4415), .A2(n4414), .ZN(n4416) );
  AND3_X1 U5500 ( .A1(n4418), .A2(n4417), .A3(n4416), .ZN(n6490) );
  INV_X1 U5501 ( .A(n6490), .ZN(n4419) );
  NAND2_X1 U5502 ( .A1(n5941), .A2(n4419), .ZN(n4420) );
  OAI21_X1 U5503 ( .B1(n5941), .B2(n4421), .A(n4420), .ZN(U3471) );
  INV_X1 U5504 ( .A(n6611), .ZN(n4424) );
  NOR2_X1 U5505 ( .A1(n5733), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5263) );
  OAI21_X1 U5506 ( .B1(n5263), .B2(READREQUEST_REG_SCAN_IN), .A(n4424), .ZN(
        n4422) );
  OAI21_X1 U5507 ( .B1(n4424), .B2(n4423), .A(n4422), .ZN(U3474) );
  INV_X1 U5508 ( .A(n4532), .ZN(n4533) );
  AOI211_X1 U5509 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4425), .A(n5263), .B(
        n4533), .ZN(n4426) );
  INV_X1 U5510 ( .A(n4426), .ZN(U2788) );
  NOR2_X1 U5511 ( .A1(n5456), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4427)
         );
  OR2_X1 U5512 ( .A1(n4428), .A2(n4427), .ZN(n5721) );
  NAND2_X1 U5513 ( .A1(n4489), .A2(n4429), .ZN(n4491) );
  INV_X1 U5514 ( .A(n3284), .ZN(n4432) );
  NOR2_X1 U5515 ( .A1(n4648), .A2(n4688), .ZN(n4430) );
  NAND4_X1 U5516 ( .A1(n4432), .A2(n4535), .A3(n4431), .A4(n4430), .ZN(n4433)
         );
  OR2_X2 U5517 ( .A1(n5492), .A2(n4648), .ZN(n5538) );
  INV_X2 U5518 ( .A(n5492), .ZN(n5537) );
  OAI21_X1 U5519 ( .B1(n4437), .B2(n4436), .A(n4435), .ZN(n5276) );
  OR2_X2 U5520 ( .A1(n5492), .A2(n5540), .ZN(n5536) );
  OAI222_X1 U5521 ( .A1(n5721), .A2(n5538), .B1(n5537), .B2(n5271), .C1(n5276), 
        .C2(n5536), .ZN(U2859) );
  NAND2_X1 U5522 ( .A1(n5445), .A2(n6496), .ZN(n4438) );
  NAND2_X1 U5523 ( .A1(n4438), .A2(n4494), .ZN(n4439) );
  NAND2_X1 U5524 ( .A1(n6135), .A2(n4672), .ZN(n6131) );
  NAND2_X1 U5525 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4633) );
  NOR2_X1 U5526 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4633), .ZN(n6159) );
  AOI22_X1 U5527 ( .A1(DATAO_REG_29__SCAN_IN), .A2(n3133), .B1(
        UWORD_REG_13__SCAN_IN), .B2(n6614), .ZN(n4440) );
  OAI21_X1 U5528 ( .B1(n4237), .B2(n6131), .A(n4440), .ZN(U2894) );
  INV_X1 U5529 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6923) );
  AOI22_X1 U5530 ( .A1(DATAO_REG_17__SCAN_IN), .A2(n3133), .B1(n6159), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n4441) );
  OAI21_X1 U5531 ( .B1(n6923), .B2(n6131), .A(n4441), .ZN(U2906) );
  AOI22_X1 U5532 ( .A1(DATAO_REG_24__SCAN_IN), .A2(n3133), .B1(n6159), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n4442) );
  OAI21_X1 U5533 ( .B1(n3840), .B2(n6131), .A(n4442), .ZN(U2899) );
  INV_X1 U5534 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6890) );
  AOI22_X1 U5535 ( .A1(DATAO_REG_18__SCAN_IN), .A2(n3133), .B1(n6159), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n4443) );
  OAI21_X1 U5536 ( .B1(n6890), .B2(n6131), .A(n4443), .ZN(U2905) );
  INV_X1 U5537 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4547) );
  AOI22_X1 U5538 ( .A1(DATAO_REG_28__SCAN_IN), .A2(n3133), .B1(n6614), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n4444) );
  OAI21_X1 U5539 ( .B1(n4547), .B2(n6131), .A(n4444), .ZN(U2895) );
  INV_X1 U5540 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4551) );
  AOI22_X1 U5541 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6159), .B1(n3133), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4445) );
  OAI21_X1 U5542 ( .B1(n4551), .B2(n6131), .A(n4445), .ZN(U2897) );
  INV_X1 U5543 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6765) );
  AOI22_X1 U5544 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6159), .B1(n3133), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4446) );
  OAI21_X1 U5545 ( .B1(n6765), .B2(n6131), .A(n4446), .ZN(U2900) );
  INV_X1 U5546 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6919) );
  AOI22_X1 U5547 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6159), .B1(n3133), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4447) );
  OAI21_X1 U5548 ( .B1(n6919), .B2(n6131), .A(n4447), .ZN(U2896) );
  INV_X1 U5549 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4449) );
  AOI22_X1 U5550 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6614), .B1(n3133), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4448) );
  OAI21_X1 U5551 ( .B1(n4449), .B2(n6131), .A(n4448), .ZN(U2904) );
  INV_X1 U5552 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4451) );
  AOI22_X1 U5553 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6614), .B1(n3133), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4450) );
  OAI21_X1 U5554 ( .B1(n4451), .B2(n6131), .A(n4450), .ZN(U2907) );
  INV_X1 U5555 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4453) );
  AOI22_X1 U5556 ( .A1(n6614), .A2(UWORD_REG_9__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4452) );
  OAI21_X1 U5557 ( .B1(n4453), .B2(n6131), .A(n4452), .ZN(U2898) );
  AOI22_X1 U5558 ( .A1(n6614), .A2(UWORD_REG_6__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4454) );
  OAI21_X1 U5559 ( .B1(n4455), .B2(n6131), .A(n4454), .ZN(U2901) );
  INV_X1 U5560 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4457) );
  AOI22_X1 U5561 ( .A1(n6614), .A2(UWORD_REG_5__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4456) );
  OAI21_X1 U5562 ( .B1(n4457), .B2(n6131), .A(n4456), .ZN(U2902) );
  INV_X1 U5563 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4544) );
  AOI22_X1 U5564 ( .A1(n6614), .A2(UWORD_REG_14__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4458) );
  OAI21_X1 U5565 ( .B1(n4544), .B2(n6131), .A(n4458), .ZN(U2893) );
  OR2_X1 U5566 ( .A1(n4460), .A2(n4459), .ZN(n4461) );
  NAND2_X1 U5567 ( .A1(n4462), .A2(n4461), .ZN(n6285) );
  INV_X1 U5568 ( .A(n5538), .ZN(n5493) );
  XNOR2_X1 U5569 ( .A(n4463), .B(n5455), .ZN(n4529) );
  AOI22_X1 U5570 ( .A1(n5493), .A2(n4529), .B1(n5492), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4464) );
  OAI21_X1 U5571 ( .B1(n5536), .B2(n6285), .A(n4464), .ZN(U2858) );
  XNOR2_X1 U5572 ( .A(n4465), .B(n6594), .ZN(n5723) );
  NAND2_X1 U5573 ( .A1(n6272), .A2(n5723), .ZN(n4470) );
  NAND2_X1 U5574 ( .A1(n4466), .A2(n5588), .ZN(n4468) );
  NAND2_X1 U5575 ( .A1(n6325), .A2(REIP_REG_0__SCAN_IN), .ZN(n5720) );
  INV_X1 U5576 ( .A(n5720), .ZN(n4467) );
  AOI21_X1 U5577 ( .B1(PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4468), .A(n4467), 
        .ZN(n4469) );
  OAI211_X1 U5578 ( .C1(n5276), .C2(n6286), .A(n4470), .B(n4469), .ZN(U2986)
         );
  NAND2_X1 U5579 ( .A1(n4572), .A2(n4537), .ZN(n4472) );
  NOR2_X1 U5580 ( .A1(n5929), .A2(n4472), .ZN(n4475) );
  INV_X1 U5581 ( .A(n4473), .ZN(n4474) );
  AND2_X1 U5582 ( .A1(n4475), .A2(n4474), .ZN(n5442) );
  INV_X1 U5583 ( .A(n5445), .ZN(n6476) );
  NAND2_X1 U5584 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4476) );
  INV_X1 U5585 ( .A(n4476), .ZN(n4477) );
  MUX2_X1 U5586 ( .A(n4477), .B(n4476), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4481) );
  AOI21_X1 U5587 ( .B1(n4508), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4479) );
  NOR2_X1 U5588 ( .A1(n3358), .A2(n4479), .ZN(n4490) );
  AOI22_X1 U5589 ( .A1(n6476), .A2(n4481), .B1(n4480), .B2(n4490), .ZN(n4488)
         );
  NAND2_X1 U5590 ( .A1(n4482), .A2(n4565), .ZN(n4516) );
  INV_X1 U5591 ( .A(n4483), .ZN(n4587) );
  INV_X1 U5592 ( .A(n4484), .ZN(n4485) );
  MUX2_X1 U5593 ( .A(n4485), .B(n4506), .S(n4508), .Z(n4486) );
  NAND3_X1 U5594 ( .A1(n4516), .A2(n4587), .A3(n4486), .ZN(n4487) );
  OAI211_X1 U5595 ( .C1(n5077), .C2(n5442), .A(n4488), .B(n4487), .ZN(n4586)
         );
  INV_X1 U5596 ( .A(n6600), .ZN(n5928) );
  AOI22_X1 U5597 ( .A1(n4586), .A2(n5928), .B1(n4490), .B2(n6592), .ZN(n4505)
         );
  INV_X1 U5598 ( .A(n4565), .ZN(n4503) );
  INV_X1 U5599 ( .A(n4491), .ZN(n4501) );
  OAI21_X1 U5600 ( .B1(n5445), .B2(READY_N), .A(n4492), .ZN(n4493) );
  OAI211_X1 U5601 ( .C1(n4495), .C2(n4494), .A(n4502), .B(n4493), .ZN(n4499)
         );
  NAND2_X1 U5602 ( .A1(n5929), .A2(n4563), .ZN(n4496) );
  NAND4_X1 U5603 ( .A1(n4499), .A2(n4498), .A3(n4497), .A4(n4496), .ZN(n4500)
         );
  INV_X1 U5604 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5940) );
  OR2_X1 U5605 ( .A1(n3350), .A2(n4633), .ZN(n6589) );
  OAI22_X1 U5606 ( .A1(n6510), .A2(n6479), .B1(n5940), .B2(n6589), .ZN(n4504)
         );
  INV_X1 U5607 ( .A(n4504), .ZN(n5932) );
  NAND2_X1 U5608 ( .A1(n3350), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U5609 ( .A1(n5932), .A2(n6590), .ZN(n6598) );
  MUX2_X1 U5610 ( .A(n4506), .B(n4505), .S(n6598), .Z(n4507) );
  INV_X1 U5611 ( .A(n4507), .ZN(U3456) );
  INV_X1 U5612 ( .A(n4508), .ZN(n4518) );
  INV_X1 U5613 ( .A(n6598), .ZN(n4522) );
  AOI21_X1 U5614 ( .B1(n6592), .B2(n4518), .A(n4522), .ZN(n4524) );
  INV_X1 U5615 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4584) );
  XNOR2_X1 U5616 ( .A(n4508), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4515)
         );
  XNOR2_X1 U5617 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4510) );
  OAI22_X1 U5618 ( .A1(n5445), .A2(n4510), .B1(n4509), .B2(n4515), .ZN(n4514)
         );
  NOR2_X1 U5619 ( .A1(n4512), .A2(n5442), .ZN(n4513) );
  AOI211_X1 U5620 ( .C1(n4516), .C2(n4515), .A(n4514), .B(n4513), .ZN(n4585)
         );
  INV_X1 U5621 ( .A(n4585), .ZN(n4521) );
  INV_X1 U5622 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5613) );
  AOI22_X1 U5623 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5613), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4657), .ZN(n5448) );
  NOR3_X1 U5624 ( .A1(n6501), .A2(n6594), .A3(n5448), .ZN(n4520) );
  INV_X1 U5625 ( .A(n6592), .ZN(n4517) );
  NOR3_X1 U5626 ( .A1(n4518), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4517), 
        .ZN(n4519) );
  AOI211_X1 U5627 ( .C1(n4521), .C2(n5928), .A(n4520), .B(n4519), .ZN(n4523)
         );
  OAI22_X1 U5628 ( .A1(n4524), .A2(n4584), .B1(n4523), .B2(n4522), .ZN(U3459)
         );
  XNOR2_X1 U5629 ( .A(n4525), .B(n4526), .ZN(n6279) );
  NAND3_X1 U5630 ( .A1(n5608), .A2(n4527), .A3(n4657), .ZN(n4531) );
  OAI21_X1 U5631 ( .B1(n5911), .B2(n6353), .A(n6594), .ZN(n5728) );
  AOI21_X1 U5632 ( .B1(n5724), .B2(n5728), .A(n4657), .ZN(n4528) );
  INV_X1 U5633 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6602) );
  NOR2_X1 U5634 ( .A1(n6349), .A2(n6602), .ZN(n6282) );
  AOI211_X1 U5635 ( .C1(n6323), .C2(n4529), .A(n4528), .B(n6282), .ZN(n4530)
         );
  OAI211_X1 U5636 ( .C1(n6279), .C2(n5913), .A(n4531), .B(n4530), .ZN(U3017)
         );
  INV_X1 U5637 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6149) );
  INV_X1 U5638 ( .A(READY_N), .ZN(n6613) );
  NAND2_X1 U5639 ( .A1(n6202), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U5640 ( .A1(n4535), .A2(n6613), .ZN(n4536) );
  NOR2_X1 U5641 ( .A1(n4537), .A2(n4536), .ZN(n4538) );
  NAND2_X1 U5642 ( .A1(n6203), .A2(DATAI_8_), .ZN(n4541) );
  OAI211_X1 U5643 ( .C1(n6149), .C2(n6166), .A(n4540), .B(n4541), .ZN(U2947)
         );
  NAND2_X1 U5644 ( .A1(n6202), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4542) );
  OAI211_X1 U5645 ( .C1(n3840), .C2(n6166), .A(n4542), .B(n4541), .ZN(U2932)
         );
  AOI22_X1 U5646 ( .A1(n6202), .A2(UWORD_REG_14__SCAN_IN), .B1(n6203), .B2(
        DATAI_14_), .ZN(n4543) );
  OAI21_X1 U5647 ( .B1(n4544), .B2(n6166), .A(n4543), .ZN(U2938) );
  INV_X1 U5648 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6137) );
  AOI22_X1 U5649 ( .A1(n6202), .A2(LWORD_REG_15__SCAN_IN), .B1(n6203), .B2(
        DATAI_15_), .ZN(n4545) );
  OAI21_X1 U5650 ( .B1(n6137), .B2(n6166), .A(n4545), .ZN(U2954) );
  AOI22_X1 U5651 ( .A1(n6202), .A2(UWORD_REG_12__SCAN_IN), .B1(n6203), .B2(
        DATAI_12_), .ZN(n4546) );
  OAI21_X1 U5652 ( .B1(n4547), .B2(n6166), .A(n4546), .ZN(U2936) );
  AOI22_X1 U5653 ( .A1(n6202), .A2(UWORD_REG_13__SCAN_IN), .B1(n6203), .B2(
        DATAI_13_), .ZN(n4548) );
  OAI21_X1 U5654 ( .B1(n4237), .B2(n6166), .A(n4548), .ZN(U2937) );
  AOI22_X1 U5655 ( .A1(n6202), .A2(UWORD_REG_11__SCAN_IN), .B1(n6203), .B2(
        DATAI_11_), .ZN(n4549) );
  OAI21_X1 U5656 ( .B1(n6919), .B2(n6166), .A(n4549), .ZN(U2935) );
  INV_X1 U5657 ( .A(DATAI_10_), .ZN(n5245) );
  NOR2_X1 U5658 ( .A1(n6194), .A2(n5245), .ZN(n4552) );
  AOI21_X1 U5659 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6202), .A(n4552), .ZN(
        n4550) );
  OAI21_X1 U5660 ( .B1(n4551), .B2(n6166), .A(n4550), .ZN(U2934) );
  INV_X1 U5661 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6875) );
  AOI21_X1 U5662 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6202), .A(n4552), .ZN(
        n4553) );
  OAI21_X1 U5663 ( .B1(n6875), .B2(n6166), .A(n4553), .ZN(U2949) );
  INV_X1 U5664 ( .A(n4605), .ZN(n4554) );
  OAI21_X1 U5665 ( .B1(n4556), .B2(n4555), .A(n4554), .ZN(n5261) );
  INV_X1 U5666 ( .A(n5261), .ZN(n6274) );
  INV_X1 U5667 ( .A(n5536), .ZN(n5505) );
  NAND2_X1 U5668 ( .A1(n4558), .A2(n4557), .ZN(n4559) );
  NAND2_X1 U5669 ( .A1(n4607), .A2(n4559), .ZN(n6350) );
  OAI22_X1 U5670 ( .A1(n6350), .A2(n5538), .B1(n5537), .B2(n4560), .ZN(n4561)
         );
  AOI21_X1 U5671 ( .B1(n6274), .B2(n5505), .A(n4561), .ZN(n4562) );
  INV_X1 U5672 ( .A(n4562), .ZN(U2857) );
  NAND3_X1 U5673 ( .A1(n5929), .A2(n4569), .A3(n4563), .ZN(n4564) );
  OAI21_X1 U5674 ( .B1(n4566), .B2(n4565), .A(n4564), .ZN(n4567) );
  INV_X1 U5675 ( .A(n4567), .ZN(n4568) );
  NAND4_X1 U5676 ( .A1(n5540), .A2(n4570), .A3(n4569), .A4(n3303), .ZN(n4571)
         );
  NOR2_X1 U5677 ( .A1(n4572), .A2(n4571), .ZN(n4573) );
  INV_X1 U5678 ( .A(n4574), .ZN(n4575) );
  NAND2_X2 U5679 ( .A1(n5539), .A2(n4575), .ZN(n5855) );
  INV_X1 U5680 ( .A(n5373), .ZN(n4576) );
  INV_X1 U5681 ( .A(DATAI_1_), .ZN(n6179) );
  INV_X1 U5682 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6704) );
  OAI222_X1 U5683 ( .A1(n6285), .A2(n5855), .B1(n5246), .B2(n6179), .C1(n5539), 
        .C2(n6704), .ZN(U2890) );
  INV_X1 U5684 ( .A(DATAI_2_), .ZN(n6181) );
  INV_X1 U5685 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6161) );
  OAI222_X1 U5686 ( .A1(n5261), .A2(n5855), .B1(n5246), .B2(n6181), .C1(n5539), 
        .C2(n6161), .ZN(U2889) );
  INV_X1 U5687 ( .A(DATAI_0_), .ZN(n6177) );
  INV_X1 U5688 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6165) );
  OAI222_X1 U5689 ( .A1(n5276), .A2(n5855), .B1(n5246), .B2(n6177), .C1(n5539), 
        .C2(n6165), .ZN(U2891) );
  AND2_X1 U5690 ( .A1(n4605), .A2(n4604), .ZN(n4578) );
  NOR2_X1 U5691 ( .A1(n4578), .A2(n4577), .ZN(n4579) );
  OR2_X1 U5692 ( .A1(n4613), .A2(n4579), .ZN(n6260) );
  INV_X1 U5693 ( .A(DATAI_4_), .ZN(n6186) );
  INV_X1 U5694 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6698) );
  OAI222_X1 U5695 ( .A1(n6260), .A2(n5855), .B1(n5246), .B2(n6186), .C1(n5539), 
        .C2(n6698), .ZN(U2887) );
  CLKBUF_X1 U5696 ( .A(n4580), .Z(n4615) );
  OR2_X1 U5697 ( .A1(n4582), .A2(n4581), .ZN(n4583) );
  NAND2_X1 U5698 ( .A1(n4615), .A2(n4583), .ZN(n6330) );
  INV_X1 U5699 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6841) );
  OAI222_X1 U5700 ( .A1(n6330), .A2(n5538), .B1(n5537), .B2(n6841), .C1(n6260), 
        .C2(n5536), .ZN(U2855) );
  MUX2_X1 U5701 ( .A(n4585), .B(n4584), .S(n6479), .Z(n6483) );
  MUX2_X1 U5702 ( .A(n4586), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6479), 
        .Z(n6486) );
  NAND2_X1 U5703 ( .A1(n6501), .A2(n6486), .ZN(n4588) );
  NAND2_X1 U5704 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5940), .ZN(n4594) );
  OAI22_X1 U5705 ( .A1(n6483), .A2(n4588), .B1(n4594), .B2(n4587), .ZN(n6494)
         );
  INV_X1 U5706 ( .A(n4589), .ZN(n4590) );
  NAND2_X1 U5707 ( .A1(n6494), .A2(n4590), .ZN(n4632) );
  INV_X1 U5708 ( .A(n4967), .ZN(n4643) );
  OR2_X1 U5709 ( .A1(n4591), .A2(n4643), .ZN(n4593) );
  XNOR2_X1 U5710 ( .A(n4593), .B(n4592), .ZN(n5267) );
  INV_X1 U5711 ( .A(n5267), .ZN(n5930) );
  AOI22_X1 U5712 ( .A1(n6479), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(n5929), .B2(n5930), .ZN(n4595) );
  OAI22_X1 U5713 ( .A1(n4595), .A2(STATE2_REG_1__SCAN_IN), .B1(n4592), .B2(
        n4594), .ZN(n6493) );
  INV_X1 U5714 ( .A(n6493), .ZN(n4596) );
  NAND3_X1 U5715 ( .A1(n4632), .A2(n4596), .A3(n5940), .ZN(n4599) );
  INV_X1 U5716 ( .A(n6589), .ZN(n4598) );
  AOI21_X1 U5717 ( .B1(n4599), .B2(n4598), .A(n4766), .ZN(n6362) );
  NAND2_X1 U5718 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n3296), .ZN(n4628) );
  AOI211_X1 U5719 ( .C1(n4794), .C2(n5939), .A(n5733), .B(n5731), .ZN(n4601)
         );
  AOI21_X1 U5720 ( .B1(n4628), .B2(n5447), .A(n4601), .ZN(n4603) );
  NAND2_X1 U5721 ( .A1(n6362), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4602) );
  OAI21_X1 U5722 ( .B1(n6362), .B2(n4603), .A(n4602), .ZN(U3464) );
  XOR2_X1 U5723 ( .A(n4605), .B(n4604), .Z(n6265) );
  XNOR2_X1 U5724 ( .A(n4607), .B(n4606), .ZN(n6338) );
  OAI22_X1 U5725 ( .A1(n6338), .A2(n5538), .B1(n5537), .B2(n6695), .ZN(n4608)
         );
  AOI21_X1 U5726 ( .B1(n6265), .B2(n5505), .A(n4608), .ZN(n4609) );
  INV_X1 U5727 ( .A(n4609), .ZN(U2856) );
  INV_X1 U5728 ( .A(n6265), .ZN(n4610) );
  INV_X1 U5729 ( .A(DATAI_3_), .ZN(n6183) );
  INV_X1 U5730 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6158) );
  OAI222_X1 U5731 ( .A1(n4610), .A2(n5855), .B1(n5246), .B2(n6183), .C1(n5539), 
        .C2(n6158), .ZN(U2888) );
  INV_X1 U5732 ( .A(n4611), .ZN(n4612) );
  XNOR2_X1 U5733 ( .A(n4613), .B(n4612), .ZN(n6248) );
  INV_X1 U5734 ( .A(n6248), .ZN(n4625) );
  NAND2_X1 U5735 ( .A1(n4615), .A2(n4614), .ZN(n4616) );
  AND2_X1 U5736 ( .A1(n4621), .A2(n4616), .ZN(n6322) );
  AOI22_X1 U5737 ( .A1(n5493), .A2(n6322), .B1(EBX_REG_5__SCAN_IN), .B2(n5492), 
        .ZN(n4617) );
  OAI21_X1 U5738 ( .B1(n4625), .B2(n5536), .A(n4617), .ZN(U2854) );
  XNOR2_X1 U5739 ( .A(n4619), .B(n4618), .ZN(n6243) );
  NAND2_X1 U5740 ( .A1(n4621), .A2(n4620), .ZN(n4622) );
  NAND2_X1 U5741 ( .A1(n5034), .A2(n4622), .ZN(n6075) );
  OAI22_X1 U5742 ( .A1(n6075), .A2(n5538), .B1(n5537), .B2(n6074), .ZN(n4623)
         );
  INV_X1 U5743 ( .A(n4623), .ZN(n4624) );
  OAI21_X1 U5744 ( .B1(n6243), .B2(n5536), .A(n4624), .ZN(U2853) );
  INV_X1 U5745 ( .A(DATAI_5_), .ZN(n6188) );
  INV_X1 U5746 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6155) );
  OAI222_X1 U5747 ( .A1(n5855), .A2(n4625), .B1(n5246), .B2(n6188), .C1(n5539), 
        .C2(n6155), .ZN(U2886) );
  INV_X1 U5748 ( .A(n6362), .ZN(n4637) );
  INV_X1 U5749 ( .A(n4627), .ZN(n4793) );
  NAND3_X1 U5750 ( .A1(n5730), .A2(n4794), .A3(n4793), .ZN(n4698) );
  NAND2_X1 U5751 ( .A1(n4762), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4903) );
  AND2_X1 U5752 ( .A1(n4903), .A2(n5039), .ZN(n5132) );
  NAND3_X1 U5753 ( .A1(n5731), .A2(n5730), .A3(n4627), .ZN(n4966) );
  AOI21_X1 U5754 ( .B1(n5132), .B2(n4966), .A(n5733), .ZN(n4630) );
  NAND2_X1 U5755 ( .A1(n6371), .A2(n5939), .ZN(n6373) );
  INV_X1 U5756 ( .A(n4628), .ZN(n5732) );
  OAI22_X1 U5757 ( .A1(n4110), .A2(n6373), .B1(n5077), .B2(n5732), .ZN(n4629)
         );
  OAI21_X1 U5758 ( .B1(n4630), .B2(n4629), .A(n4637), .ZN(n4631) );
  OAI21_X1 U5759 ( .B1(n4637), .B2(n6485), .A(n4631), .ZN(U3462) );
  INV_X1 U5760 ( .A(n4632), .ZN(n4634) );
  NOR3_X1 U5761 ( .A1(n4634), .A2(n4633), .A3(n6493), .ZN(n6503) );
  OAI22_X1 U5762 ( .A1(n3142), .A2(n5733), .B1(n3507), .B2(n5732), .ZN(n4635)
         );
  OAI21_X1 U5763 ( .B1(n6503), .B2(n4635), .A(n4637), .ZN(n4636) );
  OAI21_X1 U5764 ( .B1(n4637), .B2(n5179), .A(n4636), .ZN(U3465) );
  NOR2_X1 U5765 ( .A1(n4793), .A2(n4795), .ZN(n4638) );
  NAND2_X1 U5766 ( .A1(n5730), .A2(n4638), .ZN(n5188) );
  INV_X1 U5767 ( .A(n5188), .ZN(n4639) );
  NAND2_X1 U5768 ( .A1(n6273), .A2(DATAI_23_), .ZN(n6418) );
  NAND3_X1 U5769 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6485), .A3(n4790), .ZN(n5185) );
  OR2_X1 U5770 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5185), .ZN(n4998)
         );
  NOR2_X1 U5771 ( .A1(n4650), .A2(n6497), .ZN(n4767) );
  INV_X1 U5772 ( .A(n4640), .ZN(n4701) );
  INV_X1 U5773 ( .A(n5083), .ZN(n6365) );
  NOR2_X1 U5774 ( .A1(n4701), .A2(n6365), .ZN(n4741) );
  OAI21_X1 U5775 ( .B1(n4741), .B2(n6497), .A(n4766), .ZN(n4737) );
  AOI211_X1 U5776 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4998), .A(n4767), .B(
        n4737), .ZN(n4645) );
  NAND2_X1 U5777 ( .A1(n4110), .A2(n4845), .ZN(n4641) );
  INV_X1 U5778 ( .A(n6373), .ZN(n4735) );
  OR2_X1 U5779 ( .A1(n5188), .A2(n5939), .ZN(n4642) );
  OR2_X1 U5780 ( .A1(n4512), .A2(n5447), .ZN(n4649) );
  NAND2_X1 U5781 ( .A1(n4899), .A2(n4643), .ZN(n5178) );
  OAI211_X1 U5782 ( .C1(n4646), .C2(n4735), .A(n5184), .B(n5178), .ZN(n4644)
         );
  NAND2_X1 U5783 ( .A1(n4645), .A2(n4644), .ZN(n4996) );
  NAND2_X1 U5784 ( .A1(n4996), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U5785 ( .A1(n6273), .A2(DATAI_31_), .ZN(n6437) );
  INV_X1 U5786 ( .A(n6437), .ZN(n6414) );
  NAND2_X1 U5787 ( .A1(n4829), .A2(n4648), .ZN(n5108) );
  NOR2_X1 U5788 ( .A1(n4649), .A2(n5733), .ZN(n4706) );
  AND2_X1 U5789 ( .A1(n4650), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6366) );
  AOI22_X1 U5790 ( .A1(n4706), .A2(n5077), .B1(n6366), .B2(n4741), .ZN(n4997)
         );
  INV_X1 U5791 ( .A(DATAI_7_), .ZN(n6191) );
  OAI22_X1 U5792 ( .A1(n5108), .A2(n4998), .B1(n4997), .B2(n5107), .ZN(n4651)
         );
  AOI21_X1 U5793 ( .B1(n6414), .B2(n5169), .A(n4651), .ZN(n4652) );
  OAI211_X1 U5794 ( .C1(n5222), .C2(n6418), .A(n4653), .B(n4652), .ZN(U3059)
         );
  OAI21_X1 U5795 ( .B1(n4656), .B2(n4655), .A(n4654), .ZN(n6238) );
  NOR2_X1 U5796 ( .A1(n6351), .A2(n6075), .ZN(n4663) );
  NOR2_X1 U5798 ( .A1(n6360), .A2(n4657), .ZN(n4658) );
  OAI21_X1 U5799 ( .B1(n5690), .B2(n4658), .A(n5688), .ZN(n6347) );
  AOI21_X1 U5800 ( .B1(n4659), .B2(n5608), .A(n6347), .ZN(n6329) );
  AOI21_X1 U5801 ( .B1(n6346), .B2(n4658), .A(n6353), .ZN(n6333) );
  OAI33_X1 U5802 ( .A1(1'b0), .A2(n6329), .A3(n4660), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4659), .B3(n6333), .ZN(n4662) );
  AOI211_X1 U5803 ( .C1(n6325), .C2(REIP_REG_6__SCAN_IN), .A(n4663), .B(n4662), 
        .ZN(n4664) );
  OAI21_X1 U5804 ( .B1(n5913), .B2(n6238), .A(n4664), .ZN(U3012) );
  NAND3_X1 U5805 ( .A1(n5730), .A2(n4793), .A3(n4795), .ZN(n4666) );
  INV_X1 U5806 ( .A(n6418), .ZN(n6429) );
  INV_X1 U5807 ( .A(n3507), .ZN(n6475) );
  NAND2_X1 U5808 ( .A1(n6368), .A2(n6475), .ZN(n4838) );
  INV_X1 U5809 ( .A(n5447), .ZN(n6115) );
  OR2_X1 U5810 ( .A1(n6115), .A2(n4512), .ZN(n4968) );
  OAI21_X1 U5811 ( .B1(n4838), .B2(n4968), .A(n5027), .ZN(n4667) );
  AOI22_X1 U5812 ( .A1(n4667), .A2(n6371), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4760), .ZN(n5026) );
  OAI22_X1 U5813 ( .A1(n5108), .A2(n5027), .B1(n5026), .B2(n5107), .ZN(n4665)
         );
  AOI21_X1 U5814 ( .B1(n6429), .B2(n5029), .A(n4665), .ZN(n4671) );
  AOI21_X1 U5815 ( .B1(n4666), .B2(n6273), .A(n4735), .ZN(n4668) );
  OR2_X1 U5816 ( .A1(n4668), .A2(n4667), .ZN(n4669) );
  OAI211_X1 U5817 ( .C1(n6371), .C2(n4760), .A(n4669), .B(n4973), .ZN(n5030)
         );
  NAND2_X1 U5818 ( .A1(n5030), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4670)
         );
  OAI211_X1 U5819 ( .C1(n5033), .C2(n6437), .A(n4671), .B(n4670), .ZN(U3147)
         );
  NAND2_X1 U5820 ( .A1(n6273), .A2(DATAI_16_), .ZN(n6382) );
  NAND2_X1 U5821 ( .A1(n4996), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4675) );
  NAND2_X1 U5822 ( .A1(n6273), .A2(DATAI_24_), .ZN(n6443) );
  INV_X1 U5823 ( .A(n6443), .ZN(n6379) );
  NAND2_X1 U5824 ( .A1(n4829), .A2(n4672), .ZN(n5086) );
  OAI22_X1 U5825 ( .A1(n5086), .A2(n4998), .B1(n4997), .B2(n5085), .ZN(n4673)
         );
  AOI21_X1 U5826 ( .B1(n6379), .B2(n5169), .A(n4673), .ZN(n4674) );
  OAI211_X1 U5827 ( .C1(n5222), .C2(n6382), .A(n4675), .B(n4674), .ZN(U3052)
         );
  NAND2_X1 U5828 ( .A1(n6273), .A2(DATAI_19_), .ZN(n6396) );
  NAND2_X1 U5829 ( .A1(n4996), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4679) );
  NAND2_X1 U5830 ( .A1(n6273), .A2(DATAI_27_), .ZN(n6455) );
  INV_X1 U5831 ( .A(n6455), .ZN(n6393) );
  NAND2_X1 U5832 ( .A1(n4829), .A2(n4676), .ZN(n5113) );
  OAI22_X1 U5833 ( .A1(n5113), .A2(n4998), .B1(n4997), .B2(n5112), .ZN(n4677)
         );
  AOI21_X1 U5834 ( .B1(n6393), .B2(n5169), .A(n4677), .ZN(n4678) );
  OAI211_X1 U5835 ( .C1(n5222), .C2(n6396), .A(n4679), .B(n4678), .ZN(U3055)
         );
  NAND2_X1 U5836 ( .A1(n6273), .A2(DATAI_18_), .ZN(n6392) );
  NAND2_X1 U5837 ( .A1(n4996), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4683) );
  NAND2_X1 U5838 ( .A1(n6273), .A2(DATAI_26_), .ZN(n6449) );
  INV_X1 U5839 ( .A(n6449), .ZN(n6389) );
  NAND2_X1 U5840 ( .A1(n4829), .A2(n4680), .ZN(n5091) );
  OAI22_X1 U5841 ( .A1(n5091), .A2(n4998), .B1(n4997), .B2(n5090), .ZN(n4681)
         );
  AOI21_X1 U5842 ( .B1(n6389), .B2(n5169), .A(n4681), .ZN(n4682) );
  OAI211_X1 U5843 ( .C1(n5222), .C2(n6392), .A(n4683), .B(n4682), .ZN(U3054)
         );
  NAND2_X1 U5844 ( .A1(n6273), .A2(DATAI_21_), .ZN(n6404) );
  NAND2_X1 U5845 ( .A1(n4996), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4687) );
  NAND2_X1 U5846 ( .A1(n6273), .A2(DATAI_29_), .ZN(n6472) );
  INV_X1 U5847 ( .A(n6472), .ZN(n6401) );
  NAND2_X1 U5848 ( .A1(n4829), .A2(n4684), .ZN(n5126) );
  OAI22_X1 U5849 ( .A1(n5126), .A2(n4998), .B1(n4997), .B2(n5123), .ZN(n4685)
         );
  AOI21_X1 U5850 ( .B1(n6401), .B2(n5169), .A(n4685), .ZN(n4686) );
  OAI211_X1 U5851 ( .C1(n5222), .C2(n6404), .A(n4687), .B(n4686), .ZN(U3057)
         );
  NAND2_X1 U5852 ( .A1(n6273), .A2(DATAI_20_), .ZN(n6400) );
  NAND2_X1 U5853 ( .A1(n4996), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4691) );
  NAND2_X1 U5854 ( .A1(n6273), .A2(DATAI_28_), .ZN(n6461) );
  INV_X1 U5855 ( .A(n6461), .ZN(n6397) );
  NAND2_X1 U5856 ( .A1(n4829), .A2(n4688), .ZN(n5118) );
  OAI22_X1 U5857 ( .A1(n5118), .A2(n4998), .B1(n4997), .B2(n5117), .ZN(n4689)
         );
  AOI21_X1 U5858 ( .B1(n6397), .B2(n5169), .A(n4689), .ZN(n4690) );
  OAI211_X1 U5859 ( .C1(n5222), .C2(n6400), .A(n4691), .B(n4690), .ZN(U3056)
         );
  INV_X1 U5860 ( .A(n6400), .ZN(n6456) );
  OAI22_X1 U5861 ( .A1(n5118), .A2(n5027), .B1(n5026), .B2(n5117), .ZN(n4692)
         );
  AOI21_X1 U5862 ( .B1(n6456), .B2(n5029), .A(n4692), .ZN(n4694) );
  NAND2_X1 U5863 ( .A1(n5030), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4693)
         );
  OAI211_X1 U5864 ( .C1(n5033), .C2(n6461), .A(n4694), .B(n4693), .ZN(U3144)
         );
  INV_X1 U5865 ( .A(n6404), .ZN(n6462) );
  OAI22_X1 U5866 ( .A1(n5126), .A2(n5027), .B1(n5026), .B2(n5123), .ZN(n4695)
         );
  AOI21_X1 U5867 ( .B1(n6462), .B2(n5029), .A(n4695), .ZN(n4697) );
  NAND2_X1 U5868 ( .A1(n5030), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4696)
         );
  OAI211_X1 U5869 ( .C1(n5033), .C2(n6472), .A(n4697), .B(n4696), .ZN(U3145)
         );
  NOR2_X2 U5870 ( .A1(n4698), .A2(n4845), .ZN(n5020) );
  INV_X1 U5871 ( .A(n5020), .ZN(n4699) );
  AOI21_X1 U5872 ( .B1(n4699), .B2(n5046), .A(n5939), .ZN(n4700) );
  AOI211_X1 U5873 ( .C1(n4899), .C2(n4967), .A(n5733), .B(n4700), .ZN(n4703)
         );
  NOR3_X1 U5874 ( .A1(n5075), .A2(n6485), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4902) );
  INV_X1 U5875 ( .A(n4902), .ZN(n4904) );
  NOR2_X1 U5876 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4904), .ZN(n4704)
         );
  INV_X1 U5877 ( .A(n4767), .ZN(n6375) );
  NAND2_X1 U5878 ( .A1(n4701), .A2(n5083), .ZN(n4800) );
  AOI21_X1 U5879 ( .B1(n4800), .B2(STATE2_REG_2__SCAN_IN), .A(n4830), .ZN(
        n4791) );
  OAI211_X1 U5880 ( .C1(n3296), .C2(n4704), .A(n6375), .B(n4791), .ZN(n4702)
         );
  NAND2_X1 U5881 ( .A1(n5016), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4709)
         );
  INV_X1 U5882 ( .A(n4704), .ZN(n5018) );
  INV_X1 U5883 ( .A(n4800), .ZN(n4705) );
  AOI22_X1 U5884 ( .A1(n4706), .A2(n6368), .B1(n6366), .B2(n4705), .ZN(n5017)
         );
  OAI22_X1 U5885 ( .A1(n5108), .A2(n5018), .B1(n5017), .B2(n5107), .ZN(n4707)
         );
  AOI21_X1 U5886 ( .B1(n6429), .B2(n5020), .A(n4707), .ZN(n4708) );
  OAI211_X1 U5887 ( .C1(n5046), .C2(n6437), .A(n4709), .B(n4708), .ZN(U3123)
         );
  INV_X1 U5888 ( .A(n6382), .ZN(n6438) );
  OAI22_X1 U5889 ( .A1(n5086), .A2(n5027), .B1(n5026), .B2(n5085), .ZN(n4710)
         );
  AOI21_X1 U5890 ( .B1(n6438), .B2(n5029), .A(n4710), .ZN(n4712) );
  NAND2_X1 U5891 ( .A1(n5030), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4711)
         );
  OAI211_X1 U5892 ( .C1(n5033), .C2(n6443), .A(n4712), .B(n4711), .ZN(U3140)
         );
  INV_X1 U5893 ( .A(n6392), .ZN(n6444) );
  OAI22_X1 U5894 ( .A1(n5091), .A2(n5027), .B1(n5026), .B2(n5090), .ZN(n4713)
         );
  AOI21_X1 U5895 ( .B1(n6444), .B2(n5029), .A(n4713), .ZN(n4715) );
  NAND2_X1 U5896 ( .A1(n5030), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4714)
         );
  OAI211_X1 U5897 ( .C1(n5033), .C2(n6449), .A(n4715), .B(n4714), .ZN(U3142)
         );
  INV_X1 U5898 ( .A(n6396), .ZN(n6450) );
  OAI22_X1 U5899 ( .A1(n5113), .A2(n5027), .B1(n5026), .B2(n5112), .ZN(n4716)
         );
  AOI21_X1 U5900 ( .B1(n6450), .B2(n5029), .A(n4716), .ZN(n4718) );
  NAND2_X1 U5901 ( .A1(n5030), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4717)
         );
  OAI211_X1 U5902 ( .C1(n5033), .C2(n6455), .A(n4718), .B(n4717), .ZN(U3143)
         );
  NAND2_X1 U5903 ( .A1(n5016), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4721)
         );
  OAI22_X1 U5904 ( .A1(n5126), .A2(n5018), .B1(n5017), .B2(n5123), .ZN(n4719)
         );
  AOI21_X1 U5905 ( .B1(n6462), .B2(n5020), .A(n4719), .ZN(n4720) );
  OAI211_X1 U5906 ( .C1(n5046), .C2(n6472), .A(n4721), .B(n4720), .ZN(U3121)
         );
  NAND2_X1 U5907 ( .A1(n5016), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4724)
         );
  OAI22_X1 U5908 ( .A1(n5118), .A2(n5018), .B1(n5017), .B2(n5117), .ZN(n4722)
         );
  AOI21_X1 U5909 ( .B1(n6456), .B2(n5020), .A(n4722), .ZN(n4723) );
  OAI211_X1 U5910 ( .C1(n5046), .C2(n6461), .A(n4724), .B(n4723), .ZN(U3120)
         );
  NAND2_X1 U5911 ( .A1(n5016), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4727)
         );
  OAI22_X1 U5912 ( .A1(n5086), .A2(n5018), .B1(n5017), .B2(n5085), .ZN(n4725)
         );
  AOI21_X1 U5913 ( .B1(n6438), .B2(n5020), .A(n4725), .ZN(n4726) );
  OAI211_X1 U5914 ( .C1(n5046), .C2(n6443), .A(n4727), .B(n4726), .ZN(U3116)
         );
  NAND2_X1 U5915 ( .A1(n5016), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4730)
         );
  OAI22_X1 U5916 ( .A1(n5113), .A2(n5018), .B1(n5017), .B2(n5112), .ZN(n4728)
         );
  AOI21_X1 U5917 ( .B1(n6450), .B2(n5020), .A(n4728), .ZN(n4729) );
  OAI211_X1 U5918 ( .C1(n5046), .C2(n6455), .A(n4730), .B(n4729), .ZN(U3119)
         );
  NAND2_X1 U5919 ( .A1(n5016), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4733)
         );
  OAI22_X1 U5920 ( .A1(n5091), .A2(n5018), .B1(n5017), .B2(n5090), .ZN(n4731)
         );
  AOI21_X1 U5921 ( .B1(n6444), .B2(n5020), .A(n4731), .ZN(n4732) );
  OAI211_X1 U5922 ( .C1(n5046), .C2(n6449), .A(n4733), .B(n4732), .ZN(U3118)
         );
  NAND3_X1 U5923 ( .A1(n5131), .A2(n4794), .A3(n4110), .ZN(n4856) );
  INV_X1 U5924 ( .A(n4856), .ZN(n4734) );
  NOR3_X1 U5925 ( .A1(n5009), .A2(n5029), .A3(n5733), .ZN(n4736) );
  INV_X1 U5926 ( .A(n4512), .ZN(n5252) );
  NOR2_X1 U5927 ( .A1(n5252), .A2(n5447), .ZN(n4839) );
  NAND2_X1 U5928 ( .A1(n4839), .A2(n5077), .ZN(n4740) );
  OAI21_X1 U5929 ( .B1(n4736), .B2(n4735), .A(n4740), .ZN(n4739) );
  NAND3_X1 U5930 ( .A1(n6485), .A2(n5075), .A3(n4790), .ZN(n4853) );
  OR2_X1 U5931 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4853), .ZN(n5007)
         );
  AOI211_X1 U5932 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5007), .A(n6366), .B(
        n4737), .ZN(n4738) );
  NAND2_X1 U5933 ( .A1(n4739), .A2(n4738), .ZN(n5005) );
  NAND2_X1 U5934 ( .A1(n5005), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4744) );
  INV_X1 U5935 ( .A(n4740), .ZN(n4849) );
  AOI22_X1 U5936 ( .A1(n4849), .A2(n6371), .B1(n4767), .B2(n4741), .ZN(n5006)
         );
  OAI22_X1 U5937 ( .A1(n5108), .A2(n5007), .B1(n5006), .B2(n5107), .ZN(n4742)
         );
  AOI21_X1 U5938 ( .B1(n6429), .B2(n5009), .A(n4742), .ZN(n4743) );
  OAI211_X1 U5939 ( .C1(n5012), .C2(n6437), .A(n4744), .B(n4743), .ZN(U3027)
         );
  NAND2_X1 U5940 ( .A1(n5005), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4747) );
  OAI22_X1 U5941 ( .A1(n5091), .A2(n5007), .B1(n5006), .B2(n5090), .ZN(n4745)
         );
  AOI21_X1 U5942 ( .B1(n6444), .B2(n5009), .A(n4745), .ZN(n4746) );
  OAI211_X1 U5943 ( .C1(n5012), .C2(n6449), .A(n4747), .B(n4746), .ZN(U3022)
         );
  NAND2_X1 U5944 ( .A1(n5005), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4750) );
  OAI22_X1 U5945 ( .A1(n5086), .A2(n5007), .B1(n5006), .B2(n5085), .ZN(n4748)
         );
  AOI21_X1 U5946 ( .B1(n6438), .B2(n5009), .A(n4748), .ZN(n4749) );
  OAI211_X1 U5947 ( .C1(n5012), .C2(n6443), .A(n4750), .B(n4749), .ZN(U3020)
         );
  NAND2_X1 U5948 ( .A1(n5005), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4753) );
  OAI22_X1 U5949 ( .A1(n5113), .A2(n5007), .B1(n5006), .B2(n5112), .ZN(n4751)
         );
  AOI21_X1 U5950 ( .B1(n6450), .B2(n5009), .A(n4751), .ZN(n4752) );
  OAI211_X1 U5951 ( .C1(n5012), .C2(n6455), .A(n4753), .B(n4752), .ZN(U3023)
         );
  NAND2_X1 U5952 ( .A1(n5005), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4756) );
  OAI22_X1 U5953 ( .A1(n5118), .A2(n5007), .B1(n5006), .B2(n5117), .ZN(n4754)
         );
  AOI21_X1 U5954 ( .B1(n6456), .B2(n5009), .A(n4754), .ZN(n4755) );
  OAI211_X1 U5955 ( .C1(n5012), .C2(n6461), .A(n4756), .B(n4755), .ZN(U3024)
         );
  NAND2_X1 U5956 ( .A1(n5005), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4759) );
  OAI22_X1 U5957 ( .A1(n5126), .A2(n5007), .B1(n5006), .B2(n5123), .ZN(n4757)
         );
  AOI21_X1 U5958 ( .B1(n6462), .B2(n5009), .A(n4757), .ZN(n4758) );
  OAI211_X1 U5959 ( .C1(n5012), .C2(n6472), .A(n4759), .B(n4758), .ZN(U3025)
         );
  INV_X1 U5960 ( .A(n4760), .ZN(n4761) );
  NOR2_X1 U5961 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4761), .ZN(n4770)
         );
  OAI21_X1 U5962 ( .B1(n4990), .B2(n4763), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4764) );
  NAND3_X1 U5963 ( .A1(n4968), .A2(n6371), .A3(n4764), .ZN(n4769) );
  NAND2_X1 U5964 ( .A1(n5083), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4765) );
  NAND2_X1 U5965 ( .A1(n4766), .A2(n4765), .ZN(n6377) );
  NOR3_X1 U5966 ( .A1(n6377), .A2(n6485), .A3(n4767), .ZN(n4768) );
  NAND2_X1 U5967 ( .A1(n4986), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4774)
         );
  INV_X1 U5968 ( .A(n4770), .ZN(n4988) );
  NOR2_X1 U5969 ( .A1(n4968), .A2(n5733), .ZN(n6364) );
  INV_X1 U5970 ( .A(n6366), .ZN(n4792) );
  NOR3_X1 U5971 ( .A1(n4792), .A2(n6485), .A3(n5083), .ZN(n4771) );
  AOI21_X1 U5972 ( .B1(n6364), .B2(n6368), .A(n4771), .ZN(n4987) );
  OAI22_X1 U5973 ( .A1(n5113), .A2(n4988), .B1(n4987), .B2(n5112), .ZN(n4772)
         );
  AOI21_X1 U5974 ( .B1(n6393), .B2(n4990), .A(n4772), .ZN(n4773) );
  OAI211_X1 U5975 ( .C1(n5033), .C2(n6396), .A(n4774), .B(n4773), .ZN(U3135)
         );
  NAND2_X1 U5976 ( .A1(n4986), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4777)
         );
  OAI22_X1 U5977 ( .A1(n5108), .A2(n4988), .B1(n4987), .B2(n5107), .ZN(n4775)
         );
  AOI21_X1 U5978 ( .B1(n6414), .B2(n4990), .A(n4775), .ZN(n4776) );
  OAI211_X1 U5979 ( .C1(n5033), .C2(n6418), .A(n4777), .B(n4776), .ZN(U3139)
         );
  NAND2_X1 U5980 ( .A1(n4986), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4780)
         );
  OAI22_X1 U5981 ( .A1(n5091), .A2(n4988), .B1(n4987), .B2(n5090), .ZN(n4778)
         );
  AOI21_X1 U5982 ( .B1(n6389), .B2(n4990), .A(n4778), .ZN(n4779) );
  OAI211_X1 U5983 ( .C1(n5033), .C2(n6392), .A(n4780), .B(n4779), .ZN(U3134)
         );
  NAND2_X1 U5984 ( .A1(n4986), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4783)
         );
  OAI22_X1 U5985 ( .A1(n5086), .A2(n4988), .B1(n4987), .B2(n5085), .ZN(n4781)
         );
  AOI21_X1 U5986 ( .B1(n6379), .B2(n4990), .A(n4781), .ZN(n4782) );
  OAI211_X1 U5987 ( .C1(n5033), .C2(n6382), .A(n4783), .B(n4782), .ZN(U3132)
         );
  NAND2_X1 U5988 ( .A1(n4986), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4786)
         );
  OAI22_X1 U5989 ( .A1(n5118), .A2(n4988), .B1(n4987), .B2(n5117), .ZN(n4784)
         );
  AOI21_X1 U5990 ( .B1(n6397), .B2(n4990), .A(n4784), .ZN(n4785) );
  OAI211_X1 U5991 ( .C1(n5033), .C2(n6400), .A(n4786), .B(n4785), .ZN(U3136)
         );
  NAND2_X1 U5992 ( .A1(n4986), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4789)
         );
  OAI22_X1 U5993 ( .A1(n5126), .A2(n4988), .B1(n4987), .B2(n5123), .ZN(n4787)
         );
  AOI21_X1 U5994 ( .B1(n6401), .B2(n4990), .A(n4787), .ZN(n4788) );
  OAI211_X1 U5995 ( .C1(n5033), .C2(n6404), .A(n4789), .B(n4788), .ZN(U3137)
         );
  NAND3_X1 U5996 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5075), .A3(n4790), .ZN(n4842) );
  NOR2_X1 U5997 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4842), .ZN(n4832)
         );
  OAI211_X1 U5998 ( .C1(n3296), .C2(n4832), .A(n4792), .B(n4791), .ZN(n4799)
         );
  NAND3_X1 U5999 ( .A1(n6419), .A2(n6371), .A3(n4889), .ZN(n4797) );
  NAND2_X1 U6000 ( .A1(n4839), .A2(n6368), .ZN(n4801) );
  INV_X1 U6001 ( .A(n4801), .ZN(n4796) );
  AOI21_X1 U6002 ( .B1(n4797), .B2(n6373), .A(n4796), .ZN(n4798) );
  OAI22_X1 U6003 ( .A1(n4801), .A2(n5733), .B1(n6375), .B2(n4800), .ZN(n4831)
         );
  AOI22_X1 U6004 ( .A1(n6451), .A2(n4832), .B1(n6452), .B2(n4831), .ZN(n4802)
         );
  OAI21_X1 U6005 ( .B1(n6455), .B2(n6419), .A(n4802), .ZN(n4803) );
  AOI21_X1 U6006 ( .B1(n6450), .B2(n4835), .A(n4803), .ZN(n4804) );
  OAI21_X1 U6007 ( .B1(n4837), .B2(n6746), .A(n4804), .ZN(U3087) );
  INV_X1 U6008 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4808) );
  AOI22_X1 U6009 ( .A1(n6445), .A2(n4832), .B1(n6446), .B2(n4831), .ZN(n4805)
         );
  OAI21_X1 U6010 ( .B1(n6449), .B2(n6419), .A(n4805), .ZN(n4806) );
  AOI21_X1 U6011 ( .B1(n6444), .B2(n4835), .A(n4806), .ZN(n4807) );
  OAI21_X1 U6012 ( .B1(n4837), .B2(n4808), .A(n4807), .ZN(U3086) );
  INV_X1 U6013 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4812) );
  AOI22_X1 U6014 ( .A1(n6465), .A2(n4832), .B1(n6467), .B2(n4831), .ZN(n4809)
         );
  OAI21_X1 U6015 ( .B1(n6472), .B2(n6419), .A(n4809), .ZN(n4810) );
  AOI21_X1 U6016 ( .B1(n6462), .B2(n4835), .A(n4810), .ZN(n4811) );
  OAI21_X1 U6017 ( .B1(n4837), .B2(n4812), .A(n4811), .ZN(U3089) );
  INV_X1 U6018 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4816) );
  AOI22_X1 U6019 ( .A1(n6428), .A2(n4832), .B1(n6432), .B2(n4831), .ZN(n4813)
         );
  OAI21_X1 U6020 ( .B1(n6437), .B2(n6419), .A(n4813), .ZN(n4814) );
  AOI21_X1 U6021 ( .B1(n6429), .B2(n4835), .A(n4814), .ZN(n4815) );
  OAI21_X1 U6022 ( .B1(n4837), .B2(n4816), .A(n4815), .ZN(U3091) );
  INV_X1 U6023 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4820) );
  AOI22_X1 U6024 ( .A1(n6457), .A2(n4832), .B1(n6458), .B2(n4831), .ZN(n4817)
         );
  OAI21_X1 U6025 ( .B1(n6461), .B2(n6419), .A(n4817), .ZN(n4818) );
  AOI21_X1 U6026 ( .B1(n6456), .B2(n4835), .A(n4818), .ZN(n4819) );
  OAI21_X1 U6027 ( .B1(n4837), .B2(n4820), .A(n4819), .ZN(U3088) );
  INV_X1 U6028 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4824) );
  AOI22_X1 U6029 ( .A1(n6439), .A2(n4832), .B1(n6440), .B2(n4831), .ZN(n4821)
         );
  OAI21_X1 U6030 ( .B1(n6443), .B2(n6419), .A(n4821), .ZN(n4822) );
  AOI21_X1 U6031 ( .B1(n6438), .B2(n4835), .A(n4822), .ZN(n4823) );
  OAI21_X1 U6032 ( .B1(n4837), .B2(n4824), .A(n4823), .ZN(U3084) );
  INV_X1 U6033 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4828) );
  NAND2_X1 U6034 ( .A1(n6273), .A2(DATAI_22_), .ZN(n6410) );
  INV_X1 U6035 ( .A(n6410), .ZN(n5205) );
  NAND2_X1 U6036 ( .A1(n6273), .A2(DATAI_30_), .ZN(n5207) );
  NAND2_X1 U6037 ( .A1(n4829), .A2(n3303), .ZN(n5101) );
  INV_X1 U6038 ( .A(DATAI_6_), .ZN(n6815) );
  AOI22_X1 U6039 ( .A1(n6406), .A2(n4832), .B1(n6405), .B2(n4831), .ZN(n4825)
         );
  OAI21_X1 U6040 ( .B1(n5207), .B2(n6419), .A(n4825), .ZN(n4826) );
  AOI21_X1 U6041 ( .B1(n5205), .B2(n4835), .A(n4826), .ZN(n4827) );
  OAI21_X1 U6042 ( .B1(n4837), .B2(n4828), .A(n4827), .ZN(U3090) );
  NAND2_X1 U6043 ( .A1(n6273), .A2(DATAI_17_), .ZN(n6388) );
  INV_X1 U6044 ( .A(n6388), .ZN(n5219) );
  NAND2_X1 U6045 ( .A1(n6273), .A2(DATAI_25_), .ZN(n5223) );
  NAND2_X1 U6046 ( .A1(n4829), .A2(n4361), .ZN(n5096) );
  AOI22_X1 U6047 ( .A1(n6384), .A2(n4832), .B1(n6383), .B2(n4831), .ZN(n4833)
         );
  OAI21_X1 U6048 ( .B1(n5223), .B2(n6419), .A(n4833), .ZN(n4834) );
  AOI21_X1 U6049 ( .B1(n5219), .B2(n4835), .A(n4834), .ZN(n4836) );
  OAI21_X1 U6050 ( .B1(n4837), .B2(n6820), .A(n4836), .ZN(U3085) );
  INV_X1 U6051 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6153) );
  OAI222_X1 U6052 ( .A1(n5855), .A2(n6243), .B1(n5246), .B2(n6815), .C1(n5539), 
        .C2(n6153), .ZN(U2885) );
  INV_X1 U6053 ( .A(n4838), .ZN(n4900) );
  NOR2_X1 U6054 ( .A1(n5179), .A2(n4842), .ZN(n4885) );
  AOI21_X1 U6055 ( .B1(n4839), .B2(n4900), .A(n4885), .ZN(n4843) );
  AOI21_X1 U6056 ( .B1(n4846), .B2(STATEBS16_REG_SCAN_IN), .A(n5733), .ZN(
        n4841) );
  AOI22_X1 U6057 ( .A1(n4843), .A2(n4841), .B1(n5733), .B2(n4842), .ZN(n4840)
         );
  NAND2_X1 U6058 ( .A1(n4973), .A2(n4840), .ZN(n4884) );
  INV_X1 U6059 ( .A(n4841), .ZN(n4844) );
  OAI22_X1 U6060 ( .A1(n4844), .A2(n4843), .B1(n6497), .B2(n4842), .ZN(n4883)
         );
  AOI22_X1 U6061 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4884), .B1(n6383), 
        .B2(n4883), .ZN(n4848) );
  AOI22_X1 U6062 ( .A1(n4886), .A2(n5219), .B1(n6384), .B2(n4885), .ZN(n4847)
         );
  OAI211_X1 U6063 ( .C1(n5223), .C2(n4889), .A(n4848), .B(n4847), .ZN(U3093)
         );
  NOR2_X1 U6064 ( .A1(n5179), .A2(n4853), .ZN(n4892) );
  AOI21_X1 U6065 ( .B1(n4849), .B2(n6475), .A(n4892), .ZN(n4855) );
  OR2_X1 U6066 ( .A1(n4856), .A2(n5939), .ZN(n4850) );
  AOI22_X1 U6067 ( .A1(n4855), .A2(n4852), .B1(n5733), .B2(n4853), .ZN(n4851)
         );
  NAND2_X1 U6068 ( .A1(n4973), .A2(n4851), .ZN(n4891) );
  INV_X1 U6069 ( .A(n4852), .ZN(n4854) );
  OAI22_X1 U6070 ( .A1(n4855), .A2(n4854), .B1(n6497), .B2(n4853), .ZN(n4890)
         );
  AOI22_X1 U6071 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4891), .B1(n6405), 
        .B2(n4890), .ZN(n4858) );
  AOI22_X1 U6072 ( .A1(n6406), .A2(n4892), .B1(n5205), .B2(n5128), .ZN(n4857)
         );
  OAI211_X1 U6073 ( .C1(n5207), .C2(n4895), .A(n4858), .B(n4857), .ZN(U3034)
         );
  AOI22_X1 U6074 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4884), .B1(n6440), 
        .B2(n4883), .ZN(n4860) );
  AOI22_X1 U6075 ( .A1(n4886), .A2(n6438), .B1(n6439), .B2(n4885), .ZN(n4859)
         );
  OAI211_X1 U6076 ( .C1(n6443), .C2(n4889), .A(n4860), .B(n4859), .ZN(U3092)
         );
  AOI22_X1 U6077 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4884), .B1(n6452), 
        .B2(n4883), .ZN(n4862) );
  AOI22_X1 U6078 ( .A1(n4886), .A2(n6450), .B1(n6451), .B2(n4885), .ZN(n4861)
         );
  OAI211_X1 U6079 ( .C1(n6455), .C2(n4889), .A(n4862), .B(n4861), .ZN(U3095)
         );
  AOI22_X1 U6080 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4884), .B1(n6432), 
        .B2(n4883), .ZN(n4864) );
  AOI22_X1 U6081 ( .A1(n4886), .A2(n6429), .B1(n6428), .B2(n4885), .ZN(n4863)
         );
  OAI211_X1 U6082 ( .C1(n6437), .C2(n4889), .A(n4864), .B(n4863), .ZN(U3099)
         );
  AOI22_X1 U6083 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4891), .B1(n6383), 
        .B2(n4890), .ZN(n4866) );
  AOI22_X1 U6084 ( .A1(n6384), .A2(n4892), .B1(n5219), .B2(n5128), .ZN(n4865)
         );
  OAI211_X1 U6085 ( .C1(n5223), .C2(n4895), .A(n4866), .B(n4865), .ZN(U3029)
         );
  AOI22_X1 U6086 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4891), .B1(n6432), 
        .B2(n4890), .ZN(n4868) );
  AOI22_X1 U6087 ( .A1(n6428), .A2(n4892), .B1(n6429), .B2(n5128), .ZN(n4867)
         );
  OAI211_X1 U6088 ( .C1(n6437), .C2(n4895), .A(n4868), .B(n4867), .ZN(U3035)
         );
  AOI22_X1 U6089 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4891), .B1(n6467), 
        .B2(n4890), .ZN(n4870) );
  AOI22_X1 U6090 ( .A1(n6465), .A2(n4892), .B1(n6462), .B2(n5128), .ZN(n4869)
         );
  OAI211_X1 U6091 ( .C1(n6472), .C2(n4895), .A(n4870), .B(n4869), .ZN(U3033)
         );
  AOI22_X1 U6092 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4891), .B1(n6458), 
        .B2(n4890), .ZN(n4872) );
  AOI22_X1 U6093 ( .A1(n6457), .A2(n4892), .B1(n6456), .B2(n5128), .ZN(n4871)
         );
  OAI211_X1 U6094 ( .C1(n6461), .C2(n4895), .A(n4872), .B(n4871), .ZN(U3032)
         );
  AOI22_X1 U6095 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4891), .B1(n6440), 
        .B2(n4890), .ZN(n4874) );
  AOI22_X1 U6096 ( .A1(n6439), .A2(n4892), .B1(n6438), .B2(n5128), .ZN(n4873)
         );
  OAI211_X1 U6097 ( .C1(n6443), .C2(n4895), .A(n4874), .B(n4873), .ZN(U3028)
         );
  AOI22_X1 U6098 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4884), .B1(n6467), 
        .B2(n4883), .ZN(n4876) );
  AOI22_X1 U6099 ( .A1(n4886), .A2(n6462), .B1(n6465), .B2(n4885), .ZN(n4875)
         );
  OAI211_X1 U6100 ( .C1(n6472), .C2(n4889), .A(n4876), .B(n4875), .ZN(U3097)
         );
  AOI22_X1 U6101 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4884), .B1(n6446), 
        .B2(n4883), .ZN(n4878) );
  AOI22_X1 U6102 ( .A1(n4886), .A2(n6444), .B1(n6445), .B2(n4885), .ZN(n4877)
         );
  OAI211_X1 U6103 ( .C1(n6449), .C2(n4889), .A(n4878), .B(n4877), .ZN(U3094)
         );
  AOI22_X1 U6104 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4884), .B1(n6405), 
        .B2(n4883), .ZN(n4880) );
  AOI22_X1 U6105 ( .A1(n4886), .A2(n5205), .B1(n6406), .B2(n4885), .ZN(n4879)
         );
  OAI211_X1 U6106 ( .C1(n5207), .C2(n4889), .A(n4880), .B(n4879), .ZN(U3098)
         );
  AOI22_X1 U6107 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4891), .B1(n6452), 
        .B2(n4890), .ZN(n4882) );
  AOI22_X1 U6108 ( .A1(n6451), .A2(n4892), .B1(n6450), .B2(n5128), .ZN(n4881)
         );
  OAI211_X1 U6109 ( .C1(n6455), .C2(n4895), .A(n4882), .B(n4881), .ZN(U3031)
         );
  AOI22_X1 U6110 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4884), .B1(n6458), 
        .B2(n4883), .ZN(n4888) );
  AOI22_X1 U6111 ( .A1(n4886), .A2(n6456), .B1(n6457), .B2(n4885), .ZN(n4887)
         );
  OAI211_X1 U6112 ( .C1(n6461), .C2(n4889), .A(n4888), .B(n4887), .ZN(U3096)
         );
  AOI22_X1 U6113 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4891), .B1(n6446), 
        .B2(n4890), .ZN(n4894) );
  AOI22_X1 U6114 ( .A1(n6445), .A2(n4892), .B1(n6444), .B2(n5128), .ZN(n4893)
         );
  OAI211_X1 U6115 ( .C1(n6449), .C2(n4895), .A(n4894), .B(n4893), .ZN(U3030)
         );
  XNOR2_X1 U6116 ( .A(n4897), .B(n4896), .ZN(n6229) );
  AOI22_X1 U6117 ( .A1(n5340), .A2(DATAI_8_), .B1(n6947), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4898) );
  OAI21_X1 U6118 ( .B1(n5855), .B2(n6229), .A(n4898), .ZN(U2883) );
  NOR2_X1 U6119 ( .A1(n5179), .A2(n4904), .ZN(n4923) );
  AOI21_X1 U6120 ( .B1(n4900), .B2(n4899), .A(n4923), .ZN(n4906) );
  NAND3_X1 U6121 ( .A1(n6371), .A2(n4906), .A3(n4903), .ZN(n4901) );
  OAI211_X1 U6122 ( .C1(n6371), .C2(n4902), .A(n4973), .B(n4901), .ZN(n4922)
         );
  NAND2_X1 U6123 ( .A1(n6371), .A2(n4903), .ZN(n4905) );
  OAI22_X1 U6124 ( .A1(n4906), .A2(n4905), .B1(n6497), .B2(n4904), .ZN(n4921)
         );
  AOI22_X1 U6125 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4922), .B1(n6383), 
        .B2(n4921), .ZN(n4908) );
  INV_X1 U6126 ( .A(n5223), .ZN(n6385) );
  AOI22_X1 U6127 ( .A1(n6384), .A2(n4923), .B1(n6385), .B2(n5020), .ZN(n4907)
         );
  OAI211_X1 U6128 ( .C1(n6388), .C2(n4926), .A(n4908), .B(n4907), .ZN(U3125)
         );
  AOI22_X1 U6129 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4922), .B1(n6432), 
        .B2(n4921), .ZN(n4910) );
  AOI22_X1 U6130 ( .A1(n6428), .A2(n4923), .B1(n6414), .B2(n5020), .ZN(n4909)
         );
  OAI211_X1 U6131 ( .C1(n6418), .C2(n4926), .A(n4910), .B(n4909), .ZN(U3131)
         );
  AOI22_X1 U6132 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4922), .B1(n6446), 
        .B2(n4921), .ZN(n4912) );
  AOI22_X1 U6133 ( .A1(n6445), .A2(n4923), .B1(n6389), .B2(n5020), .ZN(n4911)
         );
  OAI211_X1 U6134 ( .C1(n6392), .C2(n4926), .A(n4912), .B(n4911), .ZN(U3126)
         );
  AOI22_X1 U6135 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4922), .B1(n6440), 
        .B2(n4921), .ZN(n4914) );
  AOI22_X1 U6136 ( .A1(n6439), .A2(n4923), .B1(n6379), .B2(n5020), .ZN(n4913)
         );
  OAI211_X1 U6137 ( .C1(n6382), .C2(n4926), .A(n4914), .B(n4913), .ZN(U3124)
         );
  AOI22_X1 U6138 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4922), .B1(n6458), 
        .B2(n4921), .ZN(n4916) );
  AOI22_X1 U6139 ( .A1(n6457), .A2(n4923), .B1(n6397), .B2(n5020), .ZN(n4915)
         );
  OAI211_X1 U6140 ( .C1(n6400), .C2(n4926), .A(n4916), .B(n4915), .ZN(U3128)
         );
  AOI22_X1 U6141 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4922), .B1(n6405), 
        .B2(n4921), .ZN(n4918) );
  INV_X1 U6142 ( .A(n5207), .ZN(n6407) );
  AOI22_X1 U6143 ( .A1(n6406), .A2(n4923), .B1(n6407), .B2(n5020), .ZN(n4917)
         );
  OAI211_X1 U6144 ( .C1(n6410), .C2(n4926), .A(n4918), .B(n4917), .ZN(U3130)
         );
  AOI22_X1 U6145 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4922), .B1(n6467), 
        .B2(n4921), .ZN(n4920) );
  AOI22_X1 U6146 ( .A1(n6465), .A2(n4923), .B1(n6401), .B2(n5020), .ZN(n4919)
         );
  OAI211_X1 U6147 ( .C1(n6404), .C2(n4926), .A(n4920), .B(n4919), .ZN(U3129)
         );
  AOI22_X1 U6148 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4922), .B1(n6452), 
        .B2(n4921), .ZN(n4925) );
  AOI22_X1 U6149 ( .A1(n6451), .A2(n4923), .B1(n6393), .B2(n5020), .ZN(n4924)
         );
  OAI211_X1 U6150 ( .C1(n6396), .C2(n4926), .A(n4925), .B(n4924), .ZN(U3127)
         );
  NAND2_X1 U6151 ( .A1(n4958), .A2(n6471), .ZN(n4928) );
  AOI21_X1 U6152 ( .B1(n4928), .B2(STATEBS16_REG_SCAN_IN), .A(n5733), .ZN(
        n4932) );
  AND2_X1 U6153 ( .A1(n4512), .A2(n5447), .ZN(n5076) );
  NOR3_X1 U6154 ( .A1(n6375), .A2(n6485), .A3(n5083), .ZN(n4929) );
  NOR2_X1 U6155 ( .A1(n6366), .A2(n6377), .ZN(n5080) );
  INV_X1 U6156 ( .A(n5040), .ZN(n4931) );
  NAND3_X1 U6157 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5075), .ZN(n5042) );
  NOR2_X1 U6158 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5042), .ZN(n4934)
         );
  NOR2_X1 U6159 ( .A1(n4934), .A2(n3296), .ZN(n4930) );
  AOI21_X1 U6160 ( .B1(n4932), .B2(n4931), .A(n4930), .ZN(n4933) );
  OAI211_X1 U6161 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6497), .A(n5080), .B(n4933), .ZN(n4956) );
  NAND2_X1 U6162 ( .A1(n4956), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4937)
         );
  INV_X1 U6163 ( .A(n4934), .ZN(n4957) );
  OAI22_X1 U6164 ( .A1(n4958), .A2(n6461), .B1(n5118), .B2(n4957), .ZN(n4935)
         );
  AOI21_X1 U6165 ( .B1(n4960), .B2(n6456), .A(n4935), .ZN(n4936) );
  OAI211_X1 U6166 ( .C1(n4963), .C2(n5117), .A(n4937), .B(n4936), .ZN(U3104)
         );
  NAND2_X1 U6167 ( .A1(n4956), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4940)
         );
  OAI22_X1 U6168 ( .A1(n4958), .A2(n6443), .B1(n5086), .B2(n4957), .ZN(n4938)
         );
  AOI21_X1 U6169 ( .B1(n4960), .B2(n6438), .A(n4938), .ZN(n4939) );
  OAI211_X1 U6170 ( .C1(n4963), .C2(n5085), .A(n4940), .B(n4939), .ZN(U3100)
         );
  NAND2_X1 U6171 ( .A1(n4956), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4943)
         );
  OAI22_X1 U6172 ( .A1(n4958), .A2(n6455), .B1(n5113), .B2(n4957), .ZN(n4941)
         );
  AOI21_X1 U6173 ( .B1(n4960), .B2(n6450), .A(n4941), .ZN(n4942) );
  OAI211_X1 U6174 ( .C1(n4963), .C2(n5112), .A(n4943), .B(n4942), .ZN(U3103)
         );
  NAND2_X1 U6175 ( .A1(n4956), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4946)
         );
  OAI22_X1 U6176 ( .A1(n4958), .A2(n5223), .B1(n5096), .B2(n4957), .ZN(n4944)
         );
  AOI21_X1 U6177 ( .B1(n4960), .B2(n5219), .A(n4944), .ZN(n4945) );
  OAI211_X1 U6178 ( .C1(n4963), .C2(n5095), .A(n4946), .B(n4945), .ZN(U3101)
         );
  NAND2_X1 U6179 ( .A1(n4956), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4949)
         );
  OAI22_X1 U6180 ( .A1(n4958), .A2(n5207), .B1(n5101), .B2(n4957), .ZN(n4947)
         );
  AOI21_X1 U6181 ( .B1(n4960), .B2(n5205), .A(n4947), .ZN(n4948) );
  OAI211_X1 U6182 ( .C1(n4963), .C2(n5100), .A(n4949), .B(n4948), .ZN(U3106)
         );
  NAND2_X1 U6183 ( .A1(n4956), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4952)
         );
  OAI22_X1 U6184 ( .A1(n4958), .A2(n6437), .B1(n5108), .B2(n4957), .ZN(n4950)
         );
  AOI21_X1 U6185 ( .B1(n4960), .B2(n6429), .A(n4950), .ZN(n4951) );
  OAI211_X1 U6186 ( .C1(n4963), .C2(n5107), .A(n4952), .B(n4951), .ZN(U3107)
         );
  NAND2_X1 U6187 ( .A1(n4956), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4955)
         );
  OAI22_X1 U6188 ( .A1(n4958), .A2(n6472), .B1(n5126), .B2(n4957), .ZN(n4953)
         );
  AOI21_X1 U6189 ( .B1(n4960), .B2(n6462), .A(n4953), .ZN(n4954) );
  OAI211_X1 U6190 ( .C1(n4963), .C2(n5123), .A(n4955), .B(n4954), .ZN(U3105)
         );
  NAND2_X1 U6191 ( .A1(n4956), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4962)
         );
  OAI22_X1 U6192 ( .A1(n4958), .A2(n6449), .B1(n5091), .B2(n4957), .ZN(n4959)
         );
  AOI21_X1 U6193 ( .B1(n4960), .B2(n6444), .A(n4959), .ZN(n4961) );
  OAI211_X1 U6194 ( .C1(n4963), .C2(n5090), .A(n4962), .B(n4961), .ZN(U3102)
         );
  XOR2_X1 U6195 ( .A(n4965), .B(n4964), .Z(n6234) );
  INV_X1 U6196 ( .A(n6234), .ZN(n5036) );
  INV_X1 U6197 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6151) );
  OAI222_X1 U6198 ( .A1(n5855), .A2(n5036), .B1(n5246), .B2(n6191), .C1(n5539), 
        .C2(n6151), .ZN(U2884) );
  NAND2_X1 U6199 ( .A1(n4966), .A2(n6371), .ZN(n4976) );
  NOR2_X1 U6200 ( .A1(n4968), .A2(n4967), .ZN(n6372) );
  NAND2_X1 U6201 ( .A1(n6372), .A2(n6475), .ZN(n4969) );
  NAND2_X1 U6202 ( .A1(n4969), .A2(n6420), .ZN(n4975) );
  INV_X1 U6203 ( .A(n4975), .ZN(n4970) );
  OAI22_X1 U6204 ( .A1(n4976), .A2(n4970), .B1(n6363), .B2(n6497), .ZN(n6431)
         );
  INV_X1 U6205 ( .A(n6431), .ZN(n5067) );
  INV_X1 U6206 ( .A(n6436), .ZN(n4980) );
  OAI22_X1 U6207 ( .A1(n6419), .A2(n6400), .B1(n5118), .B2(n6420), .ZN(n4972)
         );
  AOI21_X1 U6208 ( .B1(n6397), .B2(n4980), .A(n4972), .ZN(n4978) );
  AOI21_X1 U6209 ( .B1(n5733), .B2(n6363), .A(n5183), .ZN(n4974) );
  OAI21_X1 U6210 ( .B1(n4976), .B2(n4975), .A(n4974), .ZN(n6433) );
  NAND2_X1 U6211 ( .A1(n6433), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4977) );
  OAI211_X1 U6212 ( .C1(n5067), .C2(n5117), .A(n4978), .B(n4977), .ZN(U3080)
         );
  OAI22_X1 U6213 ( .A1(n6419), .A2(n6404), .B1(n5126), .B2(n6420), .ZN(n4979)
         );
  AOI21_X1 U6214 ( .B1(n6401), .B2(n4980), .A(n4979), .ZN(n4982) );
  NAND2_X1 U6215 ( .A1(n6433), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4981) );
  OAI211_X1 U6216 ( .C1(n5067), .C2(n5123), .A(n4982), .B(n4981), .ZN(U3081)
         );
  NAND2_X1 U6217 ( .A1(n4986), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4985)
         );
  OAI22_X1 U6218 ( .A1(n5101), .A2(n4988), .B1(n4987), .B2(n5100), .ZN(n4983)
         );
  AOI21_X1 U6219 ( .B1(n6407), .B2(n4990), .A(n4983), .ZN(n4984) );
  OAI211_X1 U6220 ( .C1(n5033), .C2(n6410), .A(n4985), .B(n4984), .ZN(U3138)
         );
  NAND2_X1 U6221 ( .A1(n4986), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4992)
         );
  OAI22_X1 U6222 ( .A1(n5096), .A2(n4988), .B1(n4987), .B2(n5095), .ZN(n4989)
         );
  AOI21_X1 U6223 ( .B1(n6385), .B2(n4990), .A(n4989), .ZN(n4991) );
  OAI211_X1 U6224 ( .C1(n5033), .C2(n6388), .A(n4992), .B(n4991), .ZN(U3133)
         );
  NAND2_X1 U6225 ( .A1(n4996), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4995) );
  OAI22_X1 U6226 ( .A1(n5096), .A2(n4998), .B1(n4997), .B2(n5095), .ZN(n4993)
         );
  AOI21_X1 U6227 ( .B1(n6385), .B2(n5169), .A(n4993), .ZN(n4994) );
  OAI211_X1 U6228 ( .C1(n5222), .C2(n6388), .A(n4995), .B(n4994), .ZN(U3053)
         );
  NAND2_X1 U6229 ( .A1(n4996), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5001) );
  OAI22_X1 U6230 ( .A1(n5101), .A2(n4998), .B1(n4997), .B2(n5100), .ZN(n4999)
         );
  AOI21_X1 U6231 ( .B1(n6407), .B2(n5169), .A(n4999), .ZN(n5000) );
  OAI211_X1 U6232 ( .C1(n5222), .C2(n6410), .A(n5001), .B(n5000), .ZN(U3058)
         );
  NAND2_X1 U6233 ( .A1(n5005), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5004) );
  OAI22_X1 U6234 ( .A1(n5096), .A2(n5007), .B1(n5006), .B2(n5095), .ZN(n5002)
         );
  AOI21_X1 U6235 ( .B1(n5219), .B2(n5009), .A(n5002), .ZN(n5003) );
  OAI211_X1 U6236 ( .C1(n5012), .C2(n5223), .A(n5004), .B(n5003), .ZN(U3021)
         );
  NAND2_X1 U6237 ( .A1(n5005), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5011) );
  OAI22_X1 U6238 ( .A1(n5101), .A2(n5007), .B1(n5006), .B2(n5100), .ZN(n5008)
         );
  AOI21_X1 U6239 ( .B1(n5205), .B2(n5009), .A(n5008), .ZN(n5010) );
  OAI211_X1 U6240 ( .C1(n5012), .C2(n5207), .A(n5011), .B(n5010), .ZN(U3026)
         );
  NAND2_X1 U6241 ( .A1(n5016), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5015)
         );
  OAI22_X1 U6242 ( .A1(n5096), .A2(n5018), .B1(n5017), .B2(n5095), .ZN(n5013)
         );
  AOI21_X1 U6243 ( .B1(n5219), .B2(n5020), .A(n5013), .ZN(n5014) );
  OAI211_X1 U6244 ( .C1(n5046), .C2(n5223), .A(n5015), .B(n5014), .ZN(U3117)
         );
  NAND2_X1 U6245 ( .A1(n5016), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5022)
         );
  OAI22_X1 U6246 ( .A1(n5101), .A2(n5018), .B1(n5017), .B2(n5100), .ZN(n5019)
         );
  AOI21_X1 U6247 ( .B1(n5205), .B2(n5020), .A(n5019), .ZN(n5021) );
  OAI211_X1 U6248 ( .C1(n5046), .C2(n5207), .A(n5022), .B(n5021), .ZN(U3122)
         );
  OAI22_X1 U6249 ( .A1(n5101), .A2(n5027), .B1(n5026), .B2(n5100), .ZN(n5023)
         );
  AOI21_X1 U6250 ( .B1(n5205), .B2(n5029), .A(n5023), .ZN(n5025) );
  NAND2_X1 U6251 ( .A1(n5030), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5024)
         );
  OAI211_X1 U6252 ( .C1(n5033), .C2(n5207), .A(n5025), .B(n5024), .ZN(U3146)
         );
  OAI22_X1 U6253 ( .A1(n5096), .A2(n5027), .B1(n5026), .B2(n5095), .ZN(n5028)
         );
  AOI21_X1 U6254 ( .B1(n5219), .B2(n5029), .A(n5028), .ZN(n5032) );
  NAND2_X1 U6255 ( .A1(n5030), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5031)
         );
  OAI211_X1 U6256 ( .C1(n5033), .C2(n5223), .A(n5032), .B(n5031), .ZN(U3141)
         );
  AOI21_X1 U6257 ( .B1(n5035), .B2(n5034), .A(n5070), .ZN(n6312) );
  INV_X1 U6258 ( .A(n6312), .ZN(n6067) );
  INV_X1 U6259 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5037) );
  OAI222_X1 U6260 ( .A1(n6067), .A2(n5538), .B1(n5037), .B2(n5537), .C1(n5536), 
        .C2(n5036), .ZN(U2852) );
  INV_X1 U6261 ( .A(n5731), .ZN(n5038) );
  OAI21_X1 U6262 ( .B1(n5039), .B2(n5038), .A(n6371), .ZN(n5045) );
  NOR2_X1 U6263 ( .A1(n5134), .A2(n6485), .ZN(n6464) );
  AOI21_X1 U6264 ( .B1(n5040), .B2(n6475), .A(n6464), .ZN(n5041) );
  OAI22_X1 U6265 ( .A1(n5045), .A2(n5041), .B1(n5042), .B2(n6497), .ZN(n6466)
         );
  INV_X1 U6266 ( .A(n6466), .ZN(n5056) );
  INV_X1 U6267 ( .A(n5041), .ZN(n5044) );
  AOI21_X1 U6268 ( .B1(n5733), .B2(n5042), .A(n5183), .ZN(n5043) );
  OAI21_X1 U6269 ( .B1(n5045), .B2(n5044), .A(n5043), .ZN(n6468) );
  AOI22_X1 U6270 ( .A1(n6384), .A2(n6464), .B1(n6463), .B2(n5219), .ZN(n5047)
         );
  OAI21_X1 U6271 ( .B1(n6471), .B2(n5223), .A(n5047), .ZN(n5048) );
  AOI21_X1 U6272 ( .B1(INSTQUEUE_REG_11__1__SCAN_IN), .B2(n6468), .A(n5048), 
        .ZN(n5049) );
  OAI21_X1 U6273 ( .B1(n5056), .B2(n5095), .A(n5049), .ZN(U3109) );
  AOI22_X1 U6274 ( .A1(n6406), .A2(n6464), .B1(n6463), .B2(n5205), .ZN(n5050)
         );
  OAI21_X1 U6275 ( .B1(n6471), .B2(n5207), .A(n5050), .ZN(n5051) );
  AOI21_X1 U6276 ( .B1(INSTQUEUE_REG_11__6__SCAN_IN), .B2(n6468), .A(n5051), 
        .ZN(n5052) );
  OAI21_X1 U6277 ( .B1(n5056), .B2(n5100), .A(n5052), .ZN(U3114) );
  AOI22_X1 U6278 ( .A1(n6428), .A2(n6464), .B1(n6463), .B2(n6429), .ZN(n5053)
         );
  OAI21_X1 U6279 ( .B1(n6471), .B2(n6437), .A(n5053), .ZN(n5054) );
  AOI21_X1 U6280 ( .B1(INSTQUEUE_REG_11__7__SCAN_IN), .B2(n6468), .A(n5054), 
        .ZN(n5055) );
  OAI21_X1 U6281 ( .B1(n5056), .B2(n5107), .A(n5055), .ZN(U3115) );
  OAI21_X1 U6282 ( .B1(n5058), .B2(n5057), .A(n5234), .ZN(n6221) );
  INV_X1 U6283 ( .A(DATAI_9_), .ZN(n6193) );
  INV_X1 U6284 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6678) );
  OAI222_X1 U6285 ( .A1(n5855), .A2(n6221), .B1(n5246), .B2(n6193), .C1(n5539), 
        .C2(n6678), .ZN(U2882) );
  NAND2_X1 U6286 ( .A1(n5068), .A2(n5059), .ZN(n5060) );
  NAND2_X1 U6287 ( .A1(n3132), .A2(n5060), .ZN(n6296) );
  OAI222_X1 U6288 ( .A1(n6296), .A2(n5538), .B1(n5537), .B2(n6042), .C1(n5536), 
        .C2(n6221), .ZN(U2850) );
  NOR2_X1 U6289 ( .A1(n6436), .A2(n5223), .ZN(n5062) );
  OAI22_X1 U6290 ( .A1(n6419), .A2(n6388), .B1(n5096), .B2(n6420), .ZN(n5061)
         );
  AOI211_X1 U6291 ( .C1(INSTQUEUE_REG_7__1__SCAN_IN), .C2(n6433), .A(n5062), 
        .B(n5061), .ZN(n5063) );
  OAI21_X1 U6292 ( .B1(n5067), .B2(n5095), .A(n5063), .ZN(U3077) );
  NOR2_X1 U6293 ( .A1(n6436), .A2(n5207), .ZN(n5065) );
  OAI22_X1 U6294 ( .A1(n6419), .A2(n6410), .B1(n5101), .B2(n6420), .ZN(n5064)
         );
  AOI211_X1 U6295 ( .C1(INSTQUEUE_REG_7__6__SCAN_IN), .C2(n6433), .A(n5065), 
        .B(n5064), .ZN(n5066) );
  OAI21_X1 U6296 ( .B1(n5067), .B2(n5100), .A(n5066), .ZN(U3082) );
  OAI21_X1 U6297 ( .B1(n5070), .B2(n5069), .A(n5068), .ZN(n6305) );
  INV_X1 U6298 ( .A(n6229), .ZN(n5071) );
  AOI22_X1 U6299 ( .A1(n5505), .A2(n5071), .B1(n5492), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5072) );
  OAI21_X1 U6300 ( .B1(n5538), .B2(n6305), .A(n5072), .ZN(U2851) );
  NAND2_X1 U6301 ( .A1(n4110), .A2(n4090), .ZN(n5074) );
  NAND3_X1 U6302 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6485), .A3(n5075), .ZN(n5139) );
  NOR2_X1 U6303 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5139), .ZN(n5082)
         );
  INV_X1 U6304 ( .A(n5172), .ZN(n5103) );
  OAI21_X1 U6305 ( .B1(n5128), .B2(n5103), .A(n6373), .ZN(n5079) );
  INV_X1 U6306 ( .A(n5135), .ZN(n5078) );
  NAND2_X1 U6307 ( .A1(n5079), .A2(n5078), .ZN(n5081) );
  NAND2_X1 U6308 ( .A1(n5122), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5089) );
  INV_X1 U6309 ( .A(n5082), .ZN(n5125) );
  NOR3_X1 U6310 ( .A1(n6375), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5083), 
        .ZN(n5084) );
  AOI21_X1 U6311 ( .B1(n5135), .B2(n6371), .A(n5084), .ZN(n5124) );
  OAI22_X1 U6312 ( .A1(n5086), .A2(n5125), .B1(n5124), .B2(n5085), .ZN(n5087)
         );
  AOI21_X1 U6313 ( .B1(n6379), .B2(n5128), .A(n5087), .ZN(n5088) );
  OAI211_X1 U6314 ( .C1(n6382), .C2(n5172), .A(n5089), .B(n5088), .ZN(U3036)
         );
  NAND2_X1 U6315 ( .A1(n5122), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5094) );
  OAI22_X1 U6316 ( .A1(n5091), .A2(n5125), .B1(n5124), .B2(n5090), .ZN(n5092)
         );
  AOI21_X1 U6317 ( .B1(n6389), .B2(n5128), .A(n5092), .ZN(n5093) );
  OAI211_X1 U6318 ( .C1(n5172), .C2(n6392), .A(n5094), .B(n5093), .ZN(U3038)
         );
  NAND2_X1 U6319 ( .A1(n5122), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5099) );
  OAI22_X1 U6320 ( .A1(n5096), .A2(n5125), .B1(n5124), .B2(n5095), .ZN(n5097)
         );
  AOI21_X1 U6321 ( .B1(n5219), .B2(n5103), .A(n5097), .ZN(n5098) );
  OAI211_X1 U6322 ( .C1(n5106), .C2(n5223), .A(n5099), .B(n5098), .ZN(U3037)
         );
  NAND2_X1 U6323 ( .A1(n5122), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5105) );
  OAI22_X1 U6324 ( .A1(n5101), .A2(n5125), .B1(n5124), .B2(n5100), .ZN(n5102)
         );
  AOI21_X1 U6325 ( .B1(n5205), .B2(n5103), .A(n5102), .ZN(n5104) );
  OAI211_X1 U6326 ( .C1(n5106), .C2(n5207), .A(n5105), .B(n5104), .ZN(U3042)
         );
  NAND2_X1 U6327 ( .A1(n5122), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5111) );
  OAI22_X1 U6328 ( .A1(n5108), .A2(n5125), .B1(n5124), .B2(n5107), .ZN(n5109)
         );
  AOI21_X1 U6329 ( .B1(n6414), .B2(n5128), .A(n5109), .ZN(n5110) );
  OAI211_X1 U6330 ( .C1(n5172), .C2(n6418), .A(n5111), .B(n5110), .ZN(U3043)
         );
  NAND2_X1 U6331 ( .A1(n5122), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5116) );
  OAI22_X1 U6332 ( .A1(n5113), .A2(n5125), .B1(n5124), .B2(n5112), .ZN(n5114)
         );
  AOI21_X1 U6333 ( .B1(n6393), .B2(n5128), .A(n5114), .ZN(n5115) );
  OAI211_X1 U6334 ( .C1(n5172), .C2(n6396), .A(n5116), .B(n5115), .ZN(U3039)
         );
  NAND2_X1 U6335 ( .A1(n5122), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5121) );
  OAI22_X1 U6336 ( .A1(n5118), .A2(n5125), .B1(n5124), .B2(n5117), .ZN(n5119)
         );
  AOI21_X1 U6337 ( .B1(n6397), .B2(n5128), .A(n5119), .ZN(n5120) );
  OAI211_X1 U6338 ( .C1(n5172), .C2(n6400), .A(n5121), .B(n5120), .ZN(U3040)
         );
  NAND2_X1 U6339 ( .A1(n5122), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5130) );
  OAI22_X1 U6340 ( .A1(n5126), .A2(n5125), .B1(n5124), .B2(n5123), .ZN(n5127)
         );
  AOI21_X1 U6341 ( .B1(n6401), .B2(n5128), .A(n5127), .ZN(n5129) );
  OAI211_X1 U6342 ( .C1(n5172), .C2(n6404), .A(n5130), .B(n5129), .ZN(U3041)
         );
  NAND3_X1 U6343 ( .A1(n5132), .A2(n5131), .A3(n5731), .ZN(n5133) );
  NAND2_X1 U6344 ( .A1(n5133), .A2(n6371), .ZN(n5141) );
  INV_X1 U6345 ( .A(n5141), .ZN(n5138) );
  NOR2_X1 U6346 ( .A1(n5134), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5170)
         );
  AOI21_X1 U6347 ( .B1(n5135), .B2(n6475), .A(n5170), .ZN(n5140) );
  INV_X1 U6348 ( .A(n5139), .ZN(n5136) );
  NOR2_X1 U6349 ( .A1(n6371), .A2(n5136), .ZN(n5137) );
  AOI211_X2 U6350 ( .C1(n5138), .C2(n5140), .A(n5137), .B(n5183), .ZN(n5177)
         );
  INV_X1 U6351 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5145) );
  OAI22_X1 U6352 ( .A1(n5141), .A2(n5140), .B1(n5139), .B2(n6497), .ZN(n5174)
         );
  AOI22_X1 U6353 ( .A1(n6451), .A2(n5170), .B1(n6450), .B2(n5169), .ZN(n5142)
         );
  OAI21_X1 U6354 ( .B1(n6455), .B2(n5172), .A(n5142), .ZN(n5143) );
  AOI21_X1 U6355 ( .B1(n5174), .B2(n6452), .A(n5143), .ZN(n5144) );
  OAI21_X1 U6356 ( .B1(n5177), .B2(n5145), .A(n5144), .ZN(U3047) );
  AOI22_X1 U6357 ( .A1(n6465), .A2(n5170), .B1(n6462), .B2(n5169), .ZN(n5146)
         );
  OAI21_X1 U6358 ( .B1(n6472), .B2(n5172), .A(n5146), .ZN(n5147) );
  AOI21_X1 U6359 ( .B1(n5174), .B2(n6467), .A(n5147), .ZN(n5148) );
  OAI21_X1 U6360 ( .B1(n5177), .B2(n3455), .A(n5148), .ZN(U3049) );
  INV_X1 U6361 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5152) );
  AOI22_X1 U6362 ( .A1(n6457), .A2(n5170), .B1(n6456), .B2(n5169), .ZN(n5149)
         );
  OAI21_X1 U6363 ( .B1(n6461), .B2(n5172), .A(n5149), .ZN(n5150) );
  AOI21_X1 U6364 ( .B1(n5174), .B2(n6458), .A(n5150), .ZN(n5151) );
  OAI21_X1 U6365 ( .B1(n5177), .B2(n5152), .A(n5151), .ZN(U3048) );
  INV_X1 U6366 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5156) );
  AOI22_X1 U6367 ( .A1(n6445), .A2(n5170), .B1(n6444), .B2(n5169), .ZN(n5153)
         );
  OAI21_X1 U6368 ( .B1(n6449), .B2(n5172), .A(n5153), .ZN(n5154) );
  AOI21_X1 U6369 ( .B1(n5174), .B2(n6446), .A(n5154), .ZN(n5155) );
  OAI21_X1 U6370 ( .B1(n5177), .B2(n5156), .A(n5155), .ZN(U3046) );
  INV_X1 U6371 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5160) );
  AOI22_X1 U6372 ( .A1(n6406), .A2(n5170), .B1(n5205), .B2(n5169), .ZN(n5157)
         );
  OAI21_X1 U6373 ( .B1(n5207), .B2(n5172), .A(n5157), .ZN(n5158) );
  AOI21_X1 U6374 ( .B1(n5174), .B2(n6405), .A(n5158), .ZN(n5159) );
  OAI21_X1 U6375 ( .B1(n5177), .B2(n5160), .A(n5159), .ZN(U3050) );
  INV_X1 U6376 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5164) );
  AOI22_X1 U6377 ( .A1(n6384), .A2(n5170), .B1(n5219), .B2(n5169), .ZN(n5161)
         );
  OAI21_X1 U6378 ( .B1(n5223), .B2(n5172), .A(n5161), .ZN(n5162) );
  AOI21_X1 U6379 ( .B1(n5174), .B2(n6383), .A(n5162), .ZN(n5163) );
  OAI21_X1 U6380 ( .B1(n5177), .B2(n5164), .A(n5163), .ZN(U3045) );
  INV_X1 U6381 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5168) );
  AOI22_X1 U6382 ( .A1(n6439), .A2(n5170), .B1(n6438), .B2(n5169), .ZN(n5165)
         );
  OAI21_X1 U6383 ( .B1(n6443), .B2(n5172), .A(n5165), .ZN(n5166) );
  AOI21_X1 U6384 ( .B1(n5174), .B2(n6440), .A(n5166), .ZN(n5167) );
  OAI21_X1 U6385 ( .B1(n5177), .B2(n5168), .A(n5167), .ZN(U3044) );
  INV_X1 U6386 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5176) );
  AOI22_X1 U6387 ( .A1(n6428), .A2(n5170), .B1(n6429), .B2(n5169), .ZN(n5171)
         );
  OAI21_X1 U6388 ( .B1(n6437), .B2(n5172), .A(n5171), .ZN(n5173) );
  AOI21_X1 U6389 ( .B1(n5174), .B2(n6432), .A(n5173), .ZN(n5175) );
  OAI21_X1 U6390 ( .B1(n5177), .B2(n5176), .A(n5175), .ZN(U3051) );
  INV_X1 U6391 ( .A(n5178), .ZN(n5180) );
  NOR2_X1 U6392 ( .A1(n5179), .A2(n5185), .ZN(n5220) );
  AOI21_X1 U6393 ( .B1(n5180), .B2(n6475), .A(n5220), .ZN(n5186) );
  INV_X1 U6394 ( .A(n5185), .ZN(n5181) );
  NOR2_X1 U6395 ( .A1(n6371), .A2(n5181), .ZN(n5182) );
  AOI211_X2 U6396 ( .C1(n5184), .C2(n5186), .A(n5183), .B(n5182), .ZN(n5228)
         );
  INV_X1 U6397 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5192) );
  INV_X1 U6398 ( .A(n5184), .ZN(n5187) );
  OAI22_X1 U6399 ( .A1(n5187), .A2(n5186), .B1(n5185), .B2(n6497), .ZN(n5225)
         );
  AOI22_X1 U6400 ( .A1(n6465), .A2(n5220), .B1(n6462), .B2(n6413), .ZN(n5189)
         );
  OAI21_X1 U6401 ( .B1(n6472), .B2(n5222), .A(n5189), .ZN(n5190) );
  AOI21_X1 U6402 ( .B1(n6467), .B2(n5225), .A(n5190), .ZN(n5191) );
  OAI21_X1 U6403 ( .B1(n5228), .B2(n5192), .A(n5191), .ZN(U3065) );
  INV_X1 U6404 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5196) );
  AOI22_X1 U6405 ( .A1(n6445), .A2(n5220), .B1(n6444), .B2(n6413), .ZN(n5193)
         );
  OAI21_X1 U6406 ( .B1(n6449), .B2(n5222), .A(n5193), .ZN(n5194) );
  AOI21_X1 U6407 ( .B1(n6446), .B2(n5225), .A(n5194), .ZN(n5195) );
  OAI21_X1 U6408 ( .B1(n5228), .B2(n5196), .A(n5195), .ZN(U3062) );
  INV_X1 U6409 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5200) );
  AOI22_X1 U6410 ( .A1(n6428), .A2(n5220), .B1(n6429), .B2(n6413), .ZN(n5197)
         );
  OAI21_X1 U6411 ( .B1(n6437), .B2(n5222), .A(n5197), .ZN(n5198) );
  AOI21_X1 U6412 ( .B1(n6432), .B2(n5225), .A(n5198), .ZN(n5199) );
  OAI21_X1 U6413 ( .B1(n5228), .B2(n5200), .A(n5199), .ZN(U3067) );
  INV_X1 U6414 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5204) );
  AOI22_X1 U6415 ( .A1(n6451), .A2(n5220), .B1(n6450), .B2(n6413), .ZN(n5201)
         );
  OAI21_X1 U6416 ( .B1(n6455), .B2(n5222), .A(n5201), .ZN(n5202) );
  AOI21_X1 U6417 ( .B1(n6452), .B2(n5225), .A(n5202), .ZN(n5203) );
  OAI21_X1 U6418 ( .B1(n5228), .B2(n5204), .A(n5203), .ZN(U3063) );
  INV_X1 U6419 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5210) );
  AOI22_X1 U6420 ( .A1(n6406), .A2(n5220), .B1(n5205), .B2(n6413), .ZN(n5206)
         );
  OAI21_X1 U6421 ( .B1(n5207), .B2(n5222), .A(n5206), .ZN(n5208) );
  AOI21_X1 U6422 ( .B1(n6405), .B2(n5225), .A(n5208), .ZN(n5209) );
  OAI21_X1 U6423 ( .B1(n5228), .B2(n5210), .A(n5209), .ZN(U3066) );
  INV_X1 U6424 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5214) );
  AOI22_X1 U6425 ( .A1(n6439), .A2(n5220), .B1(n6438), .B2(n6413), .ZN(n5211)
         );
  OAI21_X1 U6426 ( .B1(n6443), .B2(n5222), .A(n5211), .ZN(n5212) );
  AOI21_X1 U6427 ( .B1(n6440), .B2(n5225), .A(n5212), .ZN(n5213) );
  OAI21_X1 U6428 ( .B1(n5228), .B2(n5214), .A(n5213), .ZN(U3060) );
  INV_X1 U6429 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5218) );
  AOI22_X1 U6430 ( .A1(n6457), .A2(n5220), .B1(n6456), .B2(n6413), .ZN(n5215)
         );
  OAI21_X1 U6431 ( .B1(n6461), .B2(n5222), .A(n5215), .ZN(n5216) );
  AOI21_X1 U6432 ( .B1(n6458), .B2(n5225), .A(n5216), .ZN(n5217) );
  OAI21_X1 U6433 ( .B1(n5228), .B2(n5218), .A(n5217), .ZN(U3064) );
  INV_X1 U6434 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5227) );
  AOI22_X1 U6435 ( .A1(n6384), .A2(n5220), .B1(n5219), .B2(n6413), .ZN(n5221)
         );
  OAI21_X1 U6436 ( .B1(n5223), .B2(n5222), .A(n5221), .ZN(n5224) );
  AOI21_X1 U6437 ( .B1(n6383), .B2(n5225), .A(n5224), .ZN(n5226) );
  OAI21_X1 U6438 ( .B1(n5228), .B2(n5227), .A(n5226), .ZN(U3061) );
  AOI21_X1 U6439 ( .B1(n5230), .B2(n3132), .A(n5239), .ZN(n5231) );
  INV_X1 U6440 ( .A(n5231), .ZN(n6034) );
  INV_X1 U6441 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5235) );
  AOI21_X1 U6442 ( .B1(n5234), .B2(n5233), .A(n5237), .ZN(n6037) );
  INV_X1 U6443 ( .A(n6037), .ZN(n5244) );
  OAI222_X1 U6444 ( .A1(n6034), .A2(n5538), .B1(n5235), .B2(n5537), .C1(n5244), 
        .C2(n5536), .ZN(U2849) );
  OAI21_X1 U6445 ( .B1(n5237), .B2(n5236), .A(n5297), .ZN(n6213) );
  NOR2_X1 U6446 ( .A1(n5239), .A2(n5238), .ZN(n5240) );
  OR2_X1 U6447 ( .A1(n5300), .A2(n5240), .ZN(n6024) );
  OAI22_X1 U6448 ( .A1(n6024), .A2(n5538), .B1(n5537), .B2(n6877), .ZN(n5241)
         );
  INV_X1 U6449 ( .A(n5241), .ZN(n5242) );
  OAI21_X1 U6450 ( .B1(n6213), .B2(n5536), .A(n5242), .ZN(U2848) );
  AOI22_X1 U6451 ( .A1(n5340), .A2(DATAI_11_), .B1(n6947), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5243) );
  OAI21_X1 U6452 ( .B1(n6213), .B2(n5855), .A(n5243), .ZN(U2880) );
  OAI222_X1 U6453 ( .A1(n5246), .A2(n5245), .B1(n5539), .B2(n6875), .C1(n5855), 
        .C2(n5244), .ZN(U2881) );
  AND2_X1 U6454 ( .A1(n5247), .A2(n5249), .ZN(n5248) );
  NOR2_X1 U6455 ( .A1(n6070), .A2(n5248), .ZN(n6116) );
  INV_X1 U6456 ( .A(n6277), .ZN(n5259) );
  INV_X1 U6457 ( .A(n5249), .ZN(n5250) );
  OR2_X1 U6458 ( .A1(n5251), .A2(n5250), .ZN(n6114) );
  INV_X1 U6459 ( .A(n6114), .ZN(n6101) );
  NAND2_X1 U6460 ( .A1(n5252), .A2(n6101), .ZN(n5254) );
  AOI22_X1 U6461 ( .A1(n6112), .A2(EBX_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6110), .ZN(n5253) );
  OAI211_X1 U6462 ( .C1(n6350), .C2(n6123), .A(n5254), .B(n5253), .ZN(n5258)
         );
  INV_X1 U6463 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6538) );
  INV_X1 U6464 ( .A(n6096), .ZN(n6111) );
  NAND2_X1 U6465 ( .A1(n6111), .A2(REIP_REG_1__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6466 ( .A1(n5262), .A2(REIP_REG_1__SCAN_IN), .ZN(n5255) );
  AOI21_X1 U6467 ( .B1(n6063), .B2(n5255), .A(n6538), .ZN(n6098) );
  AOI21_X1 U6468 ( .B1(n6538), .B2(n5256), .A(n6098), .ZN(n5257) );
  AOI211_X1 U6469 ( .C1(n6120), .C2(n5259), .A(n5258), .B(n5257), .ZN(n5260)
         );
  OAI21_X1 U6470 ( .B1(n6116), .B2(n5261), .A(n5260), .ZN(U2825) );
  NAND2_X1 U6471 ( .A1(n5263), .A2(n5262), .ZN(n6066) );
  OAI21_X1 U6472 ( .B1(n6109), .B2(n6094), .A(n6063), .ZN(n6103) );
  OAI22_X1 U6473 ( .A1(n6103), .A2(n6542), .B1(n6123), .B2(n6330), .ZN(n5264)
         );
  AOI211_X1 U6474 ( .C1(n6110), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6083), 
        .B(n5264), .ZN(n5270) );
  NOR3_X1 U6475 ( .A1(n6096), .A2(REIP_REG_4__SCAN_IN), .A3(n6094), .ZN(n5265)
         );
  AOI21_X1 U6476 ( .B1(n6112), .B2(EBX_REG_4__SCAN_IN), .A(n5265), .ZN(n5266)
         );
  OAI21_X1 U6477 ( .B1(n5267), .B2(n6114), .A(n5266), .ZN(n5268) );
  AOI21_X1 U6478 ( .B1(n6120), .B2(n6256), .A(n5268), .ZN(n5269) );
  OAI211_X1 U6479 ( .C1(n6116), .C2(n6260), .A(n5270), .B(n5269), .ZN(U2823)
         );
  NOR2_X1 U6480 ( .A1(n3507), .A2(n6114), .ZN(n5273) );
  OAI22_X1 U6481 ( .A1(n6123), .A2(n5721), .B1(n6073), .B2(n5271), .ZN(n5272)
         );
  AOI211_X1 U6482 ( .C1(n6063), .C2(REIP_REG_0__SCAN_IN), .A(n5273), .B(n5272), 
        .ZN(n5275) );
  OAI21_X1 U6483 ( .B1(n6120), .B2(n6110), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5274) );
  OAI211_X1 U6484 ( .C1(n6116), .C2(n5276), .A(n5275), .B(n5274), .ZN(U2827)
         );
  NAND2_X1 U6485 ( .A1(n6207), .A2(n5277), .ZN(n5279) );
  XOR2_X1 U6486 ( .A(n5279), .B(n3147), .Z(n5294) );
  INV_X1 U6487 ( .A(n6038), .ZN(n5281) );
  AOI22_X1 U6488 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6325), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5280) );
  OAI21_X1 U6489 ( .B1(n6280), .B2(n5281), .A(n5280), .ZN(n5282) );
  AOI21_X1 U6490 ( .B1(n6037), .B2(n6273), .A(n5282), .ZN(n5283) );
  OAI21_X1 U6491 ( .B1(n5294), .B2(n6278), .A(n5283), .ZN(U2976) );
  INV_X1 U6492 ( .A(n6333), .ZN(n5284) );
  NAND2_X1 U6493 ( .A1(n5288), .A2(n5284), .ZN(n6316) );
  NOR2_X1 U6494 ( .A1(n5285), .A2(n6316), .ZN(n6298) );
  OAI211_X1 U6495 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6298), .B(n5286), .ZN(n5293) );
  INV_X1 U6496 ( .A(n5688), .ZN(n5290) );
  OAI22_X1 U6497 ( .A1(n5288), .A2(n5317), .B1(n5690), .B2(n5287), .ZN(n5289)
         );
  NOR2_X1 U6498 ( .A1(n5290), .A2(n5289), .ZN(n6314) );
  OAI21_X1 U6499 ( .B1(n6304), .B2(n5691), .A(n6314), .ZN(n6295) );
  OAI22_X1 U6500 ( .A1(n6351), .A2(n6034), .B1(n6551), .B2(n6349), .ZN(n5291)
         );
  AOI21_X1 U6501 ( .B1(n6295), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5291), 
        .ZN(n5292) );
  OAI211_X1 U6502 ( .C1(n5294), .C2(n5913), .A(n5293), .B(n5292), .ZN(U3008)
         );
  AOI21_X1 U6503 ( .B1(n5297), .B2(n5296), .A(n5304), .ZN(n6019) );
  INV_X1 U6504 ( .A(n6019), .ZN(n5302) );
  AOI22_X1 U6505 ( .A1(n5340), .A2(DATAI_12_), .B1(n6947), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5298) );
  OAI21_X1 U6506 ( .B1(n5302), .B2(n5855), .A(n5298), .ZN(U2879) );
  OR2_X1 U6507 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  NAND2_X1 U6508 ( .A1(n5307), .A2(n5301), .ZN(n6016) );
  INV_X1 U6509 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6701) );
  OAI222_X1 U6510 ( .A1(n6016), .A2(n5538), .B1(n5537), .B2(n6701), .C1(n5302), 
        .C2(n5536), .ZN(U2847) );
  OAI21_X1 U6511 ( .B1(n5304), .B2(n5303), .A(n5336), .ZN(n6010) );
  AOI22_X1 U6512 ( .A1(n5340), .A2(DATAI_13_), .B1(n6947), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5305) );
  OAI21_X1 U6513 ( .B1(n6010), .B2(n5855), .A(n5305), .ZN(U2878) );
  NAND2_X1 U6514 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  NAND2_X1 U6515 ( .A1(n5343), .A2(n5308), .ZN(n6006) );
  OAI22_X1 U6516 ( .A1(n6006), .A2(n5538), .B1(n5537), .B2(n5309), .ZN(n5310)
         );
  INV_X1 U6517 ( .A(n5310), .ZN(n5311) );
  OAI21_X1 U6518 ( .B1(n6010), .B2(n5536), .A(n5311), .ZN(U2846) );
  INV_X1 U6519 ( .A(n5313), .ZN(n5314) );
  NOR2_X1 U6520 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  XNOR2_X1 U6521 ( .A(n3148), .B(n5316), .ZN(n5333) );
  NOR3_X1 U6522 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6288), .A3(n6293), 
        .ZN(n5326) );
  OAI21_X1 U6523 ( .B1(n5318), .B2(n5317), .A(n5688), .ZN(n5319) );
  AOI21_X1 U6524 ( .B1(n5321), .B2(n5320), .A(n5319), .ZN(n6294) );
  OAI21_X1 U6525 ( .B1(n6353), .B2(n5322), .A(n6293), .ZN(n5323) );
  AOI21_X1 U6526 ( .B1(n6294), .B2(n5323), .A(n6782), .ZN(n5325) );
  NAND2_X1 U6527 ( .A1(n6325), .A2(REIP_REG_12__SCAN_IN), .ZN(n5329) );
  OAI21_X1 U6528 ( .B1(n6351), .B2(n6016), .A(n5329), .ZN(n5324) );
  NOR3_X1 U6529 ( .A1(n5326), .A2(n5325), .A3(n5324), .ZN(n5327) );
  OAI21_X1 U6530 ( .B1(n5333), .B2(n5913), .A(n5327), .ZN(U3006) );
  INV_X1 U6531 ( .A(n6020), .ZN(n5330) );
  NAND2_X1 U6532 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5328)
         );
  OAI211_X1 U6533 ( .C1(n6280), .C2(n5330), .A(n5329), .B(n5328), .ZN(n5331)
         );
  AOI21_X1 U6534 ( .B1(n6019), .B2(n6273), .A(n5331), .ZN(n5332) );
  OAI21_X1 U6535 ( .B1(n5333), .B2(n6278), .A(n5332), .ZN(U2974) );
  AOI21_X1 U6536 ( .B1(n5336), .B2(n5335), .A(n5339), .ZN(n5359) );
  INV_X1 U6537 ( .A(n5359), .ZN(n6002) );
  AOI22_X1 U6538 ( .A1(n5340), .A2(DATAI_14_), .B1(n6947), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5337) );
  OAI21_X1 U6539 ( .B1(n6002), .B2(n5855), .A(n5337), .ZN(U2877) );
  XNOR2_X1 U6540 ( .A(n5339), .B(n5338), .ZN(n5346) );
  AOI22_X1 U6541 ( .A1(n5340), .A2(DATAI_15_), .B1(n6947), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5341) );
  OAI21_X1 U6542 ( .B1(n5346), .B2(n5855), .A(n5341), .ZN(U2876) );
  INV_X1 U6543 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5345) );
  AND2_X1 U6544 ( .A1(n5343), .A2(n5342), .ZN(n5344) );
  OR2_X1 U6545 ( .A1(n5344), .A2(n5348), .ZN(n5994) );
  OAI222_X1 U6546 ( .A1(n6002), .A2(n5536), .B1(n5537), .B2(n5345), .C1(n5994), 
        .C2(n5538), .ZN(U2845) );
  INV_X1 U6547 ( .A(n5346), .ZN(n5983) );
  NOR2_X1 U6548 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  OR2_X1 U6549 ( .A1(n5364), .A2(n5349), .ZN(n5985) );
  OAI22_X1 U6550 ( .A1(n5985), .A2(n5538), .B1(n5537), .B2(n5350), .ZN(n5351)
         );
  AOI21_X1 U6551 ( .B1(n5983), .B2(n5505), .A(n5351), .ZN(n5352) );
  INV_X1 U6552 ( .A(n5352), .ZN(U2844) );
  XNOR2_X1 U6553 ( .A(n4164), .B(n5354), .ZN(n5355) );
  XNOR2_X1 U6554 ( .A(n5598), .B(n5355), .ZN(n5914) );
  INV_X1 U6555 ( .A(n5999), .ZN(n5357) );
  AOI22_X1 U6556 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6325), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5356) );
  OAI21_X1 U6557 ( .B1(n6280), .B2(n5357), .A(n5356), .ZN(n5358) );
  AOI21_X1 U6558 ( .B1(n5359), .B2(n6273), .A(n5358), .ZN(n5360) );
  OAI21_X1 U6559 ( .B1(n6278), .B2(n5914), .A(n5360), .ZN(U2972) );
  AOI21_X1 U6560 ( .B1(n5362), .B2(n5361), .A(n5367), .ZN(n6128) );
  INV_X1 U6561 ( .A(n6128), .ZN(n5366) );
  INV_X1 U6562 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5365) );
  OAI21_X1 U6563 ( .B1(n5364), .B2(n5363), .A(n5369), .ZN(n5982) );
  OAI222_X1 U6564 ( .A1(n5366), .A2(n5536), .B1(n5365), .B2(n5537), .C1(n5982), 
        .C2(n5538), .ZN(U2843) );
  OAI21_X1 U6565 ( .B1(n5368), .B2(n5367), .A(n5533), .ZN(n5972) );
  INV_X1 U6566 ( .A(n5523), .ZN(n5531) );
  AOI21_X1 U6567 ( .B1(n5370), .B2(n5369), .A(n5531), .ZN(n5970) );
  AOI22_X1 U6568 ( .A1(n5970), .A2(n5493), .B1(EBX_REG_17__SCAN_IN), .B2(n5492), .ZN(n5371) );
  OAI21_X1 U6569 ( .B1(n5972), .B2(n5536), .A(n5371), .ZN(U2842) );
  AOI22_X1 U6570 ( .A1(n6947), .A2(EAX_REG_17__SCAN_IN), .B1(n6946), .B2(
        DATAI_1_), .ZN(n5376) );
  NAND2_X1 U6571 ( .A1(n6948), .A2(DATAI_17_), .ZN(n5375) );
  OAI211_X1 U6572 ( .C1(n5972), .C2(n5855), .A(n5376), .B(n5375), .ZN(U2874)
         );
  INV_X1 U6573 ( .A(n3138), .ZN(n5378) );
  NAND2_X1 U6574 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  XNOR2_X1 U6575 ( .A(n5379), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5625)
         );
  NOR2_X1 U6576 ( .A1(n5381), .A2(n5380), .ZN(n5383) );
  INV_X1 U6577 ( .A(n5470), .ZN(n5765) );
  NAND2_X1 U6578 ( .A1(n5759), .A2(n6257), .ZN(n5384) );
  NAND2_X1 U6579 ( .A1(n6325), .A2(REIP_REG_29__SCAN_IN), .ZN(n5620) );
  OAI211_X1 U6580 ( .C1(n5588), .C2(n5385), .A(n5384), .B(n5620), .ZN(n5386)
         );
  AOI21_X1 U6581 ( .B1(n5765), .B2(n6273), .A(n5386), .ZN(n5387) );
  OAI21_X1 U6582 ( .B1(n5625), .B2(n6278), .A(n5387), .ZN(U2957) );
  AOI22_X1 U6583 ( .A1(n6947), .A2(EAX_REG_29__SCAN_IN), .B1(n6946), .B2(
        DATAI_13_), .ZN(n5389) );
  NAND2_X1 U6584 ( .A1(n6948), .A2(DATAI_29_), .ZN(n5388) );
  OAI211_X1 U6585 ( .C1(n5470), .C2(n5855), .A(n5389), .B(n5388), .ZN(U2862)
         );
  AOI22_X1 U6586 ( .A1(n6947), .A2(EAX_REG_30__SCAN_IN), .B1(n6946), .B2(
        DATAI_14_), .ZN(n5391) );
  NAND2_X1 U6587 ( .A1(n6948), .A2(DATAI_30_), .ZN(n5390) );
  OAI211_X1 U6588 ( .C1(n5748), .C2(n5855), .A(n5391), .B(n5390), .ZN(U2861)
         );
  NAND2_X1 U6589 ( .A1(n5496), .A2(n5392), .ZN(n5481) );
  INV_X1 U6590 ( .A(n5481), .ZN(n5394) );
  AOI22_X1 U6591 ( .A1(n6947), .A2(EAX_REG_26__SCAN_IN), .B1(n6946), .B2(
        DATAI_10_), .ZN(n5398) );
  NAND2_X1 U6592 ( .A1(n6948), .A2(DATAI_26_), .ZN(n5397) );
  OAI211_X1 U6593 ( .C1(n5787), .C2(n5855), .A(n5398), .B(n5397), .ZN(U2865)
         );
  NOR2_X1 U6594 ( .A1(n5482), .A2(n5399), .ZN(n5400) );
  OR2_X1 U6595 ( .A1(n4074), .A2(n5400), .ZN(n5644) );
  INV_X1 U6596 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5401) );
  OAI222_X1 U6597 ( .A1(n5644), .A2(n5538), .B1(n5401), .B2(n5537), .C1(n5787), 
        .C2(n5536), .ZN(U2833) );
  NAND2_X1 U6598 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NOR2_X1 U6599 ( .A1(n5405), .A2(n5406), .ZN(n5710) );
  AOI21_X1 U6600 ( .B1(n5406), .B2(n5405), .A(n5710), .ZN(n5417) );
  INV_X1 U6601 ( .A(n5407), .ZN(n5408) );
  OAI21_X1 U6602 ( .B1(n5408), .B2(n5691), .A(n6294), .ZN(n5903) );
  NAND2_X1 U6603 ( .A1(n5903), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6604 ( .A1(n6325), .A2(REIP_REG_15__SCAN_IN), .ZN(n5413) );
  OAI211_X1 U6605 ( .C1(n6351), .C2(n5985), .A(n5409), .B(n5413), .ZN(n5410)
         );
  AOI21_X1 U6606 ( .B1(n5905), .B2(n6679), .A(n5410), .ZN(n5411) );
  OAI21_X1 U6607 ( .B1(n5417), .B2(n5913), .A(n5411), .ZN(U3003) );
  INV_X1 U6608 ( .A(n5984), .ZN(n5414) );
  NAND2_X1 U6609 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5412)
         );
  OAI211_X1 U6610 ( .C1(n6280), .C2(n5414), .A(n5413), .B(n5412), .ZN(n5415)
         );
  AOI21_X1 U6611 ( .B1(n5983), .B2(n6273), .A(n5415), .ZN(n5416) );
  OAI21_X1 U6612 ( .B1(n5417), .B2(n6278), .A(n5416), .ZN(U2971) );
  INV_X1 U6613 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5418) );
  OAI222_X1 U6614 ( .A1(n5536), .A2(n5748), .B1(n5538), .B2(n5749), .C1(n5418), 
        .C2(n5537), .ZN(U2829) );
  INV_X1 U6615 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5419) );
  NOR2_X2 U6616 ( .A1(n5590), .A2(n5420), .ZN(n5583) );
  AND3_X1 U6617 ( .A1(n4164), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6618 ( .A1(n5583), .A2(n5421), .ZN(n5422) );
  XNOR2_X1 U6619 ( .A(n5424), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5581)
         );
  INV_X1 U6620 ( .A(n5484), .ZN(n5425) );
  AOI21_X1 U6621 ( .B1(n5426), .B2(n5434), .A(n5425), .ZN(n5801) );
  NAND2_X1 U6622 ( .A1(n6325), .A2(REIP_REG_24__SCAN_IN), .ZN(n5575) );
  INV_X1 U6623 ( .A(n5575), .ZN(n5430) );
  INV_X1 U6624 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6859) );
  INV_X1 U6625 ( .A(n5439), .ZN(n5428) );
  AOI211_X1 U6626 ( .C1(n6859), .C2(n5428), .A(n5427), .B(n5655), .ZN(n5429)
         );
  AOI211_X1 U6627 ( .C1(n5801), .C2(n6323), .A(n5430), .B(n5429), .ZN(n5431)
         );
  OAI21_X1 U6628 ( .B1(n5581), .B2(n5913), .A(n5431), .ZN(U2994) );
  OR2_X1 U6629 ( .A1(n5502), .A2(n5432), .ZN(n5433) );
  NAND2_X1 U6630 ( .A1(n5434), .A2(n5433), .ZN(n5809) );
  NAND2_X1 U6631 ( .A1(n5435), .A2(n6356), .ZN(n5441) );
  NOR2_X1 U6632 ( .A1(n5436), .A2(n4310), .ZN(n5437) );
  AOI211_X1 U6633 ( .C1(n5439), .C2(n4310), .A(n5438), .B(n5437), .ZN(n5440)
         );
  OAI211_X1 U6634 ( .C1(n6351), .C2(n5809), .A(n5441), .B(n5440), .ZN(U2995)
         );
  INV_X1 U6635 ( .A(n5442), .ZN(n6474) );
  OAI21_X1 U6636 ( .B1(n5450), .B2(n5443), .A(n6473), .ZN(n5444) );
  OAI21_X1 U6637 ( .B1(n5445), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n5444), 
        .ZN(n5446) );
  AOI21_X1 U6638 ( .B1(n5447), .B2(n6474), .A(n5446), .ZN(n6478) );
  NOR2_X1 U6639 ( .A1(n6501), .A2(n6594), .ZN(n5449) );
  AOI22_X1 U6640 ( .A1(n5450), .A2(n6592), .B1(n5449), .B2(n5448), .ZN(n5451)
         );
  OAI21_X1 U6641 ( .B1(n6478), .B2(n6600), .A(n5451), .ZN(n5452) );
  AOI22_X1 U6642 ( .A1(n6598), .A2(n5452), .B1(n5443), .B2(n6592), .ZN(n5453)
         );
  OAI21_X1 U6643 ( .B1(n6598), .B2(n5454), .A(n5453), .ZN(U3460) );
  OAI22_X1 U6644 ( .A1(n5456), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n5455), .B2(EBX_REG_31__SCAN_IN), .ZN(n5466) );
  INV_X1 U6645 ( .A(n5469), .ZN(n5471) );
  AOI21_X1 U6646 ( .B1(n5471), .B2(n5457), .A(n3987), .ZN(n5464) );
  INV_X1 U6647 ( .A(n5457), .ZN(n5461) );
  NOR2_X1 U6648 ( .A1(n5458), .A2(EBX_REG_29__SCAN_IN), .ZN(n5459) );
  AOI21_X1 U6649 ( .B1(n5461), .B2(n5460), .A(n5459), .ZN(n5468) );
  NOR3_X1 U6650 ( .A1(n5469), .A2(n5462), .A3(n5468), .ZN(n5463) );
  NOR2_X1 U6651 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  XOR2_X1 U6652 ( .A(n5466), .B(n5465), .Z(n5740) );
  INV_X1 U6653 ( .A(n5740), .ZN(n5467) );
  OAI22_X1 U6654 ( .A1(n5467), .A2(n5538), .B1(n5537), .B2(n6716), .ZN(U2828)
         );
  XNOR2_X1 U6655 ( .A(n5469), .B(n5468), .ZN(n5767) );
  OAI222_X1 U6656 ( .A1(n5536), .A2(n5470), .B1(n5537), .B2(n4351), .C1(n5538), 
        .C2(n5767), .ZN(U2830) );
  AOI21_X1 U6657 ( .B1(n5473), .B2(n5472), .A(n5471), .ZN(n5771) );
  AOI22_X1 U6658 ( .A1(n5771), .A2(n5493), .B1(EBX_REG_28__SCAN_IN), .B2(n5492), .ZN(n5474) );
  OAI21_X1 U6659 ( .B1(n5545), .B2(n5536), .A(n5474), .ZN(U2831) );
  OAI22_X1 U6660 ( .A1(n5635), .A2(n5538), .B1(n5537), .B2(n5475), .ZN(n5476)
         );
  INV_X1 U6661 ( .A(n5476), .ZN(n5477) );
  OAI21_X1 U6662 ( .B1(n5558), .B2(n5536), .A(n5477), .ZN(U2832) );
  NAND2_X1 U6663 ( .A1(n5481), .A2(n5480), .ZN(n6951) );
  INV_X1 U6664 ( .A(n6951), .ZN(n5792) );
  INV_X1 U6665 ( .A(n5792), .ZN(n5868) );
  INV_X1 U6666 ( .A(n5482), .ZN(n5486) );
  NAND2_X1 U6667 ( .A1(n5484), .A2(n5483), .ZN(n5485) );
  NAND2_X1 U6668 ( .A1(n5486), .A2(n5485), .ZN(n5796) );
  OAI22_X1 U6669 ( .A1(n5796), .A2(n5538), .B1(n5537), .B2(n6795), .ZN(n5487)
         );
  INV_X1 U6670 ( .A(n5487), .ZN(n5488) );
  OAI21_X1 U6671 ( .B1(n5868), .B2(n5536), .A(n5488), .ZN(U2834) );
  AOI21_X1 U6672 ( .B1(n5491), .B2(n5490), .A(n5489), .ZN(n5579) );
  INV_X1 U6673 ( .A(n5579), .ZN(n5804) );
  AOI22_X1 U6674 ( .A1(n5801), .A2(n5493), .B1(EBX_REG_24__SCAN_IN), .B2(n5492), .ZN(n5494) );
  OAI21_X1 U6675 ( .B1(n5804), .B2(n5536), .A(n5494), .ZN(U2835) );
  INV_X1 U6676 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5495) );
  OAI222_X1 U6677 ( .A1(n5807), .A2(n5536), .B1(n5537), .B2(n5495), .C1(n5809), 
        .C2(n5538), .ZN(U2836) );
  INV_X1 U6678 ( .A(n5496), .ZN(n5498) );
  AOI21_X1 U6679 ( .B1(n5499), .B2(n5498), .A(n5497), .ZN(n5856) );
  AOI21_X1 U6680 ( .B1(n5508), .B2(n5509), .A(n5500), .ZN(n5501) );
  OR2_X1 U6681 ( .A1(n5502), .A2(n5501), .ZN(n5669) );
  OAI22_X1 U6682 ( .A1(n5669), .A2(n5538), .B1(n5537), .B2(n5503), .ZN(n5504)
         );
  AOI21_X1 U6683 ( .B1(n5856), .B2(n5505), .A(n5504), .ZN(n5506) );
  INV_X1 U6684 ( .A(n5506), .ZN(U2837) );
  XOR2_X1 U6685 ( .A(n5516), .B(n5507), .Z(n5859) );
  INV_X1 U6686 ( .A(n5859), .ZN(n5596) );
  INV_X1 U6687 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6713) );
  XOR2_X1 U6688 ( .A(n5509), .B(n5508), .Z(n5830) );
  INV_X1 U6689 ( .A(n5830), .ZN(n5680) );
  OAI222_X1 U6690 ( .A1(n5596), .A2(n5536), .B1(n5537), .B2(n6713), .C1(n5538), 
        .C2(n5680), .ZN(U2838) );
  MUX2_X1 U6691 ( .A(n5512), .B(n5511), .S(n5510), .Z(n5514) );
  XNOR2_X1 U6692 ( .A(n5514), .B(n5513), .ZN(n5833) );
  AOI21_X1 U6693 ( .B1(n5517), .B2(n5519), .A(n5516), .ZN(n5870) );
  INV_X1 U6694 ( .A(n5870), .ZN(n5835) );
  OAI222_X1 U6695 ( .A1(n5538), .A2(n5833), .B1(n5536), .B2(n5835), .C1(n5834), 
        .C2(n5537), .ZN(U2839) );
  OAI21_X1 U6696 ( .B1(n5520), .B2(n5532), .A(n5519), .ZN(n5880) );
  AND2_X1 U6697 ( .A1(n5522), .A2(n5521), .ZN(n5528) );
  OR2_X1 U6698 ( .A1(n5523), .A2(n5528), .ZN(n5529) );
  XNOR2_X1 U6699 ( .A(n5529), .B(n5524), .ZN(n5848) );
  OAI22_X1 U6700 ( .A1(n5848), .A2(n5538), .B1(n5537), .B2(n5525), .ZN(n5526)
         );
  INV_X1 U6701 ( .A(n5526), .ZN(n5527) );
  OAI21_X1 U6702 ( .B1(n5880), .B2(n5536), .A(n5527), .ZN(U2840) );
  INV_X1 U6703 ( .A(n5528), .ZN(n5530) );
  OAI21_X1 U6704 ( .B1(n5531), .B2(n5530), .A(n5529), .ZN(n5963) );
  INV_X1 U6705 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6730) );
  AOI21_X1 U6706 ( .B1(n5534), .B2(n5533), .A(n5532), .ZN(n6124) );
  INV_X1 U6707 ( .A(n6124), .ZN(n5535) );
  OAI222_X1 U6708 ( .A1(n5538), .A2(n5963), .B1(n5537), .B2(n6730), .C1(n5536), 
        .C2(n5535), .ZN(U2841) );
  NAND3_X1 U6709 ( .A1(n5739), .A2(n5540), .A3(n5539), .ZN(n5542) );
  AOI22_X1 U6710 ( .A1(n6948), .A2(DATAI_31_), .B1(n6947), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U6711 ( .A1(n5542), .A2(n5541), .ZN(U2860) );
  AOI22_X1 U6712 ( .A1(n6947), .A2(EAX_REG_28__SCAN_IN), .B1(n6946), .B2(
        DATAI_12_), .ZN(n5544) );
  NAND2_X1 U6713 ( .A1(n6948), .A2(DATAI_28_), .ZN(n5543) );
  OAI211_X1 U6714 ( .C1(n5545), .C2(n5855), .A(n5544), .B(n5543), .ZN(U2863)
         );
  AOI22_X1 U6715 ( .A1(n6947), .A2(EAX_REG_27__SCAN_IN), .B1(n6946), .B2(
        DATAI_11_), .ZN(n5547) );
  NAND2_X1 U6716 ( .A1(n6948), .A2(DATAI_27_), .ZN(n5546) );
  OAI211_X1 U6717 ( .C1(n5558), .C2(n5855), .A(n5547), .B(n5546), .ZN(U2864)
         );
  AOI22_X1 U6718 ( .A1(n6947), .A2(EAX_REG_24__SCAN_IN), .B1(n6946), .B2(
        DATAI_8_), .ZN(n5549) );
  NAND2_X1 U6719 ( .A1(n6948), .A2(DATAI_24_), .ZN(n5548) );
  OAI211_X1 U6720 ( .C1(n5804), .C2(n5855), .A(n5549), .B(n5548), .ZN(U2867)
         );
  AOI22_X1 U6721 ( .A1(n6947), .A2(EAX_REG_23__SCAN_IN), .B1(n6946), .B2(
        DATAI_7_), .ZN(n5551) );
  NAND2_X1 U6722 ( .A1(n6948), .A2(DATAI_23_), .ZN(n5550) );
  OAI211_X1 U6723 ( .C1(n5807), .C2(n5855), .A(n5551), .B(n5550), .ZN(U2868)
         );
  AOI22_X1 U6724 ( .A1(n6947), .A2(EAX_REG_19__SCAN_IN), .B1(n6946), .B2(
        DATAI_3_), .ZN(n5553) );
  NAND2_X1 U6725 ( .A1(n6948), .A2(DATAI_19_), .ZN(n5552) );
  OAI211_X1 U6726 ( .C1(n5880), .C2(n5855), .A(n5553), .B(n5552), .ZN(U2872)
         );
  INV_X1 U6727 ( .A(n5554), .ZN(n5555) );
  NAND2_X1 U6728 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  XNOR2_X1 U6729 ( .A(n5557), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5643)
         );
  INV_X1 U6730 ( .A(n5558), .ZN(n5563) );
  NAND2_X1 U6731 ( .A1(n5559), .A2(n6257), .ZN(n5560) );
  NAND2_X1 U6732 ( .A1(n6325), .A2(REIP_REG_27__SCAN_IN), .ZN(n5636) );
  OAI211_X1 U6733 ( .C1(n5588), .C2(n5561), .A(n5560), .B(n5636), .ZN(n5562)
         );
  AOI21_X1 U6734 ( .B1(n5563), .B2(n6273), .A(n5562), .ZN(n5564) );
  OAI21_X1 U6735 ( .B1(n5643), .B2(n6278), .A(n5564), .ZN(U2959) );
  INV_X1 U6736 ( .A(n5565), .ZN(n5566) );
  NOR2_X1 U6737 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  XNOR2_X1 U6738 ( .A(n5569), .B(n5568), .ZN(n5652) );
  NAND2_X1 U6739 ( .A1(n6325), .A2(REIP_REG_26__SCAN_IN), .ZN(n5648) );
  OAI21_X1 U6740 ( .B1(n5588), .B2(n5570), .A(n5648), .ZN(n5573) );
  NOR2_X1 U6741 ( .A1(n5571), .A2(n6286), .ZN(n5572) );
  OAI21_X1 U6742 ( .B1(n5652), .B2(n6278), .A(n5574), .ZN(U2960) );
  NAND2_X1 U6743 ( .A1(n6257), .A2(n5799), .ZN(n5576) );
  OAI211_X1 U6744 ( .C1(n5588), .C2(n5577), .A(n5576), .B(n5575), .ZN(n5578)
         );
  AOI21_X1 U6745 ( .B1(n5579), .B2(n6273), .A(n5578), .ZN(n5580) );
  OAI21_X1 U6746 ( .B1(n5581), .B2(n6278), .A(n5580), .ZN(U2962) );
  AOI21_X1 U6747 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4164), .A(n5582), 
        .ZN(n5584) );
  XOR2_X1 U6748 ( .A(n5584), .B(n5583), .Z(n5672) );
  NAND2_X1 U6749 ( .A1(n6325), .A2(REIP_REG_22__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U6750 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5585)
         );
  OAI211_X1 U6751 ( .C1(n6280), .C2(n5816), .A(n5663), .B(n5585), .ZN(n5586)
         );
  AOI21_X1 U6752 ( .B1(n5856), .B2(n6273), .A(n5586), .ZN(n5587) );
  OAI21_X1 U6753 ( .B1(n5672), .B2(n6278), .A(n5587), .ZN(U2964) );
  NAND2_X1 U6754 ( .A1(n6325), .A2(REIP_REG_21__SCAN_IN), .ZN(n5674) );
  OAI21_X1 U6755 ( .B1(n5588), .B2(n5826), .A(n5674), .ZN(n5589) );
  AOI21_X1 U6756 ( .B1(n6257), .B2(n5824), .A(n5589), .ZN(n5595) );
  INV_X1 U6757 ( .A(n5590), .ZN(n5591) );
  OAI21_X1 U6758 ( .B1(n5593), .B2(n3149), .A(n5591), .ZN(n5673) );
  NAND2_X1 U6759 ( .A1(n5673), .A2(n6272), .ZN(n5594) );
  OAI211_X1 U6760 ( .C1(n5596), .C2(n6286), .A(n5595), .B(n5594), .ZN(U2965)
         );
  NOR2_X1 U6761 ( .A1(n4164), .A2(n4176), .ZN(n5886) );
  AOI21_X1 U6762 ( .B1(n4176), .B2(n4164), .A(n5886), .ZN(n5602) );
  OR2_X1 U6763 ( .A1(n5598), .A2(n5597), .ZN(n5600) );
  AND2_X1 U6764 ( .A1(n5600), .A2(n5599), .ZN(n5601) );
  XOR2_X1 U6765 ( .A(n5602), .B(n5601), .Z(n5901) );
  INV_X1 U6766 ( .A(n5973), .ZN(n5604) );
  AOI22_X1 U6767 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6325), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5603) );
  OAI21_X1 U6768 ( .B1(n6280), .B2(n5604), .A(n5603), .ZN(n5605) );
  AOI21_X1 U6769 ( .B1(n6128), .B2(n6273), .A(n5605), .ZN(n5606) );
  OAI21_X1 U6770 ( .B1(n6278), .B2(n5901), .A(n5606), .ZN(U2970) );
  AOI21_X1 U6771 ( .B1(n5609), .B2(n5608), .A(n5607), .ZN(n5614) );
  INV_X1 U6772 ( .A(n5610), .ZN(n5618) );
  NAND4_X1 U6773 ( .A1(n5618), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n5613), .ZN(n5611) );
  OAI211_X1 U6774 ( .C1(n5614), .C2(n5613), .A(n5612), .B(n5611), .ZN(n5615)
         );
  AOI21_X1 U6775 ( .B1(n5740), .B2(n6323), .A(n5615), .ZN(n5616) );
  OAI21_X1 U6776 ( .B1(n5617), .B2(n5913), .A(n5616), .ZN(U2987) );
  INV_X1 U6777 ( .A(n5767), .ZN(n5623) );
  NAND2_X1 U6778 ( .A1(n5618), .A2(n6714), .ZN(n5619) );
  OAI211_X1 U6779 ( .C1(n5621), .C2(n6714), .A(n5620), .B(n5619), .ZN(n5622)
         );
  AOI21_X1 U6780 ( .B1(n5623), .B2(n6323), .A(n5622), .ZN(n5624) );
  OAI21_X1 U6781 ( .B1(n5625), .B2(n5913), .A(n5624), .ZN(U2989) );
  NOR2_X1 U6782 ( .A1(n5638), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5630)
         );
  INV_X1 U6783 ( .A(n5626), .ZN(n5639) );
  NAND2_X1 U6784 ( .A1(n5631), .A2(n5638), .ZN(n5637) );
  AOI21_X1 U6785 ( .B1(n5639), .B2(n5637), .A(n5627), .ZN(n5628) );
  AOI211_X1 U6786 ( .C1(n5631), .C2(n5630), .A(n5629), .B(n5628), .ZN(n5633)
         );
  NAND2_X1 U6787 ( .A1(n5771), .A2(n6323), .ZN(n5632) );
  OAI211_X1 U6788 ( .C1(n5634), .C2(n5913), .A(n5633), .B(n5632), .ZN(U2990)
         );
  INV_X1 U6789 ( .A(n5635), .ZN(n5641) );
  OAI211_X1 U6790 ( .C1(n5639), .C2(n5638), .A(n5637), .B(n5636), .ZN(n5640)
         );
  AOI21_X1 U6791 ( .B1(n5641), .B2(n6323), .A(n5640), .ZN(n5642) );
  OAI21_X1 U6792 ( .B1(n5643), .B2(n5913), .A(n5642), .ZN(U2991) );
  INV_X1 U6793 ( .A(n5644), .ZN(n5784) );
  XNOR2_X1 U6794 ( .A(n5645), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5646)
         );
  NAND2_X1 U6795 ( .A1(n5656), .A2(n5646), .ZN(n5647) );
  OAI211_X1 U6796 ( .C1(n5655), .C2(n5649), .A(n5648), .B(n5647), .ZN(n5650)
         );
  AOI21_X1 U6797 ( .B1(n5784), .B2(n6323), .A(n5650), .ZN(n5651) );
  OAI21_X1 U6798 ( .B1(n5652), .B2(n5913), .A(n5651), .ZN(U2992) );
  INV_X1 U6799 ( .A(n4292), .ZN(n5654) );
  OAI21_X1 U6800 ( .B1(n5654), .B2(n3161), .A(n5653), .ZN(n5865) );
  NAND2_X1 U6801 ( .A1(n5865), .A2(n6356), .ZN(n5662) );
  INV_X1 U6802 ( .A(n5655), .ZN(n5660) );
  INV_X1 U6803 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5658) );
  INV_X1 U6804 ( .A(n5656), .ZN(n5657) );
  OAI22_X1 U6805 ( .A1(n6349), .A2(n5658), .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5657), .ZN(n5659) );
  AOI21_X1 U6806 ( .B1(n5660), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5659), 
        .ZN(n5661) );
  OAI211_X1 U6807 ( .C1(n5796), .C2(n6351), .A(n5662), .B(n5661), .ZN(U2993)
         );
  INV_X1 U6808 ( .A(n5663), .ZN(n5668) );
  INV_X1 U6809 ( .A(n5664), .ZN(n5665) );
  NOR3_X1 U6810 ( .A1(n5666), .A2(n5665), .A3(n5675), .ZN(n5667) );
  AOI211_X1 U6811 ( .C1(n5677), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5668), .B(n5667), .ZN(n5671) );
  INV_X1 U6812 ( .A(n5669), .ZN(n5818) );
  NAND2_X1 U6813 ( .A1(n5818), .A2(n6323), .ZN(n5670) );
  OAI211_X1 U6814 ( .C1(n5672), .C2(n5913), .A(n5671), .B(n5670), .ZN(U2996)
         );
  NAND2_X1 U6815 ( .A1(n5673), .A2(n6356), .ZN(n5679) );
  OAI21_X1 U6816 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5675), .A(n5674), 
        .ZN(n5676) );
  AOI21_X1 U6817 ( .B1(n5677), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5676), 
        .ZN(n5678) );
  OAI211_X1 U6818 ( .C1(n5680), .C2(n6351), .A(n5679), .B(n5678), .ZN(U2997)
         );
  INV_X1 U6819 ( .A(n5682), .ZN(n5684) );
  NAND2_X1 U6820 ( .A1(n5684), .A2(n5683), .ZN(n5685) );
  XNOR2_X1 U6821 ( .A(n5681), .B(n5685), .ZN(n5869) );
  NAND2_X1 U6822 ( .A1(n5869), .A2(n6356), .ZN(n5699) );
  OAI21_X1 U6823 ( .B1(n4177), .B2(n5686), .A(n6353), .ZN(n5687) );
  OAI211_X1 U6824 ( .C1(n5690), .C2(n5689), .A(n5688), .B(n5687), .ZN(n5896)
         );
  AOI21_X1 U6825 ( .B1(n6346), .B2(n4177), .A(n5896), .ZN(n5714) );
  OAI21_X1 U6826 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5691), .A(n5714), 
        .ZN(n5707) );
  INV_X1 U6827 ( .A(n5692), .ZN(n5695) );
  NAND4_X1 U6828 ( .A1(n5695), .A2(n5701), .A3(n5694), .A4(n5693), .ZN(n5696)
         );
  OAI21_X1 U6829 ( .B1(n6349), .B2(n6566), .A(n5696), .ZN(n5697) );
  AOI21_X1 U6830 ( .B1(n5707), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5697), 
        .ZN(n5698) );
  OAI211_X1 U6831 ( .C1(n5833), .C2(n6351), .A(n5699), .B(n5698), .ZN(U2998)
         );
  NOR2_X1 U6832 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n5900), .ZN(n5700)
         );
  AOI22_X1 U6833 ( .A1(n6325), .A2(REIP_REG_19__SCAN_IN), .B1(n5701), .B2(
        n5700), .ZN(n5702) );
  OAI21_X1 U6834 ( .B1(n5848), .B2(n6351), .A(n5702), .ZN(n5706) );
  OAI21_X1 U6835 ( .B1(n5703), .B2(n5704), .A(n4306), .ZN(n5876) );
  NOR2_X1 U6836 ( .A1(n5876), .A2(n5913), .ZN(n5705) );
  AOI211_X1 U6837 ( .C1(n5707), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5706), .B(n5705), .ZN(n5708) );
  INV_X1 U6838 ( .A(n5708), .ZN(U2999) );
  AND3_X1 U6839 ( .A1(n4187), .A2(n4177), .A3(n4176), .ZN(n5709) );
  INV_X1 U6840 ( .A(n5709), .ZN(n5711) );
  AOI22_X1 U6841 ( .A1(n5710), .A2(n5709), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n4164), .ZN(n5888) );
  AOI21_X1 U6842 ( .B1(n3139), .B2(n5711), .A(n5888), .ZN(n5713) );
  XNOR2_X1 U6843 ( .A(n5713), .B(n4175), .ZN(n5881) );
  INV_X1 U6844 ( .A(n5881), .ZN(n5719) );
  INV_X1 U6845 ( .A(n5963), .ZN(n5717) );
  NOR3_X1 U6846 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n4177), .A3(n5900), 
        .ZN(n5716) );
  OAI22_X1 U6847 ( .A1(n5714), .A2(n4175), .B1(n6349), .B2(n6563), .ZN(n5715)
         );
  AOI211_X1 U6848 ( .C1(n5717), .C2(n6323), .A(n5716), .B(n5715), .ZN(n5718)
         );
  OAI21_X1 U6849 ( .B1(n5719), .B2(n5913), .A(n5718), .ZN(U3000) );
  OAI21_X1 U6850 ( .B1(n6351), .B2(n5721), .A(n5720), .ZN(n5722) );
  AOI21_X1 U6851 ( .B1(n6356), .B2(n5723), .A(n5722), .ZN(n5729) );
  INV_X1 U6852 ( .A(n5910), .ZN(n5726) );
  INV_X1 U6853 ( .A(n5724), .ZN(n5725) );
  OAI21_X1 U6854 ( .B1(n5726), .B2(n5725), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5727) );
  NAND3_X1 U6855 ( .A1(n5729), .A2(n5728), .A3(n5727), .ZN(U3018) );
  XNOR2_X1 U6856 ( .A(n5731), .B(n5730), .ZN(n5734) );
  OAI22_X1 U6857 ( .A1(n5734), .A2(n5733), .B1(n4512), .B2(n5732), .ZN(n5735)
         );
  MUX2_X1 U6858 ( .A(n5735), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(n6362), 
        .Z(U3463) );
  AND2_X1 U6859 ( .A1(n3133), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OAI22_X1 U6860 ( .A1(n5737), .A2(n6716), .B1(n6099), .B2(n5736), .ZN(n5738)
         );
  INV_X1 U6861 ( .A(n5738), .ZN(n5745) );
  AOI22_X1 U6862 ( .A1(n6087), .A2(n5740), .B1(n6070), .B2(n5739), .ZN(n5744)
         );
  INV_X1 U6863 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6578) );
  NAND3_X1 U6864 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5773), .ZN(n5763) );
  NOR2_X1 U6865 ( .A1(n6578), .A2(n5763), .ZN(n5746) );
  INV_X1 U6866 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6582) );
  NAND3_X1 U6867 ( .A1(REIP_REG_30__SCAN_IN), .A2(n5746), .A3(n6582), .ZN(
        n5743) );
  NAND2_X1 U6868 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5741) );
  OAI21_X1 U6869 ( .B1(n5741), .B2(n5783), .A(n6063), .ZN(n5768) );
  OAI211_X1 U6870 ( .C1(REIP_REG_29__SCAN_IN), .C2(n6004), .A(
        REIP_REG_30__SCAN_IN), .B(n5768), .ZN(n5747) );
  NAND3_X1 U6871 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6063), .A3(n5747), .ZN(
        n5742) );
  NAND4_X1 U6872 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(U2796)
         );
  AOI22_X1 U6873 ( .A1(n6112), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6110), .ZN(n5757) );
  INV_X1 U6874 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5754) );
  INV_X1 U6875 ( .A(n5747), .ZN(n5753) );
  INV_X1 U6876 ( .A(n5746), .ZN(n5752) );
  OAI22_X1 U6877 ( .A1(n5749), .A2(n6123), .B1(n6081), .B2(n5748), .ZN(n5750)
         );
  INV_X1 U6878 ( .A(n5750), .ZN(n5751) );
  OAI221_X1 U6879 ( .B1(n5754), .B2(n5753), .C1(n5752), .C2(n5753), .A(n5751), 
        .ZN(n5755) );
  INV_X1 U6880 ( .A(n5755), .ZN(n5756) );
  OAI211_X1 U6881 ( .C1(n5758), .C2(n6108), .A(n5757), .B(n5756), .ZN(U2797)
         );
  AOI22_X1 U6882 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6110), .B1(n5759), 
        .B2(n6120), .ZN(n5760) );
  OAI21_X1 U6883 ( .B1(n6578), .B2(n5768), .A(n5760), .ZN(n5761) );
  AOI21_X1 U6884 ( .B1(EBX_REG_29__SCAN_IN), .B2(n6112), .A(n5761), .ZN(n5762)
         );
  OAI21_X1 U6885 ( .B1(n5763), .B2(REIP_REG_29__SCAN_IN), .A(n5762), .ZN(n5764) );
  AOI21_X1 U6886 ( .B1(n5765), .B2(n6070), .A(n5764), .ZN(n5766) );
  OAI21_X1 U6887 ( .B1(n5767), .B2(n6123), .A(n5766), .ZN(U2798) );
  AOI22_X1 U6888 ( .A1(n6112), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6110), .ZN(n5777) );
  OAI22_X1 U6889 ( .A1(n5769), .A2(n6108), .B1(n6862), .B2(n5768), .ZN(n5770)
         );
  INV_X1 U6890 ( .A(n5770), .ZN(n5776) );
  AOI22_X1 U6891 ( .A1(n5772), .A2(n6070), .B1(n5771), .B2(n6087), .ZN(n5775)
         );
  NAND3_X1 U6892 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5773), .A3(n6862), .ZN(
        n5774) );
  NAND4_X1 U6893 ( .A1(n5777), .A2(n5776), .A3(n5775), .A4(n5774), .ZN(U2799)
         );
  INV_X1 U6894 ( .A(n5778), .ZN(n5779) );
  OAI22_X1 U6895 ( .A1(n5779), .A2(n6108), .B1(n6073), .B2(n5401), .ZN(n5780)
         );
  AOI21_X1 U6896 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6110), .A(n5780), 
        .ZN(n5786) );
  NAND2_X1 U6897 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5793) );
  OAI21_X1 U6898 ( .B1(n5781), .B2(n5793), .A(n6857), .ZN(n5782) );
  AOI22_X1 U6899 ( .A1(n5784), .A2(n6087), .B1(n5783), .B2(n5782), .ZN(n5785)
         );
  OAI211_X1 U6900 ( .C1(n5787), .C2(n6081), .A(n5786), .B(n5785), .ZN(U2801)
         );
  OAI22_X1 U6901 ( .A1(n6073), .A2(n6795), .B1(n6099), .B2(n5788), .ZN(n5791)
         );
  INV_X1 U6902 ( .A(n5864), .ZN(n5789) );
  OAI22_X1 U6903 ( .A1(n5811), .A2(n5658), .B1(n5789), .B2(n6108), .ZN(n5790)
         );
  AOI211_X1 U6904 ( .C1(n5792), .C2(n6070), .A(n5791), .B(n5790), .ZN(n5795)
         );
  OAI211_X1 U6905 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5800), .B(n5793), .ZN(n5794) );
  OAI211_X1 U6906 ( .C1(n6123), .C2(n5796), .A(n5795), .B(n5794), .ZN(U2802)
         );
  AOI22_X1 U6907 ( .A1(n6112), .A2(EBX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6110), .ZN(n5797) );
  OAI21_X1 U6908 ( .B1(n5811), .B2(n6703), .A(n5797), .ZN(n5798) );
  AOI21_X1 U6909 ( .B1(n5799), .B2(n6120), .A(n5798), .ZN(n5803) );
  AOI22_X1 U6910 ( .A1(n6087), .A2(n5801), .B1(n5800), .B2(n6703), .ZN(n5802)
         );
  OAI211_X1 U6911 ( .C1(n5804), .C2(n6081), .A(n5803), .B(n5802), .ZN(U2803)
         );
  INV_X1 U6912 ( .A(n5805), .ZN(n5806) );
  AOI22_X1 U6913 ( .A1(n6120), .A2(n5806), .B1(EBX_REG_23__SCAN_IN), .B2(n6112), .ZN(n5815) );
  INV_X1 U6914 ( .A(n5807), .ZN(n5813) );
  NAND2_X1 U6915 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5819) );
  INV_X1 U6916 ( .A(n5819), .ZN(n5808) );
  AOI21_X1 U6917 ( .B1(n5829), .B2(n5808), .A(REIP_REG_23__SCAN_IN), .ZN(n5810) );
  OAI22_X1 U6918 ( .A1(n5811), .A2(n5810), .B1(n5809), .B2(n6123), .ZN(n5812)
         );
  AOI21_X1 U6919 ( .B1(n5813), .B2(n6070), .A(n5812), .ZN(n5814) );
  OAI211_X1 U6920 ( .C1(n6785), .C2(n6099), .A(n5815), .B(n5814), .ZN(U2804)
         );
  AOI22_X1 U6921 ( .A1(n6112), .A2(EBX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6110), .ZN(n5823) );
  INV_X1 U6922 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6901) );
  OAI22_X1 U6923 ( .A1(n5816), .A2(n6108), .B1(n6901), .B2(n5842), .ZN(n5817)
         );
  INV_X1 U6924 ( .A(n5817), .ZN(n5822) );
  AOI22_X1 U6925 ( .A1(n5856), .A2(n6070), .B1(n5818), .B2(n6087), .ZN(n5821)
         );
  OAI211_X1 U6926 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5829), .B(n5819), .ZN(n5820) );
  NAND4_X1 U6927 ( .A1(n5823), .A2(n5822), .A3(n5821), .A4(n5820), .ZN(U2805)
         );
  INV_X1 U6928 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6568) );
  AOI22_X1 U6929 ( .A1(n6120), .A2(n5824), .B1(EBX_REG_21__SCAN_IN), .B2(n6112), .ZN(n5825) );
  OAI21_X1 U6930 ( .B1(n5826), .B2(n6099), .A(n5825), .ZN(n5827) );
  AOI221_X1 U6931 ( .B1(n5829), .B2(n6568), .C1(n5828), .C2(
        REIP_REG_21__SCAN_IN), .A(n5827), .ZN(n5832) );
  AOI22_X1 U6932 ( .A1(n5859), .A2(n6070), .B1(n5830), .B2(n6087), .ZN(n5831)
         );
  NAND2_X1 U6933 ( .A1(n5832), .A2(n5831), .ZN(U2806) );
  INV_X1 U6934 ( .A(n5833), .ZN(n5839) );
  OAI22_X1 U6935 ( .A1(n6081), .A2(n5835), .B1(n6073), .B2(n5834), .ZN(n5838)
         );
  INV_X1 U6936 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5836) );
  OAI22_X1 U6937 ( .A1(n5836), .A2(n6099), .B1(n5873), .B2(n6108), .ZN(n5837)
         );
  AOI211_X1 U6938 ( .C1(n6087), .C2(n5839), .A(n5838), .B(n5837), .ZN(n5840)
         );
  OAI221_X1 U6939 ( .B1(n5842), .B2(n6566), .C1(n5842), .C2(n5841), .A(n5840), 
        .ZN(U2807) );
  INV_X1 U6940 ( .A(n5843), .ZN(n5964) );
  NAND2_X1 U6941 ( .A1(n5845), .A2(n6563), .ZN(n5961) );
  NOR2_X1 U6942 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6563), .ZN(n5844) );
  AOI22_X1 U6943 ( .A1(n5874), .A2(n6120), .B1(n5845), .B2(n5844), .ZN(n5846)
         );
  OAI211_X1 U6944 ( .C1(n6099), .C2(n5847), .A(n5846), .B(n6066), .ZN(n5850)
         );
  OAI22_X1 U6945 ( .A1(n5848), .A2(n6123), .B1(n6073), .B2(n5525), .ZN(n5849)
         );
  NOR2_X1 U6946 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  OAI21_X1 U6947 ( .B1(n5880), .B2(n6081), .A(n5851), .ZN(n5852) );
  INV_X1 U6948 ( .A(n5852), .ZN(n5853) );
  OAI221_X1 U6949 ( .B1(n5854), .B2(n5964), .C1(n5854), .C2(n5961), .A(n5853), 
        .ZN(U2808) );
  INV_X1 U6950 ( .A(n5855), .ZN(n6127) );
  AOI22_X1 U6951 ( .A1(n5856), .A2(n6127), .B1(n6948), .B2(DATAI_22_), .ZN(
        n5858) );
  AOI22_X1 U6952 ( .A1(n6947), .A2(EAX_REG_22__SCAN_IN), .B1(n6946), .B2(
        DATAI_6_), .ZN(n5857) );
  NAND2_X1 U6953 ( .A1(n5858), .A2(n5857), .ZN(U2869) );
  AOI22_X1 U6954 ( .A1(n5859), .A2(n6127), .B1(n6948), .B2(DATAI_21_), .ZN(
        n5861) );
  AOI22_X1 U6955 ( .A1(n6947), .A2(EAX_REG_21__SCAN_IN), .B1(n6946), .B2(
        DATAI_5_), .ZN(n5860) );
  NAND2_X1 U6956 ( .A1(n5861), .A2(n5860), .ZN(U2870) );
  AOI22_X1 U6957 ( .A1(n5870), .A2(n6127), .B1(n6948), .B2(DATAI_20_), .ZN(
        n5863) );
  AOI22_X1 U6958 ( .A1(n6947), .A2(EAX_REG_20__SCAN_IN), .B1(n6946), .B2(
        DATAI_4_), .ZN(n5862) );
  NAND2_X1 U6959 ( .A1(n5863), .A2(n5862), .ZN(U2871) );
  AOI22_X1 U6960 ( .A1(n6325), .A2(REIP_REG_25__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5867) );
  AOI22_X1 U6961 ( .A1(n5865), .A2(n6272), .B1(n5864), .B2(n6257), .ZN(n5866)
         );
  OAI211_X1 U6962 ( .C1(n6286), .C2(n5868), .A(n5867), .B(n5866), .ZN(U2961)
         );
  AOI22_X1 U6963 ( .A1(n6325), .A2(REIP_REG_20__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5872) );
  AOI22_X1 U6964 ( .A1(n5870), .A2(n6273), .B1(n6272), .B2(n5869), .ZN(n5871)
         );
  OAI211_X1 U6965 ( .C1(n6280), .C2(n5873), .A(n5872), .B(n5871), .ZN(U2966)
         );
  AOI22_X1 U6966 ( .A1(n6325), .A2(REIP_REG_19__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5879) );
  INV_X1 U6967 ( .A(n5874), .ZN(n5875) );
  OAI22_X1 U6968 ( .A1(n5876), .A2(n6278), .B1(n6280), .B2(n5875), .ZN(n5877)
         );
  INV_X1 U6969 ( .A(n5877), .ZN(n5878) );
  OAI211_X1 U6970 ( .C1(n6286), .C2(n5880), .A(n5879), .B(n5878), .ZN(U2967)
         );
  AOI22_X1 U6971 ( .A1(n6325), .A2(REIP_REG_18__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5883) );
  AOI22_X1 U6972 ( .A1(n6272), .A2(n5881), .B1(n6273), .B2(n6124), .ZN(n5882)
         );
  OAI211_X1 U6973 ( .C1(n6280), .C2(n5958), .A(n5883), .B(n5882), .ZN(U2968)
         );
  AOI22_X1 U6974 ( .A1(n6325), .A2(REIP_REG_17__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5891) );
  MUX2_X1 U6975 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .B(n4177), .S(n4164), 
        .Z(n5885) );
  OAI21_X1 U6976 ( .B1(n5889), .B2(n5886), .A(n5885), .ZN(n5887) );
  OAI21_X1 U6977 ( .B1(n5889), .B2(n5888), .A(n5887), .ZN(n5897) );
  AOI22_X1 U6978 ( .A1(n5897), .A2(n6272), .B1(n6257), .B2(n5966), .ZN(n5890)
         );
  OAI211_X1 U6979 ( .C1(n6286), .C2(n5972), .A(n5891), .B(n5890), .ZN(U2969)
         );
  AOI22_X1 U6980 ( .A1(n6325), .A2(REIP_REG_13__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5895) );
  XNOR2_X1 U6981 ( .A(n5892), .B(n5893), .ZN(n5924) );
  AOI22_X1 U6982 ( .A1(n5924), .A2(n6272), .B1(n6257), .B2(n6012), .ZN(n5894)
         );
  OAI211_X1 U6983 ( .C1(n6286), .C2(n6010), .A(n5895), .B(n5894), .ZN(U2973)
         );
  AOI22_X1 U6984 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5896), .B1(n6325), .B2(REIP_REG_17__SCAN_IN), .ZN(n5899) );
  AOI22_X1 U6985 ( .A1(n5897), .A2(n6356), .B1(n6323), .B2(n5970), .ZN(n5898)
         );
  OAI211_X1 U6986 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5900), .A(n5899), .B(n5898), .ZN(U3001) );
  INV_X1 U6987 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5977) );
  OAI22_X1 U6988 ( .A1(n5901), .A2(n5913), .B1(n6351), .B2(n5982), .ZN(n5902)
         );
  AOI21_X1 U6989 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n5903), .A(n5902), 
        .ZN(n5907) );
  OAI211_X1 U6990 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5905), .B(n5904), .ZN(n5906) );
  OAI211_X1 U6991 ( .C1(n5977), .C2(n6349), .A(n5907), .B(n5906), .ZN(U3002)
         );
  NOR2_X1 U6992 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5908), .ZN(n5921)
         );
  OAI21_X1 U6993 ( .B1(n6353), .B2(n5911), .A(n5908), .ZN(n5909) );
  OAI211_X1 U6994 ( .C1(n5918), .C2(n5910), .A(n6294), .B(n5909), .ZN(n5923)
         );
  AOI221_X1 U6995 ( .B1(n5912), .B2(n5921), .C1(n5911), .C2(n5921), .A(n5923), 
        .ZN(n5920) );
  NOR2_X1 U6996 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6288), .ZN(n5917)
         );
  NOR2_X1 U6997 ( .A1(n6349), .A2(n6819), .ZN(n5916) );
  OAI22_X1 U6998 ( .A1(n5914), .A2(n5913), .B1(n6351), .B2(n5994), .ZN(n5915)
         );
  AOI211_X1 U6999 ( .C1(n5918), .C2(n5917), .A(n5916), .B(n5915), .ZN(n5919)
         );
  OAI21_X1 U7000 ( .B1(n5920), .B2(n5354), .A(n5919), .ZN(U3004) );
  INV_X1 U7001 ( .A(n5921), .ZN(n5927) );
  OAI22_X1 U7002 ( .A1(n6351), .A2(n6006), .B1(n6349), .B2(n6920), .ZN(n5922)
         );
  INV_X1 U7003 ( .A(n5922), .ZN(n5926) );
  AOI22_X1 U7004 ( .A1(n5924), .A2(n6356), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5923), .ZN(n5925) );
  OAI211_X1 U7005 ( .C1(n6288), .C2(n5927), .A(n5926), .B(n5925), .ZN(U3005)
         );
  NAND3_X1 U7006 ( .A1(n5930), .A2(n5929), .A3(n5928), .ZN(n5931) );
  OAI22_X1 U7007 ( .A1(n5932), .A2(n5931), .B1(n4592), .B2(n6598), .ZN(U3455)
         );
  INV_X1 U7008 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6535) );
  AOI21_X1 U7009 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6535), .A(n6529), .ZN(n5937) );
  INV_X1 U7010 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5933) );
  NAND2_X2 U7011 ( .A1(n6529), .A2(STATE_REG_1__SCAN_IN), .ZN(n6623) );
  INV_X1 U7012 ( .A(n6623), .ZN(n6622) );
  AOI21_X1 U7013 ( .B1(n5937), .B2(n5933), .A(n6622), .ZN(U2789) );
  OAI21_X1 U7014 ( .B1(n5934), .B2(n6510), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5935) );
  OAI21_X1 U7015 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6511), .A(n5935), .ZN(
        U2790) );
  NOR2_X1 U7016 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5938) );
  OAI21_X1 U7017 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5938), .A(n6623), .ZN(n5936)
         );
  OAI21_X1 U7018 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6623), .A(n5936), .ZN(
        U2791) );
  NOR2_X1 U7019 ( .A1(n6622), .A2(n5937), .ZN(n6588) );
  OAI21_X1 U7020 ( .B1(n5938), .B2(BS16_N), .A(n6588), .ZN(n6586) );
  OAI21_X1 U7021 ( .B1(n6588), .B2(n5939), .A(n6586), .ZN(U2792) );
  OAI21_X1 U7022 ( .B1(n5941), .B2(n5940), .A(n6278), .ZN(U2793) );
  NOR4_X1 U7023 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5945) );
  NOR4_X1 U7024 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(
        n5944) );
  NOR4_X1 U7025 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5943) );
  NOR4_X1 U7026 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n5942) );
  NAND4_X1 U7027 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n5951)
         );
  NOR4_X1 U7028 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_8__SCAN_IN), .ZN(n5949) );
  AOI211_X1 U7029 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_13__SCAN_IN), .B(
        DATAWIDTH_REG_4__SCAN_IN), .ZN(n5948) );
  NOR4_X1 U7030 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n5947) );
  NOR4_X1 U7031 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5946) );
  NAND4_X1 U7032 ( .A1(n5949), .A2(n5948), .A3(n5947), .A4(n5946), .ZN(n5950)
         );
  NOR2_X1 U7033 ( .A1(n5951), .A2(n5950), .ZN(n6609) );
  INV_X1 U7034 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5953) );
  NOR3_X1 U7035 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5954) );
  OAI21_X1 U7036 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5954), .A(n6609), .ZN(n5952)
         );
  OAI21_X1 U7037 ( .B1(n6609), .B2(n5953), .A(n5952), .ZN(U2794) );
  INV_X1 U7038 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6587) );
  AOI21_X1 U7039 ( .B1(n6602), .B2(n6587), .A(n5954), .ZN(n5956) );
  INV_X1 U7040 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5955) );
  INV_X1 U7041 ( .A(n6609), .ZN(n6604) );
  AOI22_X1 U7042 ( .A1(n6609), .A2(n5956), .B1(n5955), .B2(n6604), .ZN(U2795)
         );
  NAND2_X1 U7043 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n6110), .ZN(n5957)
         );
  OAI211_X1 U7044 ( .C1(n6108), .C2(n5958), .A(n6066), .B(n5957), .ZN(n5960)
         );
  OAI22_X1 U7045 ( .A1(n5964), .A2(n6563), .B1(n6073), .B2(n6730), .ZN(n5959)
         );
  AOI211_X1 U7046 ( .C1(n6070), .C2(n6124), .A(n5960), .B(n5959), .ZN(n5962)
         );
  OAI211_X1 U7047 ( .C1(n5963), .C2(n6123), .A(n5962), .B(n5961), .ZN(U2809)
         );
  AOI21_X1 U7048 ( .B1(n6561), .B2(n5965), .A(n5964), .ZN(n5969) );
  AOI22_X1 U7049 ( .A1(n6120), .A2(n5966), .B1(EBX_REG_17__SCAN_IN), .B2(n6112), .ZN(n5967) );
  OAI211_X1 U7050 ( .C1(n6099), .C2(n6904), .A(n5967), .B(n6066), .ZN(n5968)
         );
  AOI211_X1 U7051 ( .C1(n5970), .C2(n6087), .A(n5969), .B(n5968), .ZN(n5971)
         );
  OAI21_X1 U7052 ( .B1(n6081), .B2(n5972), .A(n5971), .ZN(U2810) );
  INV_X1 U7053 ( .A(n5998), .ZN(n5976) );
  AOI21_X1 U7054 ( .B1(n6110), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6083), 
        .ZN(n5975) );
  AOI22_X1 U7055 ( .A1(n6120), .A2(n5973), .B1(EBX_REG_16__SCAN_IN), .B2(n6112), .ZN(n5974) );
  OAI211_X1 U7056 ( .C1(n5977), .C2(n5976), .A(n5975), .B(n5974), .ZN(n5978)
         );
  AOI21_X1 U7057 ( .B1(n6070), .B2(n6128), .A(n5978), .ZN(n5981) );
  OAI211_X1 U7058 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n5990), .B(n5979), .ZN(n5980) );
  OAI211_X1 U7059 ( .C1(n5982), .C2(n6123), .A(n5981), .B(n5980), .ZN(U2811)
         );
  AOI22_X1 U7060 ( .A1(n5984), .A2(n6120), .B1(n6070), .B2(n5983), .ZN(n5992)
         );
  INV_X1 U7061 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6558) );
  INV_X1 U7062 ( .A(n5985), .ZN(n5986) );
  AOI22_X1 U7063 ( .A1(n5986), .A2(n6087), .B1(EBX_REG_15__SCAN_IN), .B2(n6112), .ZN(n5987) );
  OAI211_X1 U7064 ( .C1(n6099), .C2(n5988), .A(n5987), .B(n6066), .ZN(n5989)
         );
  AOI221_X1 U7065 ( .B1(n5990), .B2(n6558), .C1(n5998), .C2(
        REIP_REG_15__SCAN_IN), .A(n5989), .ZN(n5991) );
  NAND2_X1 U7066 ( .A1(n5992), .A2(n5991), .ZN(U2812) );
  OAI21_X1 U7067 ( .B1(n6099), .B2(n5993), .A(n6066), .ZN(n5996) );
  NOR2_X1 U7068 ( .A1(n5994), .A2(n6123), .ZN(n5995) );
  AOI211_X1 U7069 ( .C1(EBX_REG_14__SCAN_IN), .C2(n6112), .A(n5996), .B(n5995), 
        .ZN(n6001) );
  OAI21_X1 U7070 ( .B1(n6920), .B2(n6014), .A(n6819), .ZN(n5997) );
  AOI22_X1 U7071 ( .A1(n5999), .A2(n6120), .B1(n5998), .B2(n5997), .ZN(n6000)
         );
  OAI211_X1 U7072 ( .C1(n6081), .C2(n6002), .A(n6001), .B(n6000), .ZN(U2813)
         );
  NOR3_X1 U7073 ( .A1(n6004), .A2(n6003), .A3(n6920), .ZN(n6005) );
  AOI211_X1 U7074 ( .C1(n6110), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6083), 
        .B(n6005), .ZN(n6009) );
  INV_X1 U7075 ( .A(n6006), .ZN(n6007) );
  AOI22_X1 U7076 ( .A1(n6007), .A2(n6087), .B1(EBX_REG_13__SCAN_IN), .B2(n6112), .ZN(n6008) );
  OAI211_X1 U7077 ( .C1(n6081), .C2(n6010), .A(n6009), .B(n6008), .ZN(n6011)
         );
  AOI21_X1 U7078 ( .B1(n6012), .B2(n6120), .A(n6011), .ZN(n6013) );
  OAI21_X1 U7079 ( .B1(REIP_REG_13__SCAN_IN), .B2(n6014), .A(n6013), .ZN(U2814) );
  AND2_X1 U7080 ( .A1(n6015), .A2(n6063), .ZN(n6029) );
  AOI22_X1 U7081 ( .A1(n6029), .A2(REIP_REG_12__SCAN_IN), .B1(
        EBX_REG_12__SCAN_IN), .B2(n6112), .ZN(n6023) );
  OAI22_X1 U7082 ( .A1(n6842), .A2(n6099), .B1(n6123), .B2(n6016), .ZN(n6017)
         );
  AOI211_X1 U7083 ( .C1(n6018), .C2(n6694), .A(n6083), .B(n6017), .ZN(n6022)
         );
  AOI22_X1 U7084 ( .A1(n6020), .A2(n6120), .B1(n6070), .B2(n6019), .ZN(n6021)
         );
  NAND3_X1 U7085 ( .A1(n6023), .A2(n6022), .A3(n6021), .ZN(U2815) );
  INV_X1 U7086 ( .A(n6024), .ZN(n6287) );
  OAI22_X1 U7087 ( .A1(n6073), .A2(n6877), .B1(n6099), .B2(n6025), .ZN(n6026)
         );
  AOI211_X1 U7088 ( .C1(n6087), .C2(n6287), .A(n6083), .B(n6026), .ZN(n6031)
         );
  INV_X1 U7089 ( .A(n6032), .ZN(n6027) );
  OAI21_X1 U7090 ( .B1(n6027), .B2(n6551), .A(n6553), .ZN(n6028) );
  AOI22_X1 U7091 ( .A1(n6210), .A2(n6120), .B1(n6029), .B2(n6028), .ZN(n6030)
         );
  OAI211_X1 U7092 ( .C1(n6081), .C2(n6213), .A(n6031), .B(n6030), .ZN(U2816)
         );
  AOI22_X1 U7093 ( .A1(n6032), .A2(n6551), .B1(EBX_REG_10__SCAN_IN), .B2(n6112), .ZN(n6041) );
  INV_X1 U7094 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6549) );
  NOR2_X1 U7095 ( .A1(n6096), .A2(n6033), .ZN(n6050) );
  OR2_X1 U7096 ( .A1(n6109), .A2(n6050), .ZN(n6052) );
  AOI21_X1 U7097 ( .B1(n6044), .B2(n6549), .A(n6052), .ZN(n6035) );
  OAI22_X1 U7098 ( .A1(n6035), .A2(n6551), .B1(n6123), .B2(n6034), .ZN(n6036)
         );
  AOI211_X1 U7099 ( .C1(n6110), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6083), 
        .B(n6036), .ZN(n6040) );
  AOI22_X1 U7100 ( .A1(n6038), .A2(n6120), .B1(n6070), .B2(n6037), .ZN(n6039)
         );
  NAND3_X1 U7101 ( .A1(n6041), .A2(n6040), .A3(n6039), .ZN(U2817) );
  INV_X1 U7102 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6047) );
  INV_X1 U7103 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6042) );
  OAI22_X1 U7104 ( .A1(n6296), .A2(n6123), .B1(n6073), .B2(n6042), .ZN(n6043)
         );
  INV_X1 U7105 ( .A(n6043), .ZN(n6046) );
  AOI221_X1 U7106 ( .B1(n6044), .B2(n6549), .C1(n6052), .C2(
        REIP_REG_9__SCAN_IN), .A(n6083), .ZN(n6045) );
  OAI211_X1 U7107 ( .C1(n6047), .C2(n6099), .A(n6046), .B(n6045), .ZN(n6048)
         );
  AOI21_X1 U7108 ( .B1(n6218), .B2(n6120), .A(n6048), .ZN(n6049) );
  OAI21_X1 U7109 ( .B1(n6081), .B2(n6221), .A(n6049), .ZN(U2818) );
  AOI22_X1 U7110 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6052), .B1(n6051), .B2(n6050), .ZN(n6056) );
  AOI22_X1 U7111 ( .A1(n6112), .A2(EBX_REG_8__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n6110), .ZN(n6053) );
  OAI211_X1 U7112 ( .C1(n6123), .C2(n6305), .A(n6053), .B(n6066), .ZN(n6054)
         );
  AOI21_X1 U7113 ( .B1(n6226), .B2(n6120), .A(n6054), .ZN(n6055) );
  OAI211_X1 U7114 ( .C1(n6081), .C2(n6229), .A(n6056), .B(n6055), .ZN(U2819)
         );
  AND2_X1 U7115 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6082), .ZN(n6057) );
  NAND2_X1 U7116 ( .A1(n6111), .A2(n6057), .ZN(n6078) );
  INV_X1 U7117 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6910) );
  INV_X1 U7118 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U7119 ( .A1(n6910), .A2(n6545), .ZN(n6059) );
  NAND2_X1 U7120 ( .A1(n6059), .A2(n6058), .ZN(n6061) );
  NAND2_X1 U7121 ( .A1(n6112), .A2(EBX_REG_7__SCAN_IN), .ZN(n6060) );
  OAI21_X1 U7122 ( .B1(n6078), .B2(n6061), .A(n6060), .ZN(n6062) );
  INV_X1 U7123 ( .A(n6062), .ZN(n6072) );
  INV_X1 U7124 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6065) );
  OAI21_X1 U7125 ( .B1(n6109), .B2(n6064), .A(n6063), .ZN(n6091) );
  OAI22_X1 U7126 ( .A1(n6065), .A2(n6099), .B1(n6910), .B2(n6091), .ZN(n6069)
         );
  OAI21_X1 U7127 ( .B1(n6123), .B2(n6067), .A(n6066), .ZN(n6068) );
  AOI211_X1 U7128 ( .C1(n6070), .C2(n6234), .A(n6069), .B(n6068), .ZN(n6071)
         );
  OAI211_X1 U7129 ( .C1(n6237), .C2(n6108), .A(n6072), .B(n6071), .ZN(U2820)
         );
  OAI22_X1 U7130 ( .A1(n6075), .A2(n6123), .B1(n6074), .B2(n6073), .ZN(n6076)
         );
  AOI211_X1 U7131 ( .C1(n6110), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6083), 
        .B(n6076), .ZN(n6077) );
  OAI221_X1 U7132 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6078), .C1(n6545), .C2(
        n6091), .A(n6077), .ZN(n6079) );
  AOI21_X1 U7133 ( .B1(n6239), .B2(n6120), .A(n6079), .ZN(n6080) );
  OAI21_X1 U7134 ( .B1(n6081), .B2(n6243), .A(n6080), .ZN(U2821) );
  AOI21_X1 U7135 ( .B1(n6111), .B2(n6082), .A(REIP_REG_5__SCAN_IN), .ZN(n6090)
         );
  NAND2_X1 U7136 ( .A1(n6112), .A2(EBX_REG_5__SCAN_IN), .ZN(n6085) );
  AOI21_X1 U7137 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n6110), .A(n6083), 
        .ZN(n6084) );
  NAND2_X1 U7138 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  AOI21_X1 U7139 ( .B1(n6322), .B2(n6087), .A(n6086), .ZN(n6089) );
  INV_X1 U7140 ( .A(n6116), .ZN(n6105) );
  NAND2_X1 U7141 ( .A1(n6248), .A2(n6105), .ZN(n6088) );
  OAI211_X1 U7142 ( .C1(n6091), .C2(n6090), .A(n6089), .B(n6088), .ZN(n6092)
         );
  INV_X1 U7143 ( .A(n6092), .ZN(n6093) );
  OAI21_X1 U7144 ( .B1(n6251), .B2(n6108), .A(n6093), .ZN(U2822) );
  INV_X1 U7145 ( .A(n6094), .ZN(n6095) );
  NOR2_X1 U7146 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  AOI22_X1 U7147 ( .A1(n6098), .A2(n6097), .B1(EBX_REG_3__SCAN_IN), .B2(n6112), 
        .ZN(n6107) );
  INV_X1 U7148 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6540) );
  INV_X1 U7149 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6895) );
  OAI22_X1 U7150 ( .A1(n6338), .A2(n6123), .B1(n6099), .B2(n6895), .ZN(n6100)
         );
  AOI21_X1 U7151 ( .B1(n6368), .B2(n6101), .A(n6100), .ZN(n6102) );
  OAI21_X1 U7152 ( .B1(n6103), .B2(n6540), .A(n6102), .ZN(n6104) );
  AOI21_X1 U7153 ( .B1(n6265), .B2(n6105), .A(n6104), .ZN(n6106) );
  OAI211_X1 U7154 ( .C1(n6268), .C2(n6108), .A(n6107), .B(n6106), .ZN(U2824)
         );
  AOI22_X1 U7155 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6110), .B1(n6109), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6122) );
  INV_X1 U7156 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6119) );
  AOI22_X1 U7157 ( .A1(n6112), .A2(EBX_REG_1__SCAN_IN), .B1(n6111), .B2(n6602), 
        .ZN(n6113) );
  OAI21_X1 U7158 ( .B1(n6115), .B2(n6114), .A(n6113), .ZN(n6118) );
  NOR2_X1 U7159 ( .A1(n6116), .A2(n6285), .ZN(n6117) );
  AOI211_X1 U7160 ( .C1(n6120), .C2(n6119), .A(n6118), .B(n6117), .ZN(n6121)
         );
  OAI211_X1 U7161 ( .C1(n4463), .C2(n6123), .A(n6122), .B(n6121), .ZN(U2826)
         );
  AOI22_X1 U7162 ( .A1(n6124), .A2(n6127), .B1(n6948), .B2(DATAI_18_), .ZN(
        n6126) );
  AOI22_X1 U7163 ( .A1(n6947), .A2(EAX_REG_18__SCAN_IN), .B1(n6946), .B2(
        DATAI_2_), .ZN(n6125) );
  NAND2_X1 U7164 ( .A1(n6126), .A2(n6125), .ZN(U2873) );
  AOI22_X1 U7165 ( .A1(n6128), .A2(n6127), .B1(n6948), .B2(DATAI_16_), .ZN(
        n6130) );
  AOI22_X1 U7166 ( .A1(n6947), .A2(EAX_REG_16__SCAN_IN), .B1(n6946), .B2(
        DATAI_0_), .ZN(n6129) );
  NAND2_X1 U7167 ( .A1(n6130), .A2(n6129), .ZN(U2875) );
  INV_X1 U7168 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6719) );
  INV_X1 U7169 ( .A(n6131), .ZN(n6132) );
  AOI22_X1 U7170 ( .A1(n6132), .A2(EAX_REG_20__SCAN_IN), .B1(
        UWORD_REG_4__SCAN_IN), .B2(n6614), .ZN(n6133) );
  OAI21_X1 U7171 ( .B1(n6719), .B2(n6134), .A(n6133), .ZN(U2903) );
  AOI22_X1 U7172 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n6614), .B1(n3133), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6136) );
  OAI21_X1 U7173 ( .B1(n6137), .B2(n6164), .A(n6136), .ZN(U2908) );
  INV_X1 U7174 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6139) );
  AOI22_X1 U7175 ( .A1(n6614), .A2(LWORD_REG_14__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6138) );
  OAI21_X1 U7176 ( .B1(n6139), .B2(n6164), .A(n6138), .ZN(U2909) );
  INV_X1 U7177 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6141) );
  AOI22_X1 U7178 ( .A1(n6614), .A2(LWORD_REG_13__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7179 ( .B1(n6141), .B2(n6164), .A(n6140), .ZN(U2910) );
  INV_X1 U7180 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6143) );
  AOI22_X1 U7181 ( .A1(DATAO_REG_12__SCAN_IN), .A2(n3133), .B1(n6159), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6142) );
  OAI21_X1 U7182 ( .B1(n6143), .B2(n6164), .A(n6142), .ZN(U2911) );
  INV_X1 U7183 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6145) );
  AOI22_X1 U7184 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6614), .B1(n3133), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6144) );
  OAI21_X1 U7185 ( .B1(n6145), .B2(n6164), .A(n6144), .ZN(U2912) );
  AOI22_X1 U7186 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6614), .B1(n3133), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6146) );
  OAI21_X1 U7187 ( .B1(n6875), .B2(n6164), .A(n6146), .ZN(U2913) );
  AOI22_X1 U7188 ( .A1(DATAO_REG_9__SCAN_IN), .A2(n3133), .B1(
        LWORD_REG_9__SCAN_IN), .B2(n6159), .ZN(n6147) );
  OAI21_X1 U7189 ( .B1(n6678), .B2(n6164), .A(n6147), .ZN(U2914) );
  AOI22_X1 U7190 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6614), .B1(n3133), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6148) );
  OAI21_X1 U7191 ( .B1(n6149), .B2(n6164), .A(n6148), .ZN(U2915) );
  AOI22_X1 U7192 ( .A1(n6614), .A2(LWORD_REG_7__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6150) );
  OAI21_X1 U7193 ( .B1(n6151), .B2(n6164), .A(n6150), .ZN(U2916) );
  AOI22_X1 U7194 ( .A1(DATAO_REG_6__SCAN_IN), .A2(n3133), .B1(
        LWORD_REG_6__SCAN_IN), .B2(n6159), .ZN(n6152) );
  OAI21_X1 U7195 ( .B1(n6153), .B2(n6164), .A(n6152), .ZN(U2917) );
  AOI22_X1 U7196 ( .A1(n6614), .A2(LWORD_REG_5__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6154) );
  OAI21_X1 U7197 ( .B1(n6155), .B2(n6164), .A(n6154), .ZN(U2918) );
  AOI22_X1 U7198 ( .A1(n6614), .A2(LWORD_REG_4__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6156) );
  OAI21_X1 U7199 ( .B1(n6698), .B2(n6164), .A(n6156), .ZN(U2919) );
  AOI22_X1 U7200 ( .A1(n6614), .A2(LWORD_REG_3__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6157) );
  OAI21_X1 U7201 ( .B1(n6158), .B2(n6164), .A(n6157), .ZN(U2920) );
  AOI22_X1 U7202 ( .A1(DATAO_REG_2__SCAN_IN), .A2(n3133), .B1(n6159), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n6160) );
  OAI21_X1 U7203 ( .B1(n6161), .B2(n6164), .A(n6160), .ZN(U2921) );
  AOI22_X1 U7204 ( .A1(n6614), .A2(LWORD_REG_1__SCAN_IN), .B1(n3133), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6162) );
  OAI21_X1 U7205 ( .B1(n6704), .B2(n6164), .A(n6162), .ZN(U2922) );
  AOI22_X1 U7206 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6614), .B1(
        DATAO_REG_0__SCAN_IN), .B2(n3133), .ZN(n6163) );
  OAI21_X1 U7207 ( .B1(n6165), .B2(n6164), .A(n6163), .ZN(U2923) );
  AOI22_X1 U7208 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6167) );
  OAI21_X1 U7209 ( .B1(n6194), .B2(n6177), .A(n6167), .ZN(U2924) );
  AOI22_X1 U7210 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6168) );
  OAI21_X1 U7211 ( .B1(n6194), .B2(n6179), .A(n6168), .ZN(U2925) );
  AOI22_X1 U7212 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6169) );
  OAI21_X1 U7213 ( .B1(n6194), .B2(n6181), .A(n6169), .ZN(U2926) );
  AOI22_X1 U7214 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6170) );
  OAI21_X1 U7215 ( .B1(n6194), .B2(n6183), .A(n6170), .ZN(U2927) );
  AOI22_X1 U7216 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6171) );
  OAI21_X1 U7217 ( .B1(n6194), .B2(n6186), .A(n6171), .ZN(U2928) );
  AOI22_X1 U7218 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6172) );
  OAI21_X1 U7219 ( .B1(n6194), .B2(n6188), .A(n6172), .ZN(U2929) );
  AOI22_X1 U7220 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6173) );
  OAI21_X1 U7221 ( .B1(n6194), .B2(n6815), .A(n6173), .ZN(U2930) );
  AOI22_X1 U7222 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6174) );
  OAI21_X1 U7223 ( .B1(n6194), .B2(n6191), .A(n6174), .ZN(U2931) );
  AOI22_X1 U7224 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6175) );
  OAI21_X1 U7225 ( .B1(n6194), .B2(n6193), .A(n6175), .ZN(U2933) );
  AOI22_X1 U7226 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6184), .B1(n6201), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n6176) );
  OAI21_X1 U7227 ( .B1(n6194), .B2(n6177), .A(n6176), .ZN(U2939) );
  AOI22_X1 U7228 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6184), .B1(n6201), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n6178) );
  OAI21_X1 U7229 ( .B1(n6194), .B2(n6179), .A(n6178), .ZN(U2940) );
  AOI22_X1 U7230 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6184), .B1(n6201), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n6180) );
  OAI21_X1 U7231 ( .B1(n6194), .B2(n6181), .A(n6180), .ZN(U2941) );
  AOI22_X1 U7232 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6184), .B1(n6201), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n6182) );
  OAI21_X1 U7233 ( .B1(n6194), .B2(n6183), .A(n6182), .ZN(U2942) );
  AOI22_X1 U7234 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6184), .B1(n6201), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n6185) );
  OAI21_X1 U7235 ( .B1(n6194), .B2(n6186), .A(n6185), .ZN(U2943) );
  AOI22_X1 U7236 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n6187) );
  OAI21_X1 U7237 ( .B1(n6194), .B2(n6188), .A(n6187), .ZN(U2944) );
  AOI22_X1 U7238 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n6189) );
  OAI21_X1 U7239 ( .B1(n6194), .B2(n6815), .A(n6189), .ZN(U2945) );
  AOI22_X1 U7240 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n6190) );
  OAI21_X1 U7241 ( .B1(n6194), .B2(n6191), .A(n6190), .ZN(U2946) );
  AOI22_X1 U7242 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n6192) );
  OAI21_X1 U7243 ( .B1(n6194), .B2(n6193), .A(n6192), .ZN(U2948) );
  AOI22_X1 U7244 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7245 ( .A1(n6203), .A2(DATAI_11_), .ZN(n6195) );
  NAND2_X1 U7246 ( .A1(n6196), .A2(n6195), .ZN(U2950) );
  AOI22_X1 U7247 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7248 ( .A1(n6203), .A2(DATAI_12_), .ZN(n6197) );
  NAND2_X1 U7249 ( .A1(n6198), .A2(n6197), .ZN(U2951) );
  AOI22_X1 U7250 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7251 ( .A1(n6203), .A2(DATAI_13_), .ZN(n6199) );
  NAND2_X1 U7252 ( .A1(n6200), .A2(n6199), .ZN(U2952) );
  AOI22_X1 U7253 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6202), .B1(n6201), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7254 ( .A1(n6203), .A2(DATAI_14_), .ZN(n6204) );
  NAND2_X1 U7255 ( .A1(n6205), .A2(n6204), .ZN(U2953) );
  AOI22_X1 U7256 ( .A1(n6325), .A2(REIP_REG_11__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7257 ( .A1(n6206), .A2(n6207), .ZN(n6209) );
  XNOR2_X1 U7258 ( .A(n4164), .B(n6293), .ZN(n6208) );
  XNOR2_X1 U7259 ( .A(n6209), .B(n6208), .ZN(n6290) );
  AOI22_X1 U7260 ( .A1(n6272), .A2(n6290), .B1(n6257), .B2(n6210), .ZN(n6211)
         );
  OAI211_X1 U7261 ( .C1(n6286), .C2(n6213), .A(n6212), .B(n6211), .ZN(U2975)
         );
  AOI22_X1 U7262 ( .A1(n6325), .A2(REIP_REG_9__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7263 ( .A1(n6216), .A2(n6215), .ZN(n6217) );
  XNOR2_X1 U7264 ( .A(n6214), .B(n6217), .ZN(n6299) );
  AOI22_X1 U7265 ( .A1(n6299), .A2(n6272), .B1(n6257), .B2(n6218), .ZN(n6219)
         );
  OAI211_X1 U7266 ( .C1(n6286), .C2(n6221), .A(n6220), .B(n6219), .ZN(U2977)
         );
  AOI22_X1 U7267 ( .A1(n6325), .A2(REIP_REG_8__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6228) );
  OAI21_X1 U7268 ( .B1(n6222), .B2(n6224), .A(n6223), .ZN(n6225) );
  INV_X1 U7269 ( .A(n6225), .ZN(n6308) );
  AOI22_X1 U7270 ( .A1(n6308), .A2(n6272), .B1(n6257), .B2(n6226), .ZN(n6227)
         );
  OAI211_X1 U7271 ( .C1(n6286), .C2(n6229), .A(n6228), .B(n6227), .ZN(U2978)
         );
  AOI22_X1 U7272 ( .A1(n6325), .A2(REIP_REG_7__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6236) );
  OR2_X1 U7273 ( .A1(n6231), .A2(n6230), .ZN(n6232) );
  AND2_X1 U7274 ( .A1(n6233), .A2(n6232), .ZN(n6311) );
  AOI22_X1 U7275 ( .A1(n6234), .A2(n6273), .B1(n6272), .B2(n6311), .ZN(n6235)
         );
  OAI211_X1 U7276 ( .C1(n6280), .C2(n6237), .A(n6236), .B(n6235), .ZN(U2979)
         );
  AOI22_X1 U7277 ( .A1(n6325), .A2(REIP_REG_6__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6242) );
  INV_X1 U7278 ( .A(n6238), .ZN(n6240) );
  AOI22_X1 U7279 ( .A1(n6240), .A2(n6272), .B1(n6257), .B2(n6239), .ZN(n6241)
         );
  OAI211_X1 U7280 ( .C1(n6286), .C2(n6243), .A(n6242), .B(n6241), .ZN(U2980)
         );
  AOI22_X1 U7281 ( .A1(n6325), .A2(REIP_REG_5__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6250) );
  OAI21_X1 U7282 ( .B1(n6246), .B2(n6245), .A(n3137), .ZN(n6247) );
  INV_X1 U7283 ( .A(n6247), .ZN(n6324) );
  AOI22_X1 U7284 ( .A1(n6324), .A2(n6272), .B1(n6273), .B2(n6248), .ZN(n6249)
         );
  OAI211_X1 U7285 ( .C1(n6280), .C2(n6251), .A(n6250), .B(n6249), .ZN(U2981)
         );
  AOI22_X1 U7286 ( .A1(n6325), .A2(REIP_REG_4__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7287 ( .B1(n6254), .B2(n6253), .A(n3136), .ZN(n6255) );
  INV_X1 U7288 ( .A(n6255), .ZN(n6332) );
  AOI22_X1 U7289 ( .A1(n6332), .A2(n6272), .B1(n6257), .B2(n6256), .ZN(n6258)
         );
  OAI211_X1 U7290 ( .C1(n6286), .C2(n6260), .A(n6259), .B(n6258), .ZN(U2982)
         );
  AOI22_X1 U7291 ( .A1(n6325), .A2(REIP_REG_3__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6267) );
  OAI21_X1 U7292 ( .B1(n6262), .B2(n6263), .A(n6261), .ZN(n6264) );
  INV_X1 U7293 ( .A(n6264), .ZN(n6340) );
  AOI22_X1 U7294 ( .A1(n6340), .A2(n6272), .B1(n6265), .B2(n6273), .ZN(n6266)
         );
  OAI211_X1 U7295 ( .C1(n6280), .C2(n6268), .A(n6267), .B(n6266), .ZN(U2983)
         );
  AOI22_X1 U7296 ( .A1(n6325), .A2(REIP_REG_2__SCAN_IN), .B1(n6283), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6276) );
  XNOR2_X1 U7297 ( .A(n6269), .B(n6360), .ZN(n6270) );
  XNOR2_X1 U7298 ( .A(n6271), .B(n6270), .ZN(n6357) );
  AOI22_X1 U7299 ( .A1(n6274), .A2(n6273), .B1(n6272), .B2(n6357), .ZN(n6275)
         );
  OAI211_X1 U7300 ( .C1(n6280), .C2(n6277), .A(n6276), .B(n6275), .ZN(U2984)
         );
  OAI22_X1 U7301 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6279), 
        .B2(n6278), .ZN(n6281) );
  AOI211_X1 U7302 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6283), .A(n6282), 
        .B(n6281), .ZN(n6284) );
  OAI21_X1 U7303 ( .B1(n6286), .B2(n6285), .A(n6284), .ZN(U2985) );
  AOI22_X1 U7304 ( .A1(n6323), .A2(n6287), .B1(n6325), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6292) );
  INV_X1 U7305 ( .A(n6288), .ZN(n6289) );
  AOI22_X1 U7306 ( .A1(n6356), .A2(n6290), .B1(n6293), .B2(n6289), .ZN(n6291)
         );
  OAI211_X1 U7307 ( .C1(n6294), .C2(n6293), .A(n6292), .B(n6291), .ZN(U3007)
         );
  INV_X1 U7308 ( .A(n6295), .ZN(n6303) );
  OAI22_X1 U7309 ( .A1(n6351), .A2(n6296), .B1(n6349), .B2(n6549), .ZN(n6297)
         );
  INV_X1 U7310 ( .A(n6297), .ZN(n6301) );
  AOI22_X1 U7311 ( .A1(n6299), .A2(n6356), .B1(n6298), .B2(n6302), .ZN(n6300)
         );
  OAI211_X1 U7312 ( .C1(n6303), .C2(n6302), .A(n6301), .B(n6300), .ZN(U3009)
         );
  AOI211_X1 U7313 ( .C1(n6315), .C2(n6310), .A(n6304), .B(n6316), .ZN(n6307)
         );
  INV_X1 U7314 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6817) );
  OAI22_X1 U7315 ( .A1(n6351), .A2(n6305), .B1(n6817), .B2(n6349), .ZN(n6306)
         );
  AOI211_X1 U7316 ( .C1(n6308), .C2(n6356), .A(n6307), .B(n6306), .ZN(n6309)
         );
  OAI21_X1 U7317 ( .B1(n6314), .B2(n6310), .A(n6309), .ZN(U3010) );
  AOI222_X1 U7318 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6325), .B1(n6323), .B2(
        n6312), .C1(n6356), .C2(n6311), .ZN(n6313) );
  OAI221_X1 U7319 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n6316), .C1(n6315), .C2(n6314), .A(n6313), .ZN(U3011) );
  OAI21_X1 U7320 ( .B1(n6319), .B2(n6318), .A(n6317), .ZN(n6320) );
  AOI21_X1 U7321 ( .B1(n6353), .B2(n6321), .A(n6320), .ZN(n6328) );
  AOI22_X1 U7322 ( .A1(n6324), .A2(n6356), .B1(n6323), .B2(n6322), .ZN(n6327)
         );
  NAND2_X1 U7323 ( .A1(n6325), .A2(REIP_REG_5__SCAN_IN), .ZN(n6326) );
  OAI211_X1 U7324 ( .C1(n6329), .C2(n6328), .A(n6327), .B(n6326), .ZN(U3013)
         );
  AOI21_X1 U7325 ( .B1(n6353), .B2(n6352), .A(n6347), .ZN(n6345) );
  OAI22_X1 U7326 ( .A1(n6351), .A2(n6330), .B1(n6542), .B2(n6349), .ZN(n6331)
         );
  AOI21_X1 U7327 ( .B1(n6332), .B2(n6356), .A(n6331), .ZN(n6336) );
  NOR2_X1 U7328 ( .A1(n6352), .A2(n6333), .ZN(n6341) );
  OAI211_X1 U7329 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6341), .B(n6334), .ZN(n6335) );
  OAI211_X1 U7330 ( .C1(n6345), .C2(n6337), .A(n6336), .B(n6335), .ZN(U3014)
         );
  OAI22_X1 U7331 ( .A1(n6351), .A2(n6338), .B1(n6349), .B2(n6540), .ZN(n6339)
         );
  INV_X1 U7332 ( .A(n6339), .ZN(n6343) );
  AOI22_X1 U7333 ( .A1(n6341), .A2(n6344), .B1(n6340), .B2(n6356), .ZN(n6342)
         );
  OAI211_X1 U7334 ( .C1(n6345), .C2(n6344), .A(n6343), .B(n6342), .ZN(U3015)
         );
  NAND2_X1 U7335 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6346), .ZN(n6361)
         );
  AOI21_X1 U7336 ( .B1(n6353), .B2(n6348), .A(n6347), .ZN(n6359) );
  OAI22_X1 U7337 ( .A1(n6351), .A2(n6350), .B1(n6538), .B2(n6349), .ZN(n6355)
         );
  AND2_X1 U7338 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  AOI211_X1 U7339 ( .C1(n6357), .C2(n6356), .A(n6355), .B(n6354), .ZN(n6358)
         );
  OAI221_X1 U7340 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6361), .C1(n6360), .C2(n6359), .A(n6358), .ZN(U3016) );
  AND2_X1 U7341 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6362), .ZN(U3019)
         );
  NOR2_X1 U7342 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6363), .ZN(n6412)
         );
  INV_X1 U7343 ( .A(n6364), .ZN(n6369) );
  NAND3_X1 U7344 ( .A1(n6366), .A2(n6365), .A3(n6485), .ZN(n6367) );
  OAI21_X1 U7345 ( .B1(n6369), .B2(n6368), .A(n6367), .ZN(n6411) );
  AOI22_X1 U7346 ( .A1(n6439), .A2(n6412), .B1(n6440), .B2(n6411), .ZN(n6381)
         );
  NAND3_X1 U7347 ( .A1(n6436), .A2(n6371), .A3(n6370), .ZN(n6374) );
  AOI21_X1 U7348 ( .B1(n6374), .B2(n6373), .A(n6372), .ZN(n6378) );
  OAI211_X1 U7349 ( .C1(n3296), .C2(n6412), .A(n6375), .B(n6485), .ZN(n6376)
         );
  AOI22_X1 U7350 ( .A1(n6415), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6379), 
        .B2(n6413), .ZN(n6380) );
  OAI211_X1 U7351 ( .C1(n6382), .C2(n6436), .A(n6381), .B(n6380), .ZN(U3068)
         );
  AOI22_X1 U7352 ( .A1(n6384), .A2(n6412), .B1(n6383), .B2(n6411), .ZN(n6387)
         );
  AOI22_X1 U7353 ( .A1(n6415), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6385), 
        .B2(n6413), .ZN(n6386) );
  OAI211_X1 U7354 ( .C1(n6388), .C2(n6436), .A(n6387), .B(n6386), .ZN(U3069)
         );
  AOI22_X1 U7355 ( .A1(n6445), .A2(n6412), .B1(n6446), .B2(n6411), .ZN(n6391)
         );
  AOI22_X1 U7356 ( .A1(n6415), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6389), 
        .B2(n6413), .ZN(n6390) );
  OAI211_X1 U7357 ( .C1(n6392), .C2(n6436), .A(n6391), .B(n6390), .ZN(U3070)
         );
  AOI22_X1 U7358 ( .A1(n6451), .A2(n6412), .B1(n6452), .B2(n6411), .ZN(n6395)
         );
  AOI22_X1 U7359 ( .A1(n6415), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6393), 
        .B2(n6413), .ZN(n6394) );
  OAI211_X1 U7360 ( .C1(n6396), .C2(n6436), .A(n6395), .B(n6394), .ZN(U3071)
         );
  AOI22_X1 U7361 ( .A1(n6457), .A2(n6412), .B1(n6458), .B2(n6411), .ZN(n6399)
         );
  AOI22_X1 U7362 ( .A1(n6415), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6397), 
        .B2(n6413), .ZN(n6398) );
  OAI211_X1 U7363 ( .C1(n6400), .C2(n6436), .A(n6399), .B(n6398), .ZN(U3072)
         );
  AOI22_X1 U7364 ( .A1(n6465), .A2(n6412), .B1(n6467), .B2(n6411), .ZN(n6403)
         );
  AOI22_X1 U7365 ( .A1(n6415), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6401), 
        .B2(n6413), .ZN(n6402) );
  OAI211_X1 U7366 ( .C1(n6404), .C2(n6436), .A(n6403), .B(n6402), .ZN(U3073)
         );
  AOI22_X1 U7367 ( .A1(n6406), .A2(n6412), .B1(n6405), .B2(n6411), .ZN(n6409)
         );
  AOI22_X1 U7368 ( .A1(n6415), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6407), 
        .B2(n6413), .ZN(n6408) );
  OAI211_X1 U7369 ( .C1(n6410), .C2(n6436), .A(n6409), .B(n6408), .ZN(U3074)
         );
  AOI22_X1 U7370 ( .A1(n6428), .A2(n6412), .B1(n6432), .B2(n6411), .ZN(n6417)
         );
  AOI22_X1 U7371 ( .A1(n6415), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6414), 
        .B2(n6413), .ZN(n6416) );
  OAI211_X1 U7372 ( .C1(n6418), .C2(n6436), .A(n6417), .B(n6416), .ZN(U3075)
         );
  INV_X1 U7373 ( .A(n6419), .ZN(n6430) );
  INV_X1 U7374 ( .A(n6420), .ZN(n6427) );
  AOI22_X1 U7375 ( .A1(n6430), .A2(n6438), .B1(n6439), .B2(n6427), .ZN(n6422)
         );
  AOI22_X1 U7376 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6433), .B1(n6440), 
        .B2(n6431), .ZN(n6421) );
  OAI211_X1 U7377 ( .C1(n6443), .C2(n6436), .A(n6422), .B(n6421), .ZN(U3076)
         );
  AOI22_X1 U7378 ( .A1(n6430), .A2(n6444), .B1(n6445), .B2(n6427), .ZN(n6424)
         );
  AOI22_X1 U7379 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6433), .B1(n6446), 
        .B2(n6431), .ZN(n6423) );
  OAI211_X1 U7380 ( .C1(n6449), .C2(n6436), .A(n6424), .B(n6423), .ZN(U3078)
         );
  AOI22_X1 U7381 ( .A1(n6430), .A2(n6450), .B1(n6451), .B2(n6427), .ZN(n6426)
         );
  AOI22_X1 U7382 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6433), .B1(n6452), 
        .B2(n6431), .ZN(n6425) );
  OAI211_X1 U7383 ( .C1(n6455), .C2(n6436), .A(n6426), .B(n6425), .ZN(U3079)
         );
  AOI22_X1 U7384 ( .A1(n6430), .A2(n6429), .B1(n6428), .B2(n6427), .ZN(n6435)
         );
  AOI22_X1 U7385 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6433), .B1(n6432), 
        .B2(n6431), .ZN(n6434) );
  OAI211_X1 U7386 ( .C1(n6437), .C2(n6436), .A(n6435), .B(n6434), .ZN(U3083)
         );
  AOI22_X1 U7387 ( .A1(n6439), .A2(n6464), .B1(n6463), .B2(n6438), .ZN(n6442)
         );
  AOI22_X1 U7388 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6468), .B1(n6440), 
        .B2(n6466), .ZN(n6441) );
  OAI211_X1 U7389 ( .C1(n6443), .C2(n6471), .A(n6442), .B(n6441), .ZN(U3108)
         );
  AOI22_X1 U7390 ( .A1(n6445), .A2(n6464), .B1(n6463), .B2(n6444), .ZN(n6448)
         );
  AOI22_X1 U7391 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6468), .B1(n6446), 
        .B2(n6466), .ZN(n6447) );
  OAI211_X1 U7392 ( .C1(n6449), .C2(n6471), .A(n6448), .B(n6447), .ZN(U3110)
         );
  AOI22_X1 U7393 ( .A1(n6451), .A2(n6464), .B1(n6463), .B2(n6450), .ZN(n6454)
         );
  AOI22_X1 U7394 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6468), .B1(n6452), 
        .B2(n6466), .ZN(n6453) );
  OAI211_X1 U7395 ( .C1(n6455), .C2(n6471), .A(n6454), .B(n6453), .ZN(U3111)
         );
  AOI22_X1 U7396 ( .A1(n6457), .A2(n6464), .B1(n6463), .B2(n6456), .ZN(n6460)
         );
  AOI22_X1 U7397 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6468), .B1(n6458), 
        .B2(n6466), .ZN(n6459) );
  OAI211_X1 U7398 ( .C1(n6461), .C2(n6471), .A(n6460), .B(n6459), .ZN(U3112)
         );
  AOI22_X1 U7399 ( .A1(n6465), .A2(n6464), .B1(n6463), .B2(n6462), .ZN(n6470)
         );
  AOI22_X1 U7400 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6468), .B1(n6467), 
        .B2(n6466), .ZN(n6469) );
  OAI211_X1 U7401 ( .C1(n6472), .C2(n6471), .A(n6470), .B(n6469), .ZN(U3113)
         );
  INV_X1 U7402 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6593) );
  AOI22_X1 U7403 ( .A1(n6475), .A2(n6474), .B1(n6473), .B2(n6593), .ZN(n6596)
         );
  NAND2_X1 U7404 ( .A1(n6476), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6601) );
  AND3_X1 U7405 ( .A1(n6596), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6601), 
        .ZN(n6477) );
  NAND2_X1 U7406 ( .A1(n6477), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6481) );
  OAI22_X1 U7407 ( .A1(n6479), .A2(n6478), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6477), .ZN(n6480) );
  NAND2_X1 U7408 ( .A1(n6481), .A2(n6480), .ZN(n6482) );
  AOI222_X1 U7409 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6483), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6482), .C1(n6483), .C2(n6482), 
        .ZN(n6484) );
  AOI222_X1 U7410 ( .A1(n6486), .A2(n6485), .B1(n6486), .B2(n6484), .C1(n6485), 
        .C2(n6484), .ZN(n6487) );
  NOR2_X1 U7411 ( .A1(n6487), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6495)
         );
  OAI21_X1 U7412 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6488), 
        .ZN(n6491) );
  NAND3_X1 U7413 ( .A1(n6491), .A2(n6490), .A3(n6489), .ZN(n6492) );
  NOR4_X1 U7414 ( .A1(n6495), .A2(n6494), .A3(n6493), .A4(n6492), .ZN(n6508)
         );
  INV_X1 U7415 ( .A(n6496), .ZN(n6500) );
  NOR3_X1 U7416 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .A3(n6524), .ZN(
        n6499) );
  AOI21_X1 U7417 ( .B1(STATE2_REG_1__SCAN_IN), .B2(READY_N), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6498) );
  AOI211_X1 U7418 ( .C1(n6500), .C2(n6499), .A(n6498), .B(n6497), .ZN(n6504)
         );
  OAI221_X1 U7419 ( .B1(n3350), .B2(n6508), .C1(n3350), .C2(n6501), .A(n6504), 
        .ZN(n6591) );
  OAI21_X1 U7420 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6613), .A(n6591), .ZN(
        n6509) );
  AOI221_X1 U7421 ( .B1(n6503), .B2(STATE2_REG_0__SCAN_IN), .C1(n6509), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6502), .ZN(n6507) );
  AOI211_X1 U7422 ( .C1(n6617), .C2(n6592), .A(STATE2_REG_0__SCAN_IN), .B(
        n6504), .ZN(n6505) );
  INV_X1 U7423 ( .A(n6505), .ZN(n6506) );
  OAI211_X1 U7424 ( .C1(n6508), .C2(n6510), .A(n6507), .B(n6506), .ZN(U3148)
         );
  OAI211_X1 U7425 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6509), .ZN(n6515) );
  OAI21_X1 U7426 ( .B1(READY_N), .B2(n6511), .A(n6510), .ZN(n6513) );
  AOI21_X1 U7427 ( .B1(n6513), .B2(n6591), .A(n6512), .ZN(n6514) );
  NAND2_X1 U7428 ( .A1(n6515), .A2(n6514), .ZN(U3149) );
  OAI221_X1 U7429 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6613), .A(n6589), .ZN(n6517) );
  OAI21_X1 U7430 ( .B1(n6617), .B2(n6517), .A(n6516), .ZN(U3150) );
  AND2_X1 U7431 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6518), .ZN(U3151) );
  INV_X1 U7432 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6823) );
  NOR2_X1 U7433 ( .A1(n6588), .A2(n6823), .ZN(U3152) );
  AND2_X1 U7434 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6518), .ZN(U3153) );
  AND2_X1 U7435 ( .A1(n6518), .A2(DATAWIDTH_REG_28__SCAN_IN), .ZN(U3154) );
  AND2_X1 U7436 ( .A1(n6518), .A2(DATAWIDTH_REG_27__SCAN_IN), .ZN(U3155) );
  AND2_X1 U7437 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6518), .ZN(U3156) );
  AND2_X1 U7438 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6518), .ZN(U3157) );
  AND2_X1 U7439 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6518), .ZN(U3158) );
  AND2_X1 U7440 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6518), .ZN(U3159) );
  INV_X1 U7441 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6748) );
  NOR2_X1 U7442 ( .A1(n6588), .A2(n6748), .ZN(U3160) );
  AND2_X1 U7443 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6518), .ZN(U3161) );
  AND2_X1 U7444 ( .A1(n6518), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  AND2_X1 U7445 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6518), .ZN(U3163) );
  AND2_X1 U7446 ( .A1(n6518), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  AND2_X1 U7447 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6518), .ZN(U3165) );
  AND2_X1 U7448 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6518), .ZN(U3166) );
  AND2_X1 U7449 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6518), .ZN(U3167) );
  AND2_X1 U7450 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6518), .ZN(U3168) );
  AND2_X1 U7451 ( .A1(n6518), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  AND2_X1 U7452 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6518), .ZN(U3170) );
  INV_X1 U7453 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6681) );
  NOR2_X1 U7454 ( .A1(n6588), .A2(n6681), .ZN(U3171) );
  AND2_X1 U7455 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6518), .ZN(U3172) );
  AND2_X1 U7456 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6518), .ZN(U3173) );
  INV_X1 U7457 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6829) );
  NOR2_X1 U7458 ( .A1(n6588), .A2(n6829), .ZN(U3174) );
  AND2_X1 U7459 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6518), .ZN(U3175) );
  AND2_X1 U7460 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6518), .ZN(U3176) );
  AND2_X1 U7461 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6518), .ZN(U3177) );
  AND2_X1 U7462 ( .A1(n6518), .A2(DATAWIDTH_REG_4__SCAN_IN), .ZN(U3178) );
  AND2_X1 U7463 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6518), .ZN(U3179) );
  AND2_X1 U7464 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6518), .ZN(U3180) );
  NOR2_X1 U7465 ( .A1(n6535), .A2(n6525), .ZN(n6526) );
  AOI22_X1 U7466 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6534) );
  AND2_X1 U7467 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6522) );
  INV_X1 U7468 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6520) );
  INV_X1 U7469 ( .A(NA_N), .ZN(n6527) );
  AOI221_X1 U7470 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6527), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6531) );
  AOI221_X1 U7471 ( .B1(n6522), .B2(n6623), .C1(n6520), .C2(n6623), .A(n6531), 
        .ZN(n6519) );
  OAI21_X1 U7472 ( .B1(n6526), .B2(n6534), .A(n6519), .ZN(U3181) );
  NOR2_X1 U7473 ( .A1(n6529), .A2(n6520), .ZN(n6528) );
  NAND2_X1 U7474 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6521) );
  OAI21_X1 U7475 ( .B1(n6528), .B2(n6522), .A(n6521), .ZN(n6523) );
  OAI211_X1 U7476 ( .C1(n6525), .C2(n6613), .A(n6524), .B(n6523), .ZN(U3182)
         );
  AOI21_X1 U7477 ( .B1(n6528), .B2(n6527), .A(n6526), .ZN(n6533) );
  AOI221_X1 U7478 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6613), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6530) );
  AOI221_X1 U7479 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6530), .C2(HOLD), .A(n6529), .ZN(n6532) );
  OAI22_X1 U7480 ( .A1(n6534), .A2(n6533), .B1(n6532), .B2(n6531), .ZN(U3183)
         );
  OR2_X1 U7481 ( .A1(n6623), .A2(STATE_REG_2__SCAN_IN), .ZN(n6581) );
  NOR2_X1 U7482 ( .A1(n6535), .A2(n6623), .ZN(n6579) );
  AOI222_X1 U7483 ( .A1(n3134), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6623), .C1(REIP_REG_1__SCAN_IN), .C2(
        n6579), .ZN(n6536) );
  INV_X1 U7484 ( .A(n6536), .ZN(U3184) );
  AOI22_X1 U7485 ( .A1(REIP_REG_3__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6623), .ZN(n6537) );
  OAI21_X1 U7486 ( .B1(n6538), .B2(n6577), .A(n6537), .ZN(U3185) );
  AOI22_X1 U7487 ( .A1(REIP_REG_4__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6623), .ZN(n6539) );
  OAI21_X1 U7488 ( .B1(n6540), .B2(n6577), .A(n6539), .ZN(U3186) );
  AOI22_X1 U7489 ( .A1(REIP_REG_5__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6623), .ZN(n6541) );
  OAI21_X1 U7490 ( .B1(n6542), .B2(n6577), .A(n6541), .ZN(U3187) );
  AOI222_X1 U7491 ( .A1(n3134), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6623), .C1(REIP_REG_5__SCAN_IN), .C2(
        n6579), .ZN(n6543) );
  INV_X1 U7492 ( .A(n6543), .ZN(U3188) );
  AOI22_X1 U7493 ( .A1(REIP_REG_7__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6623), .ZN(n6544) );
  OAI21_X1 U7494 ( .B1(n6545), .B2(n6577), .A(n6544), .ZN(U3189) );
  AOI22_X1 U7495 ( .A1(REIP_REG_8__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6623), .ZN(n6546) );
  OAI21_X1 U7496 ( .B1(n6910), .B2(n6577), .A(n6546), .ZN(U3190) );
  AOI222_X1 U7497 ( .A1(n6579), .A2(REIP_REG_8__SCAN_IN), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6623), .C1(REIP_REG_9__SCAN_IN), .C2(
        n3134), .ZN(n6547) );
  INV_X1 U7498 ( .A(n6547), .ZN(U3191) );
  AOI22_X1 U7499 ( .A1(REIP_REG_10__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6623), .ZN(n6548) );
  OAI21_X1 U7500 ( .B1(n6549), .B2(n6577), .A(n6548), .ZN(U3192) );
  AOI22_X1 U7501 ( .A1(REIP_REG_11__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6623), .ZN(n6550) );
  OAI21_X1 U7502 ( .B1(n6551), .B2(n6577), .A(n6550), .ZN(U3193) );
  AOI22_X1 U7503 ( .A1(REIP_REG_12__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6623), .ZN(n6552) );
  OAI21_X1 U7504 ( .B1(n6553), .B2(n6577), .A(n6552), .ZN(U3194) );
  AOI22_X1 U7505 ( .A1(REIP_REG_13__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6623), .ZN(n6554) );
  OAI21_X1 U7506 ( .B1(n6694), .B2(n6577), .A(n6554), .ZN(U3195) );
  AOI22_X1 U7507 ( .A1(REIP_REG_14__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6623), .ZN(n6555) );
  OAI21_X1 U7508 ( .B1(n6920), .B2(n6577), .A(n6555), .ZN(U3196) );
  AOI22_X1 U7509 ( .A1(REIP_REG_15__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6623), .ZN(n6556) );
  OAI21_X1 U7510 ( .B1(n6819), .B2(n6577), .A(n6556), .ZN(U3197) );
  AOI22_X1 U7511 ( .A1(REIP_REG_16__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6623), .ZN(n6557) );
  OAI21_X1 U7512 ( .B1(n6558), .B2(n6577), .A(n6557), .ZN(U3198) );
  AOI222_X1 U7513 ( .A1(n6579), .A2(REIP_REG_16__SCAN_IN), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6623), .C1(REIP_REG_17__SCAN_IN), .C2(
        n3134), .ZN(n6559) );
  INV_X1 U7514 ( .A(n6559), .ZN(U3199) );
  AOI22_X1 U7515 ( .A1(REIP_REG_18__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6623), .ZN(n6560) );
  OAI21_X1 U7516 ( .B1(n6561), .B2(n6577), .A(n6560), .ZN(U3200) );
  AOI22_X1 U7517 ( .A1(REIP_REG_19__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6623), .ZN(n6562) );
  OAI21_X1 U7518 ( .B1(n6563), .B2(n6577), .A(n6562), .ZN(U3201) );
  AOI222_X1 U7519 ( .A1(n6579), .A2(REIP_REG_19__SCAN_IN), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6623), .C1(REIP_REG_20__SCAN_IN), .C2(
        n3134), .ZN(n6564) );
  INV_X1 U7520 ( .A(n6564), .ZN(U3202) );
  AOI22_X1 U7521 ( .A1(REIP_REG_21__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6623), .ZN(n6565) );
  OAI21_X1 U7522 ( .B1(n6566), .B2(n6577), .A(n6565), .ZN(U3203) );
  AOI22_X1 U7523 ( .A1(REIP_REG_22__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6623), .ZN(n6567) );
  OAI21_X1 U7524 ( .B1(n6568), .B2(n6577), .A(n6567), .ZN(U3204) );
  AOI22_X1 U7525 ( .A1(REIP_REG_23__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6623), .ZN(n6569) );
  OAI21_X1 U7526 ( .B1(n6901), .B2(n6577), .A(n6569), .ZN(U3205) );
  AOI22_X1 U7527 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6579), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6623), .ZN(n6570) );
  OAI21_X1 U7528 ( .B1(n6703), .B2(n6581), .A(n6570), .ZN(U3206) );
  AOI222_X1 U7529 ( .A1(n3134), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6623), .C1(REIP_REG_24__SCAN_IN), .C2(
        n6579), .ZN(n6571) );
  INV_X1 U7530 ( .A(n6571), .ZN(U3207) );
  AOI22_X1 U7531 ( .A1(REIP_REG_26__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6623), .ZN(n6572) );
  OAI21_X1 U7532 ( .B1(n5658), .B2(n6577), .A(n6572), .ZN(U3208) );
  AOI222_X1 U7533 ( .A1(n6579), .A2(REIP_REG_26__SCAN_IN), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6623), .C1(REIP_REG_27__SCAN_IN), .C2(
        n3134), .ZN(n6573) );
  INV_X1 U7534 ( .A(n6573), .ZN(U3209) );
  AOI222_X1 U7535 ( .A1(n6579), .A2(REIP_REG_27__SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6623), .C1(REIP_REG_28__SCAN_IN), .C2(
        n3134), .ZN(n6574) );
  INV_X1 U7536 ( .A(n6574), .ZN(U3210) );
  AOI22_X1 U7537 ( .A1(REIP_REG_29__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6623), .ZN(n6575) );
  OAI21_X1 U7538 ( .B1(n6862), .B2(n6577), .A(n6575), .ZN(U3211) );
  AOI22_X1 U7539 ( .A1(REIP_REG_30__SCAN_IN), .A2(n3134), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6623), .ZN(n6576) );
  OAI21_X1 U7540 ( .B1(n6578), .B2(n6577), .A(n6576), .ZN(U3212) );
  AOI22_X1 U7541 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6579), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6623), .ZN(n6580) );
  OAI21_X1 U7542 ( .B1(n6582), .B2(n6581), .A(n6580), .ZN(U3213) );
  MUX2_X1 U7543 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6623), .Z(U3445) );
  OAI22_X1 U7544 ( .A1(n6623), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        BE_N_REG_2__SCAN_IN), .B2(n6622), .ZN(n6583) );
  INV_X1 U7545 ( .A(n6583), .ZN(U3446) );
  MUX2_X1 U7546 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6623), .Z(U3447) );
  OAI22_X1 U7547 ( .A1(n6623), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        BE_N_REG_0__SCAN_IN), .B2(n6622), .ZN(n6584) );
  INV_X1 U7548 ( .A(n6584), .ZN(U3448) );
  OAI21_X1 U7549 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6588), .A(n6586), .ZN(
        n6585) );
  INV_X1 U7550 ( .A(n6585), .ZN(U3451) );
  OAI21_X1 U7551 ( .B1(n6588), .B2(n6587), .A(n6586), .ZN(U3452) );
  OAI211_X1 U7552 ( .C1(n3296), .C2(n6591), .A(n6590), .B(n6589), .ZN(U3453)
         );
  AOI22_X1 U7553 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6594), .B1(n6593), .B2(
        n6592), .ZN(n6595) );
  OAI211_X1 U7554 ( .C1(n6596), .C2(n6600), .A(n6598), .B(n6595), .ZN(n6597)
         );
  OAI21_X1 U7555 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6598), .A(n6597), 
        .ZN(n6599) );
  OAI21_X1 U7556 ( .B1(n6601), .B2(n6600), .A(n6599), .ZN(U3461) );
  AOI21_X1 U7557 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6603) );
  AOI22_X1 U7558 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6603), .B2(n6602), .ZN(n6606) );
  INV_X1 U7559 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6605) );
  AOI22_X1 U7560 ( .A1(n6609), .A2(n6606), .B1(n6605), .B2(n6604), .ZN(U3468)
         );
  INV_X1 U7561 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6608) );
  OAI21_X1 U7562 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6609), .ZN(n6607) );
  OAI21_X1 U7563 ( .B1(n6609), .B2(n6608), .A(n6607), .ZN(U3469) );
  NAND2_X1 U7564 ( .A1(n6623), .A2(W_R_N_REG_SCAN_IN), .ZN(n6610) );
  OAI21_X1 U7565 ( .B1(n6623), .B2(READREQUEST_REG_SCAN_IN), .A(n6610), .ZN(
        U3470) );
  AOI211_X1 U7566 ( .C1(n6614), .C2(n6613), .A(n6612), .B(n6611), .ZN(n6621)
         );
  OAI211_X1 U7567 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6616), .A(n6615), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6618) );
  AOI21_X1 U7568 ( .B1(n6618), .B2(STATE2_REG_0__SCAN_IN), .A(n6617), .ZN(
        n6620) );
  NAND2_X1 U7569 ( .A1(n6621), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6619) );
  OAI21_X1 U7570 ( .B1(n6621), .B2(n6620), .A(n6619), .ZN(U3472) );
  OAI22_X1 U7571 ( .A1(n6623), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n6622), .ZN(n6624) );
  INV_X1 U7572 ( .A(n6624), .ZN(U3473) );
  INV_X1 U7573 ( .A(keyinput126), .ZN(n6625) );
  NAND4_X1 U7574 ( .A1(keyinput32), .A2(keyinput109), .A3(keyinput74), .A4(
        n6625), .ZN(n6626) );
  NOR3_X1 U7575 ( .A1(keyinput17), .A2(keyinput14), .A3(n6626), .ZN(n6638) );
  NAND2_X1 U7576 ( .A1(keyinput115), .A2(keyinput56), .ZN(n6627) );
  NOR3_X1 U7577 ( .A1(keyinput119), .A2(keyinput28), .A3(n6627), .ZN(n6628) );
  NAND3_X1 U7578 ( .A1(keyinput107), .A2(keyinput81), .A3(n6628), .ZN(n6636)
         );
  NAND2_X1 U7579 ( .A1(keyinput54), .A2(keyinput0), .ZN(n6629) );
  NOR3_X1 U7580 ( .A1(keyinput11), .A2(keyinput34), .A3(n6629), .ZN(n6634) );
  NOR4_X1 U7581 ( .A1(keyinput36), .A2(keyinput125), .A3(keyinput9), .A4(
        keyinput117), .ZN(n6633) );
  INV_X1 U7582 ( .A(keyinput73), .ZN(n6811) );
  NOR4_X1 U7583 ( .A1(keyinput48), .A2(keyinput19), .A3(keyinput93), .A4(n6811), .ZN(n6632) );
  NAND2_X1 U7584 ( .A1(keyinput40), .A2(keyinput64), .ZN(n6630) );
  NOR3_X1 U7585 ( .A1(keyinput102), .A2(keyinput99), .A3(n6630), .ZN(n6631) );
  NAND4_X1 U7586 ( .A1(n6634), .A2(n6633), .A3(n6632), .A4(n6631), .ZN(n6635)
         );
  NOR4_X1 U7587 ( .A1(keyinput39), .A2(keyinput27), .A3(n6636), .A4(n6635), 
        .ZN(n6637) );
  NAND4_X1 U7588 ( .A1(keyinput35), .A2(keyinput75), .A3(n6638), .A4(n6637), 
        .ZN(n6676) );
  NOR4_X1 U7589 ( .A1(keyinput105), .A2(keyinput60), .A3(keyinput68), .A4(
        keyinput20), .ZN(n6643) );
  NOR4_X1 U7590 ( .A1(keyinput57), .A2(keyinput49), .A3(keyinput21), .A4(
        keyinput69), .ZN(n6642) );
  NAND2_X1 U7591 ( .A1(keyinput98), .A2(keyinput118), .ZN(n6639) );
  NOR3_X1 U7592 ( .A1(keyinput80), .A2(keyinput100), .A3(n6639), .ZN(n6641) );
  NOR4_X1 U7593 ( .A1(keyinput24), .A2(keyinput116), .A3(keyinput76), .A4(
        keyinput108), .ZN(n6640) );
  NAND4_X1 U7594 ( .A1(n6643), .A2(n6642), .A3(n6641), .A4(n6640), .ZN(n6675)
         );
  NOR4_X1 U7595 ( .A1(keyinput79), .A2(keyinput70), .A3(keyinput67), .A4(
        keyinput62), .ZN(n6647) );
  NOR4_X1 U7596 ( .A1(keyinput110), .A2(keyinput103), .A3(keyinput87), .A4(
        keyinput78), .ZN(n6646) );
  NOR4_X1 U7597 ( .A1(keyinput18), .A2(keyinput3), .A3(keyinput45), .A4(
        keyinput41), .ZN(n6645) );
  NOR4_X1 U7598 ( .A1(keyinput58), .A2(keyinput46), .A3(keyinput30), .A4(
        keyinput31), .ZN(n6644) );
  NAND4_X1 U7599 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6674)
         );
  INV_X1 U7600 ( .A(keyinput92), .ZN(n6894) );
  NAND4_X1 U7601 ( .A1(keyinput90), .A2(keyinput96), .A3(keyinput51), .A4(
        n6894), .ZN(n6652) );
  OR4_X1 U7602 ( .A1(keyinput114), .A2(keyinput97), .A3(keyinput91), .A4(
        keyinput33), .ZN(n6651) );
  INV_X1 U7603 ( .A(keyinput1), .ZN(n6880) );
  NAND4_X1 U7604 ( .A1(keyinput77), .A2(keyinput2), .A3(keyinput50), .A4(n6880), .ZN(n6650) );
  NOR2_X1 U7605 ( .A1(keyinput66), .A2(keyinput38), .ZN(n6648) );
  NAND3_X1 U7606 ( .A1(keyinput88), .A2(keyinput7), .A3(n6648), .ZN(n6649) );
  NOR4_X1 U7607 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n6672)
         );
  NOR2_X1 U7608 ( .A1(keyinput43), .A2(keyinput52), .ZN(n6653) );
  NAND3_X1 U7609 ( .A1(keyinput106), .A2(keyinput72), .A3(n6653), .ZN(n6660)
         );
  NOR2_X1 U7610 ( .A1(keyinput121), .A2(keyinput61), .ZN(n6654) );
  NAND3_X1 U7611 ( .A1(keyinput123), .A2(keyinput55), .A3(n6654), .ZN(n6659)
         );
  NOR2_X1 U7612 ( .A1(keyinput85), .A2(keyinput127), .ZN(n6655) );
  NAND3_X1 U7613 ( .A1(keyinput10), .A2(keyinput83), .A3(n6655), .ZN(n6658) );
  NOR2_X1 U7614 ( .A1(keyinput23), .A2(keyinput26), .ZN(n6656) );
  NAND3_X1 U7615 ( .A1(keyinput122), .A2(keyinput111), .A3(n6656), .ZN(n6657)
         );
  NOR4_X1 U7616 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(n6671)
         );
  NAND4_X1 U7617 ( .A1(keyinput89), .A2(keyinput101), .A3(keyinput44), .A4(
        keyinput4), .ZN(n6664) );
  NAND4_X1 U7618 ( .A1(keyinput25), .A2(keyinput29), .A3(keyinput65), .A4(
        keyinput113), .ZN(n6663) );
  NAND4_X1 U7619 ( .A1(keyinput124), .A2(keyinput104), .A3(keyinput112), .A4(
        keyinput84), .ZN(n6662) );
  NAND4_X1 U7620 ( .A1(keyinput12), .A2(keyinput16), .A3(keyinput8), .A4(
        keyinput120), .ZN(n6661) );
  NOR4_X1 U7621 ( .A1(n6664), .A2(n6663), .A3(n6662), .A4(n6661), .ZN(n6670)
         );
  NAND4_X1 U7622 ( .A1(keyinput63), .A2(keyinput71), .A3(keyinput59), .A4(
        keyinput47), .ZN(n6668) );
  NAND4_X1 U7623 ( .A1(keyinput94), .A2(keyinput95), .A3(keyinput86), .A4(
        keyinput82), .ZN(n6667) );
  NAND4_X1 U7624 ( .A1(keyinput53), .A2(keyinput37), .A3(keyinput13), .A4(
        keyinput5), .ZN(n6666) );
  NAND4_X1 U7625 ( .A1(keyinput42), .A2(keyinput15), .A3(keyinput22), .A4(
        keyinput6), .ZN(n6665) );
  NOR4_X1 U7626 ( .A1(n6668), .A2(n6667), .A3(n6666), .A4(n6665), .ZN(n6669)
         );
  NAND4_X1 U7627 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n6673)
         );
  NOR4_X1 U7628 ( .A1(n6676), .A2(n6675), .A3(n6674), .A4(n6673), .ZN(n6945)
         );
  AOI22_X1 U7629 ( .A1(n6679), .A2(keyinput59), .B1(keyinput22), .B2(n6678), 
        .ZN(n6677) );
  OAI221_X1 U7630 ( .B1(n6679), .B2(keyinput59), .C1(n6678), .C2(keyinput22), 
        .A(n6677), .ZN(n6692) );
  INV_X1 U7631 ( .A(keyinput70), .ZN(n6682) );
  AOI22_X1 U7632 ( .A1(n6682), .A2(ADDRESS_REG_25__SCAN_IN), .B1(keyinput100), 
        .B2(n6681), .ZN(n6680) );
  OAI221_X1 U7633 ( .B1(n6682), .B2(ADDRESS_REG_25__SCAN_IN), .C1(n6681), .C2(
        keyinput100), .A(n6680), .ZN(n6691) );
  INV_X1 U7634 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6685) );
  AOI22_X1 U7635 ( .A1(n6685), .A2(keyinput20), .B1(keyinput5), .B2(n6684), 
        .ZN(n6683) );
  OAI221_X1 U7636 ( .B1(n6685), .B2(keyinput20), .C1(n6684), .C2(keyinput5), 
        .A(n6683), .ZN(n6690) );
  INV_X1 U7637 ( .A(keyinput6), .ZN(n6688) );
  INV_X1 U7638 ( .A(keyinput13), .ZN(n6687) );
  AOI22_X1 U7639 ( .A1(n6688), .A2(ADDRESS_REG_15__SCAN_IN), .B1(
        DATAO_REG_24__SCAN_IN), .B2(n6687), .ZN(n6686) );
  OAI221_X1 U7640 ( .B1(n6688), .B2(ADDRESS_REG_15__SCAN_IN), .C1(n6687), .C2(
        DATAO_REG_24__SCAN_IN), .A(n6686), .ZN(n6689) );
  NOR4_X1 U7641 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n6744)
         );
  AOI22_X1 U7642 ( .A1(n6695), .A2(keyinput110), .B1(keyinput82), .B2(n6694), 
        .ZN(n6693) );
  OAI221_X1 U7643 ( .B1(n6695), .B2(keyinput110), .C1(n6694), .C2(keyinput82), 
        .A(n6693), .ZN(n6708) );
  INV_X1 U7644 ( .A(keyinput4), .ZN(n6697) );
  AOI22_X1 U7645 ( .A1(n6698), .A2(keyinput84), .B1(DATAI_2_), .B2(n6697), 
        .ZN(n6696) );
  OAI221_X1 U7646 ( .B1(n6698), .B2(keyinput84), .C1(n6697), .C2(DATAI_2_), 
        .A(n6696), .ZN(n6707) );
  INV_X1 U7647 ( .A(keyinput30), .ZN(n6700) );
  AOI22_X1 U7648 ( .A1(n6701), .A2(keyinput49), .B1(DATAO_REG_29__SCAN_IN), 
        .B2(n6700), .ZN(n6699) );
  OAI221_X1 U7649 ( .B1(n6701), .B2(keyinput49), .C1(n6700), .C2(
        DATAO_REG_29__SCAN_IN), .A(n6699), .ZN(n6706) );
  AOI22_X1 U7650 ( .A1(n6704), .A2(keyinput63), .B1(n6703), .B2(keyinput47), 
        .ZN(n6702) );
  OAI221_X1 U7651 ( .B1(n6704), .B2(keyinput63), .C1(n6703), .C2(keyinput47), 
        .A(n6702), .ZN(n6705) );
  NOR4_X1 U7652 ( .A1(n6708), .A2(n6707), .A3(n6706), .A4(n6705), .ZN(n6743)
         );
  INV_X1 U7653 ( .A(keyinput57), .ZN(n6711) );
  INV_X1 U7654 ( .A(keyinput69), .ZN(n6710) );
  AOI22_X1 U7655 ( .A1(n6711), .A2(ADDRESS_REG_22__SCAN_IN), .B1(
        DATAWIDTH_REG_18__SCAN_IN), .B2(n6710), .ZN(n6709) );
  OAI221_X1 U7656 ( .B1(n6711), .B2(ADDRESS_REG_22__SCAN_IN), .C1(n6710), .C2(
        DATAWIDTH_REG_18__SCAN_IN), .A(n6709), .ZN(n6724) );
  AOI22_X1 U7657 ( .A1(n6714), .A2(keyinput41), .B1(keyinput94), .B2(n6713), 
        .ZN(n6712) );
  OAI221_X1 U7658 ( .B1(n6714), .B2(keyinput41), .C1(n6713), .C2(keyinput94), 
        .A(n6712), .ZN(n6723) );
  INV_X1 U7659 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6717) );
  AOI22_X1 U7660 ( .A1(n6717), .A2(keyinput60), .B1(keyinput89), .B2(n6716), 
        .ZN(n6715) );
  OAI221_X1 U7661 ( .B1(n6717), .B2(keyinput60), .C1(n6716), .C2(keyinput89), 
        .A(n6715), .ZN(n6722) );
  INV_X1 U7662 ( .A(keyinput21), .ZN(n6720) );
  AOI22_X1 U7663 ( .A1(n6720), .A2(LWORD_REG_11__SCAN_IN), .B1(keyinput118), 
        .B2(n6719), .ZN(n6718) );
  OAI221_X1 U7664 ( .B1(n6720), .B2(LWORD_REG_11__SCAN_IN), .C1(n6719), .C2(
        keyinput118), .A(n6718), .ZN(n6721) );
  NOR4_X1 U7665 ( .A1(n6724), .A2(n6723), .A3(n6722), .A4(n6721), .ZN(n6742)
         );
  INV_X1 U7666 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6727) );
  INV_X1 U7667 ( .A(keyinput108), .ZN(n6726) );
  AOI22_X1 U7668 ( .A1(n6727), .A2(keyinput62), .B1(UWORD_REG_3__SCAN_IN), 
        .B2(n6726), .ZN(n6725) );
  OAI221_X1 U7669 ( .B1(n6727), .B2(keyinput62), .C1(n6726), .C2(
        UWORD_REG_3__SCAN_IN), .A(n6725), .ZN(n6740) );
  INV_X1 U7670 ( .A(keyinput3), .ZN(n6729) );
  AOI22_X1 U7671 ( .A1(n6730), .A2(keyinput113), .B1(UWORD_REG_4__SCAN_IN), 
        .B2(n6729), .ZN(n6728) );
  OAI221_X1 U7672 ( .B1(n6730), .B2(keyinput113), .C1(n6729), .C2(
        UWORD_REG_4__SCAN_IN), .A(n6728), .ZN(n6739) );
  INV_X1 U7673 ( .A(DATAI_30_), .ZN(n6733) );
  INV_X1 U7674 ( .A(keyinput12), .ZN(n6732) );
  AOI22_X1 U7675 ( .A1(n6733), .A2(keyinput37), .B1(UWORD_REG_10__SCAN_IN), 
        .B2(n6732), .ZN(n6731) );
  OAI221_X1 U7676 ( .B1(n6733), .B2(keyinput37), .C1(n6732), .C2(
        UWORD_REG_10__SCAN_IN), .A(n6731), .ZN(n6738) );
  INV_X1 U7677 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6736) );
  INV_X1 U7678 ( .A(keyinput16), .ZN(n6735) );
  AOI22_X1 U7679 ( .A1(n6736), .A2(keyinput25), .B1(DATAI_7_), .B2(n6735), 
        .ZN(n6734) );
  OAI221_X1 U7680 ( .B1(n6736), .B2(keyinput25), .C1(n6735), .C2(DATAI_7_), 
        .A(n6734), .ZN(n6737) );
  NOR4_X1 U7681 ( .A1(n6740), .A2(n6739), .A3(n6738), .A4(n6737), .ZN(n6741)
         );
  NAND4_X1 U7682 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n6944)
         );
  AOI22_X1 U7683 ( .A1(n3350), .A2(keyinput31), .B1(keyinput116), .B2(n6746), 
        .ZN(n6745) );
  OAI221_X1 U7684 ( .B1(n3350), .B2(keyinput31), .C1(n6746), .C2(keyinput116), 
        .A(n6745), .ZN(n6759) );
  INV_X1 U7685 ( .A(keyinput45), .ZN(n6749) );
  AOI22_X1 U7686 ( .A1(n6749), .A2(DATAO_REG_6__SCAN_IN), .B1(keyinput112), 
        .B2(n6748), .ZN(n6747) );
  OAI221_X1 U7687 ( .B1(n6749), .B2(DATAO_REG_6__SCAN_IN), .C1(n6748), .C2(
        keyinput112), .A(n6747), .ZN(n6758) );
  INV_X1 U7688 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6752) );
  INV_X1 U7689 ( .A(keyinput124), .ZN(n6751) );
  AOI22_X1 U7690 ( .A1(n6752), .A2(keyinput76), .B1(LWORD_REG_8__SCAN_IN), 
        .B2(n6751), .ZN(n6750) );
  OAI221_X1 U7691 ( .B1(n6752), .B2(keyinput76), .C1(n6751), .C2(
        LWORD_REG_8__SCAN_IN), .A(n6750), .ZN(n6757) );
  INV_X1 U7692 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6755) );
  INV_X1 U7693 ( .A(keyinput44), .ZN(n6754) );
  AOI22_X1 U7694 ( .A1(n6755), .A2(keyinput120), .B1(DATAWIDTH_REG_20__SCAN_IN), .B2(n6754), .ZN(n6753) );
  OAI221_X1 U7695 ( .B1(n6755), .B2(keyinput120), .C1(n6754), .C2(
        DATAWIDTH_REG_20__SCAN_IN), .A(n6753), .ZN(n6756) );
  NOR4_X1 U7696 ( .A1(n6759), .A2(n6758), .A3(n6757), .A4(n6756), .ZN(n6809)
         );
  INV_X1 U7697 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6762) );
  INV_X1 U7698 ( .A(keyinput58), .ZN(n6761) );
  AOI22_X1 U7699 ( .A1(n6762), .A2(keyinput103), .B1(ADDRESS_REG_23__SCAN_IN), 
        .B2(n6761), .ZN(n6760) );
  OAI221_X1 U7700 ( .B1(n6762), .B2(keyinput103), .C1(n6761), .C2(
        ADDRESS_REG_23__SCAN_IN), .A(n6760), .ZN(n6774) );
  INV_X1 U7701 ( .A(keyinput71), .ZN(n6764) );
  AOI22_X1 U7702 ( .A1(n6765), .A2(keyinput79), .B1(DATAO_REG_17__SCAN_IN), 
        .B2(n6764), .ZN(n6763) );
  OAI221_X1 U7703 ( .B1(n6765), .B2(keyinput79), .C1(n6764), .C2(
        DATAO_REG_17__SCAN_IN), .A(n6763), .ZN(n6773) );
  INV_X1 U7704 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6768) );
  INV_X1 U7705 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6767) );
  AOI22_X1 U7706 ( .A1(n6768), .A2(keyinput18), .B1(keyinput65), .B2(n6767), 
        .ZN(n6766) );
  OAI221_X1 U7707 ( .B1(n6768), .B2(keyinput18), .C1(n6767), .C2(keyinput65), 
        .A(n6766), .ZN(n6772) );
  INV_X1 U7708 ( .A(keyinput98), .ZN(n6770) );
  AOI22_X1 U7709 ( .A1(n6594), .A2(keyinput86), .B1(DATAO_REG_18__SCAN_IN), 
        .B2(n6770), .ZN(n6769) );
  OAI221_X1 U7710 ( .B1(n6594), .B2(keyinput86), .C1(n6770), .C2(
        DATAO_REG_18__SCAN_IN), .A(n6769), .ZN(n6771) );
  NOR4_X1 U7711 ( .A1(n6774), .A2(n6773), .A3(n6772), .A4(n6771), .ZN(n6808)
         );
  INV_X1 U7712 ( .A(keyinput68), .ZN(n6777) );
  INV_X1 U7713 ( .A(keyinput95), .ZN(n6776) );
  AOI22_X1 U7714 ( .A1(n6777), .A2(READREQUEST_REG_SCAN_IN), .B1(
        DATAWIDTH_REG_27__SCAN_IN), .B2(n6776), .ZN(n6775) );
  OAI221_X1 U7715 ( .B1(n6777), .B2(READREQUEST_REG_SCAN_IN), .C1(n6776), .C2(
        DATAWIDTH_REG_27__SCAN_IN), .A(n6775), .ZN(n6789) );
  AOI22_X1 U7716 ( .A1(n6042), .A2(keyinput78), .B1(keyinput80), .B2(n6779), 
        .ZN(n6778) );
  OAI221_X1 U7717 ( .B1(n6042), .B2(keyinput78), .C1(n6779), .C2(keyinput80), 
        .A(n6778), .ZN(n6788) );
  INV_X1 U7718 ( .A(keyinput46), .ZN(n6781) );
  AOI22_X1 U7719 ( .A1(n6782), .A2(keyinput105), .B1(ADDRESS_REG_0__SCAN_IN), 
        .B2(n6781), .ZN(n6780) );
  OAI221_X1 U7720 ( .B1(n6782), .B2(keyinput105), .C1(n6781), .C2(
        ADDRESS_REG_0__SCAN_IN), .A(n6780), .ZN(n6787) );
  INV_X1 U7721 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6784) );
  AOI22_X1 U7722 ( .A1(n6785), .A2(keyinput53), .B1(n6784), .B2(keyinput8), 
        .ZN(n6783) );
  OAI221_X1 U7723 ( .B1(n6785), .B2(keyinput53), .C1(n6784), .C2(keyinput8), 
        .A(n6783), .ZN(n6786) );
  NOR4_X1 U7724 ( .A1(n6789), .A2(n6788), .A3(n6787), .A4(n6786), .ZN(n6807)
         );
  INV_X1 U7725 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6792) );
  INV_X1 U7726 ( .A(keyinput29), .ZN(n6791) );
  AOI22_X1 U7727 ( .A1(n6792), .A2(keyinput15), .B1(DATAO_REG_12__SCAN_IN), 
        .B2(n6791), .ZN(n6790) );
  OAI221_X1 U7728 ( .B1(n6792), .B2(keyinput15), .C1(n6791), .C2(
        DATAO_REG_12__SCAN_IN), .A(n6790), .ZN(n6805) );
  INV_X1 U7729 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n6794) );
  AOI22_X1 U7730 ( .A1(n6795), .A2(keyinput67), .B1(n6794), .B2(keyinput42), 
        .ZN(n6793) );
  OAI221_X1 U7731 ( .B1(n6795), .B2(keyinput67), .C1(n6794), .C2(keyinput42), 
        .A(n6793), .ZN(n6804) );
  INV_X1 U7732 ( .A(keyinput101), .ZN(n6798) );
  INV_X1 U7733 ( .A(keyinput104), .ZN(n6797) );
  AOI22_X1 U7734 ( .A1(n6798), .A2(FLUSH_REG_SCAN_IN), .B1(
        BYTEENABLE_REG_1__SCAN_IN), .B2(n6797), .ZN(n6796) );
  OAI221_X1 U7735 ( .B1(n6798), .B2(FLUSH_REG_SCAN_IN), .C1(n6797), .C2(
        BYTEENABLE_REG_1__SCAN_IN), .A(n6796), .ZN(n6803) );
  INV_X1 U7736 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6801) );
  AOI22_X1 U7737 ( .A1(n6801), .A2(keyinput87), .B1(n6800), .B2(keyinput24), 
        .ZN(n6799) );
  OAI221_X1 U7738 ( .B1(n6801), .B2(keyinput87), .C1(n6800), .C2(keyinput24), 
        .A(n6799), .ZN(n6802) );
  NOR4_X1 U7739 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n6806)
         );
  NAND4_X1 U7740 ( .A1(n6809), .A2(n6808), .A3(n6807), .A4(n6806), .ZN(n6943)
         );
  INV_X1 U7741 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n6812) );
  OAI22_X1 U7742 ( .A1(n6812), .A2(keyinput93), .B1(n6811), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6810) );
  AOI221_X1 U7743 ( .B1(n6812), .B2(keyinput93), .C1(UWORD_REG_11__SCAN_IN), 
        .C2(n6811), .A(n6810), .ZN(n6941) );
  INV_X1 U7744 ( .A(keyinput19), .ZN(n6814) );
  OAI22_X1 U7745 ( .A1(keyinput48), .A2(n6815), .B1(n6814), .B2(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n6813) );
  AOI221_X1 U7746 ( .B1(n6815), .B2(keyinput48), .C1(n6814), .C2(
        DATAWIDTH_REG_28__SCAN_IN), .A(n6813), .ZN(n6940) );
  AOI22_X1 U7747 ( .A1(n6817), .A2(keyinput40), .B1(n5271), .B2(keyinput99), 
        .ZN(n6816) );
  OAI221_X1 U7748 ( .B1(n6817), .B2(keyinput40), .C1(n5271), .C2(keyinput99), 
        .A(n6816), .ZN(n6839) );
  INV_X1 U7749 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6820) );
  AOI22_X1 U7750 ( .A1(n6820), .A2(keyinput64), .B1(keyinput102), .B2(n6819), 
        .ZN(n6818) );
  OAI221_X1 U7751 ( .B1(n6820), .B2(keyinput64), .C1(n6819), .C2(keyinput102), 
        .A(n6818), .ZN(n6838) );
  INV_X1 U7752 ( .A(keyinput119), .ZN(n6822) );
  OAI22_X1 U7753 ( .A1(keyinput56), .A2(n6823), .B1(n6822), .B2(
        BE_N_REG_2__SCAN_IN), .ZN(n6821) );
  AOI221_X1 U7754 ( .B1(n6823), .B2(keyinput56), .C1(n6822), .C2(
        BE_N_REG_2__SCAN_IN), .A(n6821), .ZN(n6836) );
  INV_X1 U7755 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6826) );
  INV_X1 U7756 ( .A(keyinput39), .ZN(n6825) );
  OAI22_X1 U7757 ( .A1(n6826), .A2(keyinput27), .B1(n6825), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6824) );
  AOI221_X1 U7758 ( .B1(n6826), .B2(keyinput27), .C1(LWORD_REG_9__SCAN_IN), 
        .C2(n6825), .A(n6824), .ZN(n6835) );
  INV_X1 U7759 ( .A(keyinput81), .ZN(n6828) );
  OAI22_X1 U7760 ( .A1(keyinput107), .A2(n6829), .B1(n6828), .B2(
        MEMORYFETCH_REG_SCAN_IN), .ZN(n6827) );
  AOI221_X1 U7761 ( .B1(n6829), .B2(keyinput107), .C1(n6828), .C2(
        MEMORYFETCH_REG_SCAN_IN), .A(n6827), .ZN(n6834) );
  INV_X1 U7762 ( .A(keyinput115), .ZN(n6832) );
  INV_X1 U7763 ( .A(keyinput28), .ZN(n6831) );
  OAI22_X1 U7764 ( .A1(n6832), .A2(BE_N_REG_0__SCAN_IN), .B1(n6831), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n6830) );
  AOI221_X1 U7765 ( .B1(n6832), .B2(BE_N_REG_0__SCAN_IN), .C1(
        DATAO_REG_28__SCAN_IN), .C2(n6831), .A(n6830), .ZN(n6833) );
  NAND4_X1 U7766 ( .A1(n6836), .A2(n6835), .A3(n6834), .A4(n6833), .ZN(n6837)
         );
  NOR3_X1 U7767 ( .A1(n6839), .A2(n6838), .A3(n6837), .ZN(n6939) );
  INV_X1 U7768 ( .A(keyinput106), .ZN(n6845) );
  INV_X1 U7769 ( .A(keyinput52), .ZN(n6844) );
  AOI22_X1 U7770 ( .A1(n6845), .A2(DATAO_REG_0__SCAN_IN), .B1(
        DATAWIDTH_REG_13__SCAN_IN), .B2(n6844), .ZN(n6843) );
  OAI221_X1 U7771 ( .B1(n6845), .B2(DATAO_REG_0__SCAN_IN), .C1(n6844), .C2(
        DATAWIDTH_REG_13__SCAN_IN), .A(n6843), .ZN(n6936) );
  INV_X1 U7772 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6848) );
  INV_X1 U7773 ( .A(keyinput55), .ZN(n6847) );
  OAI22_X1 U7774 ( .A1(keyinput123), .A2(n6848), .B1(n6847), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n6846) );
  AOI221_X1 U7775 ( .B1(n6848), .B2(keyinput123), .C1(n6847), .C2(
        LWORD_REG_6__SCAN_IN), .A(n6846), .ZN(n6869) );
  INV_X1 U7776 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6851) );
  INV_X1 U7777 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6850) );
  OAI22_X1 U7778 ( .A1(n6851), .A2(keyinput121), .B1(n6850), .B2(keyinput61), 
        .ZN(n6849) );
  AOI221_X1 U7779 ( .B1(n6851), .B2(keyinput121), .C1(keyinput61), .C2(n6850), 
        .A(n6849), .ZN(n6868) );
  INV_X1 U7780 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n6854) );
  INV_X1 U7781 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6853) );
  AOI22_X1 U7782 ( .A1(n6854), .A2(keyinput26), .B1(n6853), .B2(keyinput111), 
        .ZN(n6852) );
  OAI221_X1 U7783 ( .B1(n6854), .B2(keyinput26), .C1(n6853), .C2(keyinput111), 
        .A(n6852), .ZN(n6866) );
  INV_X1 U7784 ( .A(keyinput23), .ZN(n6856) );
  AOI22_X1 U7785 ( .A1(n6857), .A2(keyinput122), .B1(DATAO_REG_9__SCAN_IN), 
        .B2(n6856), .ZN(n6855) );
  OAI221_X1 U7786 ( .B1(n6857), .B2(keyinput122), .C1(n6856), .C2(
        DATAO_REG_9__SCAN_IN), .A(n6855), .ZN(n6865) );
  AOI22_X1 U7787 ( .A1(n4310), .A2(keyinput83), .B1(n6859), .B2(keyinput127), 
        .ZN(n6858) );
  OAI221_X1 U7788 ( .B1(n4310), .B2(keyinput83), .C1(n6859), .C2(keyinput127), 
        .A(n6858), .ZN(n6864) );
  INV_X1 U7789 ( .A(keyinput85), .ZN(n6861) );
  AOI22_X1 U7790 ( .A1(n6862), .A2(keyinput10), .B1(UWORD_REG_7__SCAN_IN), 
        .B2(n6861), .ZN(n6860) );
  OAI221_X1 U7791 ( .B1(n6862), .B2(keyinput10), .C1(n6861), .C2(
        UWORD_REG_7__SCAN_IN), .A(n6860), .ZN(n6863) );
  NOR4_X1 U7792 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6867)
         );
  NAND3_X1 U7793 ( .A1(n6869), .A2(n6868), .A3(n6867), .ZN(n6935) );
  INV_X1 U7794 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6872) );
  INV_X1 U7795 ( .A(keyinput38), .ZN(n6871) );
  AOI22_X1 U7796 ( .A1(n6872), .A2(keyinput7), .B1(LWORD_REG_10__SCAN_IN), 
        .B2(n6871), .ZN(n6870) );
  OAI221_X1 U7797 ( .B1(n6872), .B2(keyinput7), .C1(n6871), .C2(
        LWORD_REG_10__SCAN_IN), .A(n6870), .ZN(n6885) );
  INV_X1 U7798 ( .A(keyinput66), .ZN(n6874) );
  AOI22_X1 U7799 ( .A1(n6875), .A2(keyinput88), .B1(UWORD_REG_0__SCAN_IN), 
        .B2(n6874), .ZN(n6873) );
  OAI221_X1 U7800 ( .B1(n6875), .B2(keyinput88), .C1(n6874), .C2(
        UWORD_REG_0__SCAN_IN), .A(n6873), .ZN(n6884) );
  INV_X1 U7801 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6878) );
  AOI22_X1 U7802 ( .A1(n6878), .A2(keyinput2), .B1(n6877), .B2(keyinput50), 
        .ZN(n6876) );
  OAI221_X1 U7803 ( .B1(n6878), .B2(keyinput2), .C1(n6877), .C2(keyinput50), 
        .A(n6876), .ZN(n6883) );
  INV_X1 U7804 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6881) );
  AOI22_X1 U7805 ( .A1(n6881), .A2(keyinput77), .B1(DATAI_9_), .B2(n6880), 
        .ZN(n6879) );
  OAI221_X1 U7806 ( .B1(n6881), .B2(keyinput77), .C1(n6880), .C2(DATAI_9_), 
        .A(n6879), .ZN(n6882) );
  NOR4_X1 U7807 ( .A1(n6885), .A2(n6884), .A3(n6883), .A4(n6882), .ZN(n6933)
         );
  INV_X1 U7808 ( .A(keyinput33), .ZN(n6887) );
  AOI22_X1 U7809 ( .A1(n5401), .A2(keyinput91), .B1(M_IO_N_REG_SCAN_IN), .B2(
        n6887), .ZN(n6886) );
  OAI221_X1 U7810 ( .B1(n5401), .B2(keyinput91), .C1(n6887), .C2(
        M_IO_N_REG_SCAN_IN), .A(n6886), .ZN(n6899) );
  INV_X1 U7811 ( .A(keyinput97), .ZN(n6889) );
  AOI22_X1 U7812 ( .A1(n6890), .A2(keyinput114), .B1(ADDRESS_REG_4__SCAN_IN), 
        .B2(n6889), .ZN(n6888) );
  OAI221_X1 U7813 ( .B1(n6890), .B2(keyinput114), .C1(n6889), .C2(
        ADDRESS_REG_4__SCAN_IN), .A(n6888), .ZN(n6898) );
  INV_X1 U7814 ( .A(keyinput51), .ZN(n6892) );
  AOI22_X1 U7815 ( .A1(n5164), .A2(keyinput96), .B1(LWORD_REG_15__SCAN_IN), 
        .B2(n6892), .ZN(n6891) );
  OAI221_X1 U7816 ( .B1(n5164), .B2(keyinput96), .C1(n6892), .C2(
        LWORD_REG_15__SCAN_IN), .A(n6891), .ZN(n6897) );
  AOI22_X1 U7817 ( .A1(n6895), .A2(keyinput90), .B1(DATAO_REG_2__SCAN_IN), 
        .B2(n6894), .ZN(n6893) );
  OAI221_X1 U7818 ( .B1(n6895), .B2(keyinput90), .C1(n6894), .C2(
        DATAO_REG_2__SCAN_IN), .A(n6893), .ZN(n6896) );
  NOR4_X1 U7819 ( .A1(n6899), .A2(n6898), .A3(n6897), .A4(n6896), .ZN(n6932)
         );
  AOI22_X1 U7820 ( .A1(n3840), .A2(keyinput0), .B1(keyinput11), .B2(n6901), 
        .ZN(n6900) );
  OAI221_X1 U7821 ( .B1(n3840), .B2(keyinput0), .C1(n6901), .C2(keyinput11), 
        .A(n6900), .ZN(n6914) );
  INV_X1 U7822 ( .A(keyinput125), .ZN(n6903) );
  INV_X1 U7823 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6907) );
  INV_X1 U7824 ( .A(keyinput9), .ZN(n6906) );
  AOI22_X1 U7825 ( .A1(n6907), .A2(keyinput117), .B1(ADDRESS_REG_26__SCAN_IN), 
        .B2(n6906), .ZN(n6905) );
  OAI221_X1 U7826 ( .B1(n6907), .B2(keyinput117), .C1(n6906), .C2(
        ADDRESS_REG_26__SCAN_IN), .A(n6905), .ZN(n6912) );
  INV_X1 U7827 ( .A(keyinput54), .ZN(n6909) );
  AOI22_X1 U7828 ( .A1(n6910), .A2(keyinput34), .B1(ADDRESS_REG_21__SCAN_IN), 
        .B2(n6909), .ZN(n6908) );
  OAI221_X1 U7829 ( .B1(n6910), .B2(keyinput34), .C1(n6909), .C2(
        ADDRESS_REG_21__SCAN_IN), .A(n6908), .ZN(n6911) );
  NOR4_X1 U7830 ( .A1(n6914), .A2(n6913), .A3(n6912), .A4(n6911), .ZN(n6931)
         );
  INV_X1 U7831 ( .A(keyinput109), .ZN(n6917) );
  INV_X1 U7832 ( .A(keyinput74), .ZN(n6916) );
  AOI22_X1 U7833 ( .A1(n6917), .A2(DATAWIDTH_REG_4__SCAN_IN), .B1(
        UWORD_REG_13__SCAN_IN), .B2(n6916), .ZN(n6915) );
  OAI221_X1 U7834 ( .B1(n6917), .B2(DATAWIDTH_REG_4__SCAN_IN), .C1(n6916), 
        .C2(UWORD_REG_13__SCAN_IN), .A(n6915), .ZN(n6929) );
  AOI22_X1 U7835 ( .A1(n6920), .A2(keyinput17), .B1(n6919), .B2(keyinput14), 
        .ZN(n6918) );
  OAI221_X1 U7836 ( .B1(n6920), .B2(keyinput17), .C1(n6919), .C2(keyinput14), 
        .A(n6918), .ZN(n6928) );
  INV_X1 U7837 ( .A(keyinput75), .ZN(n6922) );
  AOI22_X1 U7838 ( .A1(n6923), .A2(keyinput35), .B1(ADDRESS_REG_7__SCAN_IN), 
        .B2(n6922), .ZN(n6921) );
  OAI221_X1 U7839 ( .B1(n6923), .B2(keyinput35), .C1(n6922), .C2(
        ADDRESS_REG_7__SCAN_IN), .A(n6921), .ZN(n6927) );
  XNOR2_X1 U7840 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput32), .ZN(
        n6925) );
  XNOR2_X1 U7841 ( .A(keyinput126), .B(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U7842 ( .A1(n6925), .A2(n6924), .ZN(n6926) );
  NOR4_X1 U7843 ( .A1(n6929), .A2(n6928), .A3(n6927), .A4(n6926), .ZN(n6930)
         );
  NAND4_X1 U7844 ( .A1(n6933), .A2(n6932), .A3(n6931), .A4(n6930), .ZN(n6934)
         );
  NOR4_X1 U7845 ( .A1(n6937), .A2(n6936), .A3(n6935), .A4(n6934), .ZN(n6938)
         );
  NAND4_X1 U7846 ( .A1(n6941), .A2(n6940), .A3(n6939), .A4(n6938), .ZN(n6942)
         );
  NOR4_X1 U7847 ( .A1(n6945), .A2(n6944), .A3(n6943), .A4(n6942), .ZN(n6954)
         );
  AOI22_X1 U7848 ( .A1(n6947), .A2(EAX_REG_25__SCAN_IN), .B1(n6946), .B2(
        DATAI_9_), .ZN(n6950) );
  NAND2_X1 U7849 ( .A1(n6948), .A2(DATAI_25_), .ZN(n6949) );
  OAI211_X1 U7850 ( .C1(n6951), .C2(n5855), .A(n6950), .B(n6949), .ZN(n6952)
         );
  INV_X1 U7851 ( .A(n6952), .ZN(n6953) );
  XNOR2_X1 U7852 ( .A(n6954), .B(n6953), .ZN(U2866) );
  AND4_X1 U4196 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n3252)
         );
  INV_X1 U4235 ( .A(n4676), .ZN(n3976) );
  CLKBUF_X2 U4286 ( .A(n3258), .Z(n4202) );
  BUF_X1 U3634 ( .A(n3412), .Z(n3352) );
  AND2_X1 U3756 ( .A1(n3936), .A2(n3935), .ZN(n4489) );
  CLKBUF_X2 U3587 ( .A(n3746), .Z(n3864) );
  AND3_X1 U3619 ( .A1(n3310), .A2(n3289), .A3(n4648), .ZN(n3290) );
  AND2_X1 U3707 ( .A1(n3300), .A2(n4672), .ZN(n3984) );
  CLKBUF_X1 U3903 ( .A(n3986), .Z(n5458) );
  CLKBUF_X2 U4005 ( .A(n3987), .Z(n4023) );
  AND2_X2 U4205 ( .A1(n3892), .A2(n4672), .ZN(n4534) );
  CLKBUF_X1 U4966 ( .A(n6159), .Z(n6614) );
endmodule

