

module b20_C_AntiSAT_k_128_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208;

  NAND2_X1 U4838 ( .A1(n9567), .A2(n7531), .ZN(n9568) );
  OR2_X1 U4839 ( .A1(n9645), .A2(n8820), .ZN(n9071) );
  NAND2_X1 U4840 ( .A1(n9645), .A2(n8820), .ZN(n9076) );
  NAND2_X2 U4841 ( .A1(n7516), .A2(n7515), .ZN(n9645) );
  INV_X2 U4842 ( .A(n5725), .ZN(n5748) );
  INV_X1 U4843 ( .A(n4339), .ZN(n5529) );
  CLKBUF_X2 U4844 ( .A(n5020), .Z(n5532) );
  INV_X1 U4845 ( .A(n8640), .ZN(n8541) );
  BUF_X1 U4846 ( .A(n6383), .Z(n6440) );
  CLKBUF_X2 U4847 ( .A(n6113), .Z(n4333) );
  INV_X1 U4848 ( .A(n8864), .ZN(n7575) );
  NOR2_X1 U4849 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4552) );
  NAND2_X1 U4850 ( .A1(n4978), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4977) );
  NAND2_X1 U4851 ( .A1(n8176), .A2(n7245), .ZN(n8163) );
  NAND3_X1 U4852 ( .A1(n4932), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4934) );
  OR2_X2 U4853 ( .A1(n5981), .A2(n6197), .ZN(n8565) );
  AND2_X1 U4854 ( .A1(n9460), .A2(n8912), .ZN(n9448) );
  INV_X1 U4855 ( .A(n6263), .ZN(n7574) );
  OAI21_X1 U4856 ( .B1(n7700), .B2(n7702), .A(n7701), .ZN(n7699) );
  INV_X2 U4857 ( .A(n5327), .ZN(n5312) );
  INV_X1 U4858 ( .A(n5528), .ZN(n7401) );
  NAND2_X1 U4859 ( .A1(n4840), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5840) );
  OAI211_X1 U4860 ( .C1(n5082), .C2(n4988), .A(n4991), .B(n4671), .ZN(n6380)
         );
  AOI21_X1 U4861 ( .B1(n4689), .B2(n4347), .A(n4690), .ZN(n7835) );
  OR2_X1 U4862 ( .A1(n7422), .A2(n4608), .ZN(n4607) );
  NOR2_X1 U4863 ( .A1(n8004), .A2(n8003), .ZN(n8006) );
  NAND2_X1 U4865 ( .A1(n9071), .A2(n9076), .ZN(n9474) );
  MUX2_X1 U4866 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9686), .S(n9816), .Z(n9592)
         );
  NAND2_X1 U4867 ( .A1(n7600), .A2(n7599), .ZN(n9404) );
  XNOR2_X1 U4868 ( .A(n5840), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9109) );
  CLKBUF_X2 U4869 ( .A(n5030), .Z(n5787) );
  AOI211_X1 U4870 ( .C1(n8027), .C2(n9901), .A(n8026), .B(n8025), .ZN(n8028)
         );
  BUF_X1 U4871 ( .A(n6384), .Z(n9142) );
  XNOR2_X1 U4872 ( .A(n5864), .B(n5863), .ZN(n5865) );
  NOR2_X2 U4873 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4676) );
  NOR2_X2 U4874 ( .A1(n7940), .A2(n4426), .ZN(n7956) );
  OR2_X2 U4875 ( .A1(n6882), .A2(n6877), .ZN(n4760) );
  NOR2_X2 U4876 ( .A1(n7938), .A2(n4427), .ZN(n7971) );
  NAND2_X2 U4877 ( .A1(n5170), .A2(n5169), .ZN(n5192) );
  AOI21_X2 U4878 ( .B1(n5164), .B2(n5163), .A(n5162), .ZN(n5170) );
  INV_X2 U4879 ( .A(n5980), .ZN(n6196) );
  OR2_X1 U4880 ( .A1(n5981), .A2(n6197), .ZN(n4332) );
  AOI21_X2 U4881 ( .B1(n4820), .B2(n4816), .A(n4813), .ZN(n9365) );
  NOR2_X2 U4882 ( .A1(n9870), .A2(n5068), .ZN(n9869) );
  NAND2_X2 U4883 ( .A1(n6350), .A2(n4483), .ZN(n9870) );
  NAND2_X2 U4884 ( .A1(n5614), .A2(n5613), .ZN(n5662) );
  OAI21_X2 U4885 ( .B1(n5322), .B2(n4785), .A(n4782), .ZN(n8176) );
  OAI21_X2 U4886 ( .B1(n5280), .B2(SI_15_), .A(n5281), .ZN(n5301) );
  BUF_X4 U4887 ( .A(n4940), .Z(n4443) );
  INV_X1 U4888 ( .A(n7885), .ZN(n6924) );
  NAND4_X2 U4889 ( .A1(n5128), .A2(n5127), .A3(n5126), .A4(n5125), .ZN(n7885)
         );
  OAI21_X2 U4890 ( .B1(n7835), .B2(n7717), .A(n7716), .ZN(n7784) );
  XNOR2_X2 U4891 ( .A(n4444), .B(n6384), .ZN(n6434) );
  NAND4_X2 U4892 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n6384)
         );
  OAI21_X2 U4893 ( .B1(n9315), .B2(n9321), .A(n9092), .ZN(n9303) );
  NAND2_X2 U4894 ( .A1(n9332), .A2(n8989), .ZN(n9315) );
  OAI21_X2 U4895 ( .B1(n6294), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6360) );
  OAI21_X2 U4896 ( .B1(n8256), .B2(n7451), .A(n7449), .ZN(n8246) );
  OAI21_X2 U4897 ( .B1(n7130), .B2(n4659), .A(n4655), .ZN(n8256) );
  CLKBUF_X3 U4898 ( .A(n7591), .Z(n8867) );
  NAND2_X2 U4899 ( .A1(n7584), .A2(n4413), .ZN(n4820) );
  XNOR2_X2 U4900 ( .A(n5843), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9025) );
  NAND2_X2 U4901 ( .A1(n5842), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5843) );
  NOR2_X2 U4902 ( .A1(n7986), .A2(n7985), .ZN(n8009) );
  NAND2_X2 U4903 ( .A1(n7550), .A2(n7549), .ZN(n9657) );
  XNOR2_X2 U4904 ( .A(n4977), .B(n4976), .ZN(n6307) );
  OAI21_X2 U4905 ( .B1(n5375), .B2(n5374), .A(n5373), .ZN(n5377) );
  OAI21_X2 U4906 ( .B1(n5363), .B2(n5362), .A(n5361), .ZN(n5375) );
  OAI22_X2 U4907 ( .A1(n8195), .A2(n5568), .B1(n8212), .B2(n8201), .ZN(n8182)
         );
  NAND2_X1 U4908 ( .A1(n7639), .A2(n7638), .ZN(n9331) );
  OAI21_X1 U4909 ( .B1(n8820), .B2(n9479), .A(n9473), .ZN(n9457) );
  NAND2_X1 U4910 ( .A1(n8597), .A2(n8598), .ZN(n8596) );
  AND2_X1 U4911 ( .A1(n4450), .A2(n4469), .ZN(n8597) );
  OR2_X1 U4912 ( .A1(n8481), .A2(n8480), .ZN(n4450) );
  NAND2_X1 U4913 ( .A1(n9525), .A2(n7673), .ZN(n7674) );
  NAND2_X1 U4914 ( .A1(n5557), .A2(n5556), .ZN(n7130) );
  AND2_X1 U4915 ( .A1(n9068), .A2(n8960), .ZN(n9505) );
  NOR3_X1 U4916 ( .A1(n6881), .A2(n6880), .A3(n6879), .ZN(n4943) );
  INV_X2 U4917 ( .A(n8935), .ZN(n6985) );
  OAI21_X1 U4918 ( .B1(n6677), .B2(n5550), .A(n5549), .ZN(n6763) );
  NAND2_X1 U4919 ( .A1(n8918), .A2(n8922), .ZN(n8840) );
  NAND2_X1 U4920 ( .A1(n7284), .A2(n7276), .ZN(n7429) );
  CLKBUF_X2 U4921 ( .A(n6107), .Z(n8641) );
  INV_X4 U4922 ( .A(n8565), .ZN(n8644) );
  NAND2_X1 U4923 ( .A1(n9025), .A2(n9038), .ZN(n5980) );
  NAND2_X2 U4924 ( .A1(n8429), .A2(n8432), .ZN(n5063) );
  INV_X1 U4925 ( .A(n5002), .ZN(n5030) );
  NAND2_X1 U4926 ( .A1(n8429), .A2(n4975), .ZN(n5020) );
  CLKBUF_X3 U4927 ( .A(n5005), .Z(n4339) );
  NAND2_X1 U4928 ( .A1(n6307), .A2(n8041), .ZN(n5002) );
  NAND2_X1 U4929 ( .A1(n4974), .A2(n4975), .ZN(n5338) );
  INV_X1 U4930 ( .A(n6345), .ZN(n4335) );
  OR2_X1 U4931 ( .A1(n4609), .A2(n8046), .ZN(n4473) );
  OR2_X1 U4932 ( .A1(n8540), .A2(n8769), .ZN(n4842) );
  NAND2_X1 U4933 ( .A1(n8539), .A2(n8538), .ZN(n8606) );
  OR2_X1 U4934 ( .A1(n8371), .A2(n9966), .ZN(n4627) );
  NAND2_X1 U4935 ( .A1(n4836), .A2(n4832), .ZN(n4834) );
  NAND2_X1 U4936 ( .A1(n5522), .A2(n5521), .ZN(n7413) );
  AND2_X1 U4937 ( .A1(n7381), .A2(n7380), .ZN(n8370) );
  NAND2_X1 U4938 ( .A1(n4793), .A2(n4390), .ZN(n9430) );
  NAND2_X1 U4939 ( .A1(n7802), .A2(n7806), .ZN(n5729) );
  NAND2_X1 U4940 ( .A1(n7725), .A2(n4678), .ZN(n7802) );
  CLKBUF_X1 U4941 ( .A(n4856), .Z(n4470) );
  NAND2_X1 U4942 ( .A1(n7483), .A2(n7482), .ZN(n9593) );
  NOR2_X1 U4943 ( .A1(n9355), .A2(n9339), .ZN(n4459) );
  NAND2_X1 U4944 ( .A1(n8485), .A2(n8484), .ZN(n8486) );
  AND2_X1 U4945 ( .A1(n4492), .A2(n4491), .ZN(n8002) );
  AND2_X1 U4946 ( .A1(n7358), .A2(n7362), .ZN(n8107) );
  NAND2_X1 U4947 ( .A1(n5453), .A2(n5452), .ZN(n7743) );
  OAI21_X1 U4948 ( .B1(n5704), .B2(n7878), .A(n7699), .ZN(n7862) );
  OR2_X1 U4949 ( .A1(n7941), .A2(n8242), .ZN(n4452) );
  XNOR2_X1 U4950 ( .A(n5466), .B(n5465), .ZN(n7640) );
  NAND2_X1 U4951 ( .A1(n7621), .A2(n7620), .ZN(n9372) );
  NAND2_X1 U4952 ( .A1(n7609), .A2(n7608), .ZN(n9387) );
  AND2_X1 U4953 ( .A1(n4496), .A2(n4495), .ZN(n7940) );
  NAND2_X1 U4954 ( .A1(n4702), .A2(n4701), .ZN(n7793) );
  NOR2_X1 U4955 ( .A1(n9464), .A2(n9634), .ZN(n4874) );
  AND2_X1 U4956 ( .A1(n6995), .A2(n5691), .ZN(n7026) );
  NAND2_X1 U4957 ( .A1(n6875), .A2(n6886), .ZN(n7526) );
  AOI21_X1 U4958 ( .B1(n4845), .B2(n4850), .A(n4369), .ZN(n4844) );
  AND2_X1 U4959 ( .A1(n4849), .A2(n4846), .ZN(n4845) );
  NAND2_X1 U4960 ( .A1(n6883), .A2(n8848), .ZN(n9557) );
  OR2_X1 U4961 ( .A1(n4852), .A2(n4851), .ZN(n4849) );
  OAI21_X1 U4962 ( .B1(n6878), .B2(n4760), .A(n9056), .ZN(n6885) );
  NOR2_X1 U4963 ( .A1(n7207), .A2(n7147), .ZN(n7206) );
  OR2_X1 U4964 ( .A1(n7083), .A2(n5555), .ZN(n5557) );
  OR2_X1 U4965 ( .A1(n8468), .A2(n8467), .ZN(n8682) );
  AND2_X1 U4966 ( .A1(n6702), .A2(n5684), .ZN(n6728) );
  NAND2_X1 U4967 ( .A1(n7562), .A2(n7561), .ZN(n9649) );
  OR2_X1 U4968 ( .A1(n9657), .A2(n8818), .ZN(n9068) );
  XNOR2_X1 U4969 ( .A(n7163), .B(n7171), .ZN(n7207) );
  NAND2_X1 U4970 ( .A1(n7536), .A2(n7535), .ZN(n9729) );
  NAND2_X1 U4971 ( .A1(n4675), .A2(n5551), .ZN(n6809) );
  NOR2_X1 U4972 ( .A1(n7003), .A2(n7002), .ZN(n7162) );
  NAND2_X1 U4973 ( .A1(n7530), .A2(n7529), .ZN(n9733) );
  NAND2_X1 U4974 ( .A1(n6874), .A2(n6873), .ZN(n8624) );
  NAND2_X1 U4975 ( .A1(n4504), .A2(n4503), .ZN(n4502) );
  NAND2_X1 U4976 ( .A1(n9877), .A2(n4382), .ZN(n4501) );
  NAND2_X1 U4977 ( .A1(n6737), .A2(n8861), .ZN(n4438) );
  NAND2_X1 U4978 ( .A1(n6836), .A2(n6835), .ZN(n8450) );
  NAND2_X1 U4979 ( .A1(n5120), .A2(n5119), .ZN(n6960) );
  AND2_X1 U4980 ( .A1(n6638), .A2(n9898), .ZN(n9877) );
  XNOR2_X1 U4981 ( .A(n5146), .B(n5145), .ZN(n6737) );
  NAND2_X1 U4982 ( .A1(n5100), .A2(n5099), .ZN(n5110) );
  NAND2_X1 U4983 ( .A1(n4727), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4514) );
  OR2_X1 U4984 ( .A1(n7889), .A2(n6952), .ZN(n7284) );
  NAND2_X1 U4985 ( .A1(n7264), .A2(n7268), .ZN(n7431) );
  INV_X1 U4986 ( .A(n6256), .ZN(n9927) );
  OR2_X1 U4987 ( .A1(n5270), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5293) );
  INV_X1 U4988 ( .A(n7890), .ZN(n6376) );
  OR2_X1 U4989 ( .A1(n7502), .A2(n7493), .ZN(n7579) );
  NAND2_X1 U4990 ( .A1(n4332), .A2(n6107), .ZN(n6105) );
  AND4_X1 U4991 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(n6390)
         );
  AOI21_X1 U4992 ( .B1(n4888), .B2(n4891), .A(n4405), .ZN(n4887) );
  NAND2_X1 U4993 ( .A1(n5234), .A2(n5233), .ZN(n5256) );
  INV_X1 U4994 ( .A(n5235), .ZN(n5234) );
  NAND2_X1 U4995 ( .A1(n4487), .A2(n4488), .ZN(n4486) );
  AOI21_X1 U4996 ( .B1(n4912), .B2(n4913), .A(n4911), .ZN(n4910) );
  AND2_X1 U4997 ( .A1(n4892), .A2(n4889), .ZN(n4888) );
  AND2_X1 U4998 ( .A1(n5867), .A2(n9744), .ZN(n6113) );
  OR2_X1 U4999 ( .A1(n5199), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5235) );
  INV_X1 U5000 ( .A(n5082), .ZN(n5492) );
  OR2_X1 U5001 ( .A1(n5606), .A2(n5605), .ZN(n5608) );
  AND2_X1 U5002 ( .A1(n5129), .A2(n5114), .ZN(n5115) );
  OR2_X1 U5003 ( .A1(n5185), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5199) );
  INV_X1 U5004 ( .A(n5866), .ZN(n9744) );
  AND2_X1 U5005 ( .A1(n9035), .A2(n9038), .ZN(n9037) );
  CLKBUF_X1 U5006 ( .A(n5002), .Z(n4448) );
  NOR2_X1 U5007 ( .A1(n5145), .A2(n4893), .ZN(n4892) );
  AND2_X1 U5008 ( .A1(n5094), .A2(n5078), .ZN(n5079) );
  AND2_X1 U5009 ( .A1(n5866), .A2(n5867), .ZN(n4940) );
  AND2_X1 U5010 ( .A1(n5866), .A2(n5865), .ZN(n7591) );
  AND2_X1 U5011 ( .A1(n5861), .A2(n5862), .ZN(n5866) );
  NAND2_X1 U5012 ( .A1(n4974), .A2(n8432), .ZN(n5005) );
  INV_X1 U5013 ( .A(n4975), .ZN(n8432) );
  XNOR2_X1 U5014 ( .A(n4970), .B(n4969), .ZN(n4974) );
  OR2_X1 U5015 ( .A1(n5136), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U5016 ( .A1(n5862), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5864) );
  XNOR2_X1 U5017 ( .A(n5142), .B(SI_8_), .ZN(n5145) );
  NAND2_X1 U5018 ( .A1(n5095), .A2(SI_6_), .ZN(n5109) );
  MUX2_X1 U5019 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4635), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n4634) );
  NAND2_X1 U5020 ( .A1(n8426), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4970) );
  XNOR2_X1 U5021 ( .A(n4973), .B(n4972), .ZN(n4975) );
  NOR2_X1 U5022 ( .A1(n5972), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5841) );
  MUX2_X1 U5023 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5846), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5847) );
  XNOR2_X1 U5024 ( .A(n5850), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5886) );
  OR2_X1 U5025 ( .A1(n5603), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4978) );
  AND2_X1 U5026 ( .A1(n5287), .A2(n4414), .ZN(n5596) );
  CLKBUF_X1 U5027 ( .A(n7396), .Z(n4337) );
  NOR2_X1 U5028 ( .A1(n6749), .A2(n6748), .ZN(n6840) );
  CLKBUF_X1 U5029 ( .A(n5286), .Z(n5287) );
  NAND2_X2 U5030 ( .A1(n6050), .A2(P2_U3151), .ZN(n7151) );
  INV_X1 U5031 ( .A(n4737), .ZN(n6573) );
  AND3_X1 U5032 ( .A1(n4950), .A2(n4945), .A3(n4774), .ZN(n5286) );
  INV_X4 U5033 ( .A(n5012), .ZN(n6050) );
  NOR2_X1 U5034 ( .A1(n4966), .A2(n4965), .ZN(n4967) );
  AND2_X1 U5035 ( .A1(n4377), .A2(n4775), .ZN(n4774) );
  CLKBUF_X1 U5036 ( .A(n4676), .Z(n4471) );
  AND4_X1 U5037 ( .A1(n4949), .A2(n4948), .A3(n4947), .A4(n4946), .ZN(n4950)
         );
  INV_X1 U5038 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5803) );
  NOR2_X1 U5039 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5788) );
  INV_X1 U5040 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4944) );
  NOR2_X1 U5041 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4673) );
  NOR2_X1 U5042 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4674) );
  NOR2_X1 U5043 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5789) );
  NOR2_X1 U5044 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4946) );
  NOR2_X1 U5045 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5790) );
  INV_X1 U5046 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5973) );
  INV_X4 U5047 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X2 U5048 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10063) );
  INV_X1 U5049 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4932) );
  INV_X2 U5050 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4739) );
  INV_X1 U5051 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7205) );
  INV_X2 U5052 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U5053 ( .A1(n4990), .A2(n6314), .ZN(n4737) );
  OAI21_X2 U5054 ( .B1(n7129), .B2(n7300), .A(n7315), .ZN(n7140) );
  OR2_X1 U5055 ( .A1(n4943), .A2(n6882), .ZN(n9056) );
  NOR2_X4 U5056 ( .A1(n6894), .A2(n8624), .ZN(n9567) );
  OAI21_X2 U5057 ( .B1(n6809), .B2(n5552), .A(n5553), .ZN(n6922) );
  INV_X2 U5058 ( .A(n8929), .ZN(n8932) );
  OAI21_X1 U5059 ( .B1(n5662), .B2(n7432), .A(n5661), .ZN(n4336) );
  OAI21_X1 U5060 ( .B1(n5662), .B2(n7432), .A(n5661), .ZN(n5666) );
  BUF_X8 U5061 ( .A(n7396), .Z(n4338) );
  INV_X2 U5062 ( .A(n6050), .ZN(n7396) );
  OR2_X2 U5063 ( .A1(n6424), .A2(n6475), .ZN(n6482) );
  AOI21_X2 U5064 ( .B1(n9305), .B2(n9526), .A(n9304), .ZN(n9590) );
  OAI21_X2 U5065 ( .B1(n5205), .B2(n4367), .A(n4789), .ZN(n8252) );
  XNOR2_X2 U5066 ( .A(n6344), .B(n4335), .ZN(n6347) );
  NOR2_X2 U5067 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5816) );
  NOR2_X4 U5068 ( .A1(n9442), .A2(n9432), .ZN(n9431) );
  INV_X4 U5071 ( .A(n6166), .ZN(n8496) );
  OAI222_X1 U5072 ( .A1(n8278), .A2(n6721), .B1(n8276), .B2(n4992), .C1(n8358), 
        .C2(n6720), .ZN(n9929) );
  AND4_X2 U5073 ( .A1(n4996), .A2(n4995), .A3(n4994), .A4(n4993), .ZN(n4992)
         );
  OAI21_X2 U5074 ( .B1(n7786), .B2(n7727), .A(n7726), .ZN(n7725) );
  AOI21_X2 U5075 ( .B1(n7784), .B2(n7783), .A(n7782), .ZN(n7786) );
  NAND2_X1 U5076 ( .A1(n8429), .A2(n8432), .ZN(n4340) );
  NAND2_X1 U5077 ( .A1(n5886), .A2(n9748), .ZN(n4341) );
  OAI21_X2 U5078 ( .B1(n8206), .B2(n5567), .A(n5566), .ZN(n8195) );
  INV_X1 U5079 ( .A(n4618), .ZN(n4617) );
  OAI22_X1 U5080 ( .A1(n4620), .A2(n4621), .B1(n4623), .B2(n4624), .ZN(n4618)
         );
  AND2_X1 U5081 ( .A1(n7359), .A2(n7360), .ZN(n4624) );
  NOR2_X1 U5082 ( .A1(n8112), .A2(n4399), .ZN(n4621) );
  NAND2_X1 U5083 ( .A1(n4616), .A2(n4374), .ZN(n4615) );
  AND2_X1 U5084 ( .A1(n4620), .A2(n4623), .ZN(n4619) );
  AND2_X1 U5085 ( .A1(n7317), .A2(n7316), .ZN(n7141) );
  NAND2_X1 U5086 ( .A1(n9744), .A2(n5865), .ZN(n7487) );
  AOI21_X1 U5087 ( .B1(n4613), .B2(n4615), .A(n4404), .ZN(n4612) );
  INV_X1 U5088 ( .A(n4614), .ZN(n4613) );
  NOR2_X1 U5089 ( .A1(n4708), .A2(n7817), .ZN(n4707) );
  NAND2_X1 U5090 ( .A1(n4407), .A2(n5694), .ZN(n4708) );
  NOR2_X1 U5091 ( .A1(n7416), .A2(n7415), .ZN(n7420) );
  OR2_X1 U5092 ( .A1(n7467), .A2(n7468), .ZN(n7423) );
  AND2_X1 U5093 ( .A1(n9852), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4488) );
  INV_X1 U5094 ( .A(n4714), .ZN(n4490) );
  NAND2_X1 U5095 ( .A1(n9835), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4713) );
  NAND2_X1 U5096 ( .A1(n7367), .A2(n7368), .ZN(n8081) );
  OR2_X1 U5097 ( .A1(n7771), .A2(n8134), .ZN(n7360) );
  AOI21_X1 U5098 ( .B1(n4644), .B2(n4646), .A(n4393), .ZN(n4643) );
  OR2_X1 U5099 ( .A1(n7724), .A2(n8174), .ZN(n7247) );
  OR2_X1 U5100 ( .A1(n8411), .A2(n8240), .ZN(n7342) );
  INV_X1 U5101 ( .A(n7322), .ZN(n4791) );
  NAND2_X1 U5102 ( .A1(n4661), .A2(n4365), .ZN(n4657) );
  OAI21_X1 U5103 ( .B1(n8117), .B2(n4670), .A(n4668), .ZN(n8082) );
  INV_X1 U5104 ( .A(n4669), .ZN(n4668) );
  OAI22_X1 U5105 ( .A1(n4366), .A2(n4670), .B1(n8109), .B2(n7854), .ZN(n4669)
         );
  NAND2_X1 U5106 ( .A1(n4403), .A2(n5578), .ZN(n4670) );
  CLKBUF_X1 U5107 ( .A(n5082), .Z(n5327) );
  NAND2_X1 U5108 ( .A1(n4588), .A2(n4587), .ZN(n4586) );
  NAND2_X1 U5109 ( .A1(n6971), .A2(n6972), .ZN(n4587) );
  INV_X1 U5110 ( .A(n6970), .ZN(n4588) );
  INV_X1 U5111 ( .A(n9019), .ZN(n4540) );
  NAND2_X1 U5112 ( .A1(n4815), .A2(n7617), .ZN(n4814) );
  INV_X1 U5113 ( .A(n4817), .ZN(n4815) );
  NAND2_X1 U5114 ( .A1(n9712), .A2(n8771), .ZN(n4824) );
  NAND2_X1 U5115 ( .A1(n9412), .A2(n8911), .ZN(n9396) );
  AND2_X1 U5116 ( .A1(n4807), .A2(n4805), .ZN(n4802) );
  OR2_X1 U5117 ( .A1(n9733), .A2(n8689), .ZN(n8948) );
  OR2_X1 U5118 ( .A1(n8935), .A2(n4758), .ZN(n6852) );
  INV_X1 U5119 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5807) );
  AND2_X1 U5120 ( .A1(n5726), .A2(n5724), .ZN(n4678) );
  OR2_X1 U5121 ( .A1(n7801), .A2(n7873), .ZN(n5726) );
  OR2_X1 U5122 ( .A1(n5382), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5399) );
  AND2_X1 U5123 ( .A1(n5520), .A2(n5519), .ZN(n8083) );
  INV_X1 U5124 ( .A(n5063), .ZN(n5515) );
  NAND2_X1 U5125 ( .A1(n4494), .A2(n4493), .ZN(n4492) );
  INV_X1 U5126 ( .A(n7960), .ZN(n4493) );
  OR2_X1 U5127 ( .A1(n8316), .A2(n8161), .ZN(n7249) );
  NAND2_X1 U5128 ( .A1(n4651), .A2(n4650), .ZN(n8171) );
  OR2_X1 U5129 ( .A1(n8201), .A2(n8184), .ZN(n8187) );
  OR2_X1 U5130 ( .A1(n9963), .A2(n8258), .ZN(n7322) );
  AOI21_X1 U5131 ( .B1(n4662), .B2(n5558), .A(n4348), .ZN(n4660) );
  NAND2_X1 U5132 ( .A1(n4666), .A2(n4665), .ZN(n4664) );
  INV_X1 U5133 ( .A(n7130), .ZN(n4666) );
  INV_X1 U5134 ( .A(n8209), .ZN(n8276) );
  INV_X1 U5135 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5635) );
  AND2_X1 U5136 ( .A1(n7644), .A2(n6214), .ZN(n7656) );
  NOR2_X1 U5137 ( .A1(n6509), .A2(n6510), .ZN(n6655) );
  AND2_X1 U5138 ( .A1(n8573), .A2(n4578), .ZN(n4577) );
  NAND2_X1 U5139 ( .A1(n4857), .A2(n4579), .ZN(n4578) );
  INV_X1 U5140 ( .A(n4581), .ZN(n4579) );
  AOI21_X1 U5141 ( .B1(n9309), .B2(n4443), .A(n7488), .ZN(n8803) );
  AND4_X1 U5142 ( .A1(n7557), .A2(n7556), .A3(n7555), .A4(n7554), .ZN(n8818)
         );
  AND2_X1 U5143 ( .A1(n8876), .A2(n8838), .ZN(n9272) );
  OR2_X1 U5144 ( .A1(n9339), .A2(n9118), .ZN(n4835) );
  AND2_X1 U5145 ( .A1(n4824), .A2(n4819), .ZN(n4818) );
  NAND2_X1 U5146 ( .A1(n9432), .A2(n9124), .ZN(n7583) );
  OR2_X1 U5147 ( .A1(n9729), .A2(n8762), .ZN(n9524) );
  AOI21_X1 U5148 ( .B1(n4344), .B2(n4800), .A(n9542), .ZN(n4797) );
  NAND2_X1 U5149 ( .A1(n8842), .A2(n6395), .ZN(n4544) );
  OR2_X1 U5150 ( .A1(n6440), .A2(n9142), .ZN(n6386) );
  INV_X1 U5151 ( .A(n6434), .ZN(n8842) );
  NAND2_X2 U5152 ( .A1(n5886), .A2(n9748), .ZN(n6263) );
  NOR2_X1 U5153 ( .A1(n5408), .A2(n4916), .ZN(n4915) );
  INV_X1 U5154 ( .A(n5389), .ZN(n4916) );
  INV_X1 U5155 ( .A(n7915), .ZN(n4495) );
  NOR2_X1 U5156 ( .A1(n8920), .A2(n4351), .ZN(n4517) );
  NAND2_X1 U5157 ( .A1(n8917), .A2(n4349), .ZN(n4522) );
  INV_X1 U5158 ( .A(n8921), .ZN(n4521) );
  NAND2_X1 U5159 ( .A1(n8928), .A2(n4428), .ZN(n4518) );
  INV_X1 U5160 ( .A(n8928), .ZN(n4519) );
  NAND2_X1 U5161 ( .A1(n7314), .A2(n7316), .ZN(n4602) );
  OR3_X1 U5162 ( .A1(n4529), .A2(n8968), .A3(n4527), .ZN(n8969) );
  AOI21_X1 U5163 ( .B1(n4531), .B2(n4530), .A(n9030), .ZN(n4529) );
  OAI21_X1 U5164 ( .B1(n7350), .B2(n7386), .A(n7427), .ZN(n4599) );
  NAND2_X1 U5165 ( .A1(n8983), .A2(n4551), .ZN(n4549) );
  NAND2_X1 U5166 ( .A1(n8973), .A2(n9030), .ZN(n4551) );
  INV_X1 U5167 ( .A(n8984), .ZN(n4550) );
  INV_X1 U5168 ( .A(n8983), .ZN(n4547) );
  NAND2_X1 U5169 ( .A1(n4595), .A2(n7353), .ZN(n4594) );
  OAI21_X1 U5170 ( .B1(n7349), .B2(n7388), .A(n4596), .ZN(n4595) );
  NAND2_X1 U5171 ( .A1(n7354), .A2(n7386), .ZN(n4593) );
  INV_X1 U5172 ( .A(n5129), .ZN(n4893) );
  NOR2_X1 U5173 ( .A1(n7372), .A2(n7371), .ZN(n7374) );
  NAND2_X1 U5174 ( .A1(n9841), .A2(n6338), .ZN(n6339) );
  INV_X1 U5175 ( .A(n8377), .ZN(n5579) );
  AND2_X1 U5176 ( .A1(n8457), .A2(n8456), .ZN(n4851) );
  INV_X1 U5177 ( .A(n5303), .ZN(n4907) );
  NAND2_X1 U5178 ( .A1(n5306), .A2(n5305), .ZN(n5323) );
  INV_X1 U5179 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4738) );
  NAND2_X1 U5180 ( .A1(n4471), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U5181 ( .A1(n6320), .A2(n9820), .ZN(n6321) );
  NAND2_X1 U5182 ( .A1(n4728), .A2(n4485), .ZN(n4727) );
  INV_X1 U5183 ( .A(n6339), .ZN(n4728) );
  NAND2_X1 U5184 ( .A1(n4482), .A2(n9858), .ZN(n6350) );
  NAND2_X1 U5185 ( .A1(n6643), .A2(n4420), .ZN(n6645) );
  OR2_X1 U5186 ( .A1(n5579), .A2(n8072), .ZN(n7367) );
  INV_X1 U5187 ( .A(n8156), .ZN(n4649) );
  OR2_X1 U5188 ( .A1(n7781), .A2(n8185), .ZN(n7245) );
  AND2_X1 U5189 ( .A1(n8198), .A2(n7257), .ZN(n4786) );
  OR2_X1 U5190 ( .A1(n8346), .A2(n8248), .ZN(n7337) );
  INV_X1 U5191 ( .A(n4660), .ZN(n4658) );
  NAND2_X1 U5192 ( .A1(n7889), .A2(n6952), .ZN(n7276) );
  INV_X1 U5193 ( .A(SI_9_), .ZN(n10076) );
  NAND2_X1 U5194 ( .A1(n4761), .A2(n4762), .ZN(n7087) );
  AOI21_X1 U5195 ( .B1(n4764), .B2(n4767), .A(n4763), .ZN(n4762) );
  INV_X1 U5196 ( .A(n7304), .ZN(n4763) );
  OR2_X1 U5197 ( .A1(n7266), .A2(n6938), .ZN(n7432) );
  NAND2_X1 U5198 ( .A1(n5617), .A2(n7241), .ZN(n5633) );
  INV_X1 U5199 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5595) );
  INV_X1 U5200 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4775) );
  NOR2_X1 U5201 ( .A1(n4952), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4712) );
  INV_X1 U5202 ( .A(n4471), .ZN(n6314) );
  OAI21_X1 U5203 ( .B1(n8478), .B2(n8477), .A(n8758), .ZN(n8481) );
  INV_X1 U5204 ( .A(n8814), .ZN(n4572) );
  OR2_X1 U5205 ( .A1(n4360), .A2(n4851), .ZN(n4850) );
  XNOR2_X1 U5206 ( .A(n6507), .B(n8644), .ZN(n6509) );
  NOR2_X1 U5207 ( .A1(n4860), .A2(n4582), .ZN(n4581) );
  INV_X1 U5208 ( .A(n8558), .ZN(n4860) );
  INV_X1 U5209 ( .A(n8728), .ZN(n4582) );
  NAND2_X1 U5210 ( .A1(n8596), .A2(n4469), .ZN(n8485) );
  OR2_X1 U5211 ( .A1(n9593), .A2(n8803), .ZN(n9007) );
  AND2_X1 U5212 ( .A1(n9587), .A2(n8837), .ZN(n9016) );
  OR2_X1 U5213 ( .A1(n9269), .A2(n9280), .ZN(n9006) );
  OR2_X1 U5214 ( .A1(n9323), .A2(n8999), .ZN(n8990) );
  NOR2_X1 U5215 ( .A1(n9337), .A2(n9323), .ZN(n4863) );
  NAND2_X1 U5216 ( .A1(n9367), .A2(n8879), .ZN(n4744) );
  INV_X1 U5217 ( .A(n4744), .ZN(n4743) );
  AND2_X1 U5218 ( .A1(n9649), .A2(n9129), .ZN(n7571) );
  AND2_X1 U5219 ( .A1(n8624), .A2(n8461), .ZN(n8945) );
  NAND2_X1 U5220 ( .A1(n7379), .A2(n7378), .ZN(n7395) );
  OR2_X1 U5221 ( .A1(n7377), .A2(n7376), .ZN(n7378) );
  NAND2_X1 U5222 ( .A1(n4923), .A2(SI_29_), .ZN(n7379) );
  NAND2_X1 U5223 ( .A1(n4881), .A2(n4879), .ZN(n5524) );
  AOI21_X1 U5224 ( .B1(n4883), .B2(n4885), .A(n4880), .ZN(n4879) );
  INV_X1 U5225 ( .A(n5504), .ZN(n4880) );
  AND2_X1 U5226 ( .A1(n5504), .A2(n5491), .ZN(n5502) );
  AND2_X1 U5227 ( .A1(n5486), .A2(n5473), .ZN(n5484) );
  NAND2_X1 U5228 ( .A1(n5468), .A2(n5467), .ZN(n5485) );
  NAND2_X1 U5229 ( .A1(n5466), .A2(n5465), .ZN(n5468) );
  AOI21_X1 U5230 ( .B1(n4906), .B2(n5300), .A(n4905), .ZN(n4904) );
  INV_X1 U5231 ( .A(n5323), .ZN(n4905) );
  NAND2_X1 U5232 ( .A1(n5301), .A2(n4906), .ZN(n4903) );
  AND2_X1 U5233 ( .A1(n4927), .A2(n4924), .ZN(n5280) );
  INV_X1 U5234 ( .A(n4928), .ZN(n4924) );
  NAND2_X1 U5235 ( .A1(n5209), .A2(SI_12_), .ZN(n5221) );
  NOR2_X1 U5236 ( .A1(n5207), .A2(n4901), .ZN(n4900) );
  INV_X1 U5237 ( .A(n5191), .ZN(n4901) );
  NAND2_X1 U5238 ( .A1(n5165), .A2(SI_10_), .ZN(n5191) );
  XNOR2_X1 U5239 ( .A(n5161), .B(n10076), .ZN(n5163) );
  OAI21_X1 U5240 ( .B1(n5012), .B2(n4437), .A(n4436), .ZN(n5013) );
  NAND2_X1 U5241 ( .A1(n5012), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5242 ( .A1(n5013), .A2(SI_2_), .ZN(n5022) );
  NAND2_X1 U5243 ( .A1(n5732), .A2(n7808), .ZN(n4680) );
  INV_X1 U5244 ( .A(n6051), .ZN(n4672) );
  NAND2_X1 U5245 ( .A1(n5367), .A2(n7787), .ZN(n5382) );
  INV_X1 U5246 ( .A(n5699), .ZN(n4709) );
  AND2_X1 U5247 ( .A1(n4710), .A2(n4704), .ZN(n4703) );
  INV_X1 U5248 ( .A(n5700), .ZN(n4710) );
  NAND2_X1 U5249 ( .A1(n4707), .A2(n4705), .ZN(n4704) );
  INV_X1 U5250 ( .A(n4707), .ZN(n4706) );
  XNOR2_X1 U5251 ( .A(n8316), .B(n5725), .ZN(n7801) );
  OAI21_X1 U5252 ( .B1(n7862), .B2(n4696), .A(n4693), .ZN(n7833) );
  AND2_X1 U5253 ( .A1(n5463), .A2(n5462), .ZN(n5737) );
  OAI21_X1 U5254 ( .B1(n9825), .B2(P2_REG1_REG_2__SCAN_IN), .A(n4510), .ZN(
        n9822) );
  NAND2_X1 U5255 ( .A1(n9825), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4510) );
  OR2_X1 U5256 ( .A1(n6346), .A2(n6345), .ZN(n4714) );
  XNOR2_X1 U5257 ( .A(n6645), .B(n6647), .ZN(n4717) );
  NAND2_X1 U5258 ( .A1(n4717), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9888) );
  INV_X1 U5259 ( .A(n9899), .ZN(n4503) );
  INV_X1 U5260 ( .A(n9898), .ZN(n4504) );
  NOR2_X1 U5261 ( .A1(n7014), .A2(n4391), .ZN(n7017) );
  NAND2_X1 U5262 ( .A1(n4512), .A2(n4511), .ZN(n4736) );
  INV_X1 U5263 ( .A(n7016), .ZN(n4511) );
  INV_X1 U5264 ( .A(n7017), .ZN(n4512) );
  NOR2_X1 U5265 ( .A1(n7162), .A2(n4720), .ZN(n7163) );
  NOR2_X1 U5266 ( .A1(n5181), .A2(n7135), .ZN(n4720) );
  NOR2_X1 U5267 ( .A1(n7892), .A2(n4734), .ZN(n7926) );
  NOR2_X1 U5268 ( .A1(n7177), .A2(n7158), .ZN(n4734) );
  XNOR2_X1 U5269 ( .A(n8002), .B(n8008), .ZN(n7989) );
  OR2_X1 U5270 ( .A1(n5476), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5495) );
  OR2_X1 U5271 ( .A1(n7364), .A2(n7365), .ZN(n8097) );
  NAND2_X1 U5272 ( .A1(n8117), .A2(n4366), .ZN(n8104) );
  AND2_X1 U5273 ( .A1(n7359), .A2(n7249), .ZN(n4781) );
  AND2_X1 U5274 ( .A1(n7360), .A2(n7361), .ZN(n8127) );
  OR2_X1 U5275 ( .A1(n7425), .A2(n7424), .ZN(n8135) );
  NAND2_X1 U5276 ( .A1(n5574), .A2(n5573), .ZN(n8148) );
  NAND2_X1 U5277 ( .A1(n8143), .A2(n8146), .ZN(n8142) );
  AND2_X1 U5278 ( .A1(n5406), .A2(n5405), .ZN(n8161) );
  AND3_X1 U5279 ( .A1(n5386), .A2(n5385), .A3(n5384), .ZN(n8174) );
  NAND2_X1 U5280 ( .A1(n4652), .A2(n4653), .ZN(n4651) );
  NAND2_X1 U5281 ( .A1(n5322), .A2(n4786), .ZN(n8186) );
  AND2_X1 U5282 ( .A1(n8187), .A2(n7346), .ZN(n8198) );
  AOI21_X1 U5283 ( .B1(n4639), .B2(n4637), .A(n4392), .ZN(n4636) );
  INV_X1 U5284 ( .A(n4639), .ZN(n4638) );
  INV_X1 U5285 ( .A(n5293), .ZN(n5292) );
  AND4_X1 U5286 ( .A1(n5298), .A2(n5297), .A3(n5296), .A4(n5295), .ZN(n8240)
         );
  NOR2_X1 U5287 ( .A1(n8238), .A2(n4640), .ZN(n4639) );
  INV_X1 U5288 ( .A(n5561), .ZN(n4640) );
  NAND2_X1 U5289 ( .A1(n8246), .A2(n5560), .ZN(n4641) );
  AND2_X1 U5290 ( .A1(n7337), .A2(n7340), .ZN(n8238) );
  INV_X1 U5291 ( .A(n4790), .ZN(n4789) );
  OAI21_X1 U5292 ( .B1(n4343), .B2(n4367), .A(n5241), .ZN(n4790) );
  NAND2_X1 U5293 ( .A1(n7140), .A2(n7141), .ZN(n5205) );
  NAND2_X1 U5294 ( .A1(n5205), .A2(n4343), .ZN(n8271) );
  INV_X1 U5295 ( .A(n4667), .ZN(n4663) );
  NAND2_X1 U5296 ( .A1(n4664), .A2(n4667), .ZN(n7142) );
  NAND2_X1 U5297 ( .A1(n6763), .A2(n7439), .ZN(n4675) );
  OR2_X1 U5298 ( .A1(n5088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5123) );
  OR2_X1 U5299 ( .A1(n6771), .A2(n5537), .ZN(n7134) );
  INV_X1 U5300 ( .A(n8278), .ZN(n8211) );
  NAND2_X1 U5301 ( .A1(n7403), .A2(n7402), .ZN(n7467) );
  AOI21_X1 U5302 ( .B1(n8085), .B2(n8214), .A(n8084), .ZN(n8297) );
  NAND2_X1 U5303 ( .A1(n5433), .A2(n5432), .ZN(n7771) );
  NAND2_X1 U5304 ( .A1(n5416), .A2(n5415), .ZN(n5727) );
  NAND2_X1 U5305 ( .A1(n5354), .A2(n5353), .ZN(n7715) );
  NAND2_X1 U5306 ( .A1(n5333), .A2(n5332), .ZN(n8201) );
  NAND2_X1 U5307 ( .A1(n5314), .A2(n5313), .ZN(n8336) );
  AND2_X1 U5308 ( .A1(n7152), .A2(n6676), .ZN(n9952) );
  INV_X1 U5309 ( .A(n8214), .ZN(n8358) );
  INV_X1 U5310 ( .A(n8423), .ZN(n6071) );
  NAND2_X1 U5311 ( .A1(n5597), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5606) );
  INV_X1 U5312 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5605) );
  INV_X1 U5313 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4960) );
  OR2_X1 U5314 ( .A1(n4356), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5054) );
  AND2_X1 U5315 ( .A1(n7656), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7658) );
  AND2_X1 U5316 ( .A1(n8728), .A2(n8548), .ZN(n8607) );
  XNOR2_X1 U5317 ( .A(n4862), .B(n8644), .ZN(n6160) );
  OAI21_X1 U5318 ( .B1(n6267), .B2(n6826), .A(n6132), .ZN(n4862) );
  NAND2_X1 U5319 ( .A1(n6271), .A2(n6270), .ZN(n6503) );
  NOR2_X1 U5320 ( .A1(n6271), .A2(n4564), .ZN(n4563) );
  NAND2_X1 U5321 ( .A1(n6504), .A2(n4559), .ZN(n4558) );
  INV_X1 U5322 ( .A(n4561), .ZN(n4559) );
  NAND2_X1 U5323 ( .A1(n4565), .A2(n6269), .ZN(n6504) );
  NAND2_X1 U5324 ( .A1(n4859), .A2(n8558), .ZN(n4858) );
  AND3_X1 U5325 ( .A1(n4538), .A2(n4411), .A3(n4535), .ZN(n9028) );
  NAND2_X1 U5326 ( .A1(n4540), .A2(n4383), .ZN(n4538) );
  NAND2_X1 U5327 ( .A1(n4537), .A2(n4536), .ZN(n4535) );
  AND3_X1 U5328 ( .A1(n7505), .A2(n7504), .A3(n7503), .ZN(n8709) );
  AND3_X1 U5329 ( .A1(n7512), .A2(n7511), .A3(n7510), .ZN(n8820) );
  OR2_X1 U5330 ( .A1(n5918), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6011) );
  OAI21_X1 U5331 ( .B1(n9331), .B2(n4828), .A(n4830), .ZN(n9271) );
  AOI21_X1 U5332 ( .B1(n4342), .B2(n4831), .A(n4398), .ZN(n4830) );
  NAND2_X1 U5333 ( .A1(n4342), .A2(n4829), .ZN(n4828) );
  NOR2_X1 U5334 ( .A1(n7664), .A2(n4833), .ZN(n4832) );
  INV_X1 U5335 ( .A(n4835), .ZN(n4833) );
  NOR2_X2 U5336 ( .A1(n9593), .A2(n9306), .ZN(n9307) );
  NAND2_X1 U5337 ( .A1(n8990), .A2(n9092), .ZN(n9321) );
  NAND2_X1 U5338 ( .A1(n4824), .A2(n4379), .ZN(n4817) );
  AND2_X1 U5339 ( .A1(n8879), .A2(n8886), .ZN(n9381) );
  NAND2_X1 U5340 ( .A1(n9382), .A2(n9381), .ZN(n9380) );
  OR2_X1 U5341 ( .A1(n4822), .A2(n4821), .ZN(n4819) );
  INV_X1 U5342 ( .A(n4825), .ZN(n4821) );
  AND2_X1 U5343 ( .A1(n7596), .A2(n4363), .ZN(n4822) );
  AOI21_X1 U5344 ( .B1(n4757), .B2(n8965), .A(n9474), .ZN(n4752) );
  NAND2_X1 U5345 ( .A1(n9509), .A2(n4756), .ZN(n9496) );
  INV_X1 U5346 ( .A(n4757), .ZN(n4756) );
  INV_X1 U5347 ( .A(n9509), .ZN(n4755) );
  NOR2_X1 U5348 ( .A1(n4806), .A2(n7558), .ZN(n4805) );
  INV_X1 U5349 ( .A(n4810), .ZN(n4806) );
  NAND2_X1 U5350 ( .A1(n4870), .A2(n8690), .ZN(n4810) );
  INV_X1 U5351 ( .A(n9523), .ZN(n9521) );
  NAND2_X1 U5352 ( .A1(n9558), .A2(n4799), .ZN(n4798) );
  INV_X1 U5353 ( .A(n7525), .ZN(n4799) );
  INV_X1 U5354 ( .A(n9558), .ZN(n4800) );
  OR2_X1 U5355 ( .A1(n8450), .A2(n9135), .ZN(n6869) );
  INV_X1 U5356 ( .A(n8848), .ZN(n6886) );
  INV_X1 U5357 ( .A(n6383), .ZN(n4444) );
  NOR2_X1 U5358 ( .A1(n9586), .A2(n4746), .ZN(n4745) );
  AND2_X1 U5359 ( .A1(n9587), .A2(n9658), .ZN(n4746) );
  NAND2_X1 U5360 ( .A1(n7643), .A2(n7642), .ZN(n9339) );
  NAND2_X1 U5361 ( .A1(n7640), .A2(n8861), .ZN(n7643) );
  NAND2_X1 U5362 ( .A1(n7588), .A2(n7587), .ZN(n9625) );
  NAND2_X1 U5363 ( .A1(n7577), .A2(n7576), .ZN(n9432) );
  NAND2_X1 U5364 ( .A1(n7492), .A2(n7491), .ZN(n9634) );
  INV_X1 U5365 ( .A(n9565), .ZN(n9526) );
  NOR2_X1 U5366 ( .A1(n4397), .A2(n4865), .ZN(n4864) );
  XNOR2_X1 U5367 ( .A(n5524), .B(n5523), .ZN(n8434) );
  XNOR2_X1 U5368 ( .A(n5503), .B(n5502), .ZN(n7688) );
  NAND2_X1 U5369 ( .A1(n4882), .A2(n5486), .ZN(n5503) );
  NAND2_X1 U5370 ( .A1(n5485), .A2(n5484), .ZN(n4882) );
  NAND2_X1 U5371 ( .A1(n6204), .A2(n5806), .ZN(n5813) );
  AND2_X1 U5372 ( .A1(n5427), .A2(n5414), .ZN(n5425) );
  INV_X1 U5373 ( .A(n5407), .ZN(n4914) );
  OAI21_X1 U5374 ( .B1(n5192), .B2(n4897), .A(n4894), .ZN(n5228) );
  INV_X1 U5375 ( .A(n4898), .ZN(n4897) );
  AOI21_X1 U5376 ( .B1(n4896), .B2(n4898), .A(n4895), .ZN(n4894) );
  INV_X1 U5377 ( .A(n5221), .ZN(n4895) );
  NAND2_X1 U5378 ( .A1(n5228), .A2(n5227), .ZN(n5244) );
  OAI21_X1 U5379 ( .B1(n5209), .B2(SI_12_), .A(n5221), .ZN(n5210) );
  AND2_X1 U5380 ( .A1(n4902), .A2(n4372), .ZN(n4898) );
  INV_X1 U5381 ( .A(n5210), .ZN(n4902) );
  NAND2_X1 U5382 ( .A1(n5192), .A2(n4900), .ZN(n4899) );
  AND2_X1 U5383 ( .A1(n5049), .A2(n5073), .ZN(n5050) );
  OAI21_X1 U5384 ( .B1(n5013), .B2(SI_2_), .A(n5022), .ZN(n5014) );
  AND2_X1 U5385 ( .A1(n6251), .A2(n5673), .ZN(n6288) );
  NOR2_X1 U5386 ( .A1(n4684), .A2(n7861), .ZN(n4682) );
  NOR2_X1 U5387 ( .A1(n4346), .A2(n4685), .ZN(n4684) );
  INV_X1 U5388 ( .A(n4687), .ZN(n4685) );
  NAND2_X1 U5389 ( .A1(n4687), .A2(n4688), .ZN(n4686) );
  INV_X1 U5390 ( .A(n5749), .ZN(n4688) );
  OAI21_X1 U5391 ( .B1(n8373), .B2(n7853), .A(n5781), .ZN(n5782) );
  AOI21_X1 U5392 ( .B1(n6902), .B2(n6992), .A(n4424), .ZN(n4700) );
  INV_X1 U5393 ( .A(n6374), .ZN(n5668) );
  AND2_X1 U5394 ( .A1(n5441), .A2(n5440), .ZN(n8134) );
  NAND2_X1 U5395 ( .A1(n6288), .A2(n6287), .ZN(n6286) );
  INV_X1 U5396 ( .A(n5737), .ZN(n8120) );
  INV_X1 U5397 ( .A(n8134), .ZN(n7872) );
  NAND4_X1 U5398 ( .A1(n5190), .A2(n5189), .A3(n5188), .A4(n5187), .ZN(n7882)
         );
  OR2_X1 U5399 ( .A1(n7912), .A2(n7913), .ZN(n4496) );
  NAND2_X1 U5400 ( .A1(n4452), .A2(n4371), .ZN(n4494) );
  INV_X1 U5401 ( .A(n4508), .ZN(n7978) );
  INV_X1 U5402 ( .A(n4492), .ZN(n7987) );
  NAND2_X1 U5403 ( .A1(n4730), .A2(n8011), .ZN(n4729) );
  INV_X1 U5404 ( .A(n4732), .ZN(n4730) );
  OR2_X1 U5405 ( .A1(n9891), .A2(n4433), .ZN(n4476) );
  NAND2_X1 U5406 ( .A1(n4633), .A2(n4630), .ZN(n8291) );
  NOR2_X1 U5407 ( .A1(n4632), .A2(n4631), .ZN(n4630) );
  OR2_X1 U5408 ( .A1(n8071), .A2(n8358), .ZN(n4633) );
  NOR2_X1 U5409 ( .A1(n8276), .A2(n8072), .ZN(n4631) );
  NAND2_X1 U5410 ( .A1(n5215), .A2(n5214), .ZN(n9963) );
  NOR2_X1 U5411 ( .A1(n8291), .A2(n4628), .ZN(n8371) );
  NOR2_X1 U5412 ( .A1(n4629), .A2(n9959), .ZN(n4628) );
  INV_X1 U5413 ( .A(n8292), .ZN(n4629) );
  NAND2_X1 U5414 ( .A1(n4406), .A2(n4555), .ZN(n6969) );
  NAND2_X1 U5415 ( .A1(n4560), .A2(n4557), .ZN(n4556) );
  NAND2_X1 U5416 ( .A1(n7632), .A2(n7631), .ZN(n9358) );
  OAI21_X1 U5417 ( .B1(n9340), .B2(n7663), .A(n7650), .ZN(n9118) );
  INV_X1 U5418 ( .A(n4748), .ZN(n4747) );
  OAI22_X1 U5419 ( .A1(n9280), .A2(n9281), .B1(n9279), .B2(n9278), .ZN(n4748)
         );
  OR2_X1 U5420 ( .A1(n7533), .A2(n8836), .ZN(n7536) );
  OAI211_X1 U5421 ( .C1(n5526), .C2(n4921), .A(n4919), .B(n4917), .ZN(n9743)
         );
  INV_X1 U5422 ( .A(n4922), .ZN(n4921) );
  NAND2_X1 U5423 ( .A1(n4922), .A2(n4920), .ZN(n4919) );
  NAND2_X1 U5424 ( .A1(n5526), .A2(n4918), .ZN(n4917) );
  OAI21_X1 U5425 ( .B1(n4520), .B2(n4519), .A(n4401), .ZN(n4523) );
  NAND2_X1 U5426 ( .A1(n4602), .A2(n4601), .ZN(n4600) );
  OR2_X1 U5427 ( .A1(n7321), .A2(n7388), .ZN(n4603) );
  AND2_X1 U5428 ( .A1(n7317), .A2(n7388), .ZN(n4601) );
  AND2_X1 U5429 ( .A1(n8964), .A2(n9071), .ZN(n4530) );
  AOI21_X1 U5430 ( .B1(n4528), .B2(n9076), .A(n9021), .ZN(n4527) );
  OAI22_X1 U5431 ( .A1(n8112), .A2(n4375), .B1(n7358), .B2(n7386), .ZN(n4620)
         );
  INV_X1 U5432 ( .A(n4597), .ZN(n4596) );
  OAI21_X1 U5433 ( .B1(n7351), .B2(n7352), .A(n4598), .ZN(n4597) );
  INV_X1 U5434 ( .A(n4599), .ZN(n4598) );
  AOI21_X1 U5435 ( .B1(n4368), .B2(n4548), .A(n4546), .ZN(n8994) );
  OAI21_X1 U5436 ( .B1(n4550), .B2(n4547), .A(n9381), .ZN(n4546) );
  INV_X1 U5437 ( .A(n8097), .ZN(n4622) );
  AOI21_X1 U5438 ( .B1(n4594), .B2(n4593), .A(n7355), .ZN(n7356) );
  INV_X1 U5439 ( .A(n4760), .ZN(n9060) );
  INV_X1 U5440 ( .A(n4645), .ZN(n4644) );
  OAI21_X1 U5441 ( .B1(n5573), .B2(n4646), .A(n5576), .ZN(n4645) );
  INV_X1 U5442 ( .A(n5575), .ZN(n4646) );
  OR2_X1 U5443 ( .A1(n9957), .A2(n8275), .ZN(n7317) );
  AND2_X1 U5444 ( .A1(n7302), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U5445 ( .A1(n7441), .A2(n4766), .ZN(n4765) );
  INV_X1 U5446 ( .A(n7441), .ZN(n4767) );
  INV_X1 U5447 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4776) );
  INV_X1 U5448 ( .A(n5102), .ZN(n4945) );
  AOI21_X1 U5449 ( .B1(n9018), .B2(n9272), .A(n9017), .ZN(n9020) );
  XNOR2_X1 U5450 ( .A(n7377), .B(n7375), .ZN(n4923) );
  INV_X1 U5451 ( .A(n5486), .ZN(n4885) );
  INV_X1 U5452 ( .A(n4884), .ZN(n4883) );
  OAI21_X1 U5453 ( .B1(n5484), .B2(n4885), .A(n5502), .ZN(n4884) );
  INV_X1 U5454 ( .A(n4915), .ZN(n4912) );
  INV_X1 U5455 ( .A(n5425), .ZN(n4911) );
  NOR2_X1 U5456 ( .A1(n4928), .A2(n4926), .ZN(n4925) );
  INV_X1 U5457 ( .A(SI_15_), .ZN(n4926) );
  NOR2_X1 U5458 ( .A1(n5263), .A2(SI_14_), .ZN(n4928) );
  NAND2_X1 U5459 ( .A1(n5244), .A2(n4389), .ZN(n4927) );
  NAND2_X1 U5460 ( .A1(n5263), .A2(SI_14_), .ZN(n4929) );
  INV_X1 U5461 ( .A(n5109), .ZN(n4890) );
  INV_X1 U5462 ( .A(n5115), .ZN(n4891) );
  INV_X1 U5463 ( .A(n7025), .ZN(n4705) );
  INV_X1 U5464 ( .A(n5666), .ZN(n5725) );
  INV_X1 U5465 ( .A(n7863), .ZN(n4697) );
  NOR2_X1 U5466 ( .A1(n7419), .A2(n6938), .ZN(n4771) );
  NAND2_X1 U5467 ( .A1(n7418), .A2(n7266), .ZN(n7419) );
  NAND2_X1 U5468 ( .A1(n7465), .A2(n7467), .ZN(n7418) );
  NAND2_X1 U5469 ( .A1(n4592), .A2(n4386), .ZN(n4590) );
  OR2_X1 U5470 ( .A1(n7383), .A2(n7243), .ZN(n4592) );
  NOR2_X1 U5471 ( .A1(n7465), .A2(n4773), .ZN(n4591) );
  INV_X1 U5472 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4962) );
  NAND2_X1 U5473 ( .A1(n4500), .A2(n9836), .ZN(n9841) );
  NAND2_X1 U5474 ( .A1(n9839), .A2(n9837), .ZN(n4500) );
  NAND2_X1 U5475 ( .A1(n4513), .A2(n6341), .ZN(n9859) );
  INV_X1 U5476 ( .A(n4514), .ZN(n4513) );
  NAND2_X1 U5477 ( .A1(n9877), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9900) );
  AND2_X1 U5478 ( .A1(n4736), .A2(n4735), .ZN(n7172) );
  NAND2_X1 U5479 ( .A1(n7170), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4735) );
  NAND2_X1 U5480 ( .A1(n7414), .A2(n7382), .ZN(n7372) );
  INV_X1 U5481 ( .A(n4786), .ZN(n4784) );
  INV_X1 U5482 ( .A(n5560), .ZN(n4637) );
  OR2_X1 U5483 ( .A1(n7137), .A2(n7882), .ZN(n4667) );
  NAND2_X1 U5484 ( .A1(n4456), .A2(n4455), .ZN(n7089) );
  INV_X1 U5485 ( .A(n7445), .ZN(n4455) );
  OR2_X1 U5486 ( .A1(n5633), .A2(n5612), .ZN(n5784) );
  AND2_X1 U5487 ( .A1(n4712), .A2(n4964), .ZN(n4711) );
  INV_X1 U5488 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4959) );
  NOR2_X1 U5489 ( .A1(n4571), .A2(n4572), .ZN(n4570) );
  INV_X1 U5490 ( .A(n4565), .ZN(n6271) );
  AND2_X1 U5491 ( .A1(n9115), .A2(n9114), .ZN(n4539) );
  NOR2_X1 U5492 ( .A1(n9680), .A2(n9278), .ZN(n4536) );
  INV_X1 U5493 ( .A(n4832), .ZN(n4831) );
  OR2_X1 U5494 ( .A1(n9339), .A2(n8559), .ZN(n8989) );
  NAND2_X1 U5495 ( .A1(n9625), .A2(n9123), .ZN(n4825) );
  NOR2_X1 U5496 ( .A1(n9507), .A2(n9508), .ZN(n8956) );
  AND2_X1 U5497 ( .A1(n9055), .A2(n9556), .ZN(n8848) );
  NAND2_X1 U5498 ( .A1(n6397), .A2(n9042), .ZN(n8913) );
  AND2_X1 U5499 ( .A1(n9109), .A2(n9035), .ZN(n6197) );
  AND2_X1 U5500 ( .A1(n6583), .A2(n8932), .ZN(n6740) );
  AND2_X1 U5501 ( .A1(n6553), .A2(n6393), .ZN(n4866) );
  NOR2_X1 U5502 ( .A1(n6419), .A2(n6109), .ZN(n4868) );
  NAND2_X1 U5503 ( .A1(n4869), .A2(n9796), .ZN(n6415) );
  AND2_X1 U5504 ( .A1(n5467), .A2(n5451), .ZN(n5465) );
  AND2_X1 U5505 ( .A1(n5445), .A2(n5431), .ZN(n5443) );
  INV_X1 U5506 ( .A(n4900), .ZN(n4896) );
  NAND2_X1 U5507 ( .A1(n5223), .A2(SI_13_), .ZN(n5243) );
  XNOR2_X1 U5508 ( .A(n5206), .B(SI_11_), .ZN(n5207) );
  OAI21_X1 U5509 ( .B1(n4338), .B2(n4465), .A(n4464), .ZN(n5111) );
  NAND2_X1 U5510 ( .A1(n4337), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4464) );
  OAI21_X1 U5511 ( .B1(n4338), .B2(n4435), .A(n4434), .ZN(n5075) );
  NAND2_X1 U5512 ( .A1(n4338), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4434) );
  NAND2_X1 U5513 ( .A1(n4759), .A2(n5025), .ZN(n5026) );
  INV_X1 U5514 ( .A(n5024), .ZN(n4759) );
  INV_X1 U5515 ( .A(n4934), .ZN(n4930) );
  AND2_X1 U5516 ( .A1(n7783), .A2(n5718), .ZN(n7716) );
  OR2_X1 U5517 ( .A1(n6903), .A2(n6902), .ZN(n6993) );
  AND2_X1 U5518 ( .A1(n5706), .A2(n7877), .ZN(n7755) );
  AND2_X1 U5519 ( .A1(n7832), .A2(n5711), .ZN(n7762) );
  AND2_X1 U5520 ( .A1(n7745), .A2(n5735), .ZN(n7773) );
  NAND2_X1 U5521 ( .A1(n5398), .A2(n7809), .ZN(n5417) );
  XNOR2_X1 U5522 ( .A(n4336), .B(n9927), .ZN(n5671) );
  INV_X1 U5523 ( .A(n7831), .ZN(n4691) );
  INV_X1 U5524 ( .A(n7832), .ZN(n4692) );
  AOI21_X1 U5525 ( .B1(n4695), .B2(n4698), .A(n4694), .ZN(n4693) );
  INV_X1 U5526 ( .A(n7762), .ZN(n4694) );
  INV_X1 U5527 ( .A(n7887), .ZN(n5682) );
  AND2_X1 U5528 ( .A1(n7411), .A2(n7410), .ZN(n7468) );
  OR2_X1 U5529 ( .A1(n5784), .A2(n7185), .ZN(n6304) );
  OAI21_X1 U5530 ( .B1(n4737), .B2(n4395), .A(n6319), .ZN(n6562) );
  NAND2_X1 U5531 ( .A1(n9822), .A2(n9821), .ZN(n9820) );
  AND2_X1 U5532 ( .A1(n9837), .A2(n6322), .ZN(n6323) );
  NAND2_X1 U5533 ( .A1(n6345), .A2(n4509), .ZN(n6322) );
  INV_X1 U5534 ( .A(n6321), .ZN(n4509) );
  NAND2_X1 U5535 ( .A1(n6323), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9839) );
  AND2_X1 U5536 ( .A1(n4713), .A2(n4485), .ZN(n4484) );
  NAND2_X1 U5537 ( .A1(n4515), .A2(n6340), .ZN(n6636) );
  NAND2_X1 U5538 ( .A1(n9888), .A2(n4716), .ZN(n9914) );
  OR2_X1 U5539 ( .A1(n6646), .A2(n6647), .ZN(n4716) );
  NAND2_X1 U5540 ( .A1(n9914), .A2(n9915), .ZN(n9913) );
  XNOR2_X1 U5541 ( .A(n7000), .B(n4505), .ZN(n6650) );
  NAND2_X1 U5542 ( .A1(n9913), .A2(n4498), .ZN(n7000) );
  NAND2_X1 U5543 ( .A1(n4499), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4498) );
  XNOR2_X1 U5544 ( .A(n7172), .B(n7171), .ZN(n7209) );
  NOR2_X1 U5545 ( .A1(n7209), .A2(n5198), .ZN(n7208) );
  NOR2_X1 U5546 ( .A1(n7206), .A2(n7164), .ZN(n7167) );
  XNOR2_X1 U5547 ( .A(n7911), .B(n7927), .ZN(n7901) );
  NOR2_X1 U5548 ( .A1(n7899), .A2(n4715), .ZN(n7911) );
  NOR2_X1 U5549 ( .A1(n7177), .A2(n8281), .ZN(n4715) );
  NOR2_X1 U5550 ( .A1(n7928), .A2(n7929), .ZN(n7932) );
  OR2_X1 U5551 ( .A1(n7973), .A2(n7974), .ZN(n4508) );
  AND2_X1 U5552 ( .A1(n4508), .A2(n4507), .ZN(n7984) );
  INV_X1 U5553 ( .A(n7977), .ZN(n4507) );
  NAND2_X1 U5554 ( .A1(n4516), .A2(n4733), .ZN(n4732) );
  NAND2_X1 U5555 ( .A1(n7990), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4491) );
  OR2_X1 U5556 ( .A1(n8043), .A2(n8031), .ZN(n4477) );
  NAND2_X1 U5557 ( .A1(n4479), .A2(n8043), .ZN(n4478) );
  NAND2_X1 U5558 ( .A1(n8030), .A2(n8005), .ZN(n4479) );
  OR2_X1 U5559 ( .A1(n7243), .A2(n8083), .ZN(n5521) );
  INV_X1 U5560 ( .A(n7372), .ZN(n7462) );
  NOR2_X1 U5561 ( .A1(n8073), .A2(n8278), .ZN(n4632) );
  XNOR2_X1 U5562 ( .A(n7243), .B(n7869), .ZN(n8074) );
  OR2_X1 U5563 ( .A1(n5495), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5513) );
  AOI21_X1 U5564 ( .B1(n4781), .B2(n5573), .A(n4399), .ZN(n4779) );
  INV_X1 U5565 ( .A(n4781), .ZN(n4780) );
  INV_X1 U5566 ( .A(n5456), .ZN(n5455) );
  AOI21_X1 U5567 ( .B1(n4650), .B2(n5570), .A(n4649), .ZN(n4648) );
  INV_X1 U5568 ( .A(n7350), .ZN(n4785) );
  AOI21_X1 U5569 ( .B1(n4784), .B2(n7350), .A(n4783), .ZN(n4782) );
  INV_X1 U5570 ( .A(n7427), .ZN(n4783) );
  AND2_X1 U5571 ( .A1(n7428), .A2(n7427), .ZN(n8189) );
  NAND2_X1 U5572 ( .A1(n5335), .A2(n5334), .ZN(n5355) );
  INV_X1 U5573 ( .A(n5336), .ZN(n5335) );
  AND2_X1 U5574 ( .A1(n7342), .A2(n7344), .ZN(n8223) );
  OR2_X1 U5575 ( .A1(n8206), .A2(n8223), .ZN(n8226) );
  INV_X1 U5576 ( .A(n5256), .ZN(n5255) );
  AND2_X1 U5577 ( .A1(n7332), .A2(n7333), .ZN(n8251) );
  NAND2_X1 U5578 ( .A1(n4660), .A2(n4365), .ZN(n4659) );
  INV_X1 U5579 ( .A(n4656), .ZN(n4655) );
  OAI21_X1 U5580 ( .B1(n4658), .B2(n4657), .A(n5559), .ZN(n4656) );
  NAND2_X1 U5581 ( .A1(n5153), .A2(n5152), .ZN(n5185) );
  INV_X1 U5582 ( .A(n5154), .ZN(n5153) );
  NAND2_X1 U5583 ( .A1(n5122), .A2(n5121), .ZN(n5136) );
  INV_X1 U5584 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5121) );
  INV_X1 U5585 ( .A(n5123), .ZN(n5122) );
  INV_X1 U5586 ( .A(n7884), .ZN(n7085) );
  AND2_X2 U5587 ( .A1(n6920), .A2(n7303), .ZN(n7441) );
  NAND2_X1 U5588 ( .A1(n5108), .A2(n7290), .ZN(n6807) );
  OR2_X1 U5589 ( .A1(n5087), .A2(n5086), .ZN(n6667) );
  NAND2_X1 U5590 ( .A1(n5038), .A2(n5037), .ZN(n5066) );
  INV_X1 U5591 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5038) );
  INV_X1 U5592 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5037) );
  OAI21_X1 U5593 ( .B1(n6940), .B2(n5548), .A(n5547), .ZN(n6677) );
  AND4_X1 U5594 ( .A1(n5093), .A2(n5092), .A3(n5091), .A4(n5090), .ZN(n6811)
         );
  NAND2_X1 U5595 ( .A1(n6225), .A2(n6226), .ZN(n6945) );
  NAND2_X1 U5596 ( .A1(n5475), .A2(n5474), .ZN(n8300) );
  NAND2_X1 U5597 ( .A1(n5381), .A2(n5380), .ZN(n7724) );
  NAND2_X1 U5598 ( .A1(n5366), .A2(n5365), .ZN(n7781) );
  NOR2_X1 U5599 ( .A1(n5759), .A2(n8423), .ZN(n5754) );
  AND2_X1 U5600 ( .A1(n4967), .A2(n4788), .ZN(n4787) );
  NOR2_X1 U5601 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4788) );
  AND2_X1 U5602 ( .A1(n5175), .A2(n5174), .ZN(n5179) );
  NAND2_X1 U5603 ( .A1(n4719), .A2(n5031), .ZN(n4718) );
  INV_X1 U5604 ( .A(n6658), .ZN(n4837) );
  OR2_X1 U5605 ( .A1(n6270), .A2(n4564), .ZN(n4562) );
  INV_X1 U5606 ( .A(n6655), .ZN(n4839) );
  NAND2_X1 U5607 ( .A1(n4839), .A2(n6502), .ZN(n4557) );
  NAND2_X1 U5608 ( .A1(n4839), .A2(n6269), .ZN(n4560) );
  INV_X1 U5609 ( .A(n9117), .ZN(n8999) );
  OR2_X1 U5610 ( .A1(n6486), .A2(n6485), .ZN(n6517) );
  OAI21_X1 U5611 ( .B1(n4586), .B2(n4585), .A(n4844), .ZN(n4584) );
  OR2_X1 U5612 ( .A1(n6887), .A2(n10078), .ZN(n7538) );
  INV_X1 U5613 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6179) );
  AND2_X1 U5614 ( .A1(n8492), .A2(n8491), .ZN(n8716) );
  AOI21_X1 U5615 ( .B1(n8486), .B2(n4572), .A(n4571), .ZN(n4567) );
  NAND2_X1 U5616 ( .A1(n4569), .A2(n8486), .ZN(n4568) );
  INV_X1 U5617 ( .A(n4470), .ZN(n4569) );
  AND2_X1 U5618 ( .A1(n7566), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U5619 ( .A1(n7507), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7502) );
  NOR2_X1 U5620 ( .A1(n4938), .A2(n8735), .ZN(n4852) );
  INV_X1 U5621 ( .A(n4586), .ZN(n6973) );
  OR2_X1 U5622 ( .A1(n6517), .A2(n6516), .ZN(n6749) );
  NAND2_X1 U5623 ( .A1(n4553), .A2(n8745), .ZN(n8748) );
  OR2_X1 U5624 ( .A1(n7517), .A2(n8836), .ZN(n7519) );
  NAND2_X1 U5625 ( .A1(n4847), .A2(n4849), .ZN(n8677) );
  OR2_X1 U5626 ( .A1(n6973), .A2(n4850), .ZN(n4847) );
  NOR2_X1 U5627 ( .A1(n6180), .A2(n6179), .ZN(n6274) );
  NAND2_X1 U5628 ( .A1(n4576), .A2(n4857), .ZN(n8800) );
  NOR2_X1 U5629 ( .A1(n7564), .A2(n7563), .ZN(n7566) );
  AND3_X1 U5630 ( .A1(n7497), .A2(n7496), .A3(n7495), .ZN(n8508) );
  AND4_X1 U5631 ( .A1(n6753), .A2(n6752), .A3(n6751), .A4(n6750), .ZN(n8448)
         );
  OAI21_X1 U5632 ( .B1(n9743), .B2(n8836), .A(n8835), .ZN(n9587) );
  OR2_X1 U5633 ( .A1(n7658), .A2(n7657), .ZN(n9325) );
  AND2_X1 U5634 ( .A1(n8995), .A2(n8987), .ZN(n9347) );
  AOI21_X1 U5635 ( .B1(n4743), .B2(n4742), .A(n4741), .ZN(n4740) );
  INV_X1 U5636 ( .A(n8992), .ZN(n4741) );
  INV_X1 U5637 ( .A(n9381), .ZN(n4742) );
  INV_X1 U5638 ( .A(n9347), .ZN(n9350) );
  AND2_X1 U5639 ( .A1(n4818), .A2(n7617), .ZN(n4816) );
  NAND2_X1 U5640 ( .A1(n4814), .A2(n4387), .ZN(n4813) );
  NOR2_X1 U5641 ( .A1(n7589), .A2(n8753), .ZN(n7601) );
  AND2_X1 U5642 ( .A1(n9081), .A2(n8970), .ZN(n9429) );
  AND2_X1 U5643 ( .A1(n9080), .A2(n8976), .ZN(n9449) );
  NOR2_X1 U5644 ( .A1(n7571), .A2(n4809), .ZN(n4803) );
  AND2_X1 U5645 ( .A1(n9067), .A2(n9064), .ZN(n9523) );
  INV_X1 U5646 ( .A(n7674), .ZN(n9527) );
  NAND2_X1 U5647 ( .A1(n8932), .A2(n8930), .ZN(n4454) );
  NAND2_X1 U5648 ( .A1(n6739), .A2(n6747), .ZN(n6853) );
  NOR2_X2 U5649 ( .A1(n6482), .A2(n6579), .ZN(n6583) );
  NAND2_X1 U5650 ( .A1(n6387), .A2(n9796), .ZN(n4442) );
  INV_X1 U5651 ( .A(n4526), .ZN(n4525) );
  OAI22_X1 U5652 ( .A1(n8864), .A2(n4933), .B1(n9147), .B2(n4341), .ZN(n4526)
         );
  NAND2_X1 U5653 ( .A1(n8866), .A2(n8865), .ZN(n9264) );
  NAND2_X1 U5654 ( .A1(n7655), .A2(n7654), .ZN(n9323) );
  XNOR2_X1 U5655 ( .A(n7400), .B(n7399), .ZN(n8831) );
  OAI22_X1 U5656 ( .A1(n7395), .A2(n7394), .B1(SI_30_), .B2(n7393), .ZN(n7400)
         );
  XNOR2_X1 U5657 ( .A(n7395), .B(n7394), .ZN(n8862) );
  NOR2_X1 U5658 ( .A1(n4922), .A2(n4920), .ZN(n4918) );
  INV_X1 U5659 ( .A(n5525), .ZN(n4920) );
  XNOR2_X1 U5660 ( .A(n7375), .B(SI_29_), .ZN(n4922) );
  NOR2_X1 U5661 ( .A1(n4865), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n4542) );
  XNOR2_X1 U5662 ( .A(n5485), .B(n5484), .ZN(n7652) );
  INV_X1 U5663 ( .A(n5813), .ZN(n5808) );
  NAND2_X1 U5664 ( .A1(n4903), .A2(n4904), .ZN(n5344) );
  OAI21_X1 U5665 ( .B1(n5301), .B2(n5300), .A(n5303), .ZN(n5325) );
  NAND2_X1 U5666 ( .A1(n5191), .A2(n5168), .ZN(n5171) );
  NOR2_X1 U5667 ( .A1(n5161), .A2(SI_9_), .ZN(n5162) );
  AND4_X1 U5668 ( .A1(n5275), .A2(n5274), .A3(n5273), .A4(n5272), .ZN(n8248)
         );
  INV_X1 U5669 ( .A(n4680), .ZN(n4679) );
  NAND2_X1 U5670 ( .A1(n7772), .A2(n5732), .ZN(n7709) );
  NAND2_X1 U5671 ( .A1(n5002), .A2(n4385), .ZN(n4671) );
  AND2_X1 U5672 ( .A1(n5667), .A2(n6929), .ZN(n6374) );
  AND3_X1 U5673 ( .A1(n5372), .A2(n5371), .A3(n5370), .ZN(n8185) );
  NOR2_X1 U5674 ( .A1(n7860), .A2(n4698), .ZN(n7764) );
  INV_X1 U5675 ( .A(n8212), .ZN(n8184) );
  NAND2_X1 U5676 ( .A1(n7026), .A2(n7025), .ZN(n7024) );
  OR2_X1 U5677 ( .A1(n5778), .A2(n5773), .ZN(n7810) );
  AOI21_X1 U5678 ( .B1(n4703), .B2(n4706), .A(n4352), .ZN(n4701) );
  NAND2_X1 U5679 ( .A1(n6371), .A2(n5670), .ZN(n6252) );
  NAND2_X1 U5680 ( .A1(n6728), .A2(n6727), .ZN(n6726) );
  OR2_X1 U5681 ( .A1(n5778), .A2(n5777), .ZN(n7855) );
  NOR2_X1 U5682 ( .A1(n7862), .A2(n7863), .ZN(n7860) );
  NAND2_X1 U5683 ( .A1(n4611), .A2(n5583), .ZN(n4605) );
  OR2_X1 U5684 ( .A1(n4611), .A2(n5583), .ZN(n4608) );
  XNOR2_X1 U5685 ( .A(n4954), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7472) );
  INV_X1 U5686 ( .A(n7468), .ZN(n8057) );
  INV_X1 U5687 ( .A(n8083), .ZN(n7869) );
  OR2_X1 U5688 ( .A1(n6304), .A2(P2_U3151), .ZN(n7871) );
  INV_X1 U5689 ( .A(n6811), .ZN(n7886) );
  OAI211_X1 U5690 ( .C1(n4339), .C2(n10067), .A(n5009), .B(n5008), .ZN(n4778)
         );
  AOI21_X1 U5691 ( .B1(n6573), .B2(n6315), .A(n6316), .ZN(n6571) );
  NAND2_X1 U5692 ( .A1(n9851), .A2(n9852), .ZN(n9850) );
  OAI21_X1 U5693 ( .B1(n6347), .B2(n5021), .A(n4714), .ZN(n9851) );
  INV_X1 U5694 ( .A(n4717), .ZN(n9890) );
  NAND2_X1 U5695 ( .A1(n4501), .A2(n4502), .ZN(n9903) );
  NOR2_X1 U5696 ( .A1(n6999), .A2(n4453), .ZN(n7003) );
  AND2_X1 U5697 ( .A1(n7000), .A2(n4505), .ZN(n4453) );
  INV_X1 U5698 ( .A(n4736), .ZN(n7169) );
  XNOR2_X1 U5699 ( .A(n7926), .B(n7927), .ZN(n7893) );
  NOR2_X1 U5700 ( .A1(n7893), .A2(n8355), .ZN(n7928) );
  XNOR2_X1 U5701 ( .A(n7971), .B(n7972), .ZN(n7939) );
  NOR2_X1 U5702 ( .A1(n7939), .A2(n10065), .ZN(n7973) );
  INV_X1 U5703 ( .A(n4452), .ZN(n7957) );
  NOR2_X1 U5704 ( .A1(n7999), .A2(n4724), .ZN(n4723) );
  AND2_X1 U5705 ( .A1(n9897), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n4724) );
  AND2_X1 U5706 ( .A1(n7989), .A2(n7988), .ZN(n4726) );
  OR2_X1 U5707 ( .A1(n8043), .A2(n8005), .ZN(n4480) );
  XNOR2_X1 U5708 ( .A(n7413), .B(n7462), .ZN(n8069) );
  NAND2_X1 U5709 ( .A1(n8104), .A2(n5578), .ZN(n8094) );
  NAND2_X1 U5710 ( .A1(n8117), .A2(n5577), .ZN(n8106) );
  NAND2_X1 U5711 ( .A1(n8142), .A2(n4781), .ZN(n8126) );
  NAND2_X1 U5712 ( .A1(n8148), .A2(n5575), .ZN(n8132) );
  NAND2_X1 U5713 ( .A1(n8142), .A2(n7249), .ZN(n8136) );
  NAND2_X1 U5714 ( .A1(n5397), .A2(n5396), .ZN(n8316) );
  NAND2_X1 U5715 ( .A1(n4651), .A2(n5569), .ZN(n5571) );
  AND2_X1 U5716 ( .A1(n5322), .A2(n7257), .ZN(n8199) );
  NAND2_X1 U5717 ( .A1(n4641), .A2(n5561), .ZN(n8237) );
  NAND2_X1 U5718 ( .A1(n5269), .A2(n5268), .ZN(n8346) );
  NAND2_X1 U5719 ( .A1(n5232), .A2(n5231), .ZN(n8260) );
  NAND2_X1 U5720 ( .A1(n8271), .A2(n7322), .ZN(n8262) );
  NAND2_X1 U5721 ( .A1(n4654), .A2(n4660), .ZN(n8273) );
  NAND2_X1 U5722 ( .A1(n7130), .A2(n4662), .ZN(n4654) );
  NAND2_X1 U5723 ( .A1(n4664), .A2(n4662), .ZN(n7144) );
  INV_X1 U5724 ( .A(n6667), .ZN(n9937) );
  OR2_X1 U5725 ( .A1(n6682), .A2(n8255), .ZN(n8230) );
  INV_X1 U5726 ( .A(n8230), .ZN(n8284) );
  INV_X1 U5727 ( .A(n7467), .ZN(n8367) );
  AND2_X1 U5728 ( .A1(n5494), .A2(n5493), .ZN(n8377) );
  AND2_X1 U5729 ( .A1(n8297), .A2(n8296), .ZN(n8374) );
  INV_X1 U5730 ( .A(n5727), .ZN(n8390) );
  NAND2_X1 U5731 ( .A1(n5290), .A2(n5289), .ZN(n8411) );
  INV_X1 U5732 ( .A(n6768), .ZN(n6802) );
  NAND2_X1 U5733 ( .A1(n4448), .A2(n4384), .ZN(n4589) );
  NAND2_X1 U5734 ( .A1(n6071), .A2(n6070), .ZN(n6093) );
  NAND2_X1 U5735 ( .A1(n4971), .A2(n4972), .ZN(n8426) );
  AND2_X1 U5736 ( .A1(n5604), .A2(n5603), .ZN(n7241) );
  NAND2_X1 U5737 ( .A1(n5607), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5598) );
  INV_X1 U5738 ( .A(n7472), .ZN(n7152) );
  AND2_X1 U5739 ( .A1(n5798), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6000) );
  AND2_X1 U5740 ( .A1(n7484), .A2(n7665), .ZN(n9309) );
  NAND2_X1 U5741 ( .A1(n8589), .A2(n4574), .ZN(n4573) );
  NAND2_X1 U5742 ( .A1(n8589), .A2(n4857), .ZN(n4575) );
  INV_X1 U5743 ( .A(n4577), .ZN(n4574) );
  AND2_X1 U5744 ( .A1(n8582), .A2(n8581), .ZN(n8658) );
  NAND2_X1 U5745 ( .A1(n7481), .A2(n7480), .ZN(n9269) );
  OR2_X1 U5746 ( .A1(n7656), .A2(n7645), .ZN(n9340) );
  AND2_X1 U5747 ( .A1(n6177), .A2(n6161), .ZN(n4853) );
  NAND2_X1 U5748 ( .A1(n4854), .A2(n6161), .ZN(n6175) );
  AND2_X1 U5749 ( .A1(n4848), .A2(n4852), .ZN(n8737) );
  OR2_X1 U5750 ( .A1(n6973), .A2(n4360), .ZN(n4848) );
  NAND2_X1 U5751 ( .A1(n4843), .A2(n8606), .ZN(n8768) );
  NAND2_X1 U5752 ( .A1(n6503), .A2(n6502), .ZN(n4838) );
  AND2_X1 U5753 ( .A1(n6003), .A2(n9037), .ZN(n8810) );
  AND2_X1 U5754 ( .A1(n4470), .A2(n8486), .ZN(n8815) );
  INV_X1 U5755 ( .A(n8786), .ZN(n8816) );
  NAND2_X1 U5756 ( .A1(n9026), .A2(n9035), .ZN(n4532) );
  NAND2_X1 U5757 ( .A1(n4534), .A2(n4350), .ZN(n4533) );
  AND4_X1 U5758 ( .A1(n6219), .A2(n6218), .A3(n6217), .A4(n6216), .ZN(n8837)
         );
  NAND4_X2 U5759 ( .A1(n5871), .A2(n5870), .A3(n5869), .A4(n5868), .ZN(n6385)
         );
  NAND2_X1 U5760 ( .A1(n4836), .A2(n4835), .ZN(n9320) );
  AND2_X1 U5761 ( .A1(n9380), .A2(n8879), .ZN(n9366) );
  NAND2_X1 U5762 ( .A1(n4812), .A2(n4817), .ZN(n9379) );
  NAND2_X1 U5763 ( .A1(n4811), .A2(n4818), .ZN(n4812) );
  NAND2_X1 U5764 ( .A1(n4811), .A2(n4819), .ZN(n9394) );
  NAND2_X1 U5765 ( .A1(n7584), .A2(n7583), .ZN(n4823) );
  NAND2_X1 U5766 ( .A1(n9496), .A2(n8965), .ZN(n9481) );
  INV_X1 U5767 ( .A(n9649), .ZN(n9495) );
  NOR2_X1 U5768 ( .A1(n4755), .A2(n4754), .ZN(n9497) );
  INV_X1 U5769 ( .A(n9068), .ZN(n4754) );
  NAND2_X1 U5770 ( .A1(n4804), .A2(n4808), .ZN(n9489) );
  NAND2_X1 U5771 ( .A1(n9520), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U5772 ( .A1(n9520), .A2(n4810), .ZN(n9506) );
  OAI21_X1 U5773 ( .B1(n7526), .B2(n4800), .A(n4344), .ZN(n9541) );
  NAND2_X1 U5774 ( .A1(n9555), .A2(n9558), .ZN(n9554) );
  NAND2_X1 U5775 ( .A1(n7526), .A2(n7525), .ZN(n9555) );
  NAND2_X1 U5776 ( .A1(n4544), .A2(n4358), .ZN(n4543) );
  INV_X1 U5777 ( .A(n8839), .ZN(n4545) );
  INV_X1 U5778 ( .A(n9551), .ZN(n9799) );
  NAND2_X1 U5779 ( .A1(n7688), .A2(n8861), .ZN(n7483) );
  INV_X1 U5780 ( .A(n6596), .ZN(n6475) );
  INV_X1 U5781 ( .A(n6553), .ZN(n6430) );
  INV_X1 U5782 ( .A(n9264), .ZN(n9684) );
  INV_X1 U5783 ( .A(n9585), .ZN(n4449) );
  INV_X1 U5784 ( .A(n9269), .ZN(n9295) );
  INV_X1 U5785 ( .A(n9323), .ZN(n9693) );
  INV_X1 U5786 ( .A(n9339), .ZN(n9697) );
  INV_X1 U5787 ( .A(n9358), .ZN(n9701) );
  INV_X1 U5788 ( .A(n9404), .ZN(n9712) );
  CLKBUF_X1 U5789 ( .A(n9733), .Z(n4451) );
  OR2_X1 U5790 ( .A1(n6871), .A2(n8836), .ZN(n6874) );
  INV_X1 U5791 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5859) );
  CLKBUF_X1 U5792 ( .A(n5886), .Z(n9257) );
  NAND2_X1 U5793 ( .A1(n5391), .A2(n4915), .ZN(n4909) );
  NAND2_X1 U5794 ( .A1(n4899), .A2(n4898), .ZN(n5222) );
  NAND2_X1 U5795 ( .A1(n4899), .A2(n4372), .ZN(n5211) );
  AND2_X1 U5796 ( .A1(n6089), .A2(n6014), .ZN(n7534) );
  NAND2_X1 U5797 ( .A1(n4441), .A2(n4440), .ZN(n5052) );
  INV_X1 U5798 ( .A(n5050), .ZN(n4440) );
  INV_X1 U5799 ( .A(n5051), .ZN(n4441) );
  NAND2_X1 U5800 ( .A1(n5014), .A2(n4878), .ZN(n5017) );
  INV_X1 U5801 ( .A(n5015), .ZN(n4878) );
  NAND2_X1 U5802 ( .A1(n4686), .A2(n7845), .ZN(n4683) );
  NAND2_X1 U5803 ( .A1(n6286), .A2(n5675), .ZN(n6445) );
  INV_X1 U5804 ( .A(n4496), .ZN(n7916) );
  INV_X1 U5805 ( .A(n4494), .ZN(n7961) );
  NAND2_X1 U5806 ( .A1(n4725), .A2(n4721), .ZN(P2_U3199) );
  INV_X1 U5807 ( .A(n4722), .ZN(n4721) );
  OAI21_X1 U5808 ( .B1(n8003), .B2(n4726), .A(n9916), .ZN(n4725) );
  OAI21_X1 U5809 ( .B1(n8001), .B2(n8000), .A(n4723), .ZN(n4722) );
  OAI21_X1 U5810 ( .B1(n8006), .B2(n4480), .A(n4475), .ZN(n4481) );
  AOI21_X1 U5811 ( .B1(n8065), .B2(n5656), .A(n5655), .ZN(n5657) );
  AOI21_X1 U5812 ( .B1(n8065), .B2(n5643), .A(n5642), .ZN(n5644) );
  NAND2_X1 U5813 ( .A1(n4627), .A2(n4625), .ZN(P2_U3455) );
  AOI21_X1 U5814 ( .B1(n7243), .B2(n5643), .A(n4626), .ZN(n4625) );
  NOR2_X1 U5815 ( .A1(n9965), .A2(n8372), .ZN(n4626) );
  NAND2_X1 U5816 ( .A1(n4468), .A2(n4466), .ZN(P1_U3229) );
  NOR2_X1 U5817 ( .A1(n8732), .A2(n4467), .ZN(n4466) );
  AND2_X1 U5818 ( .A1(n9358), .A2(n8784), .ZN(n4467) );
  AOI21_X1 U5819 ( .B1(n8875), .B2(n9676), .A(n4461), .ZN(n4460) );
  NOR2_X1 U5820 ( .A1(n9816), .A2(n9579), .ZN(n4461) );
  AOI21_X1 U5821 ( .B1(n8875), .B2(n9732), .A(n4463), .ZN(n4462) );
  NOR2_X1 U5822 ( .A1(n9725), .A2(n9679), .ZN(n4463) );
  AND2_X1 U5823 ( .A1(n8858), .A2(n4345), .ZN(n4342) );
  AND2_X1 U5824 ( .A1(n4792), .A2(n7316), .ZN(n4343) );
  AND2_X1 U5825 ( .A1(n4798), .A2(n7532), .ZN(n4344) );
  AOI21_X1 U5826 ( .B1(n8831), .B2(n8861), .A(n8830), .ZN(n9680) );
  INV_X2 U5827 ( .A(n6166), .ZN(n8640) );
  AND2_X1 U5828 ( .A1(n4945), .A2(n4377), .ZN(n5131) );
  INV_X1 U5829 ( .A(n8272), .ZN(n4792) );
  OR2_X1 U5830 ( .A1(n9693), .A2(n8999), .ZN(n4345) );
  CLKBUF_X1 U5831 ( .A(n6108), .Z(n6109) );
  NOR2_X1 U5832 ( .A1(n5749), .A2(n4418), .ZN(n4346) );
  AND2_X1 U5833 ( .A1(n4695), .A2(n7832), .ZN(n4347) );
  AND2_X1 U5834 ( .A1(n9957), .A2(n7881), .ZN(n4348) );
  AND4_X1 U5835 ( .A1(n6522), .A2(n6521), .A3(n6520), .A4(n6519), .ZN(n6974)
         );
  INV_X1 U5836 ( .A(n6974), .ZN(n4758) );
  AND2_X1 U5837 ( .A1(n8916), .A2(n8918), .ZN(n4349) );
  NOR2_X1 U5838 ( .A1(n9024), .A2(n9035), .ZN(n4350) );
  AND2_X1 U5839 ( .A1(n8921), .A2(n4394), .ZN(n4351) );
  AND2_X1 U5840 ( .A1(n4709), .A2(n7880), .ZN(n4352) );
  NAND2_X1 U5841 ( .A1(n5807), .A2(n5811), .ZN(n4865) );
  INV_X1 U5842 ( .A(n9387), .ZN(n4872) );
  AND2_X1 U5843 ( .A1(n4904), .A2(n5343), .ZN(n4353) );
  OR2_X1 U5844 ( .A1(n8010), .A2(n8035), .ZN(n4354) );
  AND2_X1 U5845 ( .A1(n5679), .A2(n5675), .ZN(n4355) );
  NAND2_X1 U5846 ( .A1(n4471), .A2(n4719), .ZN(n4356) );
  OR2_X1 U5847 ( .A1(n8367), .A2(n8057), .ZN(n4357) );
  NAND2_X1 U5848 ( .A1(n5483), .A2(n5482), .ZN(n7870) );
  INV_X1 U5849 ( .A(n7870), .ZN(n8109) );
  AND2_X1 U5850 ( .A1(n5511), .A2(n5510), .ZN(n8373) );
  INV_X1 U5851 ( .A(n8373), .ZN(n7243) );
  NAND2_X1 U5852 ( .A1(n7519), .A2(n7518), .ZN(n8757) );
  INV_X1 U5853 ( .A(n8757), .ZN(n4870) );
  INV_X1 U5854 ( .A(n6649), .ZN(n4499) );
  INV_X1 U5855 ( .A(n9858), .ZN(n4485) );
  OR2_X1 U5856 ( .A1(n9142), .A2(n9045), .ZN(n4358) );
  AND2_X1 U5857 ( .A1(n7260), .A2(n7261), .ZN(n4359) );
  AND2_X1 U5858 ( .A1(n8451), .A2(n8452), .ZN(n4360) );
  AND2_X1 U5859 ( .A1(n4841), .A2(n8606), .ZN(n4361) );
  AND2_X1 U5860 ( .A1(n4679), .A2(n7772), .ZN(n4362) );
  OR2_X1 U5861 ( .A1(n9432), .A2(n9124), .ZN(n4363) );
  NAND2_X1 U5862 ( .A1(n5287), .A2(n4711), .ZN(n4364) );
  NAND2_X1 U5863 ( .A1(n9963), .A2(n7880), .ZN(n4365) );
  AND2_X1 U5864 ( .A1(n8112), .A2(n5577), .ZN(n4366) );
  NAND2_X1 U5865 ( .A1(n8481), .A2(n8480), .ZN(n4469) );
  OAI21_X1 U5866 ( .B1(n4698), .B2(n4697), .A(n5708), .ZN(n4696) );
  OR2_X1 U5867 ( .A1(n5242), .A2(n4791), .ZN(n4367) );
  AND2_X1 U5868 ( .A1(n8980), .A2(n8979), .ZN(n4368) );
  NAND2_X1 U5869 ( .A1(n8469), .A2(n8683), .ZN(n4369) );
  AND2_X1 U5870 ( .A1(n4834), .A2(n4342), .ZN(n4370) );
  NAND2_X1 U5871 ( .A1(n4945), .A2(n4944), .ZN(n5104) );
  OR2_X1 U5872 ( .A1(n7972), .A2(n7956), .ZN(n4371) );
  OR2_X1 U5873 ( .A1(n5206), .A2(SI_11_), .ZN(n4372) );
  INV_X1 U5874 ( .A(n8965), .ZN(n4753) );
  AND4_X1 U5875 ( .A1(n8933), .A2(n8927), .A3(n8926), .A4(n9030), .ZN(n4373)
         );
  INV_X1 U5876 ( .A(n7290), .ZN(n4766) );
  INV_X1 U5877 ( .A(n6502), .ZN(n4564) );
  INV_X1 U5878 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5839) );
  OR2_X1 U5879 ( .A1(n7362), .A2(n7388), .ZN(n4374) );
  AND4_X1 U5880 ( .A1(n6491), .A2(n6490), .A3(n6489), .A4(n6488), .ZN(n8930)
         );
  AND2_X1 U5881 ( .A1(n7360), .A2(n7388), .ZN(n4375) );
  OR3_X1 U5882 ( .A1(n7466), .A2(n7465), .A3(n7464), .ZN(n4376) );
  NAND2_X1 U5883 ( .A1(n5287), .A2(n4951), .ZN(n4958) );
  AND2_X1 U5884 ( .A1(n4944), .A2(n4776), .ZN(n4377) );
  INV_X1 U5885 ( .A(n5573), .ZN(n8146) );
  NOR2_X1 U5886 ( .A1(n7357), .A2(n7356), .ZN(n4378) );
  AND2_X1 U5887 ( .A1(n9404), .A2(n9122), .ZN(n4379) );
  NOR2_X1 U5888 ( .A1(n8864), .A2(n6130), .ZN(n4380) );
  NOR2_X1 U5889 ( .A1(n8941), .A2(n8940), .ZN(n4381) );
  NOR2_X1 U5890 ( .A1(n9899), .A2(n6622), .ZN(n4382) );
  NOR2_X1 U5891 ( .A1(n9099), .A2(n4539), .ZN(n4383) );
  AND2_X1 U5892 ( .A1(n6129), .A2(n6050), .ZN(n4384) );
  INV_X1 U5893 ( .A(n8010), .ZN(n4733) );
  INV_X1 U5894 ( .A(n4457), .ZN(n4985) );
  OAI211_X1 U5895 ( .C1(n5012), .C2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n4458), .ZN(n4457) );
  INV_X1 U5896 ( .A(n4873), .ZN(n9403) );
  AND2_X1 U5897 ( .A1(n4672), .A2(n6050), .ZN(n4385) );
  AND2_X1 U5898 ( .A1(n7384), .A2(n4591), .ZN(n4386) );
  INV_X1 U5899 ( .A(n5558), .ZN(n4665) );
  NOR2_X1 U5900 ( .A1(n5324), .A2(n4907), .ZN(n4906) );
  OR2_X1 U5901 ( .A1(n7754), .A2(n7755), .ZN(n4698) );
  NAND2_X1 U5902 ( .A1(n9387), .A2(n9121), .ZN(n4387) );
  AND2_X1 U5903 ( .A1(n6749), .A2(n6748), .ZN(n4388) );
  AND2_X1 U5904 ( .A1(n5243), .A2(n4929), .ZN(n4389) );
  OR2_X1 U5905 ( .A1(n9446), .A2(n8508), .ZN(n4390) );
  INV_X1 U5906 ( .A(n4809), .ZN(n4808) );
  INV_X1 U5907 ( .A(n4857), .ZN(n4580) );
  AND2_X1 U5908 ( .A1(n8698), .A2(n4858), .ZN(n4857) );
  INV_X1 U5909 ( .A(n4677), .ZN(n7804) );
  NAND2_X1 U5910 ( .A1(n7725), .A2(n5724), .ZN(n4677) );
  AND2_X1 U5911 ( .A1(n4506), .A2(n4505), .ZN(n4391) );
  AND4_X1 U5912 ( .A1(n6279), .A2(n6278), .A3(n6277), .A4(n6276), .ZN(n6508)
         );
  NOR2_X1 U5913 ( .A1(n8346), .A2(n7877), .ZN(n4392) );
  NOR2_X1 U5914 ( .A1(n5727), .A2(n8150), .ZN(n4393) );
  NAND2_X1 U5915 ( .A1(n9053), .A2(n9049), .ZN(n4394) );
  AND2_X1 U5916 ( .A1(n6318), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4395) );
  OR2_X1 U5917 ( .A1(n6649), .A2(n9972), .ZN(n4396) );
  OR2_X1 U5918 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n4397) );
  NOR2_X1 U5919 ( .A1(n9593), .A2(n9116), .ZN(n4398) );
  NAND2_X1 U5920 ( .A1(n7361), .A2(n8125), .ZN(n4399) );
  NAND2_X1 U5921 ( .A1(n7500), .A2(n7499), .ZN(n9466) );
  INV_X1 U5922 ( .A(n9466), .ZN(n4875) );
  AND2_X1 U5923 ( .A1(n5033), .A2(n5054), .ZN(n6345) );
  INV_X1 U5924 ( .A(n4942), .ZN(n4807) );
  OR2_X1 U5925 ( .A1(n8836), .A2(n6051), .ZN(n4400) );
  INV_X1 U5926 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4861) );
  INV_X1 U5927 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4951) );
  AND2_X1 U5928 ( .A1(n4373), .A2(n4518), .ZN(n4401) );
  OR2_X1 U5929 ( .A1(n5338), .A2(n4997), .ZN(n4402) );
  OR2_X1 U5930 ( .A1(n8300), .A2(n7870), .ZN(n4403) );
  OAI21_X1 U5931 ( .B1(n4693), .B2(n4692), .A(n4691), .ZN(n4690) );
  INV_X1 U5932 ( .A(n8858), .ZN(n9302) );
  OR2_X1 U5933 ( .A1(n8081), .A2(n7366), .ZN(n4404) );
  AND2_X1 U5934 ( .A1(n5144), .A2(n5143), .ZN(n4405) );
  NAND2_X1 U5935 ( .A1(n4561), .A2(n4839), .ZN(n4406) );
  NAND2_X1 U5936 ( .A1(n7224), .A2(n7882), .ZN(n4407) );
  INV_X1 U5937 ( .A(n4696), .ZN(n4695) );
  AND2_X1 U5938 ( .A1(n4823), .A2(n4363), .ZN(n4408) );
  OR2_X1 U5939 ( .A1(n8065), .A2(n8073), .ZN(n7414) );
  INV_X1 U5940 ( .A(n7414), .ZN(n4773) );
  AND2_X1 U5941 ( .A1(n8916), .A2(n8922), .ZN(n4409) );
  AND2_X1 U5942 ( .A1(n7276), .A2(n4768), .ZN(n4410) );
  NAND2_X1 U5943 ( .A1(n8875), .A2(n9260), .ZN(n4411) );
  INV_X1 U5944 ( .A(n7651), .ZN(n4829) );
  AND2_X1 U5945 ( .A1(n4745), .A2(n9588), .ZN(n4412) );
  AND2_X1 U5946 ( .A1(n8390), .A2(n8150), .ZN(n7425) );
  AND2_X1 U5947 ( .A1(n4825), .A2(n7583), .ZN(n4413) );
  AND2_X1 U5948 ( .A1(n4711), .A2(n4962), .ZN(n4414) );
  AND2_X1 U5949 ( .A1(n4502), .A2(n4396), .ZN(n4415) );
  OR2_X1 U5950 ( .A1(n4803), .A2(n4942), .ZN(n4416) );
  INV_X1 U5951 ( .A(n9456), .ZN(n9459) );
  AND2_X1 U5952 ( .A1(n8912), .A2(n8975), .ZN(n9456) );
  AND2_X1 U5953 ( .A1(n7426), .A2(n5569), .ZN(n4650) );
  INV_X1 U5954 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4964) );
  INV_X1 U5955 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4719) );
  NAND2_X1 U5956 ( .A1(n4732), .A2(n4731), .ZN(n4417) );
  INV_X1 U5957 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4933) );
  INV_X1 U5958 ( .A(n7007), .ZN(n4505) );
  NAND2_X1 U5959 ( .A1(n7024), .A2(n5694), .ZN(n7222) );
  NAND2_X1 U5960 ( .A1(n4568), .A2(n4567), .ZN(n8704) );
  INV_X1 U5961 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4435) );
  AND2_X1 U5962 ( .A1(n5747), .A2(n8095), .ZN(n4418) );
  OAI21_X1 U5963 ( .B1(n9743), .B2(n5528), .A(n5527), .ZN(n8065) );
  OR2_X1 U5964 ( .A1(n9693), .A2(n8828), .ZN(n4419) );
  INV_X1 U5965 ( .A(n7880), .ZN(n8258) );
  NAND2_X1 U5966 ( .A1(n5131), .A2(n4950), .ZN(n5284) );
  NAND2_X1 U5967 ( .A1(n5792), .A2(n5793), .ZN(n6149) );
  OR2_X1 U5968 ( .A1(n6644), .A2(n6765), .ZN(n4420) );
  AND2_X1 U5969 ( .A1(n5501), .A2(n5500), .ZN(n8072) );
  INV_X1 U5970 ( .A(n8072), .ZN(n8095) );
  INV_X1 U5971 ( .A(n4662), .ZN(n4661) );
  NOR2_X1 U5972 ( .A1(n7141), .A2(n4663), .ZN(n4662) );
  AND2_X1 U5973 ( .A1(n5205), .A2(n7316), .ZN(n4421) );
  AND4_X1 U5974 ( .A1(n7544), .A2(n7543), .A3(n7542), .A4(n7541), .ZN(n8762)
         );
  AND4_X1 U5975 ( .A1(n6892), .A2(n6891), .A3(n6890), .A4(n6889), .ZN(n8689)
         );
  AND4_X1 U5976 ( .A1(n6845), .A2(n6844), .A3(n6843), .A4(n6842), .ZN(n8461)
         );
  INV_X1 U5977 ( .A(n4876), .ZN(n9476) );
  AND4_X1 U5978 ( .A1(n7524), .A2(n7523), .A3(n7522), .A4(n7521), .ZN(n8690)
         );
  AND2_X1 U5979 ( .A1(n4641), .A2(n4639), .ZN(n4422) );
  AND2_X1 U5980 ( .A1(n8558), .A2(n8556), .ZN(n8727) );
  INV_X1 U5981 ( .A(n8727), .ZN(n4859) );
  AND2_X1 U5982 ( .A1(n8486), .A2(n8814), .ZN(n4423) );
  AOI21_X1 U5983 ( .B1(n4915), .B2(n5390), .A(n4914), .ZN(n4913) );
  INV_X1 U5984 ( .A(n9573), .ZN(n6473) );
  INV_X1 U5985 ( .A(n9643), .ZN(n9676) );
  NAND2_X1 U5986 ( .A1(n5753), .A2(n5752), .ZN(n7845) );
  XNOR2_X1 U5987 ( .A(n5598), .B(P2_IR_REG_25__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U5988 ( .A1(n6807), .A2(n7441), .ZN(n6806) );
  INV_X2 U5989 ( .A(n9811), .ZN(n9725) );
  XOR2_X1 U5990 ( .A(n5690), .B(n7884), .Z(n4424) );
  AND2_X1 U5991 ( .A1(n6483), .A2(n9053), .ZN(n6878) );
  NAND2_X1 U5992 ( .A1(n6504), .A2(n4838), .ZN(n6656) );
  OR2_X1 U5993 ( .A1(n4558), .A2(n4563), .ZN(n4425) );
  AND2_X1 U5994 ( .A1(n7943), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4426) );
  AND2_X1 U5995 ( .A1(n7943), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4427) );
  NAND2_X1 U5996 ( .A1(n8924), .A2(n8923), .ZN(n4428) );
  NAND2_X1 U5997 ( .A1(n5601), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5634) );
  INV_X1 U5998 ( .A(n9933), .ZN(n9959) );
  INV_X1 U5999 ( .A(n7266), .ZN(n7417) );
  XNOR2_X1 U6000 ( .A(n5535), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7266) );
  AND2_X1 U6001 ( .A1(n7990), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4429) );
  AND2_X1 U6002 ( .A1(n8043), .A2(n8030), .ZN(n4430) );
  INV_X1 U6003 ( .A(n4867), .ZN(n6423) );
  NAND2_X1 U6004 ( .A1(n4868), .A2(n4869), .ZN(n4867) );
  AND2_X1 U6005 ( .A1(n4727), .A2(n6341), .ZN(n4431) );
  OR2_X1 U6006 ( .A1(n4731), .A2(n8035), .ZN(n4432) );
  AND2_X1 U6007 ( .A1(n4478), .A2(n4477), .ZN(n4433) );
  NAND2_X1 U6008 ( .A1(n9045), .A2(n6393), .ZN(n6435) );
  INV_X1 U6009 ( .A(n6435), .ZN(n4869) );
  XNOR2_X1 U6010 ( .A(n4961), .B(n4960), .ZN(n8046) );
  INV_X1 U6011 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4437) );
  INV_X1 U6012 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4465) );
  OAI21_X2 U6013 ( .B1(n9509), .B2(n4753), .A(n4752), .ZN(n9480) );
  AOI21_X2 U6014 ( .B1(n9303), .B2(n9302), .A(n7678), .ZN(n9276) );
  NAND2_X1 U6015 ( .A1(n5045), .A2(n5044), .ZN(n5051) );
  NAND2_X1 U6016 ( .A1(n9543), .A2(n9542), .ZN(n9525) );
  OAI21_X1 U6017 ( .B1(n9382), .B2(n4744), .A(n4740), .ZN(n9349) );
  OAI21_X1 U6018 ( .B1(n6876), .B2(n6881), .A(n8942), .ZN(n6882) );
  NAND2_X1 U6019 ( .A1(n9448), .A2(n9449), .ZN(n9447) );
  NAND2_X1 U6020 ( .A1(n7671), .A2(n8948), .ZN(n9543) );
  NAND2_X1 U6021 ( .A1(n4930), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4439) );
  NAND2_X1 U6022 ( .A1(n4449), .A2(n4412), .ZN(n9685) );
  NAND2_X1 U6023 ( .A1(n5080), .A2(n5079), .ZN(n4877) );
  XNOR2_X1 U6024 ( .A(n4750), .B(n9277), .ZN(n4749) );
  NAND2_X1 U6025 ( .A1(n5010), .A2(n4982), .ZN(n4986) );
  AOI21_X2 U6026 ( .B1(n9424), .B2(n9429), .A(n9089), .ZN(n9412) );
  NAND2_X1 U6027 ( .A1(n5074), .A2(n5073), .ZN(n5080) );
  OR2_X1 U6028 ( .A1(n6427), .A2(n6398), .ZN(n6399) );
  OAI211_X1 U6029 ( .C1(n4935), .C2(n4933), .A(n4439), .B(n4931), .ZN(n4979)
         );
  NAND2_X2 U6030 ( .A1(n4438), .A2(n6738), .ZN(n8935) );
  NAND2_X1 U6031 ( .A1(n5011), .A2(n5010), .ZN(n5015) );
  NOR2_X2 U6032 ( .A1(n6165), .A2(n6164), .ZN(n6553) );
  AOI21_X2 U6033 ( .B1(n9365), .B2(n7628), .A(n7627), .ZN(n9348) );
  NAND2_X1 U6034 ( .A1(n6870), .A2(n6869), .ZN(n6875) );
  NAND2_X1 U6035 ( .A1(n9539), .A2(n7546), .ZN(n9522) );
  NAND2_X1 U6036 ( .A1(n6406), .A2(n4442), .ZN(n6414) );
  NAND2_X1 U6037 ( .A1(n6396), .A2(n9042), .ZN(n8839) );
  OAI21_X1 U6038 ( .B1(n9139), .B2(n6430), .A(n6421), .ZN(n6392) );
  AOI21_X2 U6039 ( .B1(n9301), .B2(n9302), .A(n4370), .ZN(n9591) );
  NAND2_X1 U6040 ( .A1(n6414), .A2(n8840), .ZN(n6413) );
  NAND2_X1 U6041 ( .A1(n6582), .A2(n6743), .ZN(n6736) );
  NAND2_X1 U6042 ( .A1(n6433), .A2(n6434), .ZN(n6432) );
  NAND2_X1 U6043 ( .A1(n6853), .A2(n6852), .ZN(n6854) );
  NAND2_X1 U6044 ( .A1(n9441), .A2(n7572), .ZN(n4793) );
  NAND2_X1 U6045 ( .A1(n4446), .A2(n4445), .ZN(n6256) );
  NAND2_X1 U6046 ( .A1(n5492), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4445) );
  INV_X1 U6047 ( .A(n4447), .ZN(n4446) );
  OAI21_X1 U6048 ( .B1(n5528), .B2(n6096), .A(n5018), .ZN(n4447) );
  NAND2_X1 U6049 ( .A1(n4794), .A2(n4939), .ZN(n9441) );
  NOR2_X2 U6050 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  NAND2_X1 U6051 ( .A1(n4556), .A2(n4565), .ZN(n4555) );
  NAND2_X1 U6052 ( .A1(n4855), .A2(n8483), .ZN(n4856) );
  INV_X1 U6053 ( .A(n8731), .ZN(n4468) );
  NAND2_X1 U6054 ( .A1(n5446), .A2(n5445), .ZN(n5466) );
  NAND2_X1 U6055 ( .A1(n4617), .A2(n4619), .ZN(n4616) );
  NAND2_X1 U6056 ( .A1(n4590), .A2(n4936), .ZN(n7391) );
  NAND2_X1 U6057 ( .A1(n5428), .A2(n5427), .ZN(n5444) );
  INV_X1 U6058 ( .A(n8107), .ZN(n8112) );
  NAND2_X1 U6059 ( .A1(n9028), .A2(n9025), .ZN(n4534) );
  NAND2_X1 U6060 ( .A1(n4533), .A2(n4532), .ZN(n9027) );
  OAI21_X1 U6061 ( .B1(n5391), .B2(n5390), .A(n5389), .ZN(n5409) );
  INV_X1 U6062 ( .A(n9022), .ZN(n4537) );
  NAND2_X1 U6063 ( .A1(n4886), .A2(n4887), .ZN(n5164) );
  NAND2_X1 U6064 ( .A1(n6736), .A2(n4454), .ZN(n6739) );
  NAND2_X1 U6065 ( .A1(n9457), .A2(n4795), .ZN(n4794) );
  OR2_X1 U6066 ( .A1(n9276), .A2(n9275), .ZN(n4751) );
  OR2_X2 U6067 ( .A1(n9349), .A2(n9350), .ZN(n9352) );
  OAI21_X1 U6068 ( .B1(n8840), .B2(n8913), .A(n8918), .ZN(n6427) );
  AND3_X2 U6069 ( .A1(n5793), .A2(n4861), .A3(n5792), .ZN(n6204) );
  NAND2_X1 U6070 ( .A1(n5192), .A2(n5191), .ZN(n5208) );
  NAND2_X1 U6071 ( .A1(n8686), .A2(n8475), .ZN(n8759) );
  INV_X1 U6072 ( .A(n8470), .ZN(n4846) );
  NOR2_X1 U6073 ( .A1(n7901), .A2(n8265), .ZN(n7912) );
  NAND2_X1 U6074 ( .A1(n9818), .A2(n9819), .ZN(n9817) );
  OAI21_X1 U6075 ( .B1(n9869), .B2(n6352), .A(n6351), .ZN(n6643) );
  NAND2_X1 U6076 ( .A1(n5130), .A2(n5129), .ZN(n5146) );
  OAI21_X1 U6077 ( .B1(n4749), .B2(n9565), .A(n4747), .ZN(n9585) );
  NAND2_X1 U6078 ( .A1(n5116), .A2(n5115), .ZN(n5130) );
  INV_X1 U6079 ( .A(n4845), .ZN(n4585) );
  NAND2_X1 U6080 ( .A1(n5051), .A2(n5050), .ZN(n5074) );
  OR2_X1 U6081 ( .A1(n8836), .A2(n6096), .ZN(n6097) );
  NAND2_X2 U6082 ( .A1(n9522), .A2(n9521), .ZN(n9520) );
  NAND2_X1 U6083 ( .A1(n4834), .A2(n4345), .ZN(n9301) );
  NAND2_X2 U6084 ( .A1(n5857), .A2(n5847), .ZN(n9748) );
  NAND2_X1 U6085 ( .A1(n5387), .A2(n7247), .ZN(n8143) );
  INV_X1 U6086 ( .A(n7087), .ZN(n4456) );
  OAI21_X1 U6087 ( .B1(n8236), .B2(n5276), .A(n7337), .ZN(n8229) );
  OAI21_X2 U6088 ( .B1(n8098), .B2(n7364), .A(n7363), .ZN(n8089) );
  OAI21_X1 U6089 ( .B1(n4611), .B2(n6938), .A(n4357), .ZN(n4610) );
  OAI21_X1 U6090 ( .B1(n7413), .B2(n4773), .A(n7420), .ZN(n4772) );
  NAND2_X1 U6091 ( .A1(n5012), .A2(n5978), .ZN(n4458) );
  NAND2_X1 U6092 ( .A1(n4909), .A2(n4913), .ZN(n5426) );
  NAND4_X2 U6093 ( .A1(n5793), .A2(n5792), .A3(n4861), .A4(n5794), .ZN(n6294)
         );
  AND2_X2 U6094 ( .A1(n6261), .A2(n6260), .ZN(n4565) );
  NAND2_X1 U6095 ( .A1(n4876), .A2(n4875), .ZN(n9464) );
  NAND2_X1 U6096 ( .A1(n4873), .A2(n4872), .ZN(n9385) );
  NAND2_X1 U6097 ( .A1(n4871), .A2(n4870), .ZN(n9531) );
  INV_X1 U6098 ( .A(n4459), .ZN(n9337) );
  NAND2_X1 U6099 ( .A1(n9307), .A2(n9295), .ZN(n9283) );
  NAND2_X1 U6100 ( .A1(n5023), .A2(n5022), .ZN(n5028) );
  OAI21_X1 U6101 ( .B1(n9678), .B2(n9814), .A(n4460), .ZN(P1_U3553) );
  OAI21_X1 U6102 ( .B1(n9678), .B2(n9811), .A(n4462), .ZN(P1_U3521) );
  NAND3_X1 U6103 ( .A1(n5816), .A2(n5823), .A3(n4552), .ZN(n5830) );
  NAND2_X1 U6104 ( .A1(n4474), .A2(n9456), .ZN(n9460) );
  NAND2_X1 U6105 ( .A1(n9498), .A2(n9068), .ZN(n4757) );
  INV_X1 U6106 ( .A(n9458), .ZN(n4474) );
  NAND2_X1 U6107 ( .A1(n5115), .A2(n4890), .ZN(n4889) );
  NAND2_X1 U6108 ( .A1(n4359), .A2(n6716), .ZN(n7272) );
  NAND2_X1 U6109 ( .A1(n4609), .A2(n4605), .ZN(n4604) );
  NAND2_X1 U6110 ( .A1(n4604), .A2(n4473), .ZN(n4472) );
  OAI21_X2 U6111 ( .B1(n8697), .B2(n8698), .A(n8800), .ZN(n8699) );
  NAND2_X1 U6112 ( .A1(n8759), .A2(n8760), .ZN(n8758) );
  NAND2_X1 U6113 ( .A1(n6157), .A2(n6156), .ZN(n4854) );
  NAND2_X2 U6114 ( .A1(n8549), .A2(n8607), .ZN(n8609) );
  NAND2_X1 U6115 ( .A1(n8664), .A2(n8536), .ZN(n8539) );
  NAND2_X1 U6116 ( .A1(n4584), .A2(n8684), .ZN(n8686) );
  NAND2_X1 U6117 ( .A1(n8665), .A2(n8666), .ZN(n8664) );
  NAND2_X1 U6118 ( .A1(n4554), .A2(n8630), .ZN(n8632) );
  NAND2_X1 U6119 ( .A1(n4770), .A2(n4376), .ZN(n4611) );
  NAND2_X1 U6120 ( .A1(n6761), .A2(n7291), .ZN(n5108) );
  INV_X1 U6121 ( .A(n4610), .ZN(n4609) );
  OAI211_X1 U6122 ( .C1(n7272), .C2(n7429), .A(n4769), .B(n7284), .ZN(n5061)
         );
  NAND2_X1 U6123 ( .A1(n8075), .A2(n8074), .ZN(n5522) );
  OAI21_X1 U6124 ( .B1(n8089), .B2(n8081), .A(n7367), .ZN(n8075) );
  NAND2_X1 U6125 ( .A1(n4772), .A2(n4771), .ZN(n4770) );
  NAND3_X1 U6126 ( .A1(n4472), .A2(n4607), .A3(n4606), .ZN(n7475) );
  NAND2_X1 U6127 ( .A1(n9371), .A2(n9701), .ZN(n9355) );
  NAND2_X4 U6128 ( .A1(n6263), .A2(n6050), .ZN(n8864) );
  INV_X1 U6129 ( .A(n4874), .ZN(n9442) );
  INV_X1 U6130 ( .A(n4863), .ZN(n9306) );
  NOR2_X2 U6131 ( .A1(n9531), .A2(n9657), .ZN(n9513) );
  NOR2_X2 U6132 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  NAND2_X1 U6133 ( .A1(n4751), .A2(n9274), .ZN(n4750) );
  AOI21_X2 U6134 ( .B1(n9396), .B2(n7677), .A(n7676), .ZN(n9382) );
  AOI21_X1 U6135 ( .B1(n8006), .B2(n4430), .A(n4476), .ZN(n4475) );
  NOR2_X1 U6136 ( .A1(n8006), .A2(n8005), .ZN(n8032) );
  NAND2_X1 U6137 ( .A1(n4481), .A2(n8053), .ZN(P2_U3201) );
  NAND3_X1 U6138 ( .A1(n4486), .A2(n4489), .A3(n4713), .ZN(n4482) );
  NAND2_X1 U6139 ( .A1(n4490), .A2(n9852), .ZN(n4489) );
  INV_X1 U6140 ( .A(n6347), .ZN(n4487) );
  NAND3_X1 U6141 ( .A1(n4486), .A2(n4489), .A3(n4484), .ZN(n4483) );
  AND3_X2 U6142 ( .A1(n4356), .A2(n4718), .A3(n4497), .ZN(n9825) );
  NAND3_X1 U6143 ( .A1(n6314), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_2__SCAN_IN), .ZN(n4497) );
  NAND2_X1 U6144 ( .A1(n4501), .A2(n4415), .ZN(n4506) );
  XNOR2_X1 U6145 ( .A(n4506), .B(n4505), .ZN(n6639) );
  NOR2_X2 U6146 ( .A1(n7984), .A2(n4429), .ZN(n8007) );
  NAND2_X1 U6147 ( .A1(n4514), .A2(n6341), .ZN(n4515) );
  INV_X1 U6148 ( .A(n8009), .ZN(n4516) );
  OAI21_X1 U6149 ( .B1(n8009), .B2(n4354), .A(n4432), .ZN(n8036) );
  OAI21_X1 U6150 ( .B1(n4522), .B2(n4521), .A(n4517), .ZN(n4524) );
  NAND2_X1 U6151 ( .A1(n8917), .A2(n4409), .ZN(n4520) );
  NAND3_X1 U6152 ( .A1(n4524), .A2(n4523), .A3(n4381), .ZN(n8947) );
  NAND2_X1 U6153 ( .A1(n4400), .A2(n4525), .ZN(n6383) );
  NAND4_X1 U6154 ( .A1(n8958), .A2(n9071), .A3(n9068), .A4(n9070), .ZN(n4528)
         );
  NAND3_X1 U6155 ( .A1(n8963), .A2(n9076), .A3(n9075), .ZN(n4531) );
  NAND2_X1 U6156 ( .A1(n4541), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5849) );
  NAND4_X1 U6157 ( .A1(n5806), .A2(n4542), .A3(n5792), .A4(n5793), .ZN(n4541)
         );
  NAND2_X1 U6158 ( .A1(n5849), .A2(n5848), .ZN(n5850) );
  NAND3_X1 U6159 ( .A1(n4544), .A2(n4358), .A3(n6396), .ZN(n6397) );
  XNOR2_X1 U6160 ( .A(n4545), .B(n4543), .ZN(n6410) );
  AOI21_X1 U6161 ( .B1(n8972), .B2(n9021), .A(n4549), .ZN(n4548) );
  INV_X2 U6162 ( .A(n5830), .ZN(n5793) );
  NOR2_X2 U6163 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5823) );
  NAND2_X1 U6164 ( .A1(n8632), .A2(n8744), .ZN(n4553) );
  NAND2_X1 U6165 ( .A1(n8628), .A2(n8629), .ZN(n4554) );
  NAND2_X2 U6166 ( .A1(n4341), .A2(n4338), .ZN(n8836) );
  NAND2_X1 U6167 ( .A1(n4837), .A2(n4562), .ZN(n4561) );
  NAND2_X1 U6168 ( .A1(n4856), .A2(n4570), .ZN(n4566) );
  OAI211_X1 U6169 ( .C1(n4571), .C2(n8486), .A(n8495), .B(n4566), .ZN(n8504)
         );
  INV_X1 U6170 ( .A(n8706), .ZN(n4571) );
  NAND2_X1 U6171 ( .A1(n8813), .A2(n8486), .ZN(n8705) );
  NAND2_X1 U6172 ( .A1(n4423), .A2(n4470), .ZN(n8813) );
  OAI21_X1 U6173 ( .B1(n8609), .B2(n4580), .A(n4577), .ZN(n8590) );
  NAND2_X1 U6174 ( .A1(n8609), .A2(n4581), .ZN(n4576) );
  NAND2_X1 U6175 ( .A1(n8609), .A2(n8728), .ZN(n8557) );
  OAI21_X1 U6176 ( .B1(n8609), .B2(n4575), .A(n4573), .ZN(n8653) );
  AND2_X1 U6177 ( .A1(n5806), .A2(n4864), .ZN(n4583) );
  NAND2_X1 U6178 ( .A1(n6204), .A2(n4583), .ZN(n5845) );
  NAND2_X1 U6179 ( .A1(n5845), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5846) );
  NAND2_X2 U6180 ( .A1(n5002), .A2(n6050), .ZN(n5528) );
  AND3_X2 U6181 ( .A1(n5034), .A2(n5035), .A3(n4589), .ZN(n6952) );
  NAND3_X1 U6182 ( .A1(n4603), .A2(n4792), .A3(n4600), .ZN(n7325) );
  NAND3_X1 U6183 ( .A1(n7422), .A2(n4609), .A3(n5583), .ZN(n4606) );
  OAI21_X1 U6184 ( .B1(n4378), .B2(n4614), .A(n4612), .ZN(n7370) );
  OAI21_X2 U6185 ( .B1(n4615), .B2(n4617), .A(n4622), .ZN(n4614) );
  NAND2_X1 U6186 ( .A1(n7361), .A2(n7386), .ZN(n4623) );
  NAND2_X4 U6187 ( .A1(n4634), .A2(n4978), .ZN(n8041) );
  NAND2_X1 U6188 ( .A1(n5603), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4635) );
  NAND2_X1 U6189 ( .A1(n4968), .A2(n4967), .ZN(n5603) );
  OAI21_X1 U6190 ( .B1(n8246), .B2(n4638), .A(n4636), .ZN(n8206) );
  NAND2_X1 U6191 ( .A1(n5574), .A2(n4644), .ZN(n4642) );
  NAND2_X1 U6192 ( .A1(n4642), .A2(n4643), .ZN(n8116) );
  INV_X1 U6193 ( .A(n8182), .ZN(n4652) );
  NAND2_X1 U6194 ( .A1(n4647), .A2(n4648), .ZN(n5572) );
  NAND2_X1 U6195 ( .A1(n8182), .A2(n4650), .ZN(n4647) );
  INV_X1 U6196 ( .A(n5570), .ZN(n4653) );
  INV_X1 U6197 ( .A(n6380), .ZN(n9923) );
  NAND2_X1 U6198 ( .A1(n7891), .A2(n9923), .ZN(n7264) );
  NAND3_X1 U6199 ( .A1(n4676), .A2(n4674), .A3(n4673), .ZN(n5102) );
  INV_X1 U6200 ( .A(n5729), .ZN(n5731) );
  NAND2_X1 U6201 ( .A1(n7772), .A2(n4680), .ZN(n5736) );
  NAND2_X1 U6202 ( .A1(n7693), .A2(n4682), .ZN(n4681) );
  OAI211_X1 U6203 ( .C1(n7693), .C2(n4683), .A(n5783), .B(n4681), .ZN(P2_U3160) );
  NAND2_X1 U6204 ( .A1(n5749), .A2(n4418), .ZN(n4687) );
  NAND2_X1 U6205 ( .A1(n6286), .A2(n4355), .ZN(n6442) );
  INV_X1 U6206 ( .A(n7862), .ZN(n4689) );
  NAND2_X1 U6207 ( .A1(n6903), .A2(n6992), .ZN(n4699) );
  NAND2_X1 U6208 ( .A1(n4699), .A2(n4700), .ZN(n6995) );
  NAND2_X1 U6209 ( .A1(n7026), .A2(n4703), .ZN(n4702) );
  AND2_X1 U6210 ( .A1(n5286), .A2(n4712), .ZN(n4968) );
  NOR2_X2 U6211 ( .A1(n7793), .A2(n7792), .ZN(n7700) );
  NAND2_X1 U6212 ( .A1(n5669), .A2(n5668), .ZN(n6371) );
  NAND2_X1 U6213 ( .A1(n5731), .A2(n5730), .ZN(n7772) );
  NAND2_X1 U6214 ( .A1(n5746), .A2(n5745), .ZN(n7693) );
  NAND2_X1 U6215 ( .A1(n5742), .A2(n7841), .ZN(n7844) );
  MUX2_X1 U6216 ( .A(n6724), .B(P2_REG2_REG_2__SCAN_IN), .S(n9825), .Z(n9819)
         );
  NAND2_X1 U6217 ( .A1(n4417), .A2(n4729), .ZN(n8027) );
  INV_X1 U6218 ( .A(n8011), .ZN(n4731) );
  NAND3_X2 U6219 ( .A1(n7205), .A2(n4739), .A3(n4738), .ZN(n4935) );
  NAND2_X2 U6220 ( .A1(n6985), .A2(n4758), .ZN(n8931) );
  MUX2_X1 U6221 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6050), .Z(n5024) );
  NAND2_X1 U6222 ( .A1(n5108), .A2(n4764), .ZN(n4761) );
  NAND2_X1 U6223 ( .A1(n7284), .A2(n4410), .ZN(n4769) );
  INV_X1 U6224 ( .A(n7260), .ZN(n4768) );
  INV_X1 U6225 ( .A(n7429), .ZN(n6226) );
  NAND2_X1 U6226 ( .A1(n7272), .A2(n7260), .ZN(n6225) );
  NAND2_X1 U6227 ( .A1(n5007), .A2(n4777), .ZN(n7890) );
  INV_X1 U6228 ( .A(n4778), .ZN(n4777) );
  OAI21_X1 U6229 ( .B1(n8143), .B2(n4780), .A(n4779), .ZN(n5442) );
  AND2_X1 U6230 ( .A1(n4968), .A2(n4787), .ZN(n4971) );
  OR2_X1 U6231 ( .A1(n9466), .A2(n9126), .ZN(n4795) );
  NAND2_X1 U6232 ( .A1(n7526), .A2(n4344), .ZN(n4796) );
  NAND2_X1 U6233 ( .A1(n4796), .A2(n4797), .ZN(n9539) );
  NAND2_X1 U6234 ( .A1(n9520), .A2(n4802), .ZN(n4801) );
  NAND2_X1 U6235 ( .A1(n4801), .A2(n4416), .ZN(n9475) );
  NOR2_X1 U6236 ( .A1(n9517), .A2(n8818), .ZN(n4809) );
  CLKBUF_X1 U6237 ( .A(n4820), .Z(n4811) );
  INV_X1 U6238 ( .A(n6129), .ZN(n4826) );
  OAI21_X1 U6239 ( .B1(n4826), .B2(n8836), .A(n6131), .ZN(n4827) );
  INV_X2 U6240 ( .A(n8836), .ZN(n8861) );
  NOR2_X2 U6241 ( .A1(n4380), .A2(n4827), .ZN(n6826) );
  OR2_X2 U6242 ( .A1(n9331), .A2(n7651), .ZN(n4836) );
  NAND3_X1 U6243 ( .A1(n8812), .A2(n8811), .A3(n4419), .ZN(P1_U3240) );
  INV_X1 U6244 ( .A(n9109), .ZN(n7478) );
  NAND2_X1 U6245 ( .A1(n5841), .A2(n5803), .ZN(n4840) );
  INV_X1 U6246 ( .A(n8540), .ZN(n4843) );
  INV_X1 U6247 ( .A(n4842), .ZN(n4841) );
  NAND2_X1 U6248 ( .A1(n4842), .A2(n8606), .ZN(n8549) );
  INV_X1 U6249 ( .A(n6973), .ZN(n8455) );
  NAND2_X1 U6250 ( .A1(n4854), .A2(n4853), .ZN(n6261) );
  INV_X1 U6251 ( .A(n8485), .ZN(n4855) );
  NAND2_X1 U6252 ( .A1(n8557), .A2(n8727), .ZN(n8730) );
  NAND2_X1 U6253 ( .A1(n8730), .A2(n8558), .ZN(n8697) );
  INV_X2 U6254 ( .A(n6267), .ZN(n8646) );
  INV_X1 U6255 ( .A(n6826), .ZN(n6419) );
  NOR2_X2 U6256 ( .A1(n9283), .A2(n9587), .ZN(n9282) );
  NAND2_X1 U6257 ( .A1(n5808), .A2(n5807), .ZN(n5810) );
  NOR2_X2 U6258 ( .A1(n5845), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5860) );
  NAND4_X1 U6259 ( .A1(n6826), .A2(n9045), .A3(n9796), .A4(n4866), .ZN(n6424)
         );
  NOR2_X2 U6260 ( .A1(n9568), .A2(n9729), .ZN(n4871) );
  NOR2_X2 U6261 ( .A1(n9385), .A2(n9372), .ZN(n9371) );
  NOR2_X2 U6262 ( .A1(n9415), .A2(n9404), .ZN(n4873) );
  NOR2_X2 U6263 ( .A1(n9490), .A2(n9645), .ZN(n4876) );
  NAND2_X1 U6264 ( .A1(n4877), .A2(n5094), .ZN(n5100) );
  NAND2_X1 U6265 ( .A1(n5081), .A2(n4877), .ZN(n6262) );
  NAND2_X1 U6266 ( .A1(n5485), .A2(n4883), .ZN(n4881) );
  NAND2_X1 U6267 ( .A1(n5110), .A2(n4888), .ZN(n4886) );
  NAND2_X1 U6268 ( .A1(n5110), .A2(n5109), .ZN(n5116) );
  NAND2_X1 U6269 ( .A1(n4903), .A2(n4353), .ZN(n5348) );
  NAND2_X1 U6270 ( .A1(n5377), .A2(n5376), .ZN(n5391) );
  NAND2_X1 U6271 ( .A1(n4908), .A2(n4910), .ZN(n5428) );
  NAND3_X1 U6272 ( .A1(n5377), .A2(n4913), .A3(n5376), .ZN(n4908) );
  NAND2_X1 U6273 ( .A1(n5526), .A2(n5525), .ZN(n7377) );
  NAND2_X1 U6274 ( .A1(n4927), .A2(n4925), .ZN(n5279) );
  NAND2_X1 U6275 ( .A1(n5244), .A2(n5243), .ZN(n5264) );
  NAND3_X1 U6276 ( .A1(n4935), .A2(n4934), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n4931) );
  NAND2_X2 U6277 ( .A1(n4935), .A2(n4934), .ZN(n5012) );
  NAND2_X1 U6278 ( .A1(n5572), .A2(n8165), .ZN(n8159) );
  NAND2_X1 U6279 ( .A1(n5729), .A2(n5728), .ZN(n5732) );
  OR2_X1 U6280 ( .A1(n4971), .A2(n5031), .ZN(n4973) );
  AOI22_X1 U6281 ( .A1(n9271), .A2(n9270), .B1(n9295), .B2(n9280), .ZN(n9273)
         );
  INV_X1 U6282 ( .A(n4974), .ZN(n8429) );
  XNOR2_X1 U6283 ( .A(n5849), .B(n5809), .ZN(n7477) );
  OAI21_X1 U6284 ( .B1(n8070), .B2(n4941), .A(n5581), .ZN(n5582) );
  NAND2_X1 U6285 ( .A1(n5795), .A2(n4937), .ZN(n5972) );
  OAI222_X1 U6286 ( .A1(P1_U3086), .A2(n9038), .B1(n9747), .B2(n6939), .C1(
        n7586), .C2(n9750), .ZN(P1_U3335) );
  NAND2_X1 U6287 ( .A1(n5348), .A2(n5347), .ZN(n5363) );
  NAND2_X1 U6288 ( .A1(n5279), .A2(n5278), .ZN(n5281) );
  NAND2_X1 U6289 ( .A1(n5524), .A2(n5523), .ZN(n5526) );
  NAND2_X1 U6290 ( .A1(n5002), .A2(n4338), .ZN(n5082) );
  AND2_X2 U6291 ( .A1(n6682), .A2(n8279), .ZN(n8269) );
  AND2_X2 U6292 ( .A1(n6675), .A2(n5652), .ZN(n10192) );
  INV_X1 U6293 ( .A(n8357), .ZN(n5656) );
  NAND2_X1 U6294 ( .A1(n5775), .A2(n7388), .ZN(n8278) );
  AND2_X1 U6295 ( .A1(n5640), .A2(n5639), .ZN(n9966) );
  AND2_X1 U6296 ( .A1(n7390), .A2(n7389), .ZN(n4936) );
  INV_X1 U6297 ( .A(n8420), .ZN(n5643) );
  AND3_X1 U6298 ( .A1(n5963), .A2(n5799), .A3(n10063), .ZN(n4937) );
  INV_X2 U6299 ( .A(n9816), .ZN(n9814) );
  AND2_X1 U6300 ( .A1(n8454), .A2(n8453), .ZN(n4938) );
  OR2_X1 U6301 ( .A1(n4875), .A2(n8709), .ZN(n4939) );
  INV_X1 U6302 ( .A(n9729), .ZN(n7545) );
  INV_X1 U6303 ( .A(n4451), .ZN(n7531) );
  AND2_X1 U6304 ( .A1(n8373), .A2(n8083), .ZN(n4941) );
  INV_X1 U6305 ( .A(n9432), .ZN(n9717) );
  AND2_X1 U6306 ( .A1(n9495), .A2(n8708), .ZN(n4942) );
  OR2_X1 U6307 ( .A1(n7868), .A2(n7388), .ZN(n7389) );
  NAND2_X1 U6308 ( .A1(n7243), .A2(n7869), .ZN(n5581) );
  INV_X1 U6309 ( .A(n6105), .ZN(n6267) );
  INV_X1 U6310 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6485) );
  INV_X1 U6311 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5799) );
  INV_X1 U6312 ( .A(n6444), .ZN(n5679) );
  INV_X1 U6313 ( .A(n8370), .ZN(n7385) );
  INV_X1 U6314 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6516) );
  OR2_X1 U6315 ( .A1(n8535), .A2(n8534), .ZN(n8536) );
  OR2_X1 U6316 ( .A1(n9634), .A2(n9125), .ZN(n7572) );
  INV_X1 U6317 ( .A(n8945), .ZN(n9556) );
  NAND2_X1 U6318 ( .A1(n5743), .A2(n8109), .ZN(n5744) );
  INV_X1 U6319 ( .A(n5368), .ZN(n5367) );
  INV_X1 U6320 ( .A(n5399), .ZN(n5398) );
  INV_X1 U6321 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5064) );
  XNOR2_X1 U6322 ( .A(n5582), .B(n7462), .ZN(n5585) );
  NAND2_X1 U6323 ( .A1(n5292), .A2(n5291), .ZN(n5315) );
  NAND2_X1 U6324 ( .A1(n5255), .A2(n5254), .ZN(n5270) );
  INV_X1 U6325 ( .A(n7388), .ZN(n7386) );
  OR2_X1 U6326 ( .A1(n5648), .A2(n5632), .ZN(n5759) );
  XNOR2_X1 U6327 ( .A(n6054), .B(n8565), .ZN(n6100) );
  INV_X1 U6328 ( .A(n6270), .ZN(n6269) );
  INV_X1 U6329 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6748) );
  AND2_X1 U6330 ( .A1(n8801), .A2(n8799), .ZN(n8573) );
  NOR2_X1 U6331 ( .A1(n7622), .A2(n8615), .ZN(n7644) );
  OR2_X1 U6332 ( .A1(n7611), .A2(n7610), .ZN(n7622) );
  INV_X1 U6333 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10078) );
  OR2_X1 U6334 ( .A1(n7110), .A2(n7111), .ZN(n7194) );
  INV_X1 U6335 ( .A(n6455), .ZN(n6192) );
  OR2_X1 U6336 ( .A1(n6475), .A2(n9138), .ZN(n6476) );
  OR2_X1 U6337 ( .A1(n9140), .A2(n6419), .ZN(n6389) );
  INV_X1 U6338 ( .A(n8819), .ZN(n9259) );
  NAND2_X1 U6339 ( .A1(n5444), .A2(n5443), .ZN(n5446) );
  NAND2_X1 U6340 ( .A1(n5111), .A2(SI_7_), .ZN(n5129) );
  OR2_X1 U6341 ( .A1(n5417), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5434) );
  OR2_X1 U6342 ( .A1(n5355), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5368) );
  AND2_X1 U6343 ( .A1(n7840), .A2(n5740), .ZN(n7746) );
  INV_X1 U6344 ( .A(n6929), .ZN(n6221) );
  NAND2_X1 U6345 ( .A1(n5065), .A2(n5064), .ZN(n5088) );
  AND2_X1 U6346 ( .A1(n6310), .A2(n6309), .ZN(n9906) );
  INV_X1 U6347 ( .A(n8081), .ZN(n8088) );
  NAND2_X1 U6348 ( .A1(n5455), .A2(n5454), .ZN(n5476) );
  INV_X1 U6349 ( .A(n7875), .ZN(n8197) );
  AND2_X1 U6350 ( .A1(n9952), .A2(n7417), .ZN(n5755) );
  AND2_X1 U6351 ( .A1(n7386), .A2(n5650), .ZN(n6670) );
  INV_X1 U6352 ( .A(n7879), .ZN(n8277) );
  OR2_X1 U6353 ( .A1(n5194), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5230) );
  OR2_X1 U6354 ( .A1(n7552), .A2(n7551), .ZN(n7564) );
  NOR2_X1 U6355 ( .A1(n7538), .A2(n7537), .ZN(n7540) );
  INV_X1 U6356 ( .A(n6176), .ZN(n6177) );
  OR2_X1 U6357 ( .A1(n7579), .A2(n7578), .ZN(n7589) );
  NAND2_X1 U6358 ( .A1(n6113), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6004) );
  OR2_X1 U6359 ( .A1(n9760), .A2(n9759), .ZN(n9762) );
  INV_X1 U6360 ( .A(n8857), .ZN(n9333) );
  AND2_X1 U6361 ( .A1(n8985), .A2(n8992), .ZN(n9367) );
  OR2_X1 U6362 ( .A1(n6028), .A2(n8902), .ZN(n8819) );
  AND2_X1 U6363 ( .A1(n6201), .A2(n6200), .ZN(n9565) );
  AND2_X1 U6364 ( .A1(n5243), .A2(n5226), .ZN(n5227) );
  INV_X1 U6365 ( .A(n5171), .ZN(n5169) );
  AND2_X1 U6366 ( .A1(n5109), .A2(n5098), .ZN(n5099) );
  INV_X1 U6367 ( .A(n7810), .ZN(n7857) );
  NAND2_X1 U6368 ( .A1(n5770), .A2(n5769), .ZN(n7850) );
  OR2_X1 U6369 ( .A1(n8054), .A2(n5063), .ZN(n7411) );
  AND4_X1 U6370 ( .A1(n5321), .A2(n5320), .A3(n5319), .A4(n5318), .ZN(n8224)
         );
  AND4_X1 U6371 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n8275)
         );
  AND2_X1 U6372 ( .A1(P2_U3893), .A2(n6307), .ZN(n9867) );
  INV_X1 U6373 ( .A(n9882), .ZN(n9897) );
  OR2_X1 U6374 ( .A1(n9947), .A2(n6676), .ZN(n8255) );
  AND2_X1 U6375 ( .A1(n5772), .A2(n7388), .ZN(n8209) );
  NAND2_X1 U6376 ( .A1(n6071), .A2(n5755), .ZN(n8279) );
  INV_X1 U6377 ( .A(n8279), .ZN(n8218) );
  INV_X1 U6378 ( .A(n8287), .ZN(n8267) );
  AND2_X1 U6379 ( .A1(n5649), .A2(n5648), .ZN(n6675) );
  INV_X1 U6380 ( .A(n9947), .ZN(n9964) );
  NAND2_X1 U6381 ( .A1(n7134), .A2(n9938), .ZN(n9933) );
  NAND2_X1 U6382 ( .A1(n7152), .A2(n7417), .ZN(n9947) );
  AND2_X1 U6383 ( .A1(n5266), .A2(n5251), .ZN(n7930) );
  AND4_X1 U6384 ( .A1(n7669), .A2(n7668), .A3(n7667), .A4(n7666), .ZN(n9280)
         );
  INV_X1 U6385 ( .A(n4443), .ZN(n7663) );
  AND2_X1 U6386 ( .A1(n6236), .A2(n6235), .ZN(n9251) );
  AND2_X1 U6387 ( .A1(n5939), .A2(n9257), .ZN(n9779) );
  NAND2_X1 U6388 ( .A1(n9106), .A2(n5992), .ZN(n9433) );
  AND2_X1 U6389 ( .A1(n5976), .A2(n5975), .ZN(n9658) );
  NAND2_X1 U6390 ( .A1(n5948), .A2(n5947), .ZN(n6455) );
  INV_X1 U6391 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10014) );
  NOR2_X1 U6392 ( .A1(n9996), .A2(n9995), .ZN(n7061) );
  INV_X1 U6393 ( .A(n5782), .ZN(n5783) );
  INV_X1 U6394 ( .A(n7845), .ZN(n7861) );
  AND2_X1 U6395 ( .A1(n5756), .A2(n8279), .ZN(n7853) );
  AND2_X1 U6396 ( .A1(n7411), .A2(n5534), .ZN(n8073) );
  INV_X1 U6397 ( .A(n8161), .ZN(n7873) );
  OR2_X1 U6398 ( .A1(P2_U3150), .A2(n6308), .ZN(n9882) );
  INV_X1 U6399 ( .A(n9867), .ZN(n9911) );
  INV_X1 U6400 ( .A(n9901), .ZN(n8000) );
  OR2_X1 U6401 ( .A1(n8269), .A2(n6715), .ZN(n8287) );
  NAND2_X1 U6402 ( .A1(n10192), .A2(n9964), .ZN(n8357) );
  INV_X1 U6403 ( .A(n10192), .ZN(n10190) );
  OR2_X1 U6404 ( .A1(n9966), .A2(n9947), .ZN(n8420) );
  INV_X2 U6405 ( .A(n9966), .ZN(n9965) );
  OR2_X1 U6406 ( .A1(n5762), .A2(P2_U3151), .ZN(n8423) );
  INV_X1 U6407 ( .A(n9625), .ZN(n9421) );
  OR3_X1 U6408 ( .A1(n6002), .A2(n5977), .A3(n9658), .ZN(n8786) );
  INV_X1 U6409 ( .A(n8784), .ZN(n8828) );
  OAI21_X1 U6410 ( .B1(n9325), .B2(n7663), .A(n7662), .ZN(n9117) );
  INV_X1 U6411 ( .A(n8930), .ZN(n9136) );
  AOI21_X1 U6412 ( .B1(n7681), .B2(n9526), .A(n8654), .ZN(n9300) );
  OR2_X1 U6413 ( .A1(n9802), .A2(n6540), .ZN(n9551) );
  AND2_X1 U6414 ( .A1(n6462), .A2(n9433), .ZN(n9573) );
  INV_X1 U6415 ( .A(n6473), .ZN(n9802) );
  NAND2_X1 U6416 ( .A1(n9816), .A2(n9658), .ZN(n9643) );
  NAND2_X1 U6417 ( .A1(n9725), .A2(n9658), .ZN(n9722) );
  NOR2_X1 U6418 ( .A1(n6210), .A2(n6209), .ZN(n9813) );
  INV_X1 U6419 ( .A(n9813), .ZN(n9811) );
  NAND2_X1 U6420 ( .A1(n9106), .A2(n6455), .ZN(n9804) );
  INV_X1 U6421 ( .A(n9025), .ZN(n9044) );
  INV_X1 U6422 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U6423 ( .A1(n7062), .A2(n7061), .ZN(n9994) );
  INV_X2 U6424 ( .A(n7871), .ZN(P2_U3893) );
  NOR2_X1 U6425 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4949) );
  NOR2_X1 U6426 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4948) );
  NOR2_X1 U6427 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4947) );
  NAND2_X1 U6428 ( .A1(n4959), .A2(n4960), .ZN(n4952) );
  INV_X1 U6429 ( .A(n5596), .ZN(n4953) );
  NAND2_X1 U6430 ( .A1(n4953), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4954) );
  INV_X1 U6431 ( .A(n4968), .ZN(n4955) );
  NAND2_X1 U6432 ( .A1(n4955), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4956) );
  MUX2_X1 U6433 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4956), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n4957) );
  NAND2_X1 U6434 ( .A1(n4957), .A2(n4364), .ZN(n6938) );
  NAND2_X1 U6435 ( .A1(n4958), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6436 ( .A1(n5328), .A2(n4959), .ZN(n5330) );
  NAND2_X1 U6437 ( .A1(n5330), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4961) );
  INV_X1 U6438 ( .A(n8046), .ZN(n5583) );
  AND2_X1 U6439 ( .A1(n6938), .A2(n5583), .ZN(n6676) );
  INV_X1 U6440 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5599) );
  NAND4_X1 U6441 ( .A1(n5605), .A2(n5599), .A3(n5595), .A4(n4962), .ZN(n4966)
         );
  INV_X1 U6442 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4963) );
  NAND3_X1 U6443 ( .A1(n4964), .A2(n5635), .A3(n4963), .ZN(n4965) );
  INV_X1 U6444 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4976) );
  INV_X1 U6445 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4972) );
  INV_X1 U6446 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4969) );
  INV_X4 U6447 ( .A(n5338), .ZN(n7404) );
  NAND2_X1 U6448 ( .A1(n7404), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4996) );
  INV_X1 U6449 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6299) );
  OR2_X1 U6450 ( .A1(n4339), .A2(n6299), .ZN(n4995) );
  INV_X1 U6451 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6930) );
  OR2_X1 U6452 ( .A1(n5063), .A2(n6930), .ZN(n4994) );
  OR2_X1 U6453 ( .A1(n5020), .A2(n10089), .ZN(n4993) );
  NAND2_X1 U6454 ( .A1(n4979), .A2(SI_1_), .ZN(n5010) );
  INV_X1 U6455 ( .A(n4979), .ZN(n4981) );
  INV_X1 U6456 ( .A(SI_1_), .ZN(n4980) );
  NAND2_X1 U6457 ( .A1(n4981), .A2(n4980), .ZN(n4982) );
  INV_X1 U6458 ( .A(n4986), .ZN(n4984) );
  INV_X1 U6459 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4983) );
  INV_X1 U6460 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U6461 ( .A1(n4984), .A2(n4985), .ZN(n5011) );
  NAND2_X1 U6462 ( .A1(n4986), .A2(n4457), .ZN(n4987) );
  NAND2_X1 U6463 ( .A1(n5011), .A2(n4987), .ZN(n6051) );
  INV_X1 U6464 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U6465 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4989) );
  MUX2_X1 U6466 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4989), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n4990) );
  NAND2_X1 U6467 ( .A1(n5030), .A2(n6573), .ZN(n4991) );
  NAND2_X1 U6468 ( .A1(n4992), .A2(n6380), .ZN(n7268) );
  NAND4_X1 U6469 ( .A1(n4996), .A2(n4995), .A3(n4994), .A4(n4993), .ZN(n7891)
         );
  INV_X1 U6470 ( .A(n7431), .ZN(n5003) );
  INV_X1 U6471 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n4997) );
  INV_X1 U6472 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6362) );
  OR2_X1 U6473 ( .A1(n5005), .A2(n6362), .ZN(n5000) );
  INV_X1 U6474 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6774) );
  OR2_X1 U6475 ( .A1(n5063), .A2(n6774), .ZN(n4999) );
  INV_X1 U6476 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6363) );
  OR2_X1 U6477 ( .A1(n5020), .A2(n6363), .ZN(n4998) );
  NAND4_X1 U6478 ( .A1(n4402), .A2(n5000), .A3(n4999), .A4(n4998), .ZN(n6934)
         );
  NAND2_X1 U6479 ( .A1(n6050), .A2(SI_0_), .ZN(n5001) );
  XNOR2_X1 U6480 ( .A(n5001), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8441) );
  MUX2_X1 U6481 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8441), .S(n5002), .Z(n6777) );
  INV_X1 U6482 ( .A(n6777), .ZN(n8364) );
  OR2_X1 U6483 ( .A1(n6934), .A2(n8364), .ZN(n6929) );
  NAND2_X1 U6484 ( .A1(n5003), .A2(n6221), .ZN(n5004) );
  NAND2_X1 U6485 ( .A1(n5004), .A2(n7268), .ZN(n6716) );
  INV_X1 U6486 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5006) );
  OR2_X1 U6487 ( .A1(n5338), .A2(n5006), .ZN(n5009) );
  INV_X1 U6488 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6259) );
  OR2_X1 U6489 ( .A1(n4340), .A2(n6259), .ZN(n5008) );
  INV_X1 U6490 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6724) );
  OR2_X1 U6491 ( .A1(n5020), .A2(n6724), .ZN(n5007) );
  INV_X1 U6492 ( .A(n5014), .ZN(n5016) );
  NAND2_X1 U6493 ( .A1(n5016), .A2(n5015), .ZN(n5023) );
  NAND2_X1 U6494 ( .A1(n5017), .A2(n5023), .ZN(n6096) );
  INV_X1 U6495 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U6496 ( .A1(n5030), .A2(n9825), .ZN(n5018) );
  NAND2_X1 U6497 ( .A1(n6376), .A2(n6256), .ZN(n7260) );
  NAND2_X1 U6498 ( .A1(n7890), .A2(n9927), .ZN(n7261) );
  NAND2_X1 U6499 ( .A1(n7404), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5544) );
  INV_X1 U6500 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5019) );
  OR2_X1 U6501 ( .A1(n4339), .A2(n5019), .ZN(n5543) );
  OR2_X1 U6502 ( .A1(n5063), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5542) );
  INV_X1 U6503 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5021) );
  OR2_X1 U6504 ( .A1(n5020), .A2(n5021), .ZN(n5541) );
  NAND4_X1 U6505 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .ZN(n7889)
         );
  NAND2_X1 U6506 ( .A1(n5024), .A2(SI_3_), .ZN(n5044) );
  INV_X1 U6507 ( .A(SI_3_), .ZN(n5025) );
  AND2_X1 U6508 ( .A1(n5044), .A2(n5026), .ZN(n5027) );
  NAND2_X1 U6509 ( .A1(n5028), .A2(n5027), .ZN(n5045) );
  OR2_X1 U6510 ( .A1(n5028), .A2(n5027), .ZN(n5029) );
  AND2_X1 U6511 ( .A1(n5045), .A2(n5029), .ZN(n6129) );
  NAND2_X1 U6512 ( .A1(n5492), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U6513 ( .A1(n4356), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5032) );
  MUX2_X1 U6514 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5032), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5033) );
  NAND2_X1 U6515 ( .A1(n5787), .A2(n6345), .ZN(n5034) );
  NAND2_X1 U6516 ( .A1(n5529), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5043) );
  INV_X1 U6517 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5036) );
  OR2_X1 U6518 ( .A1(n5338), .A2(n5036), .ZN(n5042) );
  NAND2_X1 U6519 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5039) );
  AND2_X1 U6520 ( .A1(n5066), .A2(n5039), .ZN(n6446) );
  OR2_X1 U6521 ( .A1(n5063), .A2(n6446), .ZN(n5041) );
  INV_X1 U6522 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6348) );
  OR2_X1 U6523 ( .A1(n5532), .A2(n6348), .ZN(n5040) );
  NAND4_X1 U6524 ( .A1(n5043), .A2(n5042), .A3(n5041), .A4(n5040), .ZN(n7888)
         );
  MUX2_X1 U6525 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5012), .Z(n5046) );
  NAND2_X1 U6526 ( .A1(n5046), .A2(SI_4_), .ZN(n5073) );
  INV_X1 U6527 ( .A(n5046), .ZN(n5048) );
  INV_X1 U6528 ( .A(SI_4_), .ZN(n5047) );
  NAND2_X1 U6529 ( .A1(n5048), .A2(n5047), .ZN(n5049) );
  NAND2_X1 U6530 ( .A1(n5074), .A2(n5052), .ZN(n6162) );
  NAND2_X1 U6531 ( .A1(n5492), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6532 ( .A1(n5054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5053) );
  MUX2_X1 U6533 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5053), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5057) );
  INV_X1 U6534 ( .A(n5054), .ZN(n5056) );
  INV_X1 U6535 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U6536 ( .A1(n5056), .A2(n5055), .ZN(n5083) );
  NAND2_X1 U6537 ( .A1(n5057), .A2(n5083), .ZN(n9835) );
  INV_X1 U6538 ( .A(n9835), .ZN(n6349) );
  NAND2_X1 U6539 ( .A1(n5787), .A2(n6349), .ZN(n5058) );
  OAI211_X1 U6540 ( .C1(n5528), .C2(n6162), .A(n5059), .B(n5058), .ZN(n9931)
         );
  NOR2_X1 U6541 ( .A1(n7888), .A2(n9931), .ZN(n5548) );
  INV_X1 U6542 ( .A(n5548), .ZN(n5060) );
  NAND2_X1 U6543 ( .A1(n7888), .A2(n9931), .ZN(n5547) );
  NAND2_X1 U6544 ( .A1(n5060), .A2(n5547), .ZN(n7434) );
  NAND2_X1 U6545 ( .A1(n5061), .A2(n7434), .ZN(n6947) );
  INV_X1 U6546 ( .A(n7888), .ZN(n6678) );
  NAND2_X1 U6547 ( .A1(n6678), .A2(n9931), .ZN(n7277) );
  NAND2_X1 U6548 ( .A1(n6947), .A2(n7277), .ZN(n6668) );
  NAND2_X1 U6549 ( .A1(n5529), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5072) );
  INV_X1 U6550 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5062) );
  OR2_X1 U6551 ( .A1(n5338), .A2(n5062), .ZN(n5071) );
  INV_X1 U6552 ( .A(n5066), .ZN(n5065) );
  NAND2_X1 U6553 ( .A1(n5066), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5067) );
  AND2_X1 U6554 ( .A1(n5088), .A2(n5067), .ZN(n6698) );
  OR2_X1 U6555 ( .A1(n5063), .A2(n6698), .ZN(n5070) );
  INV_X1 U6556 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5068) );
  OR2_X1 U6557 ( .A1(n5532), .A2(n5068), .ZN(n5069) );
  NAND4_X1 U6558 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), .ZN(n7887)
         );
  NAND2_X1 U6559 ( .A1(n5075), .A2(SI_5_), .ZN(n5094) );
  INV_X1 U6560 ( .A(n5075), .ZN(n5077) );
  INV_X1 U6561 ( .A(SI_5_), .ZN(n5076) );
  NAND2_X1 U6562 ( .A1(n5077), .A2(n5076), .ZN(n5078) );
  OR2_X1 U6563 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  NOR2_X1 U6564 ( .A1(n6262), .A2(n5528), .ZN(n5087) );
  NAND2_X1 U6565 ( .A1(n5083), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5085) );
  INV_X1 U6566 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5084) );
  XNOR2_X1 U6567 ( .A(n5085), .B(n5084), .ZN(n9858) );
  OAI22_X1 U6568 ( .A1(n5327), .A2(n4435), .B1(n4448), .B2(n9858), .ZN(n5086)
         );
  NAND2_X1 U6569 ( .A1(n7887), .A2(n9937), .ZN(n7286) );
  NAND2_X1 U6570 ( .A1(n6668), .A2(n7286), .ZN(n6761) );
  NAND2_X1 U6571 ( .A1(n7404), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5093) );
  INV_X1 U6572 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6765) );
  OR2_X1 U6573 ( .A1(n5532), .A2(n6765), .ZN(n5092) );
  NAND2_X1 U6574 ( .A1(n5088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5089) );
  AND2_X1 U6575 ( .A1(n5123), .A2(n5089), .ZN(n6766) );
  OR2_X1 U6576 ( .A1(n5063), .A2(n6766), .ZN(n5091) );
  OR2_X1 U6577 ( .A1(n4339), .A2(n6781), .ZN(n5090) );
  MUX2_X1 U6578 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4338), .Z(n5095) );
  INV_X1 U6579 ( .A(n5095), .ZN(n5097) );
  INV_X1 U6580 ( .A(SI_6_), .ZN(n5096) );
  NAND2_X1 U6581 ( .A1(n5097), .A2(n5096), .ZN(n5098) );
  OR2_X1 U6582 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  NAND2_X1 U6583 ( .A1(n5110), .A2(n5101), .ZN(n6478) );
  OR2_X1 U6584 ( .A1(n6478), .A2(n5528), .ZN(n5107) );
  NAND2_X1 U6585 ( .A1(n5102), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5103) );
  MUX2_X1 U6586 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5103), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5105) );
  AND2_X1 U6587 ( .A1(n5105), .A2(n5104), .ZN(n6644) );
  AOI22_X1 U6588 ( .A1(n5312), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5787), .B2(
        n6644), .ZN(n5106) );
  NAND2_X1 U6589 ( .A1(n5107), .A2(n5106), .ZN(n6768) );
  NAND2_X1 U6590 ( .A1(n6811), .A2(n6768), .ZN(n7280) );
  NAND2_X1 U6591 ( .A1(n5682), .A2(n6667), .ZN(n7278) );
  AND2_X1 U6592 ( .A1(n7280), .A2(n7278), .ZN(n7291) );
  NAND2_X1 U6593 ( .A1(n7886), .A2(n6802), .ZN(n7290) );
  INV_X1 U6594 ( .A(n5111), .ZN(n5113) );
  INV_X1 U6595 ( .A(SI_7_), .ZN(n5112) );
  NAND2_X1 U6596 ( .A1(n5113), .A2(n5112), .ZN(n5114) );
  OR2_X1 U6597 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  NAND2_X1 U6598 ( .A1(n5130), .A2(n5117), .ZN(n6511) );
  OR2_X1 U6599 ( .A1(n6511), .A2(n5528), .ZN(n5120) );
  NAND2_X1 U6600 ( .A1(n5104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5118) );
  XNOR2_X1 U6601 ( .A(n5118), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6647) );
  AOI22_X1 U6602 ( .A1(n5312), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5787), .B2(
        n6647), .ZN(n5119) );
  NAND2_X1 U6603 ( .A1(n7404), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5128) );
  INV_X1 U6604 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6622) );
  OR2_X1 U6605 ( .A1(n4339), .A2(n6622), .ZN(n5127) );
  NAND2_X1 U6606 ( .A1(n5123), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5124) );
  AND2_X1 U6607 ( .A1(n5136), .A2(n5124), .ZN(n6904) );
  OR2_X1 U6608 ( .A1(n5063), .A2(n6904), .ZN(n5126) );
  INV_X1 U6609 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6623) );
  OR2_X1 U6610 ( .A1(n5532), .A2(n6623), .ZN(n5125) );
  OR2_X1 U6611 ( .A1(n6960), .A2(n6924), .ZN(n6920) );
  NAND2_X1 U6612 ( .A1(n6960), .A2(n6924), .ZN(n7303) );
  MUX2_X1 U6613 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n4337), .Z(n5142) );
  NAND2_X1 U6614 ( .A1(n6737), .A2(n7401), .ZN(n5134) );
  OR2_X1 U6615 ( .A1(n5131), .A2(n5031), .ZN(n5132) );
  XNOR2_X1 U6616 ( .A(n5132), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6649) );
  AOI22_X1 U6617 ( .A1(n5312), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5787), .B2(
        n6649), .ZN(n5133) );
  NAND2_X1 U6618 ( .A1(n5134), .A2(n5133), .ZN(n9945) );
  NAND2_X1 U6619 ( .A1(n5529), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5141) );
  INV_X1 U6620 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5135) );
  OR2_X1 U6621 ( .A1(n5338), .A2(n5135), .ZN(n5140) );
  NAND2_X1 U6622 ( .A1(n5136), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5137) );
  AND2_X1 U6623 ( .A1(n5154), .A2(n5137), .ZN(n6987) );
  OR2_X1 U6624 ( .A1(n5063), .A2(n6987), .ZN(n5139) );
  INV_X1 U6625 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6648) );
  OR2_X1 U6626 ( .A1(n5532), .A2(n6648), .ZN(n5138) );
  NAND4_X1 U6627 ( .A1(n5141), .A2(n5140), .A3(n5139), .A4(n5138), .ZN(n7884)
         );
  OR2_X1 U6628 ( .A1(n9945), .A2(n7085), .ZN(n7295) );
  AND2_X1 U6629 ( .A1(n7295), .A2(n6920), .ZN(n7302) );
  NAND2_X1 U6630 ( .A1(n9945), .A2(n7085), .ZN(n7304) );
  INV_X1 U6631 ( .A(n5142), .ZN(n5144) );
  INV_X1 U6632 ( .A(SI_8_), .ZN(n5143) );
  MUX2_X1 U6633 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n4338), .Z(n5161) );
  XNOR2_X1 U6634 ( .A(n5164), .B(n5163), .ZN(n6833) );
  NAND2_X1 U6635 ( .A1(n6833), .A2(n7401), .ZN(n5150) );
  INV_X1 U6636 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5147) );
  AND2_X1 U6637 ( .A1(n5131), .A2(n5147), .ZN(n5175) );
  OR2_X1 U6638 ( .A1(n5175), .A2(n5031), .ZN(n5148) );
  XNOR2_X1 U6639 ( .A(n5148), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7007) );
  AOI22_X1 U6640 ( .A1(n5312), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5787), .B2(
        n7007), .ZN(n5149) );
  NAND2_X1 U6641 ( .A1(n5150), .A2(n5149), .ZN(n7101) );
  NAND2_X1 U6642 ( .A1(n7404), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5160) );
  INV_X1 U6643 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5151) );
  OR2_X1 U6644 ( .A1(n4339), .A2(n5151), .ZN(n5159) );
  INV_X1 U6645 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6646 ( .A1(n5154), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5155) );
  AND2_X1 U6647 ( .A1(n5185), .A2(n5155), .ZN(n7027) );
  OR2_X1 U6648 ( .A1(n5063), .A2(n7027), .ZN(n5158) );
  INV_X1 U6649 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5156) );
  OR2_X1 U6650 ( .A1(n5532), .A2(n5156), .ZN(n5157) );
  NAND4_X1 U6651 ( .A1(n5160), .A2(n5159), .A3(n5158), .A4(n5157), .ZN(n7883)
         );
  INV_X1 U6652 ( .A(n7883), .ZN(n6925) );
  OR2_X1 U6653 ( .A1(n7101), .A2(n6925), .ZN(n7301) );
  NAND2_X1 U6654 ( .A1(n7101), .A2(n6925), .ZN(n7305) );
  NAND2_X1 U6655 ( .A1(n7301), .A2(n7305), .ZN(n7445) );
  NAND2_X1 U6656 ( .A1(n7089), .A2(n7301), .ZN(n7129) );
  MUX2_X1 U6657 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4338), .Z(n5165) );
  INV_X1 U6658 ( .A(n5165), .ZN(n5167) );
  INV_X1 U6659 ( .A(SI_10_), .ZN(n5166) );
  NAND2_X1 U6660 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  INV_X1 U6661 ( .A(n5170), .ZN(n5172) );
  NAND2_X1 U6662 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  NAND2_X1 U6663 ( .A1(n5192), .A2(n5173), .ZN(n6871) );
  OR2_X1 U6664 ( .A1(n6871), .A2(n5528), .ZN(n5183) );
  INV_X1 U6665 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5174) );
  NOR2_X1 U6666 ( .A1(n5179), .A2(n5031), .ZN(n5176) );
  MUX2_X1 U6667 ( .A(n5031), .B(n5176), .S(P2_IR_REG_10__SCAN_IN), .Z(n5177)
         );
  INV_X1 U6668 ( .A(n5177), .ZN(n5180) );
  INV_X1 U6669 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6670 ( .A1(n5179), .A2(n5178), .ZN(n5194) );
  NAND2_X1 U6671 ( .A1(n5180), .A2(n5194), .ZN(n7170) );
  INV_X1 U6672 ( .A(n7170), .ZN(n5181) );
  AOI22_X1 U6673 ( .A1(n5312), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5787), .B2(
        n5181), .ZN(n5182) );
  NAND2_X1 U6674 ( .A1(n5183), .A2(n5182), .ZN(n7137) );
  INV_X1 U6675 ( .A(n7137), .ZN(n9948) );
  NAND2_X1 U6676 ( .A1(n7404), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5190) );
  INV_X1 U6677 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5184) );
  OR2_X1 U6678 ( .A1(n4339), .A2(n5184), .ZN(n5189) );
  NAND2_X1 U6679 ( .A1(n5185), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5186) );
  AND2_X1 U6680 ( .A1(n5199), .A2(n5186), .ZN(n7225) );
  OR2_X1 U6681 ( .A1(n5063), .A2(n7225), .ZN(n5188) );
  INV_X1 U6682 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7135) );
  OR2_X1 U6683 ( .A1(n5532), .A2(n7135), .ZN(n5187) );
  AND2_X1 U6684 ( .A1(n9948), .A2(n7882), .ZN(n7300) );
  INV_X1 U6685 ( .A(n7882), .ZN(n7086) );
  NAND2_X1 U6686 ( .A1(n7137), .A2(n7086), .ZN(n7315) );
  MUX2_X1 U6687 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4338), .Z(n5206) );
  XNOR2_X1 U6688 ( .A(n5208), .B(n5207), .ZN(n7527) );
  NAND2_X1 U6689 ( .A1(n7527), .A2(n7401), .ZN(n5197) );
  NAND2_X1 U6690 ( .A1(n5194), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5193) );
  MUX2_X1 U6691 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5193), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5195) );
  AND2_X1 U6692 ( .A1(n5195), .A2(n5230), .ZN(n7171) );
  AOI22_X1 U6693 ( .A1(n5312), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5787), .B2(
        n7171), .ZN(n5196) );
  NAND2_X1 U6694 ( .A1(n5197), .A2(n5196), .ZN(n9957) );
  NAND2_X1 U6695 ( .A1(n7404), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5204) );
  INV_X1 U6696 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5198) );
  OR2_X1 U6697 ( .A1(n4339), .A2(n5198), .ZN(n5203) );
  NAND2_X1 U6698 ( .A1(n5199), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5200) );
  AND2_X1 U6699 ( .A1(n5235), .A2(n5200), .ZN(n7822) );
  OR2_X1 U6700 ( .A1(n5063), .A2(n7822), .ZN(n5202) );
  INV_X1 U6701 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7147) );
  OR2_X1 U6702 ( .A1(n5532), .A2(n7147), .ZN(n5201) );
  NAND2_X1 U6703 ( .A1(n9957), .A2(n8275), .ZN(n7316) );
  MUX2_X1 U6704 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4338), .Z(n5209) );
  NAND2_X1 U6705 ( .A1(n5211), .A2(n5210), .ZN(n5212) );
  NAND2_X1 U6706 ( .A1(n5212), .A2(n5222), .ZN(n7533) );
  OR2_X1 U6707 ( .A1(n7533), .A2(n5528), .ZN(n5215) );
  NAND2_X1 U6708 ( .A1(n5230), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5213) );
  XNOR2_X1 U6709 ( .A(n5213), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7177) );
  AOI22_X1 U6710 ( .A1(n5312), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5787), .B2(
        n7177), .ZN(n5214) );
  NAND2_X1 U6711 ( .A1(n5529), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5220) );
  INV_X1 U6712 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5216) );
  OR2_X1 U6713 ( .A1(n5338), .A2(n5216), .ZN(n5219) );
  INV_X1 U6714 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10170) );
  XNOR2_X1 U6715 ( .A(n5235), .B(n10170), .ZN(n8280) );
  OR2_X1 U6716 ( .A1(n4340), .A2(n8280), .ZN(n5218) );
  INV_X1 U6717 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8281) );
  OR2_X1 U6718 ( .A1(n5532), .A2(n8281), .ZN(n5217) );
  NAND4_X1 U6719 ( .A1(n5220), .A2(n5219), .A3(n5218), .A4(n5217), .ZN(n7880)
         );
  NAND2_X1 U6720 ( .A1(n9963), .A2(n8258), .ZN(n7323) );
  NAND2_X1 U6721 ( .A1(n7322), .A2(n7323), .ZN(n8272) );
  MUX2_X1 U6722 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4338), .Z(n5223) );
  INV_X1 U6723 ( .A(n5223), .ZN(n5225) );
  INV_X1 U6724 ( .A(SI_13_), .ZN(n5224) );
  NAND2_X1 U6725 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  OR2_X1 U6726 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  NAND2_X1 U6727 ( .A1(n5244), .A2(n5229), .ZN(n7517) );
  OR2_X1 U6728 ( .A1(n7517), .A2(n5528), .ZN(n5232) );
  OAI21_X1 U6729 ( .B1(n5230), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5247) );
  XNOR2_X1 U6730 ( .A(n5247), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7927) );
  AOI22_X1 U6731 ( .A1(n5312), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5787), .B2(
        n7927), .ZN(n5231) );
  NAND2_X1 U6732 ( .A1(n7404), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5240) );
  INV_X1 U6733 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8355) );
  OR2_X1 U6734 ( .A1(n4339), .A2(n8355), .ZN(n5239) );
  NOR2_X1 U6735 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .ZN(n5233) );
  OAI21_X1 U6736 ( .B1(n5235), .B2(P2_REG3_REG_12__SCAN_IN), .A(
        P2_REG3_REG_13__SCAN_IN), .ZN(n5236) );
  AND2_X1 U6737 ( .A1(n5256), .A2(n5236), .ZN(n8264) );
  OR2_X1 U6738 ( .A1(n4340), .A2(n8264), .ZN(n5238) );
  INV_X1 U6739 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8265) );
  OR2_X1 U6740 ( .A1(n5532), .A2(n8265), .ZN(n5237) );
  NAND4_X1 U6741 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n7879)
         );
  NOR2_X1 U6742 ( .A1(n8260), .A2(n8277), .ZN(n5242) );
  NAND2_X1 U6743 ( .A1(n8260), .A2(n8277), .ZN(n5241) );
  MUX2_X1 U6744 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4338), .Z(n5263) );
  XNOR2_X1 U6745 ( .A(n5263), .B(SI_14_), .ZN(n5245) );
  XNOR2_X1 U6746 ( .A(n5264), .B(n5245), .ZN(n7547) );
  NAND2_X1 U6747 ( .A1(n7547), .A2(n7401), .ZN(n5253) );
  INV_X1 U6748 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6749 ( .A1(n5247), .A2(n5246), .ZN(n5248) );
  NAND2_X1 U6750 ( .A1(n5248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5250) );
  INV_X1 U6751 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6752 ( .A1(n5250), .A2(n5249), .ZN(n5266) );
  OR2_X1 U6753 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  AOI22_X1 U6754 ( .A1(n5312), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5787), .B2(
        n7930), .ZN(n5252) );
  NAND2_X1 U6755 ( .A1(n5253), .A2(n5252), .ZN(n7698) );
  INV_X1 U6756 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8351) );
  OR2_X1 U6757 ( .A1(n4339), .A2(n8351), .ZN(n5261) );
  INV_X1 U6758 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10003) );
  OR2_X1 U6759 ( .A1(n5338), .A2(n10003), .ZN(n5260) );
  INV_X1 U6760 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6761 ( .A1(n5256), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5257) );
  AND2_X1 U6762 ( .A1(n5270), .A2(n5257), .ZN(n8249) );
  OR2_X1 U6763 ( .A1(n5063), .A2(n8249), .ZN(n5259) );
  INV_X1 U6764 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7914) );
  OR2_X1 U6765 ( .A1(n5532), .A2(n7914), .ZN(n5258) );
  NAND4_X1 U6766 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n7878)
         );
  INV_X1 U6767 ( .A(n7878), .ZN(n8259) );
  OR2_X1 U6768 ( .A1(n7698), .A2(n8259), .ZN(n7332) );
  NAND2_X1 U6769 ( .A1(n8252), .A2(n7332), .ZN(n5262) );
  NAND2_X1 U6770 ( .A1(n7698), .A2(n8259), .ZN(n7333) );
  NAND2_X1 U6771 ( .A1(n5262), .A2(n7333), .ZN(n8236) );
  MUX2_X1 U6772 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4338), .Z(n5277) );
  XNOR2_X1 U6773 ( .A(n5277), .B(SI_15_), .ZN(n5265) );
  XNOR2_X1 U6774 ( .A(n5280), .B(n5265), .ZN(n7559) );
  NAND2_X1 U6775 ( .A1(n7559), .A2(n7401), .ZN(n5269) );
  NAND2_X1 U6776 ( .A1(n5266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5267) );
  XNOR2_X1 U6777 ( .A(n5267), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7972) );
  AOI22_X1 U6778 ( .A1(n5312), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7972), .B2(
        n5787), .ZN(n5268) );
  NAND2_X1 U6779 ( .A1(n7404), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5275) );
  INV_X1 U6780 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8242) );
  OR2_X1 U6781 ( .A1(n5532), .A2(n8242), .ZN(n5274) );
  NAND2_X1 U6782 ( .A1(n5270), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5271) );
  AND2_X1 U6783 ( .A1(n5293), .A2(n5271), .ZN(n8241) );
  OR2_X1 U6784 ( .A1(n4340), .A2(n8241), .ZN(n5273) );
  INV_X1 U6785 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10065) );
  OR2_X1 U6786 ( .A1(n4339), .A2(n10065), .ZN(n5272) );
  NAND2_X1 U6787 ( .A1(n8346), .A2(n8248), .ZN(n7340) );
  INV_X1 U6788 ( .A(n7340), .ZN(n5276) );
  INV_X1 U6789 ( .A(n5277), .ZN(n5278) );
  MUX2_X1 U6790 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4338), .Z(n5302) );
  INV_X1 U6791 ( .A(SI_16_), .ZN(n5282) );
  XNOR2_X1 U6792 ( .A(n5302), .B(n5282), .ZN(n5283) );
  XNOR2_X1 U6793 ( .A(n5301), .B(n5283), .ZN(n7513) );
  NAND2_X1 U6794 ( .A1(n7513), .A2(n7401), .ZN(n5290) );
  NAND2_X1 U6795 ( .A1(n5284), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5285) );
  MUX2_X1 U6796 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5285), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5288) );
  INV_X1 U6797 ( .A(n5287), .ZN(n5309) );
  AND2_X1 U6798 ( .A1(n5288), .A2(n5309), .ZN(n7976) );
  AOI22_X1 U6799 ( .A1(n5312), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5787), .B2(
        n7976), .ZN(n5289) );
  NAND2_X1 U6800 ( .A1(n7404), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5298) );
  INV_X1 U6801 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7975) );
  OR2_X1 U6802 ( .A1(n4339), .A2(n7975), .ZN(n5297) );
  INV_X1 U6803 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6804 ( .A1(n5293), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5294) );
  AND2_X1 U6805 ( .A1(n5315), .A2(n5294), .ZN(n8232) );
  OR2_X1 U6806 ( .A1(n5063), .A2(n8232), .ZN(n5296) );
  OR2_X1 U6807 ( .A1(n5532), .A2(n7959), .ZN(n5295) );
  NAND2_X1 U6808 ( .A1(n8411), .A2(n8240), .ZN(n7344) );
  NAND2_X1 U6809 ( .A1(n8229), .A2(n7344), .ZN(n5299) );
  NAND2_X1 U6810 ( .A1(n5299), .A2(n7342), .ZN(n8216) );
  NOR2_X1 U6811 ( .A1(n5302), .A2(SI_16_), .ZN(n5300) );
  NAND2_X1 U6812 ( .A1(n5302), .A2(SI_16_), .ZN(n5303) );
  INV_X1 U6813 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6453) );
  INV_X1 U6814 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5304) );
  MUX2_X1 U6815 ( .A(n6453), .B(n5304), .S(n4338), .Z(n5306) );
  INV_X1 U6816 ( .A(SI_17_), .ZN(n5305) );
  INV_X1 U6817 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U6818 ( .A1(n5307), .A2(SI_17_), .ZN(n5308) );
  NAND2_X1 U6819 ( .A1(n5323), .A2(n5308), .ZN(n5324) );
  XNOR2_X1 U6820 ( .A(n5325), .B(n5324), .ZN(n7498) );
  NAND2_X1 U6821 ( .A1(n7498), .A2(n7401), .ZN(n5314) );
  NAND2_X1 U6822 ( .A1(n5309), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5310) );
  MUX2_X1 U6823 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5310), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5311) );
  NAND2_X1 U6824 ( .A1(n5311), .A2(n4958), .ZN(n8014) );
  INV_X1 U6825 ( .A(n8014), .ZN(n8008) );
  AOI22_X1 U6826 ( .A1(n5312), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5787), .B2(
        n8008), .ZN(n5313) );
  OR2_X2 U6827 ( .A1(n5315), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6828 ( .A1(n5315), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6829 ( .A1(n5336), .A2(n5316), .ZN(n8217) );
  NAND2_X1 U6830 ( .A1(n5515), .A2(n8217), .ZN(n5321) );
  INV_X1 U6831 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7986) );
  OR2_X1 U6832 ( .A1(n4339), .A2(n7986), .ZN(n5320) );
  INV_X1 U6833 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5317) );
  OR2_X1 U6834 ( .A1(n5338), .A2(n5317), .ZN(n5319) );
  INV_X1 U6835 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7988) );
  OR2_X1 U6836 ( .A1(n5532), .A2(n7988), .ZN(n5318) );
  OR2_X1 U6837 ( .A1(n8336), .A2(n8224), .ZN(n7258) );
  NAND2_X1 U6838 ( .A1(n8336), .A2(n8224), .ZN(n7257) );
  NAND2_X1 U6839 ( .A1(n7258), .A2(n7257), .ZN(n8215) );
  OR2_X2 U6840 ( .A1(n8216), .A2(n8215), .ZN(n5322) );
  INV_X1 U6841 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6713) );
  INV_X1 U6842 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5326) );
  MUX2_X1 U6843 ( .A(n6713), .B(n5326), .S(n4338), .Z(n5345) );
  XNOR2_X1 U6844 ( .A(n5345), .B(SI_18_), .ZN(n5343) );
  XNOR2_X1 U6845 ( .A(n5344), .B(n5343), .ZN(n7489) );
  NAND2_X1 U6846 ( .A1(n7489), .A2(n7401), .ZN(n5333) );
  INV_X1 U6847 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U6848 ( .A1(n5329), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5331) );
  AND2_X1 U6849 ( .A1(n5331), .A2(n5330), .ZN(n6711) );
  AOI22_X1 U6850 ( .A1(n5312), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5787), .B2(
        n6711), .ZN(n5332) );
  INV_X1 U6851 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6852 ( .A1(n5336), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6853 ( .A1(n5355), .A2(n5337), .ZN(n8200) );
  NAND2_X1 U6854 ( .A1(n5515), .A2(n8200), .ZN(n5342) );
  INV_X1 U6855 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8405) );
  OR2_X1 U6856 ( .A1(n5338), .A2(n8405), .ZN(n5341) );
  INV_X1 U6857 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8016) );
  OR2_X1 U6858 ( .A1(n5020), .A2(n8016), .ZN(n5340) );
  INV_X1 U6859 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8334) );
  OR2_X1 U6860 ( .A1(n4339), .A2(n8334), .ZN(n5339) );
  NAND4_X1 U6861 ( .A1(n5342), .A2(n5341), .A3(n5340), .A4(n5339), .ZN(n8212)
         );
  NAND2_X1 U6862 ( .A1(n8201), .A2(n8184), .ZN(n7346) );
  INV_X1 U6863 ( .A(n5345), .ZN(n5346) );
  NAND2_X1 U6864 ( .A1(n5346), .A2(SI_18_), .ZN(n5347) );
  INV_X1 U6865 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6817) );
  INV_X1 U6866 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6819) );
  MUX2_X1 U6867 ( .A(n6817), .B(n6819), .S(n4338), .Z(n5350) );
  INV_X1 U6868 ( .A(SI_19_), .ZN(n5349) );
  NAND2_X1 U6869 ( .A1(n5350), .A2(n5349), .ZN(n5361) );
  INV_X1 U6870 ( .A(n5350), .ZN(n5351) );
  NAND2_X1 U6871 ( .A1(n5351), .A2(SI_19_), .ZN(n5352) );
  NAND2_X1 U6872 ( .A1(n5361), .A2(n5352), .ZN(n5362) );
  XNOR2_X1 U6873 ( .A(n5363), .B(n5362), .ZN(n7573) );
  NAND2_X1 U6874 ( .A1(n7573), .A2(n7401), .ZN(n5354) );
  AOI22_X1 U6875 ( .A1(n5312), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5583), .B2(
        n5787), .ZN(n5353) );
  NAND2_X1 U6876 ( .A1(n5355), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6877 ( .A1(n5368), .A2(n5356), .ZN(n8190) );
  NAND2_X1 U6878 ( .A1(n8190), .A2(n5515), .ZN(n5360) );
  NAND2_X1 U6879 ( .A1(n7404), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5359) );
  INV_X1 U6880 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8033) );
  OR2_X1 U6881 ( .A1(n5020), .A2(n8033), .ZN(n5358) );
  INV_X1 U6882 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8329) );
  OR2_X1 U6883 ( .A1(n4339), .A2(n8329), .ZN(n5357) );
  NAND4_X1 U6884 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), .ZN(n7875)
         );
  OR2_X1 U6885 ( .A1(n7715), .A2(n8197), .ZN(n7428) );
  AND2_X1 U6886 ( .A1(n7428), .A2(n8187), .ZN(n7350) );
  NAND2_X1 U6887 ( .A1(n7715), .A2(n8197), .ZN(n7427) );
  INV_X1 U6888 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10075) );
  INV_X1 U6889 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7586) );
  MUX2_X1 U6890 ( .A(n10075), .B(n7586), .S(n4338), .Z(n5373) );
  XNOR2_X1 U6891 ( .A(n5373), .B(SI_20_), .ZN(n5364) );
  XNOR2_X1 U6892 ( .A(n5375), .B(n5364), .ZN(n7585) );
  NAND2_X1 U6893 ( .A1(n7585), .A2(n7401), .ZN(n5366) );
  NAND2_X1 U6894 ( .A1(n5312), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5365) );
  INV_X1 U6895 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U6896 ( .A1(n5368), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6897 ( .A1(n5382), .A2(n5369), .ZN(n8177) );
  NAND2_X1 U6898 ( .A1(n8177), .A2(n5515), .ZN(n5372) );
  AOI22_X1 U6899 ( .A1(n5529), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n7404), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5371) );
  INV_X1 U6900 ( .A(n5020), .ZN(n5587) );
  NAND2_X1 U6901 ( .A1(n5587), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5370) );
  INV_X1 U6902 ( .A(SI_20_), .ZN(n5374) );
  NAND2_X1 U6903 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  MUX2_X1 U6904 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4338), .Z(n5388) );
  INV_X1 U6905 ( .A(SI_21_), .ZN(n5378) );
  XNOR2_X1 U6906 ( .A(n5388), .B(n5378), .ZN(n5379) );
  XNOR2_X1 U6907 ( .A(n5391), .B(n5379), .ZN(n7597) );
  NAND2_X1 U6908 ( .A1(n7597), .A2(n7401), .ZN(n5381) );
  NAND2_X1 U6909 ( .A1(n5312), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6910 ( .A1(n5382), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6911 ( .A1(n5399), .A2(n5383), .ZN(n8166) );
  NAND2_X1 U6912 ( .A1(n8166), .A2(n5515), .ZN(n5386) );
  AOI22_X1 U6913 ( .A1(n5529), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n7404), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n5385) );
  INV_X1 U6914 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n10102) );
  OR2_X1 U6915 ( .A1(n5532), .A2(n10102), .ZN(n5384) );
  NAND2_X1 U6916 ( .A1(n7724), .A2(n8174), .ZN(n7246) );
  NAND2_X1 U6917 ( .A1(n7781), .A2(n8185), .ZN(n8162) );
  AND2_X1 U6918 ( .A1(n7246), .A2(n8162), .ZN(n7253) );
  NAND2_X1 U6919 ( .A1(n8163), .A2(n7253), .ZN(n5387) );
  NOR2_X1 U6920 ( .A1(n5388), .A2(SI_21_), .ZN(n5390) );
  NAND2_X1 U6921 ( .A1(n5388), .A2(SI_21_), .ZN(n5389) );
  INV_X1 U6922 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10083) );
  INV_X1 U6923 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7607) );
  MUX2_X1 U6924 ( .A(n10083), .B(n7607), .S(n4338), .Z(n5393) );
  INV_X1 U6925 ( .A(SI_22_), .ZN(n5392) );
  NAND2_X1 U6926 ( .A1(n5393), .A2(n5392), .ZN(n5407) );
  INV_X1 U6927 ( .A(n5393), .ZN(n5394) );
  NAND2_X1 U6928 ( .A1(n5394), .A2(SI_22_), .ZN(n5395) );
  NAND2_X1 U6929 ( .A1(n5407), .A2(n5395), .ZN(n5408) );
  XNOR2_X1 U6930 ( .A(n5409), .B(n5408), .ZN(n7606) );
  NAND2_X1 U6931 ( .A1(n7606), .A2(n7401), .ZN(n5397) );
  NAND2_X1 U6932 ( .A1(n5492), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5396) );
  INV_X1 U6933 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U6934 ( .A1(n5399), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6935 ( .A1(n5417), .A2(n5400), .ZN(n8144) );
  NAND2_X1 U6936 ( .A1(n8144), .A2(n5515), .ZN(n5406) );
  INV_X1 U6937 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6938 ( .A1(n5529), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6939 ( .A1(n7404), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5401) );
  OAI211_X1 U6940 ( .C1(n5403), .C2(n5532), .A(n5402), .B(n5401), .ZN(n5404)
         );
  INV_X1 U6941 ( .A(n5404), .ZN(n5405) );
  NAND2_X1 U6942 ( .A1(n8316), .A2(n8161), .ZN(n7244) );
  NAND2_X1 U6943 ( .A1(n7249), .A2(n7244), .ZN(n5573) );
  INV_X1 U6944 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5410) );
  INV_X1 U6945 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7619) );
  MUX2_X1 U6946 ( .A(n5410), .B(n7619), .S(n4338), .Z(n5412) );
  INV_X1 U6947 ( .A(SI_23_), .ZN(n5411) );
  NAND2_X1 U6948 ( .A1(n5412), .A2(n5411), .ZN(n5427) );
  INV_X1 U6949 ( .A(n5412), .ZN(n5413) );
  NAND2_X1 U6950 ( .A1(n5413), .A2(SI_23_), .ZN(n5414) );
  XNOR2_X1 U6951 ( .A(n5426), .B(n5425), .ZN(n7618) );
  NAND2_X1 U6952 ( .A1(n7618), .A2(n7401), .ZN(n5416) );
  NAND2_X1 U6953 ( .A1(n5312), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6954 ( .A1(n5417), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6955 ( .A1(n5434), .A2(n5418), .ZN(n8137) );
  NAND2_X1 U6956 ( .A1(n8137), .A2(n5515), .ZN(n5424) );
  INV_X1 U6957 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6958 ( .A1(n7404), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6959 ( .A1(n5529), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5419) );
  OAI211_X1 U6960 ( .C1(n5421), .C2(n5532), .A(n5420), .B(n5419), .ZN(n5422)
         );
  INV_X1 U6961 ( .A(n5422), .ZN(n5423) );
  NAND2_X1 U6962 ( .A1(n5424), .A2(n5423), .ZN(n8150) );
  INV_X1 U6963 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7237) );
  INV_X1 U6964 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7630) );
  MUX2_X1 U6965 ( .A(n7237), .B(n7630), .S(n4338), .Z(n5429) );
  NAND2_X1 U6966 ( .A1(n5429), .A2(n10157), .ZN(n5445) );
  INV_X1 U6967 ( .A(n5429), .ZN(n5430) );
  NAND2_X1 U6968 ( .A1(n5430), .A2(SI_24_), .ZN(n5431) );
  XNOR2_X1 U6969 ( .A(n5444), .B(n5443), .ZN(n7629) );
  NAND2_X1 U6970 ( .A1(n7629), .A2(n7401), .ZN(n5433) );
  NAND2_X1 U6971 ( .A1(n5312), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5432) );
  OR2_X2 U6972 ( .A1(n5434), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6973 ( .A1(n5434), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6974 ( .A1(n5456), .A2(n5435), .ZN(n8124) );
  NAND2_X1 U6975 ( .A1(n8124), .A2(n5515), .ZN(n5441) );
  INV_X1 U6976 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U6977 ( .A1(n7404), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6978 ( .A1(n5529), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5436) );
  OAI211_X1 U6979 ( .C1(n5532), .C2(n5438), .A(n5437), .B(n5436), .ZN(n5439)
         );
  INV_X1 U6980 ( .A(n5439), .ZN(n5440) );
  NAND2_X1 U6981 ( .A1(n7771), .A2(n8134), .ZN(n7361) );
  INV_X1 U6982 ( .A(n8150), .ZN(n7808) );
  NAND2_X1 U6983 ( .A1(n5727), .A2(n7808), .ZN(n8125) );
  NAND2_X1 U6984 ( .A1(n5442), .A2(n7360), .ZN(n8113) );
  INV_X1 U6985 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5447) );
  INV_X1 U6986 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7641) );
  MUX2_X1 U6987 ( .A(n5447), .B(n7641), .S(n4338), .Z(n5449) );
  INV_X1 U6988 ( .A(SI_25_), .ZN(n5448) );
  NAND2_X1 U6989 ( .A1(n5449), .A2(n5448), .ZN(n5467) );
  INV_X1 U6990 ( .A(n5449), .ZN(n5450) );
  NAND2_X1 U6991 ( .A1(n5450), .A2(SI_25_), .ZN(n5451) );
  NAND2_X1 U6992 ( .A1(n7640), .A2(n7401), .ZN(n5453) );
  NAND2_X1 U6993 ( .A1(n5312), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5452) );
  INV_X1 U6994 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U6995 ( .A1(n5456), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U6996 ( .A1(n5476), .A2(n5457), .ZN(n8111) );
  NAND2_X1 U6997 ( .A1(n8111), .A2(n5515), .ZN(n5463) );
  INV_X1 U6998 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6999 ( .A1(n7404), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7000 ( .A1(n5529), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5458) );
  OAI211_X1 U7001 ( .C1(n5460), .C2(n5532), .A(n5459), .B(n5458), .ZN(n5461)
         );
  INV_X1 U7002 ( .A(n5461), .ZN(n5462) );
  NAND2_X1 U7003 ( .A1(n7743), .A2(n5737), .ZN(n7362) );
  NAND2_X1 U7004 ( .A1(n8113), .A2(n7362), .ZN(n5464) );
  OR2_X2 U7005 ( .A1(n7743), .A2(n5737), .ZN(n7358) );
  NAND2_X1 U7006 ( .A1(n5464), .A2(n7358), .ZN(n8098) );
  INV_X1 U7007 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5469) );
  INV_X1 U7008 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7653) );
  MUX2_X1 U7009 ( .A(n5469), .B(n7653), .S(n4338), .Z(n5471) );
  INV_X1 U7010 ( .A(SI_26_), .ZN(n5470) );
  NAND2_X1 U7011 ( .A1(n5471), .A2(n5470), .ZN(n5486) );
  INV_X1 U7012 ( .A(n5471), .ZN(n5472) );
  NAND2_X1 U7013 ( .A1(n5472), .A2(SI_26_), .ZN(n5473) );
  NAND2_X1 U7014 ( .A1(n7652), .A2(n7401), .ZN(n5475) );
  NAND2_X1 U7015 ( .A1(n5492), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U7016 ( .A1(n5476), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U7017 ( .A1(n5495), .A2(n5477), .ZN(n8099) );
  NAND2_X1 U7018 ( .A1(n8099), .A2(n5515), .ZN(n5483) );
  INV_X1 U7019 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U7020 ( .A1(n5529), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U7021 ( .A1(n7404), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5478) );
  OAI211_X1 U7022 ( .C1(n5480), .C2(n5020), .A(n5479), .B(n5478), .ZN(n5481)
         );
  INV_X1 U7023 ( .A(n5481), .ZN(n5482) );
  NOR2_X1 U7024 ( .A1(n8300), .A2(n8109), .ZN(n7364) );
  NAND2_X1 U7025 ( .A1(n8300), .A2(n8109), .ZN(n7363) );
  INV_X1 U7026 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5487) );
  INV_X1 U7027 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7689) );
  MUX2_X1 U7028 ( .A(n5487), .B(n7689), .S(n4338), .Z(n5489) );
  INV_X1 U7029 ( .A(SI_27_), .ZN(n5488) );
  NAND2_X1 U7030 ( .A1(n5489), .A2(n5488), .ZN(n5504) );
  INV_X1 U7031 ( .A(n5489), .ZN(n5490) );
  NAND2_X1 U7032 ( .A1(n5490), .A2(SI_27_), .ZN(n5491) );
  NAND2_X1 U7033 ( .A1(n7688), .A2(n7401), .ZN(n5494) );
  NAND2_X1 U7034 ( .A1(n5492), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7035 ( .A1(n5495), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7036 ( .A1(n5513), .A2(n5496), .ZN(n8087) );
  NAND2_X1 U7037 ( .A1(n8087), .A2(n5515), .ZN(n5501) );
  INV_X1 U7038 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8090) );
  NAND2_X1 U7039 ( .A1(n5529), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7040 ( .A1(n7404), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5497) );
  OAI211_X1 U7041 ( .C1(n8090), .C2(n5020), .A(n5498), .B(n5497), .ZN(n5499)
         );
  INV_X1 U7042 ( .A(n5499), .ZN(n5500) );
  NAND2_X1 U7043 ( .A1(n5579), .A2(n8072), .ZN(n7368) );
  INV_X1 U7044 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5505) );
  INV_X1 U7045 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9749) );
  MUX2_X1 U7046 ( .A(n5505), .B(n9749), .S(n4338), .Z(n5507) );
  INV_X1 U7047 ( .A(SI_28_), .ZN(n5506) );
  NAND2_X1 U7048 ( .A1(n5507), .A2(n5506), .ZN(n5525) );
  INV_X1 U7049 ( .A(n5507), .ZN(n5508) );
  NAND2_X1 U7050 ( .A1(n5508), .A2(SI_28_), .ZN(n5509) );
  AND2_X1 U7051 ( .A1(n5525), .A2(n5509), .ZN(n5523) );
  NAND2_X1 U7052 ( .A1(n8434), .A2(n7401), .ZN(n5511) );
  NAND2_X1 U7053 ( .A1(n5312), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5510) );
  INV_X1 U7054 ( .A(n5513), .ZN(n5512) );
  INV_X1 U7055 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U7056 ( .A1(n5512), .A2(n5774), .ZN(n8054) );
  NAND2_X1 U7057 ( .A1(n5513), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7058 ( .A1(n8054), .A2(n5514), .ZN(n8076) );
  NAND2_X1 U7059 ( .A1(n8076), .A2(n5515), .ZN(n5520) );
  INV_X1 U7060 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U7061 ( .A1(n5529), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7062 ( .A1(n7404), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5516) );
  OAI211_X1 U7063 ( .C1(n10066), .C2(n5532), .A(n5517), .B(n5516), .ZN(n5518)
         );
  INV_X1 U7064 ( .A(n5518), .ZN(n5519) );
  MUX2_X1 U7065 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4338), .Z(n7375) );
  NAND2_X1 U7066 ( .A1(n5312), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5527) );
  INV_X1 U7067 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U7068 ( .A1(n7404), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7069 ( .A1(n5529), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5530) );
  OAI211_X1 U7070 ( .C1(n8063), .C2(n5532), .A(n5531), .B(n5530), .ZN(n5533)
         );
  INV_X1 U7071 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U7072 ( .A1(n8065), .A2(n8073), .ZN(n7382) );
  INV_X1 U7073 ( .A(n8069), .ZN(n5594) );
  NAND2_X1 U7074 ( .A1(n4364), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5535) );
  AND2_X2 U7075 ( .A1(n7472), .A2(n7266), .ZN(n7388) );
  NAND2_X1 U7076 ( .A1(n6938), .A2(n8046), .ZN(n5659) );
  INV_X1 U7077 ( .A(n5659), .ZN(n5536) );
  NAND2_X1 U7078 ( .A1(n7388), .A2(n5536), .ZN(n5771) );
  NAND2_X1 U7079 ( .A1(n5771), .A2(n9947), .ZN(n6771) );
  AOI21_X1 U7080 ( .B1(n7472), .B2(n8046), .A(n5536), .ZN(n5537) );
  NAND2_X1 U7081 ( .A1(n6934), .A2(n6777), .ZN(n6933) );
  NAND2_X1 U7082 ( .A1(n7431), .A2(n6933), .ZN(n6932) );
  NAND2_X1 U7083 ( .A1(n4992), .A2(n9923), .ZN(n5538) );
  NAND2_X1 U7084 ( .A1(n6932), .A2(n5538), .ZN(n6719) );
  NAND2_X1 U7085 ( .A1(n6719), .A2(n7430), .ZN(n5540) );
  NAND2_X1 U7086 ( .A1(n6376), .A2(n9927), .ZN(n5539) );
  NAND2_X1 U7087 ( .A1(n5540), .A2(n5539), .ZN(n6227) );
  NAND2_X1 U7088 ( .A1(n6227), .A2(n7429), .ZN(n5546) );
  AND4_X1 U7089 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .ZN(n6721)
         );
  NAND2_X1 U7090 ( .A1(n6721), .A2(n6952), .ZN(n5545) );
  NAND2_X1 U7091 ( .A1(n5546), .A2(n5545), .ZN(n6940) );
  AND2_X1 U7092 ( .A1(n7887), .A2(n6667), .ZN(n5550) );
  NAND2_X1 U7093 ( .A1(n5682), .A2(n9937), .ZN(n5549) );
  NAND2_X1 U7094 ( .A1(n7280), .A2(n7290), .ZN(n7439) );
  NAND2_X1 U7095 ( .A1(n6811), .A2(n6802), .ZN(n5551) );
  NOR2_X1 U7096 ( .A1(n6960), .A2(n7885), .ZN(n5552) );
  NAND2_X1 U7097 ( .A1(n6960), .A2(n7885), .ZN(n5553) );
  AND2_X1 U7098 ( .A1(n9945), .A2(n7884), .ZN(n5554) );
  OAI22_X1 U7099 ( .A1(n6922), .A2(n5554), .B1(n9945), .B2(n7884), .ZN(n7083)
         );
  NOR2_X1 U7100 ( .A1(n7101), .A2(n7883), .ZN(n5555) );
  NAND2_X1 U7101 ( .A1(n7101), .A2(n7883), .ZN(n5556) );
  AND2_X1 U7102 ( .A1(n7137), .A2(n7882), .ZN(n5558) );
  INV_X1 U7103 ( .A(n8275), .ZN(n7881) );
  OR2_X1 U7104 ( .A1(n9963), .A2(n7880), .ZN(n5559) );
  NOR2_X1 U7105 ( .A1(n8260), .A2(n7879), .ZN(n7451) );
  NAND2_X1 U7106 ( .A1(n8260), .A2(n7879), .ZN(n7449) );
  OR2_X1 U7107 ( .A1(n7698), .A2(n7878), .ZN(n5560) );
  NAND2_X1 U7108 ( .A1(n7698), .A2(n7878), .ZN(n5561) );
  INV_X1 U7109 ( .A(n8248), .ZN(n7877) );
  INV_X1 U7110 ( .A(n8224), .ZN(n7876) );
  NAND2_X1 U7111 ( .A1(n8336), .A2(n7876), .ZN(n5563) );
  INV_X1 U7112 ( .A(n5563), .ZN(n5562) );
  NOR2_X1 U7113 ( .A1(n5562), .A2(n8215), .ZN(n5565) );
  OR2_X1 U7114 ( .A1(n8223), .A2(n5565), .ZN(n5567) );
  INV_X1 U7115 ( .A(n8240), .ZN(n8210) );
  NAND2_X1 U7116 ( .A1(n8411), .A2(n8210), .ZN(n8207) );
  AND2_X1 U7117 ( .A1(n8207), .A2(n5563), .ZN(n5564) );
  OR2_X1 U7118 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  AND2_X1 U7119 ( .A1(n8201), .A2(n8212), .ZN(n5568) );
  NOR2_X1 U7120 ( .A1(n7715), .A2(n7875), .ZN(n5570) );
  NAND2_X1 U7121 ( .A1(n7715), .A2(n7875), .ZN(n5569) );
  NAND2_X1 U7122 ( .A1(n7245), .A2(n8162), .ZN(n7426) );
  INV_X1 U7123 ( .A(n8185), .ZN(n7874) );
  OR2_X1 U7124 ( .A1(n7781), .A2(n7874), .ZN(n8156) );
  NAND2_X1 U7125 ( .A1(n7247), .A2(n7246), .ZN(n8165) );
  INV_X1 U7126 ( .A(n8174), .ZN(n8149) );
  OR2_X1 U7127 ( .A1(n7724), .A2(n8149), .ZN(n8145) );
  NAND2_X1 U7128 ( .A1(n8159), .A2(n8145), .ZN(n5574) );
  OR2_X1 U7129 ( .A1(n8316), .A2(n7873), .ZN(n5575) );
  NAND2_X1 U7130 ( .A1(n5727), .A2(n8150), .ZN(n5576) );
  OR2_X2 U7131 ( .A1(n8116), .A2(n8127), .ZN(n8117) );
  NAND2_X1 U7132 ( .A1(n7771), .A2(n7872), .ZN(n5577) );
  OR2_X1 U7133 ( .A1(n7743), .A2(n8120), .ZN(n5578) );
  INV_X1 U7134 ( .A(n8300), .ZN(n7854) );
  NOR2_X1 U7135 ( .A1(n8377), .A2(n8072), .ZN(n5580) );
  OAI22_X1 U7136 ( .A1(n8082), .A2(n5580), .B1(n8095), .B2(n5579), .ZN(n8070)
         );
  NAND2_X1 U7137 ( .A1(n7472), .A2(n5583), .ZN(n5636) );
  INV_X1 U7138 ( .A(n6938), .ZN(n7421) );
  NAND2_X1 U7139 ( .A1(n7266), .A2(n7421), .ZN(n5584) );
  NAND2_X1 U7140 ( .A1(n5636), .A2(n5584), .ZN(n8214) );
  NAND2_X1 U7141 ( .A1(n5585), .A2(n8214), .ZN(n5593) );
  INV_X1 U7142 ( .A(n6307), .ZN(n7469) );
  INV_X1 U7143 ( .A(n8041), .ZN(n6313) );
  NAND2_X1 U7144 ( .A1(n7469), .A2(n6313), .ZN(n5586) );
  NAND2_X1 U7145 ( .A1(n4448), .A2(n5586), .ZN(n5775) );
  INV_X1 U7146 ( .A(n5775), .ZN(n5772) );
  INV_X1 U7147 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U7148 ( .A1(n5587), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7149 ( .A1(n7404), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5588) );
  OAI211_X1 U7150 ( .C1(n4339), .C2(n10132), .A(n5589), .B(n5588), .ZN(n5590)
         );
  INV_X1 U7151 ( .A(n5590), .ZN(n5591) );
  NAND2_X1 U7152 ( .A1(n7411), .A2(n5591), .ZN(n7868) );
  AOI21_X1 U7153 ( .B1(P2_B_REG_SCAN_IN), .B2(n4448), .A(n8278), .ZN(n8056) );
  AOI22_X1 U7154 ( .A1(n7869), .A2(n8209), .B1(n7868), .B2(n8056), .ZN(n5592)
         );
  OAI211_X1 U7155 ( .C1(n8069), .C2(n7134), .A(n5593), .B(n5592), .ZN(n8061)
         );
  AOI21_X1 U7156 ( .B1(n9952), .B2(n5594), .A(n8061), .ZN(n5653) );
  NAND2_X1 U7157 ( .A1(n5596), .A2(n5595), .ZN(n5601) );
  NAND2_X1 U7158 ( .A1(n5634), .A2(n5635), .ZN(n5597) );
  NAND2_X1 U7159 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  NAND3_X1 U7160 ( .A1(n5605), .A2(n5599), .A3(n5635), .ZN(n5600) );
  OAI21_X1 U7161 ( .B1(n5601), .B2(n5600), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5602) );
  MUX2_X1 U7162 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5602), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5604) );
  NAND2_X1 U7163 ( .A1(n5608), .A2(n5607), .ZN(n5612) );
  INV_X1 U7164 ( .A(P2_B_REG_SCAN_IN), .ZN(n10091) );
  XNOR2_X1 U7165 ( .A(n5612), .B(n10091), .ZN(n5609) );
  NAND2_X1 U7166 ( .A1(n5609), .A2(n7241), .ZN(n5610) );
  NAND2_X1 U7167 ( .A1(n5633), .A2(n5610), .ZN(n5615) );
  INV_X1 U7168 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7169 ( .A1(n5615), .A2(n5611), .ZN(n5614) );
  INV_X1 U7170 ( .A(n7241), .ZN(n5618) );
  NAND2_X1 U7171 ( .A1(n5612), .A2(n5618), .ZN(n5613) );
  INV_X1 U7172 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7173 ( .A1(n5615), .A2(n5616), .ZN(n5621) );
  INV_X1 U7174 ( .A(n5617), .ZN(n5619) );
  NAND2_X1 U7175 ( .A1(n5619), .A2(n5618), .ZN(n5620) );
  NAND2_X1 U7176 ( .A1(n5621), .A2(n5620), .ZN(n6671) );
  OR2_X1 U7177 ( .A1(n5662), .A2(n6671), .ZN(n5648) );
  NOR2_X1 U7178 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5625) );
  NOR4_X1 U7179 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n5624) );
  NOR4_X1 U7180 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5623) );
  NOR4_X1 U7181 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5622) );
  NAND4_X1 U7182 ( .A1(n5625), .A2(n5624), .A3(n5623), .A4(n5622), .ZN(n5631)
         );
  NOR4_X1 U7183 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5629) );
  NOR4_X1 U7184 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5628) );
  NOR4_X1 U7185 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5627) );
  NOR4_X1 U7186 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5626) );
  NAND4_X1 U7187 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), .ZN(n5630)
         );
  OAI21_X1 U7188 ( .B1(n5631), .B2(n5630), .A(n5615), .ZN(n5646) );
  INV_X1 U7189 ( .A(n5646), .ZN(n5632) );
  XNOR2_X1 U7190 ( .A(n5634), .B(n5635), .ZN(n5785) );
  NAND2_X1 U7191 ( .A1(n5784), .A2(n5785), .ZN(n5762) );
  OR2_X1 U7192 ( .A1(n5636), .A2(n7432), .ZN(n5765) );
  NAND2_X1 U7193 ( .A1(n5771), .A2(n5765), .ZN(n5637) );
  NAND2_X1 U7194 ( .A1(n5754), .A2(n5637), .ZN(n5640) );
  AND3_X1 U7195 ( .A1(n5662), .A2(n6671), .A3(n5646), .ZN(n5767) );
  NAND2_X1 U7196 ( .A1(n5767), .A2(n6071), .ZN(n5778) );
  OR2_X1 U7197 ( .A1(n8046), .A2(n6938), .ZN(n5638) );
  OAI211_X1 U7198 ( .C1(n7152), .C2(n5638), .A(n7386), .B(n9947), .ZN(n5750)
         );
  AND2_X1 U7199 ( .A1(n5750), .A2(n8255), .ZN(n5757) );
  OR2_X1 U7200 ( .A1(n5778), .A2(n5757), .ZN(n5639) );
  OR2_X1 U7201 ( .A1(n5653), .A2(n9966), .ZN(n5645) );
  INV_X1 U7202 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5641) );
  NOR2_X1 U7203 ( .A1(n9965), .A2(n5641), .ZN(n5642) );
  NAND2_X1 U7204 ( .A1(n5645), .A2(n5644), .ZN(P2_U3456) );
  NAND2_X1 U7205 ( .A1(n7388), .A2(n5659), .ZN(n5760) );
  NAND2_X1 U7206 ( .A1(n5646), .A2(n5760), .ZN(n5647) );
  NOR2_X1 U7207 ( .A1(n8423), .A2(n5647), .ZN(n5649) );
  INV_X1 U7208 ( .A(n6671), .ZN(n8424) );
  NOR2_X1 U7209 ( .A1(n5662), .A2(n5755), .ZN(n5651) );
  NAND3_X1 U7210 ( .A1(n7472), .A2(n7421), .A3(n8046), .ZN(n5650) );
  MUX2_X1 U7211 ( .A(n8424), .B(n5651), .S(n6670), .Z(n5652) );
  OR2_X1 U7212 ( .A1(n5653), .A2(n10190), .ZN(n5658) );
  INV_X1 U7213 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5654) );
  NOR2_X1 U7214 ( .A1(n10192), .A2(n5654), .ZN(n5655) );
  NAND2_X1 U7215 ( .A1(n5658), .A2(n5657), .ZN(P2_U3488) );
  NAND2_X1 U7216 ( .A1(n7266), .A2(n6938), .ZN(n5660) );
  AND2_X1 U7217 ( .A1(n5660), .A2(n5659), .ZN(n5661) );
  XNOR2_X1 U7218 ( .A(n7698), .B(n5748), .ZN(n5703) );
  INV_X1 U7219 ( .A(n5703), .ZN(n5704) );
  XNOR2_X1 U7220 ( .A(n9948), .B(n5748), .ZN(n7224) );
  XNOR2_X1 U7221 ( .A(n7141), .B(n5725), .ZN(n7817) );
  XNOR2_X1 U7222 ( .A(n5666), .B(n6380), .ZN(n5664) );
  INV_X1 U7223 ( .A(n5664), .ZN(n5663) );
  NAND2_X1 U7224 ( .A1(n5663), .A2(n7891), .ZN(n5665) );
  NAND2_X1 U7225 ( .A1(n5664), .A2(n4992), .ZN(n5670) );
  NAND2_X1 U7226 ( .A1(n5665), .A2(n5670), .ZN(n6373) );
  INV_X1 U7227 ( .A(n6373), .ZN(n5669) );
  OR2_X1 U7228 ( .A1(n4336), .A2(n6777), .ZN(n5667) );
  XNOR2_X1 U7229 ( .A(n5671), .B(n6376), .ZN(n6253) );
  NAND2_X1 U7230 ( .A1(n6252), .A2(n6253), .ZN(n6251) );
  INV_X1 U7231 ( .A(n5671), .ZN(n5672) );
  NAND2_X1 U7232 ( .A1(n5672), .A2(n6376), .ZN(n5673) );
  XNOR2_X1 U7233 ( .A(n4336), .B(n6952), .ZN(n5674) );
  XNOR2_X1 U7234 ( .A(n5674), .B(n6721), .ZN(n6287) );
  NAND2_X1 U7235 ( .A1(n5674), .A2(n7889), .ZN(n5675) );
  XNOR2_X1 U7236 ( .A(n4336), .B(n9931), .ZN(n5676) );
  NAND2_X1 U7237 ( .A1(n5676), .A2(n6678), .ZN(n6704) );
  INV_X1 U7238 ( .A(n5676), .ZN(n5677) );
  NAND2_X1 U7239 ( .A1(n5677), .A2(n7888), .ZN(n5678) );
  NAND2_X1 U7240 ( .A1(n6704), .A2(n5678), .ZN(n6444) );
  NAND2_X1 U7241 ( .A1(n6442), .A2(n6704), .ZN(n5680) );
  XNOR2_X1 U7242 ( .A(n5748), .B(n9937), .ZN(n5681) );
  XNOR2_X1 U7243 ( .A(n5681), .B(n5682), .ZN(n6703) );
  NAND2_X1 U7244 ( .A1(n5680), .A2(n6703), .ZN(n6702) );
  INV_X1 U7245 ( .A(n5681), .ZN(n5683) );
  NAND2_X1 U7246 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  XNOR2_X1 U7247 ( .A(n5748), .B(n6802), .ZN(n5685) );
  XNOR2_X1 U7248 ( .A(n5685), .B(n6811), .ZN(n6727) );
  NAND2_X1 U7249 ( .A1(n5685), .A2(n7886), .ZN(n5686) );
  NAND2_X1 U7250 ( .A1(n6726), .A2(n5686), .ZN(n6903) );
  XNOR2_X1 U7251 ( .A(n5748), .B(n6960), .ZN(n5687) );
  NAND2_X1 U7252 ( .A1(n5687), .A2(n6924), .ZN(n6992) );
  INV_X1 U7253 ( .A(n5687), .ZN(n5688) );
  NAND2_X1 U7254 ( .A1(n5688), .A2(n7885), .ZN(n5689) );
  NAND2_X1 U7255 ( .A1(n6992), .A2(n5689), .ZN(n6902) );
  XNOR2_X1 U7256 ( .A(n5748), .B(n9945), .ZN(n5690) );
  NAND2_X1 U7257 ( .A1(n5690), .A2(n7085), .ZN(n5691) );
  XNOR2_X1 U7258 ( .A(n7101), .B(n5748), .ZN(n5692) );
  XNOR2_X1 U7259 ( .A(n5692), .B(n7883), .ZN(n7025) );
  INV_X1 U7260 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U7261 ( .A1(n5693), .A2(n7883), .ZN(n5694) );
  NOR3_X1 U7262 ( .A1(n9948), .A2(n5725), .A3(n7882), .ZN(n5695) );
  INV_X1 U7263 ( .A(n7141), .ZN(n7448) );
  AOI211_X1 U7264 ( .C1(n8275), .C2(n5725), .A(n5695), .B(n7448), .ZN(n5698)
         );
  NOR3_X1 U7265 ( .A1(n7137), .A2(n7882), .A3(n5748), .ZN(n5696) );
  AOI211_X1 U7266 ( .C1(n8275), .C2(n5748), .A(n5696), .B(n7141), .ZN(n5697)
         );
  XNOR2_X1 U7267 ( .A(n9963), .B(n5748), .ZN(n5699) );
  XNOR2_X1 U7268 ( .A(n5699), .B(n7880), .ZN(n7736) );
  OAI21_X1 U7269 ( .B1(n5698), .B2(n5697), .A(n7736), .ZN(n5700) );
  XNOR2_X1 U7270 ( .A(n8260), .B(n5748), .ZN(n5701) );
  NAND2_X1 U7271 ( .A1(n5701), .A2(n8277), .ZN(n5702) );
  OAI21_X1 U7272 ( .B1(n5701), .B2(n8277), .A(n5702), .ZN(n7792) );
  INV_X1 U7273 ( .A(n5702), .ZN(n7702) );
  XNOR2_X1 U7274 ( .A(n5703), .B(n7878), .ZN(n7701) );
  XNOR2_X1 U7275 ( .A(n8346), .B(n5748), .ZN(n5705) );
  XNOR2_X1 U7276 ( .A(n5705), .B(n8248), .ZN(n7863) );
  INV_X1 U7277 ( .A(n5705), .ZN(n5706) );
  XNOR2_X1 U7278 ( .A(n8411), .B(n5748), .ZN(n5707) );
  NAND2_X1 U7279 ( .A1(n5707), .A2(n8240), .ZN(n5708) );
  OAI21_X1 U7280 ( .B1(n5707), .B2(n8240), .A(n5708), .ZN(n7754) );
  INV_X1 U7281 ( .A(n5708), .ZN(n7763) );
  XNOR2_X1 U7282 ( .A(n8336), .B(n5748), .ZN(n5709) );
  NAND2_X1 U7283 ( .A1(n5709), .A2(n8224), .ZN(n7832) );
  INV_X1 U7284 ( .A(n5709), .ZN(n5710) );
  NAND2_X1 U7285 ( .A1(n5710), .A2(n7876), .ZN(n5711) );
  XNOR2_X1 U7286 ( .A(n8201), .B(n5748), .ZN(n5712) );
  NAND2_X1 U7287 ( .A1(n5712), .A2(n8184), .ZN(n5715) );
  INV_X1 U7288 ( .A(n5712), .ZN(n5713) );
  NAND2_X1 U7289 ( .A1(n5713), .A2(n8212), .ZN(n5714) );
  NAND2_X1 U7290 ( .A1(n5715), .A2(n5714), .ZN(n7831) );
  INV_X1 U7291 ( .A(n5715), .ZN(n7717) );
  XNOR2_X1 U7292 ( .A(n7715), .B(n5748), .ZN(n5716) );
  NAND2_X1 U7293 ( .A1(n5716), .A2(n8197), .ZN(n7783) );
  INV_X1 U7294 ( .A(n5716), .ZN(n5717) );
  NAND2_X1 U7295 ( .A1(n5717), .A2(n7875), .ZN(n5718) );
  XNOR2_X1 U7296 ( .A(n7781), .B(n5748), .ZN(n5719) );
  NAND2_X1 U7297 ( .A1(n5719), .A2(n8185), .ZN(n5722) );
  INV_X1 U7298 ( .A(n5719), .ZN(n5720) );
  NAND2_X1 U7299 ( .A1(n5720), .A2(n7874), .ZN(n5721) );
  NAND2_X1 U7300 ( .A1(n5722), .A2(n5721), .ZN(n7782) );
  INV_X1 U7301 ( .A(n5722), .ZN(n7727) );
  XNOR2_X1 U7302 ( .A(n7724), .B(n5748), .ZN(n5723) );
  XNOR2_X1 U7303 ( .A(n5723), .B(n8149), .ZN(n7726) );
  NAND2_X1 U7304 ( .A1(n5723), .A2(n8174), .ZN(n5724) );
  NAND2_X1 U7305 ( .A1(n7801), .A2(n7873), .ZN(n7806) );
  XNOR2_X1 U7306 ( .A(n5727), .B(n5748), .ZN(n5730) );
  INV_X1 U7307 ( .A(n5730), .ZN(n5728) );
  XNOR2_X1 U7308 ( .A(n7771), .B(n5748), .ZN(n5733) );
  NAND2_X1 U7309 ( .A1(n5733), .A2(n8134), .ZN(n7745) );
  INV_X1 U7310 ( .A(n5733), .ZN(n5734) );
  NAND2_X1 U7311 ( .A1(n5734), .A2(n7872), .ZN(n5735) );
  NAND2_X1 U7312 ( .A1(n5736), .A2(n7773), .ZN(n7744) );
  NAND2_X1 U7313 ( .A1(n7744), .A2(n7745), .ZN(n5741) );
  XNOR2_X1 U7314 ( .A(n7743), .B(n5748), .ZN(n5738) );
  NAND2_X1 U7315 ( .A1(n5738), .A2(n5737), .ZN(n7840) );
  INV_X1 U7316 ( .A(n5738), .ZN(n5739) );
  NAND2_X1 U7317 ( .A1(n5739), .A2(n8120), .ZN(n5740) );
  NAND2_X1 U7318 ( .A1(n5741), .A2(n7746), .ZN(n7748) );
  NAND2_X1 U7319 ( .A1(n7748), .A2(n7840), .ZN(n5742) );
  XNOR2_X1 U7320 ( .A(n8300), .B(n5748), .ZN(n5743) );
  XNOR2_X1 U7321 ( .A(n5743), .B(n7870), .ZN(n7841) );
  NAND2_X1 U7322 ( .A1(n7844), .A2(n5744), .ZN(n7691) );
  INV_X1 U7323 ( .A(n7691), .ZN(n5746) );
  XNOR2_X1 U7324 ( .A(n8377), .B(n5748), .ZN(n5747) );
  XNOR2_X1 U7325 ( .A(n5747), .B(n8095), .ZN(n7690) );
  INV_X1 U7326 ( .A(n7690), .ZN(n5745) );
  XOR2_X1 U7327 ( .A(n5748), .B(n8074), .Z(n5749) );
  INV_X1 U7328 ( .A(n5750), .ZN(n5751) );
  NAND2_X1 U7329 ( .A1(n5754), .A2(n5751), .ZN(n5753) );
  OR2_X1 U7330 ( .A1(n5778), .A2(n5765), .ZN(n5752) );
  NAND2_X1 U7331 ( .A1(n5754), .A2(n9964), .ZN(n5756) );
  INV_X1 U7332 ( .A(n5757), .ZN(n5758) );
  NAND2_X1 U7333 ( .A1(n5759), .A2(n5758), .ZN(n5764) );
  INV_X1 U7334 ( .A(n5760), .ZN(n5761) );
  NOR2_X1 U7335 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  OAI211_X1 U7336 ( .C1(n5767), .C2(n5765), .A(n5764), .B(n5763), .ZN(n5766)
         );
  NAND2_X1 U7337 ( .A1(n5766), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5770) );
  INV_X1 U7338 ( .A(n5767), .ZN(n5768) );
  NOR2_X1 U7339 ( .A1(n8423), .A2(n5771), .ZN(n7470) );
  NAND2_X1 U7340 ( .A1(n5768), .A2(n7470), .ZN(n5769) );
  INV_X1 U7341 ( .A(n5771), .ZN(n5776) );
  NAND2_X1 U7342 ( .A1(n5776), .A2(n5772), .ZN(n5773) );
  OAI22_X1 U7343 ( .A1(n8072), .A2(n7810), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5774), .ZN(n5780) );
  NAND2_X1 U7344 ( .A1(n5776), .A2(n5775), .ZN(n5777) );
  NOR2_X1 U7345 ( .A1(n8073), .A2(n7855), .ZN(n5779) );
  AOI211_X1 U7346 ( .C1(n8076), .C2(n7850), .A(n5780), .B(n5779), .ZN(n5781)
         );
  INV_X1 U7347 ( .A(n5785), .ZN(n7185) );
  NAND2_X1 U7348 ( .A1(n5785), .A2(n7388), .ZN(n5786) );
  NAND2_X1 U7349 ( .A1(n6304), .A2(n5786), .ZN(n6312) );
  OAI21_X1 U7350 ( .B1(n6312), .B2(n5787), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  NOR2_X1 U7351 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5791) );
  AND4_X2 U7352 ( .A1(n5791), .A2(n5790), .A3(n5789), .A4(n5788), .ZN(n5792)
         );
  INV_X1 U7353 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5794) );
  INV_X1 U7354 ( .A(n6294), .ZN(n5795) );
  NOR2_X1 U7355 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5963) );
  NAND2_X1 U7356 ( .A1(n5840), .A2(n5839), .ZN(n5796) );
  NAND2_X1 U7357 ( .A1(n5796), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5797) );
  XNOR2_X1 U7358 ( .A(n5797), .B(P1_IR_REG_23__SCAN_IN), .ZN(n5844) );
  INV_X1 U7359 ( .A(n5844), .ZN(n5798) );
  NOR2_X1 U7360 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5800) );
  NAND4_X1 U7361 ( .A1(n5800), .A2(n5799), .A3(n5839), .A4(n10063), .ZN(n5805)
         );
  INV_X1 U7362 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5802) );
  INV_X1 U7363 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5801) );
  NAND4_X1 U7364 ( .A1(n5973), .A2(n5803), .A3(n5802), .A4(n5801), .ZN(n5804)
         );
  INV_X1 U7365 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U7366 ( .A1(n5810), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5812) );
  INV_X1 U7367 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5811) );
  XNOR2_X1 U7368 ( .A(n5812), .B(n5811), .ZN(n7240) );
  NAND2_X1 U7369 ( .A1(n5813), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5814) );
  MUX2_X1 U7370 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5814), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5815) );
  NAND2_X1 U7371 ( .A1(n5815), .A2(n5810), .ZN(n7234) );
  OR3_X2 U7372 ( .A1(n7477), .A2(n7240), .A3(n7234), .ZN(n5995) );
  INV_X1 U7373 ( .A(n5995), .ZN(n5985) );
  AND2_X2 U7374 ( .A1(n6000), .A2(n5985), .ZN(P1_U3973) );
  AND2_X1 U7375 ( .A1(n4338), .A2(P1_U3086), .ZN(n7188) );
  INV_X2 U7376 ( .A(n7188), .ZN(n9747) );
  NOR2_X1 U7377 ( .A1(n4338), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9740) );
  INV_X1 U7378 ( .A(n9740), .ZN(n9750) );
  INV_X1 U7379 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6095) );
  OR2_X1 U7380 ( .A1(n5816), .A2(n9738), .ZN(n5825) );
  INV_X1 U7381 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5819) );
  XNOR2_X1 U7382 ( .A(n5825), .B(n5819), .ZN(n6099) );
  OAI222_X1 U7383 ( .A1(n9747), .A2(n6096), .B1(n9750), .B2(n6095), .C1(
        P1_U3086), .C2(n6099), .ZN(P1_U3353) );
  INV_X1 U7384 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7385 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5817) );
  XNOR2_X1 U7386 ( .A(n5818), .B(n5817), .ZN(n9147) );
  OAI222_X1 U7387 ( .A1(n9747), .A2(n6051), .B1(n9750), .B2(n4933), .C1(
        P1_U3086), .C2(n9147), .ZN(P1_U3354) );
  INV_X1 U7388 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7389 ( .A1(n5825), .A2(n5819), .ZN(n5820) );
  NAND2_X1 U7390 ( .A1(n5820), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5822) );
  INV_X1 U7391 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5821) );
  XNOR2_X1 U7392 ( .A(n5822), .B(n5821), .ZN(n9157) );
  OAI222_X1 U7393 ( .A1(n9750), .A2(n6130), .B1(n9747), .B2(n4826), .C1(n9157), 
        .C2(P1_U3086), .ZN(P1_U3352) );
  INV_X1 U7394 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6163) );
  INV_X1 U7395 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9738) );
  OR2_X1 U7396 ( .A1(n5823), .A2(n9738), .ZN(n5824) );
  NAND2_X1 U7397 ( .A1(n5825), .A2(n5824), .ZN(n5827) );
  XNOR2_X1 U7398 ( .A(n5827), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9175) );
  OAI222_X1 U7399 ( .A1(n9750), .A2(n6163), .B1(P1_U3086), .B2(n9175), .C1(
        n6162), .C2(n9747), .ZN(P1_U3351) );
  INV_X1 U7400 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5826) );
  AND2_X1 U7401 ( .A1(n4338), .A2(P2_U3151), .ZN(n8438) );
  INV_X1 U7402 ( .A(n8438), .ZN(n7236) );
  OAI222_X1 U7403 ( .A1(P2_U3151), .A2(n9835), .B1(n7151), .B2(n6162), .C1(
        n5826), .C2(n7236), .ZN(P2_U3291) );
  OAI21_X1 U7404 ( .B1(n5827), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5828) );
  XNOR2_X1 U7405 ( .A(n5828), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9191) );
  AOI22_X1 U7406 ( .A1(n9191), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9740), .ZN(n5829) );
  OAI21_X1 U7407 ( .B1(n6262), .B2(n9747), .A(n5829), .ZN(P1_U3350) );
  OAI222_X1 U7408 ( .A1(P2_U3151), .A2(n9858), .B1(n7151), .B2(n6262), .C1(
        n4435), .C2(n7236), .ZN(P2_U3290) );
  NAND2_X1 U7409 ( .A1(n5830), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5831) );
  MUX2_X1 U7410 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5831), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5832) );
  OR2_X1 U7411 ( .A1(n5830), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5853) );
  AND2_X1 U7412 ( .A1(n5832), .A2(n5853), .ZN(n9204) );
  AOI22_X1 U7413 ( .A1(n9204), .A2(P1_STATE_REG_SCAN_IN), .B1(n9740), .B2(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n5833) );
  OAI21_X1 U7414 ( .B1(n6478), .B2(n9747), .A(n5833), .ZN(P1_U3349) );
  AOI22_X1 U7415 ( .A1(n8438), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n6573), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n5834) );
  OAI21_X1 U7416 ( .B1(n6051), .B2(n7151), .A(n5834), .ZN(P2_U3294) );
  INV_X1 U7417 ( .A(n6644), .ZN(n6634) );
  INV_X1 U7418 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5835) );
  OAI222_X1 U7419 ( .A1(P2_U3151), .A2(n6634), .B1(n7151), .B2(n6478), .C1(
        n5835), .C2(n7236), .ZN(P2_U3289) );
  INV_X1 U7420 ( .A(n9825), .ZN(n6302) );
  OAI222_X1 U7421 ( .A1(P2_U3151), .A2(n6302), .B1(n7151), .B2(n6096), .C1(
        n4437), .C2(n7236), .ZN(P2_U3293) );
  INV_X1 U7422 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5836) );
  OAI222_X1 U7423 ( .A1(P2_U3151), .A2(n4335), .B1(n7151), .B2(n4826), .C1(
        n5836), .C2(n7236), .ZN(P2_U3292) );
  NAND2_X1 U7424 ( .A1(n5853), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5837) );
  XNOR2_X1 U7425 ( .A(n5837), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9219) );
  AOI22_X1 U7426 ( .A1(n9219), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9740), .ZN(n5838) );
  OAI21_X1 U7427 ( .B1(n6511), .B2(n9747), .A(n5838), .ZN(P1_U3348) );
  INV_X1 U7428 ( .A(n6647), .ZN(n9876) );
  OAI222_X1 U7429 ( .A1(P2_U3151), .A2(n9876), .B1(n7151), .B2(n6511), .C1(
        n4465), .C2(n7236), .ZN(P2_U3288) );
  AND2_X1 U7430 ( .A1(n6000), .A2(n5995), .ZN(n9106) );
  NAND2_X1 U7431 ( .A1(n5844), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9108) );
  INV_X1 U7432 ( .A(n9108), .ZN(n9040) );
  OR2_X1 U7433 ( .A1(n9106), .A2(n9040), .ZN(n5885) );
  INV_X1 U7434 ( .A(n5841), .ZN(n5842) );
  NAND2_X1 U7435 ( .A1(n9109), .A2(n9025), .ZN(n8902) );
  OR2_X1 U7436 ( .A1(n5844), .A2(n8902), .ZN(n5851) );
  INV_X1 U7437 ( .A(n5860), .ZN(n5857) );
  NAND2_X1 U7438 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n5848) );
  AND2_X1 U7439 ( .A1(n5851), .A2(n4341), .ZN(n5884) );
  INV_X1 U7440 ( .A(n5884), .ZN(n5852) );
  NAND2_X1 U7441 ( .A1(n5885), .A2(n5852), .ZN(n9788) );
  INV_X1 U7442 ( .A(n9788), .ZN(n9230) );
  NOR2_X1 U7443 ( .A1(n9230), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U7444 ( .A(n6737), .ZN(n5856) );
  NOR2_X1 U7445 ( .A1(n5853), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5874) );
  OR2_X1 U7446 ( .A1(n5874), .A2(n9738), .ZN(n5879) );
  XNOR2_X1 U7447 ( .A(n5879), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9231) );
  AOI22_X1 U7448 ( .A1(n9231), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9740), .ZN(n5854) );
  OAI21_X1 U7449 ( .B1(n5856), .B2(n9747), .A(n5854), .ZN(P1_U3347) );
  INV_X1 U7450 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5855) );
  OAI222_X1 U7451 ( .A1(n4499), .A2(P2_U3151), .B1(n7151), .B2(n5856), .C1(
        n5855), .C2(n7236), .ZN(P2_U3287) );
  NAND2_X1 U7452 ( .A1(n5857), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5858) );
  MUX2_X1 U7453 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5858), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5861) );
  NAND2_X1 U7454 ( .A1(n5860), .A2(n5859), .ZN(n5862) );
  INV_X1 U7455 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5863) );
  INV_X1 U7456 ( .A(n5865), .ZN(n5867) );
  NAND2_X1 U7457 ( .A1(n4940), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7458 ( .A1(n7591), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5870) );
  INV_X1 U7459 ( .A(n7487), .ZN(n6062) );
  NAND2_X1 U7460 ( .A1(n6062), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7461 ( .A1(n6113), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7462 ( .A1(n6385), .A2(P1_U3973), .ZN(n5872) );
  OAI21_X1 U7463 ( .B1(P1_U3973), .B2(n4983), .A(n5872), .ZN(P1_U3554) );
  NOR2_X1 U7464 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5873) );
  NAND2_X1 U7465 ( .A1(n5874), .A2(n5873), .ZN(n5918) );
  NAND2_X1 U7466 ( .A1(n5918), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5875) );
  XNOR2_X1 U7467 ( .A(n5875), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6872) );
  AOI22_X1 U7468 ( .A1(n6872), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9740), .ZN(n5876) );
  OAI21_X1 U7469 ( .B1(n6871), .B2(n9747), .A(n5876), .ZN(P1_U3345) );
  INV_X1 U7470 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5877) );
  OAI222_X1 U7471 ( .A1(P2_U3151), .A2(n7170), .B1(n7151), .B2(n6871), .C1(
        n5877), .C2(n7236), .ZN(P2_U3285) );
  INV_X1 U7472 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10007) );
  INV_X1 U7473 ( .A(n6833), .ZN(n5883) );
  INV_X1 U7474 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7475 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  NAND2_X1 U7476 ( .A1(n5880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5881) );
  XNOR2_X1 U7477 ( .A(n5881), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6834) );
  INV_X1 U7478 ( .A(n6834), .ZN(n9766) );
  OAI222_X1 U7479 ( .A1(n9750), .A2(n10007), .B1(n9747), .B2(n5883), .C1(n9766), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U7480 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5882) );
  OAI222_X1 U7481 ( .A1(P2_U3151), .A2(n4505), .B1(n7151), .B2(n5883), .C1(
        n5882), .C2(n7236), .ZN(P2_U3286) );
  AND2_X1 U7482 ( .A1(n5885), .A2(n5884), .ZN(n5939) );
  INV_X1 U7483 ( .A(n9748), .ZN(n6028) );
  OAI21_X1 U7484 ( .B1(n9257), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6028), .ZN(
        n6030) );
  INV_X1 U7485 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9150) );
  AOI21_X1 U7486 ( .B1(n9257), .B2(n9150), .A(n6030), .ZN(n5887) );
  INV_X1 U7487 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9149) );
  MUX2_X1 U7488 ( .A(n6030), .B(n5887), .S(n9149), .Z(n5890) );
  INV_X1 U7489 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n5888) );
  INV_X1 U7490 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6469) );
  OAI22_X1 U7491 ( .A1(n9788), .A2(n5888), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6469), .ZN(n5889) );
  AOI21_X1 U7492 ( .B1(n5939), .B2(n5890), .A(n5889), .ZN(n5892) );
  NAND3_X1 U7493 ( .A1(n9779), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9150), .ZN(
        n5891) );
  NAND2_X1 U7494 ( .A1(n5892), .A2(n5891), .ZN(P1_U3243) );
  INV_X1 U7495 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5893) );
  MUX2_X1 U7496 ( .A(n5893), .B(P1_REG1_REG_2__SCAN_IN), .S(n6099), .Z(n6019)
         );
  INV_X1 U7497 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5894) );
  MUX2_X1 U7498 ( .A(n5894), .B(P1_REG1_REG_1__SCAN_IN), .S(n9147), .Z(n5896)
         );
  AND2_X1 U7499 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n5895) );
  NAND2_X1 U7500 ( .A1(n5896), .A2(n5895), .ZN(n9152) );
  INV_X1 U7501 ( .A(n9147), .ZN(n9143) );
  NAND2_X1 U7502 ( .A1(n9143), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7503 ( .A1(n9152), .A2(n5897), .ZN(n6018) );
  NAND2_X1 U7504 ( .A1(n6019), .A2(n6018), .ZN(n5899) );
  INV_X1 U7505 ( .A(n6099), .ZN(n6027) );
  NAND2_X1 U7506 ( .A1(n6027), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7507 ( .A1(n5899), .A2(n5898), .ZN(n9163) );
  INV_X1 U7508 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5900) );
  MUX2_X1 U7509 ( .A(n5900), .B(P1_REG1_REG_3__SCAN_IN), .S(n9157), .Z(n9164)
         );
  NAND2_X1 U7510 ( .A1(n9163), .A2(n9164), .ZN(n9179) );
  INV_X1 U7511 ( .A(n9157), .ZN(n5923) );
  NAND2_X1 U7512 ( .A1(n5923), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U7513 ( .A1(n9179), .A2(n9178), .ZN(n5902) );
  MUX2_X1 U7514 ( .A(n9176), .B(P1_REG1_REG_4__SCAN_IN), .S(n9175), .Z(n5901)
         );
  NAND2_X1 U7515 ( .A1(n5902), .A2(n5901), .ZN(n9194) );
  INV_X1 U7516 ( .A(n9175), .ZN(n9171) );
  NAND2_X1 U7517 ( .A1(n9171), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U7518 ( .A1(n9194), .A2(n9193), .ZN(n5905) );
  INV_X1 U7519 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5903) );
  MUX2_X1 U7520 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n5903), .S(n9191), .Z(n5904)
         );
  NAND2_X1 U7521 ( .A1(n5905), .A2(n5904), .ZN(n9207) );
  NAND2_X1 U7522 ( .A1(n9191), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9206) );
  NAND2_X1 U7523 ( .A1(n9207), .A2(n9206), .ZN(n5908) );
  INV_X1 U7524 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5906) );
  MUX2_X1 U7525 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n5906), .S(n9204), .Z(n5907)
         );
  NAND2_X1 U7526 ( .A1(n5908), .A2(n5907), .ZN(n9222) );
  NAND2_X1 U7527 ( .A1(n9204), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U7528 ( .A1(n9222), .A2(n9221), .ZN(n5911) );
  INV_X1 U7529 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5909) );
  MUX2_X1 U7530 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n5909), .S(n9219), .Z(n5910)
         );
  NAND2_X1 U7531 ( .A1(n5911), .A2(n5910), .ZN(n9234) );
  NAND2_X1 U7532 ( .A1(n9219), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U7533 ( .A1(n9234), .A2(n9233), .ZN(n5914) );
  INV_X1 U7534 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5912) );
  MUX2_X1 U7535 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n5912), .S(n9231), .Z(n5913)
         );
  NAND2_X1 U7536 ( .A1(n5914), .A2(n5913), .ZN(n9236) );
  NAND2_X1 U7537 ( .A1(n9231), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7538 ( .A1(n9236), .A2(n5915), .ZN(n9760) );
  INV_X1 U7539 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5916) );
  MUX2_X1 U7540 ( .A(n5916), .B(P1_REG1_REG_9__SCAN_IN), .S(n6834), .Z(n9759)
         );
  OAI21_X1 U7541 ( .B1(n6834), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9762), .ZN(
        n6040) );
  INV_X1 U7542 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5917) );
  MUX2_X1 U7543 ( .A(n5917), .B(P1_REG1_REG_10__SCAN_IN), .S(n6872), .Z(n6039)
         );
  NOR2_X1 U7544 ( .A1(n6040), .A2(n6039), .ZN(n6038) );
  AOI21_X1 U7545 ( .B1(n6872), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6038), .ZN(
        n6076) );
  NAND2_X1 U7546 ( .A1(n6011), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5919) );
  XNOR2_X1 U7547 ( .A(n5919), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7528) );
  XNOR2_X1 U7548 ( .A(n7528), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n6075) );
  XNOR2_X1 U7549 ( .A(n6076), .B(n6075), .ZN(n5945) );
  INV_X1 U7550 ( .A(n9779), .ZN(n7196) );
  NAND2_X1 U7551 ( .A1(n5939), .A2(n9748), .ZN(n9767) );
  INV_X1 U7552 ( .A(n9767), .ZN(n9781) );
  INV_X1 U7553 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n5920) );
  OR2_X1 U7554 ( .A1(n10078), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8782) );
  OAI21_X1 U7555 ( .B1(n9788), .B2(n5920), .A(n8782), .ZN(n5943) );
  XNOR2_X1 U7556 ( .A(n6099), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6022) );
  XNOR2_X1 U7557 ( .A(n9147), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9146) );
  AND2_X1 U7558 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9145) );
  NAND2_X1 U7559 ( .A1(n9146), .A2(n9145), .ZN(n9144) );
  NAND2_X1 U7560 ( .A1(n9143), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7561 ( .A1(n9144), .A2(n5921), .ZN(n6021) );
  NAND2_X1 U7562 ( .A1(n6022), .A2(n6021), .ZN(n6020) );
  NAND2_X1 U7563 ( .A1(n6027), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7564 ( .A1(n6020), .A2(n5922), .ZN(n9161) );
  XNOR2_X1 U7565 ( .A(n9157), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U7566 ( .A1(n9161), .A2(n9162), .ZN(n9160) );
  NAND2_X1 U7567 ( .A1(n5923), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7568 ( .A1(n9160), .A2(n5924), .ZN(n9173) );
  INV_X1 U7569 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5925) );
  MUX2_X1 U7570 ( .A(n5925), .B(P1_REG2_REG_4__SCAN_IN), .S(n9175), .Z(n9174)
         );
  NAND2_X1 U7571 ( .A1(n9173), .A2(n9174), .ZN(n9172) );
  NAND2_X1 U7572 ( .A1(n9171), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7573 ( .A1(n9172), .A2(n5926), .ZN(n9189) );
  INV_X1 U7574 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5927) );
  XNOR2_X1 U7575 ( .A(n9191), .B(n5927), .ZN(n9190) );
  NAND2_X1 U7576 ( .A1(n9189), .A2(n9190), .ZN(n9188) );
  NAND2_X1 U7577 ( .A1(n9191), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7578 ( .A1(n9188), .A2(n5928), .ZN(n9200) );
  INV_X1 U7579 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6603) );
  MUX2_X1 U7580 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6603), .S(n9204), .Z(n9201)
         );
  NAND2_X1 U7581 ( .A1(n9200), .A2(n9201), .ZN(n9199) );
  NAND2_X1 U7582 ( .A1(n9204), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7583 ( .A1(n9199), .A2(n5929), .ZN(n9217) );
  INV_X1 U7584 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U7585 ( .A(n9219), .B(n5930), .ZN(n9218) );
  NAND2_X1 U7586 ( .A1(n9217), .A2(n9218), .ZN(n9216) );
  NAND2_X1 U7587 ( .A1(n9219), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7588 ( .A1(n9216), .A2(n5931), .ZN(n9227) );
  INV_X1 U7589 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5932) );
  MUX2_X1 U7590 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n5932), .S(n9231), .Z(n9228)
         );
  NAND2_X1 U7591 ( .A1(n9227), .A2(n9228), .ZN(n9756) );
  INV_X1 U7592 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5933) );
  XNOR2_X1 U7593 ( .A(n6834), .B(n5933), .ZN(n9754) );
  NAND2_X1 U7594 ( .A1(n9231), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9755) );
  AND2_X1 U7595 ( .A1(n9754), .A2(n9755), .ZN(n5934) );
  NAND2_X1 U7596 ( .A1(n9756), .A2(n5934), .ZN(n9753) );
  OAI21_X1 U7597 ( .B1(n6834), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9753), .ZN(
        n6042) );
  INV_X1 U7598 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5935) );
  MUX2_X1 U7599 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n5935), .S(n6872), .Z(n5936)
         );
  INV_X1 U7600 ( .A(n5936), .ZN(n6043) );
  NOR2_X1 U7601 ( .A1(n6042), .A2(n6043), .ZN(n6041) );
  AOI21_X1 U7602 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6872), .A(n6041), .ZN(
        n5941) );
  NAND2_X1 U7603 ( .A1(n7528), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5937) );
  OAI21_X1 U7604 ( .B1(n7528), .B2(P1_REG2_REG_11__SCAN_IN), .A(n5937), .ZN(
        n5940) );
  INV_X1 U7605 ( .A(n9257), .ZN(n5938) );
  AND2_X1 U7606 ( .A1(n6028), .A2(n5938), .ZN(n9105) );
  AND2_X1 U7607 ( .A1(n5939), .A2(n9105), .ZN(n9785) );
  INV_X1 U7608 ( .A(n9785), .ZN(n9241) );
  NOR2_X1 U7609 ( .A1(n5941), .A2(n5940), .ZN(n6079) );
  AOI211_X1 U7610 ( .C1(n5941), .C2(n5940), .A(n9241), .B(n6079), .ZN(n5942)
         );
  AOI211_X1 U7611 ( .C1(n9781), .C2(n7528), .A(n5943), .B(n5942), .ZN(n5944)
         );
  OAI21_X1 U7612 ( .B1(n5945), .B2(n7196), .A(n5944), .ZN(P1_U3254) );
  INV_X1 U7613 ( .A(n7477), .ZN(n5948) );
  NAND2_X1 U7614 ( .A1(n7240), .A2(P1_B_REG_SCAN_IN), .ZN(n5946) );
  MUX2_X1 U7615 ( .A(P1_B_REG_SCAN_IN), .B(n5946), .S(n7234), .Z(n5947) );
  INV_X1 U7616 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7617 ( .A1(n6192), .A2(n5949), .ZN(n5950) );
  NAND2_X1 U7618 ( .A1(n7477), .A2(n7234), .ZN(n9737) );
  NAND2_X1 U7619 ( .A1(n5950), .A2(n9737), .ZN(n6459) );
  NOR4_X1 U7620 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5954) );
  NOR4_X1 U7621 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5953) );
  NOR4_X1 U7622 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5952) );
  NOR4_X1 U7623 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5951) );
  AND4_X1 U7624 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), .ZN(n5960)
         );
  NOR2_X1 U7625 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .ZN(
        n5958) );
  NOR4_X1 U7626 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5957) );
  NOR4_X1 U7627 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5956) );
  NOR4_X1 U7628 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5955) );
  AND4_X1 U7629 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n5959)
         );
  NAND2_X1 U7630 ( .A1(n5960), .A2(n5959), .ZN(n6191) );
  INV_X1 U7631 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5961) );
  NOR2_X1 U7632 ( .A1(n6191), .A2(n5961), .ZN(n6456) );
  NAND2_X1 U7633 ( .A1(n7477), .A2(n7240), .ZN(n9736) );
  OAI21_X1 U7634 ( .B1(n6455), .B2(n6456), .A(n9736), .ZN(n5962) );
  NOR2_X1 U7635 ( .A1(n6459), .A2(n5962), .ZN(n5994) );
  NAND2_X1 U7636 ( .A1(n5994), .A2(n9106), .ZN(n6002) );
  INV_X1 U7637 ( .A(n8902), .ZN(n5977) );
  NAND2_X1 U7638 ( .A1(n7478), .A2(n9044), .ZN(n6465) );
  INV_X1 U7639 ( .A(n6465), .ZN(n5976) );
  NAND2_X1 U7640 ( .A1(n6360), .A2(n10063), .ZN(n6611) );
  INV_X1 U7641 ( .A(n6611), .ZN(n5964) );
  NAND2_X1 U7642 ( .A1(n5964), .A2(n5963), .ZN(n5971) );
  AND2_X1 U7643 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5965) );
  NAND2_X1 U7644 ( .A1(n6611), .A2(n5965), .ZN(n5970) );
  INV_X1 U7645 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7646 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n5966) );
  NAND2_X1 U7647 ( .A1(n5966), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5967) );
  OAI21_X1 U7648 ( .B1(n5968), .B2(P1_IR_REG_31__SCAN_IN), .A(n5967), .ZN(
        n5969) );
  AND3_X2 U7649 ( .A1(n5971), .A2(n5970), .A3(n5969), .ZN(n9039) );
  INV_X2 U7650 ( .A(n9039), .ZN(n9035) );
  NAND2_X1 U7651 ( .A1(n5972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5974) );
  XNOR2_X1 U7652 ( .A(n5974), .B(n5973), .ZN(n9038) );
  INV_X1 U7653 ( .A(n9037), .ZN(n5975) );
  NAND2_X2 U7654 ( .A1(n6196), .A2(n5995), .ZN(n6166) );
  NAND2_X1 U7655 ( .A1(n6385), .A2(n8496), .ZN(n5984) );
  NAND2_X1 U7656 ( .A1(n4338), .A2(SI_0_), .ZN(n5979) );
  XNOR2_X1 U7657 ( .A(n5979), .B(n5978), .ZN(n9751) );
  MUX2_X1 U7658 ( .A(n9149), .B(n9751), .S(n4341), .Z(n6393) );
  INV_X1 U7659 ( .A(n6393), .ZN(n6464) );
  NAND2_X1 U7660 ( .A1(n5980), .A2(n5995), .ZN(n5981) );
  NAND2_X1 U7661 ( .A1(n6196), .A2(n9039), .ZN(n9553) );
  NAND2_X1 U7662 ( .A1(n7478), .A2(n9037), .ZN(n5982) );
  NAND3_X1 U7663 ( .A1(n9553), .A2(n5995), .A3(n5982), .ZN(n6107) );
  NAND2_X1 U7664 ( .A1(n6464), .A2(n6105), .ZN(n5983) );
  AND2_X1 U7665 ( .A1(n5984), .A2(n5983), .ZN(n6056) );
  NAND2_X1 U7666 ( .A1(n5985), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7667 ( .A1(n6056), .A2(n5986), .ZN(n5991) );
  INV_X1 U7668 ( .A(n6107), .ZN(n8567) );
  NAND2_X1 U7669 ( .A1(n6385), .A2(n8567), .ZN(n5989) );
  OAI22_X1 U7670 ( .A1(n6393), .A2(n6166), .B1(n9149), .B2(n5995), .ZN(n5987)
         );
  INV_X1 U7671 ( .A(n5987), .ZN(n5988) );
  NAND2_X1 U7672 ( .A1(n5989), .A2(n5988), .ZN(n5990) );
  NAND2_X1 U7673 ( .A1(n5991), .A2(n5990), .ZN(n6058) );
  OAI21_X1 U7674 ( .B1(n5991), .B2(n5990), .A(n6058), .ZN(n6029) );
  OR2_X1 U7675 ( .A1(n6465), .A2(n9038), .ZN(n6463) );
  OR2_X1 U7676 ( .A1(n6002), .A2(n6463), .ZN(n5993) );
  INV_X1 U7677 ( .A(n9038), .ZN(n6199) );
  OR2_X2 U7678 ( .A1(n6465), .A2(n6199), .ZN(n9570) );
  OR2_X1 U7679 ( .A1(n9570), .A2(n9035), .ZN(n6190) );
  INV_X1 U7680 ( .A(n6190), .ZN(n5992) );
  NAND2_X1 U7681 ( .A1(n5993), .A2(n9433), .ZN(n8784) );
  INV_X1 U7682 ( .A(n5994), .ZN(n5999) );
  INV_X1 U7683 ( .A(n9658), .ZN(n9805) );
  NAND2_X1 U7684 ( .A1(n5999), .A2(n9805), .ZN(n5997) );
  OR2_X1 U7685 ( .A1(n9037), .A2(n8902), .ZN(n6458) );
  AND2_X1 U7686 ( .A1(n6458), .A2(n5995), .ZN(n5996) );
  NAND2_X1 U7687 ( .A1(n5997), .A2(n5996), .ZN(n6141) );
  INV_X1 U7688 ( .A(n6141), .ZN(n6001) );
  NOR2_X1 U7689 ( .A1(n6463), .A2(P1_U3086), .ZN(n5998) );
  NAND2_X1 U7690 ( .A1(n5999), .A2(n5998), .ZN(n6142) );
  NAND3_X1 U7691 ( .A1(n6001), .A2(n6000), .A3(n6142), .ZN(n6119) );
  INV_X1 U7692 ( .A(n6119), .ZN(n6008) );
  INV_X1 U7693 ( .A(n6002), .ZN(n6003) );
  INV_X1 U7694 ( .A(n8810), .ZN(n8822) );
  NAND2_X1 U7695 ( .A1(n4940), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7696 ( .A1(n7591), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6006) );
  INV_X1 U7697 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6535) );
  OR2_X1 U7698 ( .A1(n7487), .A2(n6535), .ZN(n6005) );
  NAND2_X1 U7699 ( .A1(n9142), .A2(n9259), .ZN(n6467) );
  OAI22_X1 U7700 ( .A1(n6008), .A2(n6469), .B1(n8822), .B2(n6467), .ZN(n6009)
         );
  AOI21_X1 U7701 ( .B1(n6464), .B2(n8784), .A(n6009), .ZN(n6010) );
  OAI21_X1 U7702 ( .B1(n8786), .B2(n6029), .A(n6010), .ZN(P1_U3232) );
  OAI21_X1 U7703 ( .B1(n6011), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6013) );
  INV_X1 U7704 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7705 ( .A1(n6013), .A2(n6012), .ZN(n6089) );
  OR2_X1 U7706 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  AOI22_X1 U7707 ( .A1(n7534), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9740), .ZN(n6015) );
  OAI21_X1 U7708 ( .B1(n7533), .B2(n9747), .A(n6015), .ZN(P1_U3343) );
  INV_X1 U7709 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6017) );
  INV_X1 U7710 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6016) );
  OAI22_X1 U7711 ( .A1(n9788), .A2(n6017), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6016), .ZN(n6026) );
  XNOR2_X1 U7712 ( .A(n6019), .B(n6018), .ZN(n6024) );
  OAI211_X1 U7713 ( .C1(n6022), .C2(n6021), .A(n9785), .B(n6020), .ZN(n6023)
         );
  OAI21_X1 U7714 ( .B1(n7196), .B2(n6024), .A(n6023), .ZN(n6025) );
  AOI211_X1 U7715 ( .C1(n6027), .C2(n9781), .A(n6026), .B(n6025), .ZN(n6033)
         );
  NAND3_X1 U7716 ( .A1(n6029), .A2(n9257), .A3(n6028), .ZN(n6032) );
  AOI22_X1 U7717 ( .A1(n9149), .A2(n6030), .B1(n9105), .B2(n9145), .ZN(n6031)
         );
  NAND3_X1 U7718 ( .A1(n6032), .A2(P1_U3973), .A3(n6031), .ZN(n9184) );
  NAND2_X1 U7719 ( .A1(n6033), .A2(n9184), .ZN(P1_U3245) );
  INV_X1 U7720 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6034) );
  INV_X1 U7721 ( .A(n7527), .ZN(n6036) );
  INV_X1 U7722 ( .A(n7528), .ZN(n6074) );
  OAI222_X1 U7723 ( .A1(n9750), .A2(n6034), .B1(n9747), .B2(n6036), .C1(
        P1_U3086), .C2(n6074), .ZN(P1_U3344) );
  INV_X1 U7724 ( .A(n7171), .ZN(n7212) );
  INV_X1 U7725 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6035) );
  OAI222_X1 U7726 ( .A1(n7212), .A2(P2_U3151), .B1(n7151), .B2(n6036), .C1(
        n6035), .C2(n7236), .ZN(P2_U3284) );
  INV_X1 U7727 ( .A(n7177), .ZN(n7900) );
  INV_X1 U7728 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6037) );
  OAI222_X1 U7729 ( .A1(P2_U3151), .A2(n7900), .B1(n7151), .B2(n7533), .C1(
        n6037), .C2(n7236), .ZN(P2_U3283) );
  AOI211_X1 U7730 ( .C1(n6040), .C2(n6039), .A(n7196), .B(n6038), .ZN(n6049)
         );
  AOI211_X1 U7731 ( .C1(n6043), .C2(n6042), .A(n9241), .B(n6041), .ZN(n6048)
         );
  INV_X1 U7732 ( .A(n6872), .ZN(n6046) );
  INV_X1 U7733 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8620) );
  NOR2_X1 U7734 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8620), .ZN(n6044) );
  AOI21_X1 U7735 ( .B1(n9230), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6044), .ZN(
        n6045) );
  OAI21_X1 U7736 ( .B1(n6046), .B2(n9767), .A(n6045), .ZN(n6047) );
  OR3_X1 U7737 ( .A1(n6049), .A2(n6048), .A3(n6047), .ZN(P1_U3253) );
  INV_X2 U7738 ( .A(n6440), .ZN(n9045) );
  NAND2_X1 U7739 ( .A1(n6384), .A2(n8496), .ZN(n6053) );
  NAND2_X1 U7740 ( .A1(n6383), .A2(n6105), .ZN(n6052) );
  NAND2_X1 U7741 ( .A1(n6053), .A2(n6052), .ZN(n6054) );
  AND2_X1 U7742 ( .A1(n6383), .A2(n8496), .ZN(n6055) );
  AOI21_X1 U7743 ( .B1(n9142), .B2(n8567), .A(n6055), .ZN(n6101) );
  XNOR2_X1 U7744 ( .A(n6100), .B(n6101), .ZN(n6060) );
  NAND2_X1 U7745 ( .A1(n6056), .A2(n8644), .ZN(n6057) );
  AND2_X1 U7746 ( .A1(n6058), .A2(n6057), .ZN(n6059) );
  NAND2_X1 U7747 ( .A1(n6060), .A2(n6059), .ZN(n6104) );
  OAI21_X1 U7748 ( .B1(n6060), .B2(n6059), .A(n6104), .ZN(n6061) );
  NAND2_X1 U7749 ( .A1(n6061), .A2(n8816), .ZN(n6069) );
  INV_X1 U7750 ( .A(n6385), .ZN(n6067) );
  OR2_X1 U7751 ( .A1(n8902), .A2(n9748), .ZN(n9281) );
  NAND2_X1 U7752 ( .A1(n7591), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7753 ( .A1(n4940), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7754 ( .A1(n6062), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7755 ( .A1(n6113), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6063) );
  AND4_X2 U7756 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n6387)
         );
  OAI22_X1 U7757 ( .A1(n6067), .A2(n9281), .B1(n6387), .B2(n8819), .ZN(n6437)
         );
  AOI22_X1 U7758 ( .A1(n6437), .A2(n8810), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6119), .ZN(n6068) );
  OAI211_X1 U7759 ( .C1(n9045), .C2(n8828), .A(n6069), .B(n6068), .ZN(P1_U3222) );
  INV_X1 U7760 ( .A(n5615), .ZN(n6070) );
  INV_X1 U7761 ( .A(n5612), .ZN(n6072) );
  NOR4_X1 U7762 ( .A1(n6072), .A2(n7241), .A3(n7185), .A4(P2_U3151), .ZN(n6073) );
  AOI21_X1 U7763 ( .B1(n6093), .B2(n5611), .A(n6073), .ZN(P2_U3376) );
  AND2_X1 U7764 ( .A1(n6093), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U7765 ( .A1(n6093), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U7766 ( .A1(n6093), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7767 ( .A1(n6093), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U7768 ( .A1(n6093), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U7769 ( .A1(n6093), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U7770 ( .A1(n6093), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7771 ( .A1(n6093), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U7772 ( .A1(n6093), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7773 ( .A1(n6093), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U7774 ( .A1(n6093), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U7775 ( .A1(n6093), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7776 ( .A1(n6093), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U7777 ( .A1(n6093), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U7778 ( .A1(n6093), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U7779 ( .A1(n6093), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7780 ( .A1(n6093), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7781 ( .A1(n6093), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U7782 ( .A1(n6093), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U7783 ( .A1(n6093), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U7784 ( .A1(n6093), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U7785 ( .A1(n6093), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U7786 ( .A1(n6093), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U7787 ( .A1(n6093), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U7788 ( .A1(n6093), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U7789 ( .A1(n6093), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U7790 ( .A1(n6093), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7791 ( .A1(n6093), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  INV_X1 U7792 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10080) );
  OAI22_X1 U7793 ( .A1(n6076), .A2(n6075), .B1(n10080), .B2(n6074), .ZN(n6078)
         );
  XNOR2_X1 U7794 ( .A(n7534), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n6077) );
  NOR2_X1 U7795 ( .A1(n6078), .A2(n6077), .ZN(n6234) );
  AOI21_X1 U7796 ( .B1(n6078), .B2(n6077), .A(n6234), .ZN(n6088) );
  AOI21_X1 U7797 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7528), .A(n6079), .ZN(
        n6082) );
  NOR2_X1 U7798 ( .A1(n7534), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6080) );
  AOI21_X1 U7799 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7534), .A(n6080), .ZN(
        n6081) );
  NAND2_X1 U7800 ( .A1(n6081), .A2(n6082), .ZN(n6244) );
  AOI221_X1 U7801 ( .B1(n6082), .B2(n6244), .C1(n6081), .C2(n6244), .A(n9241), 
        .ZN(n6083) );
  INV_X1 U7802 ( .A(n6083), .ZN(n6087) );
  INV_X1 U7803 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7804 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8693) );
  OAI21_X1 U7805 ( .B1(n9788), .B2(n6084), .A(n8693), .ZN(n6085) );
  AOI21_X1 U7806 ( .B1(n9781), .B2(n7534), .A(n6085), .ZN(n6086) );
  OAI211_X1 U7807 ( .C1(n6088), .C2(n7196), .A(n6087), .B(n6086), .ZN(P1_U3255) );
  INV_X1 U7808 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7809 ( .A1(n6089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6090) );
  XNOR2_X1 U7810 ( .A(n6090), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9248) );
  INV_X1 U7811 ( .A(n9248), .ZN(n6238) );
  OAI222_X1 U7812 ( .A1(n9750), .A2(n6091), .B1(n9747), .B2(n7517), .C1(n6238), 
        .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U7813 ( .A(n7927), .ZN(n7917) );
  INV_X1 U7814 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6092) );
  OAI222_X1 U7815 ( .A1(P2_U3151), .A2(n7917), .B1(n7151), .B2(n7517), .C1(
        n6092), .C2(n7236), .ZN(P2_U3282) );
  INV_X1 U7816 ( .A(n6093), .ZN(n6094) );
  INV_X1 U7817 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10169) );
  NOR2_X1 U7818 ( .A1(n6094), .A2(n10169), .ZN(P2_U3262) );
  INV_X1 U7819 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10082) );
  NOR2_X1 U7820 ( .A1(n6094), .A2(n10082), .ZN(P2_U3248) );
  OR2_X1 U7821 ( .A1(n8864), .A2(n6095), .ZN(n6098) );
  OAI211_X1 U7822 ( .C1(n6263), .C2(n6099), .A(n6098), .B(n6097), .ZN(n6108)
         );
  INV_X1 U7823 ( .A(n6108), .ZN(n9796) );
  INV_X1 U7824 ( .A(n6100), .ZN(n6102) );
  NAND2_X1 U7825 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  NAND2_X1 U7826 ( .A1(n6104), .A2(n6103), .ZN(n6123) );
  OAI22_X1 U7827 ( .A1(n6387), .A2(n6166), .B1(n9796), .B2(n6267), .ZN(n6106)
         );
  XNOR2_X1 U7828 ( .A(n6106), .B(n8644), .ZN(n6126) );
  OR2_X1 U7829 ( .A1(n6387), .A2(n8641), .ZN(n6111) );
  NAND2_X1 U7830 ( .A1(n6109), .A2(n8640), .ZN(n6110) );
  NAND2_X1 U7831 ( .A1(n6111), .A2(n6110), .ZN(n6124) );
  XNOR2_X1 U7832 ( .A(n6126), .B(n6124), .ZN(n6122) );
  XNOR2_X1 U7833 ( .A(n6123), .B(n6122), .ZN(n6112) );
  NAND2_X1 U7834 ( .A1(n6112), .A2(n8816), .ZN(n6121) );
  INV_X1 U7835 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U7836 ( .A1(n4940), .A2(n6823), .ZN(n6117) );
  NAND2_X1 U7837 ( .A1(n7591), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7838 ( .A1(n6062), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7839 ( .A1(n6113), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6114) );
  NAND4_X1 U7840 ( .A1(n6117), .A2(n6116), .A3(n6115), .A4(n6114), .ZN(n9140)
         );
  INV_X1 U7841 ( .A(n9140), .ZN(n6388) );
  INV_X1 U7842 ( .A(n9142), .ZN(n6118) );
  OAI22_X1 U7843 ( .A1(n6388), .A2(n8819), .B1(n6118), .B2(n9281), .ZN(n6409)
         );
  AOI22_X1 U7844 ( .A1(n6409), .A2(n8810), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6119), .ZN(n6120) );
  OAI211_X1 U7845 ( .C1(n9796), .C2(n8828), .A(n6121), .B(n6120), .ZN(P1_U3237) );
  NAND2_X1 U7846 ( .A1(n6123), .A2(n6122), .ZN(n6128) );
  INV_X1 U7847 ( .A(n6124), .ZN(n6125) );
  NAND2_X1 U7848 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  NAND2_X1 U7849 ( .A1(n6128), .A2(n6127), .ZN(n6157) );
  OR2_X1 U7850 ( .A1(n4341), .A2(n9157), .ZN(n6131) );
  NAND2_X1 U7851 ( .A1(n9140), .A2(n8640), .ZN(n6132) );
  NAND2_X1 U7852 ( .A1(n9140), .A2(n8567), .ZN(n6134) );
  OR2_X1 U7853 ( .A1(n6826), .A2(n8541), .ZN(n6133) );
  NAND2_X1 U7854 ( .A1(n6134), .A2(n6133), .ZN(n6158) );
  XNOR2_X1 U7855 ( .A(n6160), .B(n6158), .ZN(n6156) );
  XOR2_X1 U7856 ( .A(n6157), .B(n6156), .Z(n6147) );
  NAND2_X1 U7857 ( .A1(n8867), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6140) );
  INV_X1 U7858 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7859 ( .A1(n6823), .A2(n6135), .ZN(n6136) );
  NAND2_X1 U7860 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6180) );
  AND2_X1 U7861 ( .A1(n6136), .A2(n6180), .ZN(n6550) );
  NAND2_X1 U7862 ( .A1(n4443), .A2(n6550), .ZN(n6139) );
  INV_X2 U7863 ( .A(n7487), .ZN(n8868) );
  NAND2_X1 U7864 ( .A1(n8868), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7865 ( .A1(n6113), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6137) );
  OAI22_X1 U7866 ( .A1(n6387), .A2(n9281), .B1(n6390), .B2(n8819), .ZN(n6416)
         );
  AOI22_X1 U7867 ( .A1(n6416), .A2(n8810), .B1(n6419), .B2(n8784), .ZN(n6146)
         );
  NAND2_X1 U7868 ( .A1(n6141), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6144) );
  AND2_X1 U7869 ( .A1(n6142), .A2(n9108), .ZN(n6143) );
  NAND2_X1 U7870 ( .A1(n6144), .A2(n6143), .ZN(n8825) );
  INV_X1 U7871 ( .A(n8825), .ZN(n8808) );
  MUX2_X1 U7872 ( .A(n8808), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6145) );
  OAI211_X1 U7873 ( .C1(n6147), .C2(n8786), .A(n6146), .B(n6145), .ZN(P1_U3218) );
  NAND2_X1 U7874 ( .A1(P2_U3893), .A2(n6934), .ZN(n6148) );
  OAI21_X1 U7875 ( .B1(P2_U3893), .B2(n5978), .A(n6148), .ZN(P2_U3491) );
  INV_X1 U7876 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6153) );
  INV_X1 U7877 ( .A(n7547), .ZN(n6155) );
  NAND2_X1 U7878 ( .A1(n6149), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6150) );
  MUX2_X1 U7879 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6150), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6151) );
  INV_X1 U7880 ( .A(n6151), .ZN(n6152) );
  NOR2_X1 U7881 ( .A1(n6152), .A2(n6204), .ZN(n7548) );
  INV_X1 U7882 ( .A(n7548), .ZN(n6687) );
  OAI222_X1 U7883 ( .A1(n9750), .A2(n6153), .B1(n9747), .B2(n6155), .C1(
        P1_U3086), .C2(n6687), .ZN(P1_U3341) );
  INV_X1 U7884 ( .A(n7930), .ZN(n7943) );
  INV_X1 U7885 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6154) );
  OAI222_X1 U7886 ( .A1(n7943), .A2(P2_U3151), .B1(n7151), .B2(n6155), .C1(
        n6154), .C2(n7236), .ZN(P2_U3281) );
  INV_X1 U7887 ( .A(n6550), .ZN(n6189) );
  INV_X1 U7888 ( .A(n6158), .ZN(n6159) );
  NAND2_X1 U7889 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  NOR2_X1 U7890 ( .A1(n6162), .A2(n8836), .ZN(n6165) );
  OAI22_X1 U7891 ( .A1(n8864), .A2(n6163), .B1(n9175), .B2(n6263), .ZN(n6164)
         );
  OAI22_X1 U7892 ( .A1(n6390), .A2(n6166), .B1(n6553), .B2(n6267), .ZN(n6167)
         );
  XNOR2_X1 U7893 ( .A(n6167), .B(n8565), .ZN(n6170) );
  OR2_X1 U7894 ( .A1(n6390), .A2(n8641), .ZN(n6169) );
  NAND2_X1 U7895 ( .A1(n6430), .A2(n8640), .ZN(n6168) );
  NAND2_X1 U7896 ( .A1(n6169), .A2(n6168), .ZN(n6171) );
  NAND2_X1 U7897 ( .A1(n6170), .A2(n6171), .ZN(n6260) );
  INV_X1 U7898 ( .A(n6170), .ZN(n6173) );
  INV_X1 U7899 ( .A(n6171), .ZN(n6172) );
  NAND2_X1 U7900 ( .A1(n6173), .A2(n6172), .ZN(n6174) );
  NAND2_X1 U7901 ( .A1(n6260), .A2(n6174), .ZN(n6176) );
  AOI21_X1 U7902 ( .B1(n6175), .B2(n6176), .A(n8786), .ZN(n6178) );
  NAND2_X1 U7903 ( .A1(n6178), .A2(n6261), .ZN(n6188) );
  INV_X1 U7904 ( .A(n9281), .ZN(n8804) );
  NAND2_X1 U7905 ( .A1(n8867), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6185) );
  AND2_X1 U7906 ( .A1(n6180), .A2(n6179), .ZN(n6181) );
  NOR2_X1 U7907 ( .A1(n6274), .A2(n6181), .ZN(n6593) );
  NAND2_X1 U7908 ( .A1(n4443), .A2(n6593), .ZN(n6184) );
  NAND2_X1 U7909 ( .A1(n8868), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7910 ( .A1(n4333), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6182) );
  NAND4_X1 U7911 ( .A1(n6185), .A2(n6184), .A3(n6183), .A4(n6182), .ZN(n9138)
         );
  AOI22_X1 U7912 ( .A1(n8804), .A2(n9140), .B1(n9138), .B2(n9259), .ZN(n6428)
         );
  NAND2_X1 U7913 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9168) );
  OAI21_X1 U7914 ( .B1(n6428), .B2(n8822), .A(n9168), .ZN(n6186) );
  AOI21_X1 U7915 ( .B1(n6430), .B2(n8784), .A(n6186), .ZN(n6187) );
  OAI211_X1 U7916 ( .C1(n8808), .C2(n6189), .A(n6188), .B(n6187), .ZN(P1_U3230) );
  AND2_X1 U7917 ( .A1(n6190), .A2(n6458), .ZN(n6195) );
  NAND2_X1 U7918 ( .A1(n6192), .A2(n6191), .ZN(n6194) );
  OAI21_X1 U7919 ( .B1(n6455), .B2(P1_D_REG_1__SCAN_IN), .A(n9736), .ZN(n6193)
         );
  NAND4_X1 U7920 ( .A1(n6195), .A2(n9106), .A3(n6194), .A4(n6193), .ZN(n6210)
         );
  NOR2_X4 U7921 ( .A1(n6210), .A2(n6459), .ZN(n9816) );
  AND2_X1 U7922 ( .A1(n6197), .A2(n6196), .ZN(n9104) );
  OAI21_X1 U7923 ( .B1(n6197), .B2(n9037), .A(n6465), .ZN(n6198) );
  OR2_X1 U7924 ( .A1(n9104), .A2(n6198), .ZN(n9560) );
  AND2_X1 U7925 ( .A1(n7478), .A2(n9039), .ZN(n9021) );
  NAND2_X1 U7926 ( .A1(n9021), .A2(n9038), .ZN(n9671) );
  NAND2_X1 U7927 ( .A1(n9560), .A2(n9671), .ZN(n9809) );
  OR2_X1 U7928 ( .A1(n9035), .A2(n7478), .ZN(n6201) );
  NAND2_X1 U7929 ( .A1(n9025), .A2(n6199), .ZN(n6200) );
  NOR2_X1 U7930 ( .A1(n6385), .A2(n6393), .ZN(n6395) );
  INV_X1 U7931 ( .A(n6395), .ZN(n6436) );
  NAND2_X1 U7932 ( .A1(n6385), .A2(n6393), .ZN(n9041) );
  NAND2_X1 U7933 ( .A1(n6436), .A2(n9041), .ZN(n8841) );
  OAI21_X1 U7934 ( .B1(n9809), .B2(n9526), .A(n8841), .ZN(n6202) );
  OAI211_X1 U7935 ( .C1(n6465), .C2(n6393), .A(n6202), .B(n6467), .ZN(n6211)
         );
  NAND2_X1 U7936 ( .A1(n6211), .A2(n9816), .ZN(n6203) );
  OAI21_X1 U7937 ( .B1(n9816), .B2(n9150), .A(n6203), .ZN(P1_U3522) );
  INV_X1 U7938 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6206) );
  INV_X1 U7939 ( .A(n7559), .ZN(n6208) );
  OR2_X1 U7940 ( .A1(n6204), .A2(n9738), .ZN(n6205) );
  XNOR2_X1 U7941 ( .A(n6205), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7560) );
  INV_X1 U7942 ( .A(n7560), .ZN(n6789) );
  OAI222_X1 U7943 ( .A1(n9750), .A2(n6206), .B1(n9747), .B2(n6208), .C1(
        P1_U3086), .C2(n6789), .ZN(P1_U3340) );
  INV_X1 U7944 ( .A(n7972), .ZN(n7962) );
  INV_X1 U7945 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6207) );
  OAI222_X1 U7946 ( .A1(n7962), .A2(P2_U3151), .B1(n7151), .B2(n6208), .C1(
        n6207), .C2(n7236), .ZN(P2_U3280) );
  INV_X1 U7947 ( .A(n6459), .ZN(n6209) );
  INV_X1 U7948 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7949 ( .A1(n6211), .A2(n9725), .ZN(n6212) );
  OAI21_X1 U7950 ( .B1(n9725), .B2(n6213), .A(n6212), .ZN(P1_U3453) );
  NAND2_X1 U7951 ( .A1(n8867), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7952 ( .A1(n6274), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U7953 ( .A1(n6840), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6887) );
  INV_X1 U7954 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7537) );
  NAND2_X1 U7955 ( .A1(n7540), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7552) );
  INV_X1 U7956 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7551) );
  INV_X1 U7957 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7563) );
  INV_X1 U7958 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7493) );
  INV_X1 U7959 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7578) );
  INV_X1 U7960 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U7961 ( .A1(n7601), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7611) );
  INV_X1 U7962 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n7610) );
  INV_X1 U7963 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8615) );
  AND2_X1 U7964 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n6214) );
  NAND2_X1 U7965 ( .A1(n7658), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n7665) );
  INV_X1 U7966 ( .A(n7665), .ZN(n6215) );
  AND2_X1 U7967 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n6215), .ZN(n9284) );
  NAND2_X1 U7968 ( .A1(n4443), .A2(n9284), .ZN(n6218) );
  NAND2_X1 U7969 ( .A1(n8868), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7970 ( .A1(n4333), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6216) );
  INV_X1 U7971 ( .A(P1_U3973), .ZN(n9128) );
  NAND2_X1 U7972 ( .A1(n9128), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6220) );
  OAI21_X1 U7973 ( .B1(n8837), .B2(n9128), .A(n6220), .ZN(P1_U3583) );
  NOR2_X1 U7974 ( .A1(n7850), .A2(P2_U3151), .ZN(n6377) );
  NAND2_X1 U7975 ( .A1(n6934), .A2(n8364), .ZN(n7265) );
  INV_X1 U7976 ( .A(n7265), .ZN(n6222) );
  OR2_X1 U7977 ( .A1(n6222), .A2(n6221), .ZN(n8360) );
  OAI22_X1 U7978 ( .A1(n7853), .A2(n8364), .B1(n4992), .B2(n7855), .ZN(n6223)
         );
  AOI21_X1 U7979 ( .B1(n8360), .B2(n7845), .A(n6223), .ZN(n6224) );
  OAI21_X1 U7980 ( .B1(n6377), .B2(n6774), .A(n6224), .ZN(P2_U3172) );
  INV_X1 U7981 ( .A(n9952), .ZN(n9938) );
  OAI21_X1 U7982 ( .B1(n6225), .B2(n6226), .A(n6945), .ZN(n6956) );
  XNOR2_X1 U7983 ( .A(n6227), .B(n6226), .ZN(n6228) );
  OAI222_X1 U7984 ( .A1(n8278), .A2(n6678), .B1(n8276), .B2(n6376), .C1(n8358), 
        .C2(n6228), .ZN(n6953) );
  AOI21_X1 U7985 ( .B1(n9933), .B2(n6956), .A(n6953), .ZN(n6233) );
  INV_X1 U7986 ( .A(n6952), .ZN(n6291) );
  AOI22_X1 U7987 ( .A1(n5656), .A2(n6291), .B1(n10190), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n6229) );
  OAI21_X1 U7988 ( .B1(n6233), .B2(n10190), .A(n6229), .ZN(P2_U3462) );
  INV_X1 U7989 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6230) );
  OAI22_X1 U7990 ( .A1(n6952), .A2(n8420), .B1(n9965), .B2(n6230), .ZN(n6231)
         );
  INV_X1 U7991 ( .A(n6231), .ZN(n6232) );
  OAI21_X1 U7992 ( .B1(n6233), .B2(n9966), .A(n6232), .ZN(P2_U3399) );
  INV_X1 U7993 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n6242) );
  XNOR2_X1 U7994 ( .A(n6687), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n6240) );
  INV_X1 U7995 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6237) );
  XNOR2_X1 U7996 ( .A(n6238), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9250) );
  OR2_X1 U7997 ( .A1(n7534), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6236) );
  INV_X1 U7998 ( .A(n6234), .ZN(n6235) );
  NAND2_X1 U7999 ( .A1(n9250), .A2(n9251), .ZN(n9249) );
  OAI21_X1 U8000 ( .B1(n6238), .B2(n6237), .A(n9249), .ZN(n6239) );
  NAND2_X1 U8001 ( .A1(n6240), .A2(n6239), .ZN(n6686) );
  OAI211_X1 U8002 ( .C1(n6240), .C2(n6239), .A(n9779), .B(n6686), .ZN(n6241)
         );
  NAND2_X1 U8003 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8602) );
  OAI211_X1 U8004 ( .C1(n9788), .C2(n6242), .A(n6241), .B(n8602), .ZN(n6249)
         );
  NAND2_X1 U8005 ( .A1(n9248), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6243) );
  OAI21_X1 U8006 ( .B1(n9248), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6243), .ZN(
        n9244) );
  OAI21_X1 U8007 ( .B1(n7534), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6244), .ZN(
        n9243) );
  NOR2_X1 U8008 ( .A1(n9244), .A2(n9243), .ZN(n9242) );
  AOI21_X1 U8009 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9248), .A(n9242), .ZN(
        n6247) );
  NAND2_X1 U8010 ( .A1(n7548), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6245) );
  OAI21_X1 U8011 ( .B1(n7548), .B2(P1_REG2_REG_14__SCAN_IN), .A(n6245), .ZN(
        n6246) );
  NOR2_X1 U8012 ( .A1(n6247), .A2(n6246), .ZN(n6692) );
  AOI211_X1 U8013 ( .C1(n6247), .C2(n6246), .A(n6692), .B(n9241), .ZN(n6248)
         );
  AOI211_X1 U8014 ( .C1(n9781), .C2(n7548), .A(n6249), .B(n6248), .ZN(n6250)
         );
  INV_X1 U8015 ( .A(n6250), .ZN(P1_U3257) );
  OAI21_X1 U8016 ( .B1(n6253), .B2(n6252), .A(n6251), .ZN(n6254) );
  NAND2_X1 U8017 ( .A1(n6254), .A2(n7845), .ZN(n6258) );
  INV_X1 U8018 ( .A(n7853), .ZN(n7866) );
  OAI22_X1 U8019 ( .A1(n4992), .A2(n7810), .B1(n7855), .B2(n6721), .ZN(n6255)
         );
  AOI21_X1 U8020 ( .B1(n7866), .B2(n6256), .A(n6255), .ZN(n6257) );
  OAI211_X1 U8021 ( .C1(n6377), .C2(n6259), .A(n6258), .B(n6257), .ZN(P2_U3177) );
  OR2_X1 U8022 ( .A1(n6262), .A2(n8836), .ZN(n6265) );
  AOI22_X1 U8023 ( .A1(n7575), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7574), .B2(
        n9191), .ZN(n6264) );
  AND2_X2 U8024 ( .A1(n6265), .A2(n6264), .ZN(n6596) );
  NAND2_X1 U8025 ( .A1(n9138), .A2(n8496), .ZN(n6266) );
  OAI21_X1 U8026 ( .B1(n6596), .B2(n6267), .A(n6266), .ZN(n6268) );
  XNOR2_X1 U8027 ( .A(n6268), .B(n8565), .ZN(n6270) );
  NAND2_X1 U8028 ( .A1(n6504), .A2(n6503), .ZN(n6273) );
  AND2_X1 U8029 ( .A1(n9138), .A2(n8567), .ZN(n6272) );
  AOI21_X1 U8030 ( .B1(n6475), .B2(n8640), .A(n6272), .ZN(n6502) );
  XNOR2_X1 U8031 ( .A(n6273), .B(n6502), .ZN(n6285) );
  NAND2_X1 U8032 ( .A1(n8867), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6279) );
  OR2_X1 U8033 ( .A1(n6274), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6275) );
  AND2_X1 U8034 ( .A1(n6486), .A2(n6275), .ZN(n6663) );
  NAND2_X1 U8035 ( .A1(n4443), .A2(n6663), .ZN(n6278) );
  NAND2_X1 U8036 ( .A1(n8868), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U8037 ( .A1(n4333), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6276) );
  OR2_X1 U8038 ( .A1(n6508), .A2(n8819), .ZN(n6281) );
  OR2_X1 U8039 ( .A1(n6390), .A2(n9281), .ZN(n6280) );
  NAND2_X1 U8040 ( .A1(n6281), .A2(n6280), .ZN(n6402) );
  NAND2_X1 U8041 ( .A1(n6402), .A2(n8810), .ZN(n6282) );
  NAND2_X1 U8042 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9185) );
  OAI211_X1 U8043 ( .C1(n8828), .C2(n6596), .A(n6282), .B(n9185), .ZN(n6283)
         );
  AOI21_X1 U8044 ( .B1(n6593), .B2(n8825), .A(n6283), .ZN(n6284) );
  OAI21_X1 U8045 ( .B1(n6285), .B2(n8786), .A(n6284), .ZN(P1_U3227) );
  OAI211_X1 U8046 ( .C1(n6288), .C2(n6287), .A(n6286), .B(n7845), .ZN(n6293)
         );
  OAI22_X1 U8047 ( .A1(n6376), .A2(n7810), .B1(n7855), .B2(n6678), .ZN(n6290)
         );
  MUX2_X1 U8048 ( .A(n7850), .B(P2_U3151), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n6289) );
  AOI211_X1 U8049 ( .C1(n6291), .C2(n7866), .A(n6290), .B(n6289), .ZN(n6292)
         );
  NAND2_X1 U8050 ( .A1(n6293), .A2(n6292), .ZN(P2_U3158) );
  INV_X1 U8051 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6296) );
  INV_X1 U8052 ( .A(n7513), .ZN(n6298) );
  NAND2_X1 U8053 ( .A1(n6294), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6295) );
  XNOR2_X1 U8054 ( .A(n6295), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7514) );
  INV_X1 U8055 ( .A(n7514), .ZN(n7105) );
  OAI222_X1 U8056 ( .A1(n9750), .A2(n6296), .B1(n9747), .B2(n6298), .C1(n7105), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U8057 ( .A(n7976), .ZN(n7990) );
  INV_X1 U8058 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6297) );
  OAI222_X1 U8059 ( .A1(P2_U3151), .A2(n7990), .B1(n7151), .B2(n6298), .C1(
        n6297), .C2(n7236), .ZN(P2_U3279) );
  MUX2_X1 U8060 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8041), .Z(n6331) );
  XNOR2_X1 U8061 ( .A(n6331), .B(n6345), .ZN(n6333) );
  MUX2_X1 U8062 ( .A(n10089), .B(n6299), .S(n8041), .Z(n6301) );
  XNOR2_X1 U8063 ( .A(n6301), .B(n6573), .ZN(n6566) );
  MUX2_X1 U8064 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n8041), .Z(n6300) );
  INV_X1 U8065 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6318) );
  NOR2_X1 U8066 ( .A1(n6300), .A2(n6318), .ZN(n6565) );
  OAI22_X1 U8067 ( .A1(n6566), .A2(n6565), .B1(n6573), .B2(n6301), .ZN(n9830)
         );
  MUX2_X1 U8068 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8041), .Z(n6303) );
  XNOR2_X1 U8069 ( .A(n6303), .B(n9825), .ZN(n9831) );
  AOI22_X1 U8070 ( .A1(n9830), .A2(n9831), .B1(n6303), .B2(n6302), .ZN(n6334)
         );
  XOR2_X1 U8071 ( .A(n6333), .B(n6334), .Z(n6330) );
  INV_X1 U8072 ( .A(n6304), .ZN(n6308) );
  INV_X1 U8073 ( .A(n6312), .ZN(n6306) );
  NOR2_X1 U8074 ( .A1(n8041), .A2(P2_U3151), .ZN(n8437) );
  AND2_X1 U8075 ( .A1(n8437), .A2(n6307), .ZN(n6305) );
  NAND2_X1 U8076 ( .A1(n6306), .A2(n6305), .ZN(n6310) );
  OR2_X1 U8077 ( .A1(n6307), .A2(P2_U3151), .ZN(n6311) );
  INV_X1 U8078 ( .A(n6311), .ZN(n8435) );
  NAND2_X1 U8079 ( .A1(n6308), .A2(n8435), .ZN(n6309) );
  NOR2_X1 U8080 ( .A1(n6312), .A2(n6311), .ZN(n6366) );
  NAND2_X1 U8081 ( .A1(n6366), .A2(n6313), .ZN(n9891) );
  INV_X1 U8082 ( .A(n9891), .ZN(n9916) );
  NAND2_X1 U8083 ( .A1(n6318), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6315) );
  NOR2_X1 U8084 ( .A1(n6314), .A2(n6363), .ZN(n6316) );
  NAND2_X1 U8085 ( .A1(n6571), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6570) );
  INV_X1 U8086 ( .A(n6316), .ZN(n6317) );
  NAND2_X1 U8087 ( .A1(n6570), .A2(n6317), .ZN(n9818) );
  OAI21_X1 U8088 ( .B1(n9825), .B2(n6724), .A(n9817), .ZN(n6344) );
  XNOR2_X1 U8089 ( .A(n6347), .B(n5021), .ZN(n6325) );
  AND2_X1 U8090 ( .A1(n6366), .A2(n8041), .ZN(n9901) );
  INV_X1 U8091 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10067) );
  OR2_X1 U8092 ( .A1(n6562), .A2(n6299), .ZN(n6563) );
  NAND2_X1 U8093 ( .A1(n6563), .A2(n6319), .ZN(n9821) );
  OR2_X1 U8094 ( .A1(n9825), .A2(n10067), .ZN(n6320) );
  NAND2_X1 U8095 ( .A1(n6321), .A2(n4335), .ZN(n9837) );
  OAI21_X1 U8096 ( .B1(n6323), .B2(P2_REG1_REG_3__SCAN_IN), .A(n9839), .ZN(
        n6324) );
  AOI22_X1 U8097 ( .A1(n9916), .A2(n6325), .B1(n9901), .B2(n6324), .ZN(n6327)
         );
  NAND2_X1 U8098 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6326) );
  OAI211_X1 U8099 ( .C1(n9906), .C2(n4335), .A(n6327), .B(n6326), .ZN(n6328)
         );
  AOI21_X1 U8100 ( .B1(n9897), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6328), .ZN(
        n6329) );
  OAI21_X1 U8101 ( .B1(n9911), .B2(n6330), .A(n6329), .ZN(P2_U3185) );
  MUX2_X1 U8102 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8041), .Z(n6624) );
  XNOR2_X1 U8103 ( .A(n6624), .B(n6644), .ZN(n6626) );
  MUX2_X1 U8104 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8041), .Z(n6335) );
  INV_X1 U8105 ( .A(n6335), .ZN(n6336) );
  INV_X1 U8106 ( .A(n6331), .ZN(n6332) );
  AOI22_X1 U8107 ( .A1(n6334), .A2(n6333), .B1(n6345), .B2(n6332), .ZN(n9849)
         );
  XNOR2_X1 U8108 ( .A(n6335), .B(n6349), .ZN(n9848) );
  NAND2_X1 U8109 ( .A1(n9849), .A2(n9848), .ZN(n9847) );
  OAI21_X1 U8110 ( .B1(n6349), .B2(n6336), .A(n9847), .ZN(n9865) );
  MUX2_X1 U8111 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8041), .Z(n6337) );
  XNOR2_X1 U8112 ( .A(n6337), .B(n4485), .ZN(n9866) );
  AOI22_X1 U8113 ( .A1(n9865), .A2(n9866), .B1(n6337), .B2(n9858), .ZN(n6627)
         );
  XOR2_X1 U8114 ( .A(n6626), .B(n6627), .Z(n6359) );
  INV_X1 U8115 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9968) );
  MUX2_X1 U8116 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9968), .S(n9835), .Z(n9836)
         );
  NAND2_X1 U8117 ( .A1(n9835), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U8118 ( .A1(n6339), .A2(n9858), .ZN(n6341) );
  XNOR2_X1 U8119 ( .A(n6644), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n6340) );
  INV_X1 U8120 ( .A(n6340), .ZN(n6342) );
  NAND3_X1 U8121 ( .A1(n9859), .A2(n6342), .A3(n6341), .ZN(n6343) );
  AOI21_X1 U8122 ( .B1(n6636), .B2(n6343), .A(n8000), .ZN(n6355) );
  INV_X1 U8123 ( .A(n6344), .ZN(n6346) );
  MUX2_X1 U8124 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6348), .S(n9835), .Z(n9852)
         );
  INV_X1 U8125 ( .A(n6350), .ZN(n6352) );
  XNOR2_X1 U8126 ( .A(n6644), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6351) );
  OR3_X1 U8127 ( .A1(n9869), .A2(n6352), .A3(n6351), .ZN(n6353) );
  AOI21_X1 U8128 ( .B1(n6643), .B2(n6353), .A(n9891), .ZN(n6354) );
  NOR2_X1 U8129 ( .A1(n6355), .A2(n6354), .ZN(n6356) );
  NAND2_X1 U8130 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6729) );
  OAI211_X1 U8131 ( .C1(n9906), .C2(n6634), .A(n6356), .B(n6729), .ZN(n6357)
         );
  AOI21_X1 U8132 ( .B1(n9897), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6357), .ZN(
        n6358) );
  OAI21_X1 U8133 ( .B1(n9911), .B2(n6359), .A(n6358), .ZN(P2_U3188) );
  INV_X1 U8134 ( .A(n7498), .ZN(n6454) );
  XNOR2_X1 U8135 ( .A(n6360), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9780) );
  AOI22_X1 U8136 ( .A1(n9780), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9740), .ZN(n6361) );
  OAI21_X1 U8137 ( .B1(n6454), .B2(n9747), .A(n6361), .ZN(P1_U3338) );
  INV_X1 U8138 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6370) );
  INV_X1 U8139 ( .A(n9906), .ZN(n9826) );
  MUX2_X1 U8140 ( .A(n6363), .B(n6362), .S(n8041), .Z(n6364) );
  NOR2_X1 U8141 ( .A1(n6364), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6365) );
  OAI22_X1 U8142 ( .A1(n9867), .A2(n6366), .B1(n6565), .B2(n6365), .ZN(n6367)
         );
  OAI21_X1 U8143 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6774), .A(n6367), .ZN(n6368) );
  AOI21_X1 U8144 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9826), .A(n6368), .ZN(n6369) );
  OAI21_X1 U8145 ( .B1(n9882), .B2(n6370), .A(n6369), .ZN(P2_U3182) );
  INV_X1 U8146 ( .A(n6371), .ZN(n6372) );
  AOI21_X1 U8147 ( .B1(n6374), .B2(n6373), .A(n6372), .ZN(n6382) );
  INV_X1 U8148 ( .A(n6934), .ZN(n6375) );
  OAI22_X1 U8149 ( .A1(n6376), .A2(n7855), .B1(n7810), .B2(n6375), .ZN(n6379)
         );
  NOR2_X1 U8150 ( .A1(n6377), .A2(n6930), .ZN(n6378) );
  AOI211_X1 U8151 ( .C1(n6380), .C2(n7866), .A(n6379), .B(n6378), .ZN(n6381)
         );
  OAI21_X1 U8152 ( .B1(n7861), .B2(n6382), .A(n6381), .ZN(P2_U3162) );
  INV_X1 U8153 ( .A(n6390), .ZN(n9139) );
  INV_X1 U8154 ( .A(n6387), .ZN(n9141) );
  NAND2_X1 U8155 ( .A1(n6385), .A2(n6464), .ZN(n6433) );
  NAND2_X1 U8156 ( .A1(n6432), .A2(n6386), .ZN(n6407) );
  NAND2_X1 U8157 ( .A1(n6387), .A2(n6109), .ZN(n6396) );
  NAND2_X1 U8158 ( .A1(n9141), .A2(n9796), .ZN(n9042) );
  NAND2_X1 U8159 ( .A1(n6407), .A2(n8839), .ZN(n6406) );
  NAND2_X1 U8160 ( .A1(n6388), .A2(n6419), .ZN(n8918) );
  NAND2_X1 U8161 ( .A1(n9140), .A2(n6826), .ZN(n8922) );
  NAND2_X1 U8162 ( .A1(n6413), .A2(n6389), .ZN(n6422) );
  NAND2_X1 U8163 ( .A1(n6390), .A2(n6430), .ZN(n8923) );
  NAND2_X1 U8164 ( .A1(n9139), .A2(n6553), .ZN(n9049) );
  AND2_X1 U8165 ( .A1(n8923), .A2(n9049), .ZN(n8916) );
  INV_X1 U8166 ( .A(n8916), .ZN(n6426) );
  NAND2_X1 U8167 ( .A1(n6422), .A2(n6426), .ZN(n6421) );
  NAND2_X1 U8168 ( .A1(n6596), .A2(n9138), .ZN(n9053) );
  INV_X1 U8169 ( .A(n9138), .ZN(n6391) );
  NAND2_X1 U8170 ( .A1(n6391), .A2(n6475), .ZN(n8924) );
  NAND2_X1 U8171 ( .A1(n9053), .A2(n8924), .ZN(n8845) );
  NAND2_X1 U8172 ( .A1(n6392), .A2(n8845), .ZN(n6477) );
  OAI21_X1 U8173 ( .B1(n6392), .B2(n8845), .A(n6477), .ZN(n6598) );
  AOI21_X1 U8174 ( .B1(n6424), .B2(n6475), .A(n9570), .ZN(n6394) );
  AND2_X1 U8175 ( .A1(n6394), .A2(n6482), .ZN(n6592) );
  INV_X1 U8176 ( .A(n8923), .ZN(n6398) );
  NAND2_X1 U8177 ( .A1(n6399), .A2(n9049), .ZN(n6401) );
  INV_X1 U8178 ( .A(n8845), .ZN(n6400) );
  NAND2_X1 U8179 ( .A1(n6401), .A2(n6400), .ZN(n6483) );
  OAI211_X1 U8180 ( .C1(n6401), .C2(n6400), .A(n6483), .B(n9526), .ZN(n6404)
         );
  INV_X1 U8181 ( .A(n6402), .ZN(n6403) );
  NAND2_X1 U8182 ( .A1(n6404), .A2(n6403), .ZN(n6591) );
  AOI211_X1 U8183 ( .C1(n6598), .C2(n9809), .A(n6592), .B(n6591), .ZN(n6497)
         );
  AOI22_X1 U8184 ( .A1(n9676), .A2(n6475), .B1(n9814), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n6405) );
  OAI21_X1 U8185 ( .B1(n6497), .B2(n9814), .A(n6405), .ZN(P1_U3527) );
  OAI21_X1 U8186 ( .B1(n6407), .B2(n8839), .A(n6406), .ZN(n9798) );
  INV_X1 U8187 ( .A(n6415), .ZN(n6408) );
  AOI211_X1 U8188 ( .C1(n6109), .C2(n6435), .A(n9570), .B(n6408), .ZN(n9791)
         );
  AOI21_X1 U8189 ( .B1(n6410), .B2(n9526), .A(n6409), .ZN(n9801) );
  INV_X1 U8190 ( .A(n9801), .ZN(n6411) );
  AOI211_X1 U8191 ( .C1(n9809), .C2(n9798), .A(n9791), .B(n6411), .ZN(n6530)
         );
  AOI22_X1 U8192 ( .A1(n9676), .A2(n6109), .B1(n9814), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6412) );
  OAI21_X1 U8193 ( .B1(n6530), .B2(n9814), .A(n6412), .ZN(P1_U3524) );
  OAI21_X1 U8194 ( .B1(n6414), .B2(n8840), .A(n6413), .ZN(n6828) );
  AOI211_X1 U8195 ( .C1(n6419), .C2(n6415), .A(n9570), .B(n6423), .ZN(n6822)
         );
  INV_X1 U8196 ( .A(n8913), .ZN(n9048) );
  XNOR2_X1 U8197 ( .A(n9048), .B(n8840), .ZN(n6418) );
  INV_X1 U8198 ( .A(n6416), .ZN(n6417) );
  OAI21_X1 U8199 ( .B1(n6418), .B2(n9565), .A(n6417), .ZN(n6820) );
  AOI211_X1 U8200 ( .C1(n9809), .C2(n6828), .A(n6822), .B(n6820), .ZN(n6534)
         );
  AOI22_X1 U8201 ( .A1(n9676), .A2(n6419), .B1(n9814), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n6420) );
  OAI21_X1 U8202 ( .B1(n6534), .B2(n9814), .A(n6420), .ZN(P1_U3525) );
  OAI21_X1 U8203 ( .B1(n6422), .B2(n6426), .A(n6421), .ZN(n6555) );
  INV_X1 U8204 ( .A(n6424), .ZN(n6425) );
  AOI211_X1 U8205 ( .C1(n6430), .C2(n4867), .A(n9570), .B(n6425), .ZN(n6549)
         );
  XNOR2_X1 U8206 ( .A(n6427), .B(n6426), .ZN(n6429) );
  OAI21_X1 U8207 ( .B1(n6429), .B2(n9565), .A(n6428), .ZN(n6548) );
  AOI211_X1 U8208 ( .C1(n9809), .C2(n6555), .A(n6549), .B(n6548), .ZN(n6501)
         );
  AOI22_X1 U8209 ( .A1(n9676), .A2(n6430), .B1(n9814), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6431) );
  OAI21_X1 U8210 ( .B1(n6501), .B2(n9814), .A(n6431), .ZN(P1_U3526) );
  OAI21_X1 U8211 ( .B1(n6434), .B2(n6433), .A(n6432), .ZN(n6545) );
  AOI211_X1 U8212 ( .C1(n6464), .C2(n6440), .A(n9570), .B(n4869), .ZN(n6541)
         );
  XNOR2_X1 U8213 ( .A(n8842), .B(n6436), .ZN(n6439) );
  INV_X1 U8214 ( .A(n6437), .ZN(n6438) );
  OAI21_X1 U8215 ( .B1(n6439), .B2(n9565), .A(n6438), .ZN(n6539) );
  AOI211_X1 U8216 ( .C1(n9809), .C2(n6545), .A(n6541), .B(n6539), .ZN(n6538)
         );
  AOI22_X1 U8217 ( .A1(n9676), .A2(n6440), .B1(n9814), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n6441) );
  OAI21_X1 U8218 ( .B1(n6538), .B2(n9814), .A(n6441), .ZN(P1_U3523) );
  INV_X1 U8219 ( .A(n6442), .ZN(n6443) );
  AOI21_X1 U8220 ( .B1(n6445), .B2(n6444), .A(n6443), .ZN(n6452) );
  INV_X1 U8221 ( .A(n6446), .ZN(n6948) );
  INV_X1 U8222 ( .A(n9931), .ZN(n7285) );
  INV_X1 U8223 ( .A(n7855), .ZN(n7796) );
  NAND2_X1 U8224 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9856) );
  INV_X1 U8225 ( .A(n9856), .ZN(n6447) );
  AOI21_X1 U8226 ( .B1(n7796), .B2(n7887), .A(n6447), .ZN(n6449) );
  NAND2_X1 U8227 ( .A1(n7857), .A2(n7889), .ZN(n6448) );
  OAI211_X1 U8228 ( .C1(n7853), .C2(n7285), .A(n6449), .B(n6448), .ZN(n6450)
         );
  AOI21_X1 U8229 ( .B1(n6948), .B2(n7850), .A(n6450), .ZN(n6451) );
  OAI21_X1 U8230 ( .B1(n6452), .B2(n7861), .A(n6451), .ZN(P2_U3170) );
  OAI222_X1 U8231 ( .A1(n8014), .A2(P2_U3151), .B1(n7151), .B2(n6454), .C1(
        n6453), .C2(n7236), .ZN(P2_U3278) );
  INV_X1 U8232 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U8233 ( .A1(n9106), .A2(n6456), .ZN(n6457) );
  NAND2_X1 U8234 ( .A1(n9804), .A2(n6457), .ZN(n6461) );
  AND3_X1 U8235 ( .A1(n6459), .A2(n9736), .A3(n6458), .ZN(n6460) );
  NAND2_X1 U8236 ( .A1(n6461), .A2(n6460), .ZN(n6462) );
  OR2_X1 U8237 ( .A1(n9802), .A2(n9039), .ZN(n9532) );
  NOR2_X1 U8238 ( .A1(n9532), .A2(n9570), .ZN(n9503) );
  OR2_X2 U8239 ( .A1(n9802), .A2(n6463), .ZN(n9795) );
  INV_X1 U8240 ( .A(n9795), .ZN(n6821) );
  OAI21_X1 U8241 ( .B1(n9503), .B2(n6821), .A(n6464), .ZN(n6472) );
  INV_X1 U8242 ( .A(n9104), .ZN(n6466) );
  NAND3_X1 U8243 ( .A1(n8841), .A2(n6466), .A3(n6465), .ZN(n6468) );
  OAI211_X1 U8244 ( .C1(n9433), .C2(n6469), .A(n6468), .B(n6467), .ZN(n6470)
         );
  NAND2_X1 U8245 ( .A1(n6470), .A2(n6473), .ZN(n6471) );
  OAI211_X1 U8246 ( .C1(n6474), .C2(n6473), .A(n6472), .B(n6471), .ZN(P1_U3293) );
  NAND2_X1 U8247 ( .A1(n6477), .A2(n6476), .ZN(n6481) );
  OR2_X1 U8248 ( .A1(n6478), .A2(n8836), .ZN(n6480) );
  AOI22_X1 U8249 ( .A1(n7575), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7574), .B2(
        n9204), .ZN(n6479) );
  NAND2_X1 U8250 ( .A1(n6480), .A2(n6479), .ZN(n6579) );
  OR2_X1 U8251 ( .A1(n6579), .A2(n6508), .ZN(n8925) );
  NAND2_X1 U8252 ( .A1(n6579), .A2(n6508), .ZN(n8927) );
  NAND2_X1 U8253 ( .A1(n8925), .A2(n8927), .ZN(n6484) );
  NAND2_X1 U8254 ( .A1(n6481), .A2(n6484), .ZN(n6581) );
  OAI21_X1 U8255 ( .B1(n6481), .B2(n6484), .A(n6581), .ZN(n6607) );
  AOI211_X1 U8256 ( .C1(n6579), .C2(n6482), .A(n9570), .B(n6583), .ZN(n6606)
         );
  XNOR2_X1 U8257 ( .A(n6878), .B(n6484), .ZN(n6492) );
  NAND2_X1 U8258 ( .A1(n6486), .A2(n6485), .ZN(n6487) );
  AND2_X1 U8259 ( .A1(n6517), .A2(n6487), .ZN(n6585) );
  NAND2_X1 U8260 ( .A1(n4443), .A2(n6585), .ZN(n6491) );
  NAND2_X1 U8261 ( .A1(n8867), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8262 ( .A1(n6062), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U8263 ( .A1(n4333), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6488) );
  AOI22_X1 U8264 ( .A1(n9136), .A2(n9259), .B1(n8804), .B2(n9138), .ZN(n6661)
         );
  OAI21_X1 U8265 ( .B1(n6492), .B2(n9565), .A(n6661), .ZN(n6601) );
  AOI211_X1 U8266 ( .C1(n9809), .C2(n6607), .A(n6606), .B(n6601), .ZN(n6561)
         );
  AOI22_X1 U8267 ( .A1(n9676), .A2(n6579), .B1(n9814), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n6493) );
  OAI21_X1 U8268 ( .B1(n6561), .B2(n9814), .A(n6493), .ZN(P1_U3528) );
  INV_X1 U8269 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6494) );
  OAI22_X1 U8270 ( .A1(n9722), .A2(n6596), .B1(n9725), .B2(n6494), .ZN(n6495)
         );
  INV_X1 U8271 ( .A(n6495), .ZN(n6496) );
  OAI21_X1 U8272 ( .B1(n6497), .B2(n9811), .A(n6496), .ZN(P1_U3468) );
  INV_X1 U8273 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6498) );
  OAI22_X1 U8274 ( .A1(n9722), .A2(n6553), .B1(n9725), .B2(n6498), .ZN(n6499)
         );
  INV_X1 U8275 ( .A(n6499), .ZN(n6500) );
  OAI21_X1 U8276 ( .B1(n6501), .B2(n9811), .A(n6500), .ZN(P1_U3465) );
  NAND2_X1 U8277 ( .A1(n6579), .A2(n8646), .ZN(n6506) );
  OR2_X1 U8278 ( .A1(n6508), .A2(n8541), .ZN(n6505) );
  NAND2_X1 U8279 ( .A1(n6506), .A2(n6505), .ZN(n6507) );
  INV_X1 U8280 ( .A(n6508), .ZN(n9137) );
  AOI22_X1 U8281 ( .A1(n6579), .A2(n8640), .B1(n9137), .B2(n8567), .ZN(n6510)
         );
  AND2_X1 U8282 ( .A1(n6509), .A2(n6510), .ZN(n6658) );
  OR2_X1 U8283 ( .A1(n6511), .A2(n8836), .ZN(n6513) );
  AOI22_X1 U8284 ( .A1(n7575), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7574), .B2(
        n9219), .ZN(n6512) );
  NAND2_X2 U8285 ( .A1(n6513), .A2(n6512), .ZN(n8929) );
  AOI22_X1 U8286 ( .A1(n8929), .A2(n8646), .B1(n8640), .B2(n9136), .ZN(n6514)
         );
  XNOR2_X1 U8287 ( .A(n6514), .B(n8565), .ZN(n6967) );
  AOI22_X1 U8288 ( .A1(n8929), .A2(n8496), .B1(n8567), .B2(n9136), .ZN(n6968)
         );
  XNOR2_X1 U8289 ( .A(n6967), .B(n6968), .ZN(n6515) );
  XNOR2_X1 U8290 ( .A(n6969), .B(n6515), .ZN(n6526) );
  NAND2_X1 U8291 ( .A1(n8867), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U8292 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  NAND2_X1 U8293 ( .A1(n6749), .A2(n6518), .ZN(n6980) );
  INV_X1 U8294 ( .A(n6980), .ZN(n6862) );
  NAND2_X1 U8295 ( .A1(n4443), .A2(n6862), .ZN(n6521) );
  NAND2_X1 U8296 ( .A1(n8868), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8297 ( .A1(n4333), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6519) );
  AOI22_X1 U8298 ( .A1(n9259), .A2(n4758), .B1(n9137), .B2(n8804), .ZN(n6577)
         );
  NAND2_X1 U8299 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9213) );
  NAND2_X1 U8300 ( .A1(n8825), .A2(n6585), .ZN(n6523) );
  OAI211_X1 U8301 ( .C1(n6577), .C2(n8822), .A(n9213), .B(n6523), .ZN(n6524)
         );
  AOI21_X1 U8302 ( .B1(n8929), .B2(n8784), .A(n6524), .ZN(n6525) );
  OAI21_X1 U8303 ( .B1(n6526), .B2(n8786), .A(n6525), .ZN(P1_U3213) );
  INV_X1 U8304 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6527) );
  OAI22_X1 U8305 ( .A1(n9722), .A2(n9796), .B1(n9725), .B2(n6527), .ZN(n6528)
         );
  INV_X1 U8306 ( .A(n6528), .ZN(n6529) );
  OAI21_X1 U8307 ( .B1(n6530), .B2(n9811), .A(n6529), .ZN(P1_U3459) );
  INV_X1 U8308 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6531) );
  OAI22_X1 U8309 ( .A1(n9722), .A2(n6826), .B1(n9725), .B2(n6531), .ZN(n6532)
         );
  INV_X1 U8310 ( .A(n6532), .ZN(n6533) );
  OAI21_X1 U8311 ( .B1(n6534), .B2(n9811), .A(n6533), .ZN(P1_U3462) );
  OAI22_X1 U8312 ( .A1(n9722), .A2(n9045), .B1(n9725), .B2(n6535), .ZN(n6536)
         );
  INV_X1 U8313 ( .A(n6536), .ZN(n6537) );
  OAI21_X1 U8314 ( .B1(n6538), .B2(n9811), .A(n6537), .ZN(P1_U3456) );
  INV_X1 U8315 ( .A(n6539), .ZN(n6547) );
  AND2_X1 U8316 ( .A1(n9560), .A2(n9553), .ZN(n6540) );
  INV_X2 U8317 ( .A(n9532), .ZN(n9790) );
  NAND2_X1 U8318 ( .A1(n6541), .A2(n9790), .ZN(n6543) );
  INV_X2 U8319 ( .A(n9433), .ZN(n9792) );
  AOI22_X1 U8320 ( .A1(n9802), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9792), .ZN(n6542) );
  OAI211_X1 U8321 ( .C1(n9045), .C2(n9795), .A(n6543), .B(n6542), .ZN(n6544)
         );
  AOI21_X1 U8322 ( .B1(n9799), .B2(n6545), .A(n6544), .ZN(n6546) );
  OAI21_X1 U8323 ( .B1(n9802), .B2(n6547), .A(n6546), .ZN(P1_U3292) );
  INV_X1 U8324 ( .A(n6548), .ZN(n6557) );
  NAND2_X1 U8325 ( .A1(n6549), .A2(n9790), .ZN(n6552) );
  AOI22_X1 U8326 ( .A1(n9802), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6550), .B2(
        n9792), .ZN(n6551) );
  OAI211_X1 U8327 ( .C1(n6553), .C2(n9795), .A(n6552), .B(n6551), .ZN(n6554)
         );
  AOI21_X1 U8328 ( .B1(n9799), .B2(n6555), .A(n6554), .ZN(n6556) );
  OAI21_X1 U8329 ( .B1(n9802), .B2(n6557), .A(n6556), .ZN(P1_U3289) );
  NAND2_X1 U8330 ( .A1(n7871), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6558) );
  OAI21_X1 U8331 ( .B1(n8073), .B2(n7871), .A(n6558), .ZN(P2_U3520) );
  INV_X1 U8332 ( .A(n6579), .ZN(n6666) );
  INV_X1 U8333 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10135) );
  OAI22_X1 U8334 ( .A1(n6666), .A2(n9722), .B1(n9725), .B2(n10135), .ZN(n6559)
         );
  INV_X1 U8335 ( .A(n6559), .ZN(n6560) );
  OAI21_X1 U8336 ( .B1(n6561), .B2(n9811), .A(n6560), .ZN(P1_U3471) );
  INV_X1 U8337 ( .A(n6562), .ZN(n6564) );
  OAI21_X1 U8338 ( .B1(n6564), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6563), .ZN(
        n6569) );
  XNOR2_X1 U8339 ( .A(n6566), .B(n6565), .ZN(n6567) );
  OAI22_X1 U8340 ( .A1(n9911), .A2(n6567), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6930), .ZN(n6568) );
  AOI21_X1 U8341 ( .B1(n9901), .B2(n6569), .A(n6568), .ZN(n6575) );
  OAI21_X1 U8342 ( .B1(n6571), .B2(P2_REG2_REG_1__SCAN_IN), .A(n6570), .ZN(
        n6572) );
  AOI22_X1 U8343 ( .A1(n6573), .A2(n9826), .B1(n9916), .B2(n6572), .ZN(n6574)
         );
  OAI211_X1 U8344 ( .C1(n9981), .C2(n9882), .A(n6575), .B(n6574), .ZN(P2_U3183) );
  NAND2_X1 U8345 ( .A1(n6878), .A2(n8925), .ZN(n6576) );
  NAND2_X1 U8346 ( .A1(n6576), .A2(n8927), .ZN(n6745) );
  XNOR2_X1 U8347 ( .A(n8929), .B(n8930), .ZN(n6743) );
  XNOR2_X1 U8348 ( .A(n6745), .B(n6743), .ZN(n6578) );
  OAI21_X1 U8349 ( .B1(n6578), .B2(n9565), .A(n6577), .ZN(n6614) );
  INV_X1 U8350 ( .A(n6614), .ZN(n6590) );
  NAND2_X1 U8351 ( .A1(n6508), .A2(n6666), .ZN(n6580) );
  NAND2_X1 U8352 ( .A1(n6581), .A2(n6580), .ZN(n6582) );
  OAI21_X1 U8353 ( .B1(n6582), .B2(n6743), .A(n6736), .ZN(n6616) );
  INV_X1 U8354 ( .A(n6583), .ZN(n6584) );
  AOI211_X1 U8355 ( .C1(n8929), .C2(n6584), .A(n9570), .B(n6740), .ZN(n6615)
         );
  NAND2_X1 U8356 ( .A1(n6615), .A2(n9790), .ZN(n6587) );
  AOI22_X1 U8357 ( .A1(n9802), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6585), .B2(
        n9792), .ZN(n6586) );
  OAI211_X1 U8358 ( .C1(n8932), .C2(n9795), .A(n6587), .B(n6586), .ZN(n6588)
         );
  AOI21_X1 U8359 ( .B1(n6616), .B2(n9799), .A(n6588), .ZN(n6589) );
  OAI21_X1 U8360 ( .B1(n9802), .B2(n6590), .A(n6589), .ZN(P1_U3286) );
  INV_X1 U8361 ( .A(n6591), .ZN(n6600) );
  NAND2_X1 U8362 ( .A1(n6592), .A2(n9790), .ZN(n6595) );
  AOI22_X1 U8363 ( .A1(n9802), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6593), .B2(
        n9792), .ZN(n6594) );
  OAI211_X1 U8364 ( .C1(n6596), .C2(n9795), .A(n6595), .B(n6594), .ZN(n6597)
         );
  AOI21_X1 U8365 ( .B1(n6598), .B2(n9799), .A(n6597), .ZN(n6599) );
  OAI21_X1 U8366 ( .B1(n9802), .B2(n6600), .A(n6599), .ZN(P1_U3288) );
  INV_X1 U8367 ( .A(n6601), .ZN(n6610) );
  NOR2_X1 U8368 ( .A1(n9795), .A2(n6666), .ZN(n6605) );
  INV_X1 U8369 ( .A(n6663), .ZN(n6602) );
  OAI22_X1 U8370 ( .A1(n6473), .A2(n6603), .B1(n6602), .B2(n9433), .ZN(n6604)
         );
  AOI211_X1 U8371 ( .C1(n6606), .C2(n9790), .A(n6605), .B(n6604), .ZN(n6609)
         );
  NAND2_X1 U8372 ( .A1(n6607), .A2(n9799), .ZN(n6608) );
  OAI211_X1 U8373 ( .C1(n6610), .C2(n9802), .A(n6609), .B(n6608), .ZN(P1_U3287) );
  INV_X1 U8374 ( .A(n7489), .ZN(n6712) );
  NAND2_X1 U8375 ( .A1(n6611), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6612) );
  XNOR2_X1 U8376 ( .A(n6612), .B(P1_IR_REG_18__SCAN_IN), .ZN(n7490) );
  AOI22_X1 U8377 ( .A1(n7490), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9740), .ZN(n6613) );
  OAI21_X1 U8378 ( .B1(n6712), .B2(n9747), .A(n6613), .ZN(P1_U3337) );
  AOI211_X1 U8379 ( .C1(n9809), .C2(n6616), .A(n6615), .B(n6614), .ZN(n6621)
         );
  AOI22_X1 U8380 ( .A1(n8929), .A2(n9676), .B1(n9814), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n6617) );
  OAI21_X1 U8381 ( .B1(n6621), .B2(n9814), .A(n6617), .ZN(P1_U3529) );
  INV_X1 U8382 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6618) );
  OAI22_X1 U8383 ( .A1(n8932), .A2(n9722), .B1(n9725), .B2(n6618), .ZN(n6619)
         );
  INV_X1 U8384 ( .A(n6619), .ZN(n6620) );
  OAI21_X1 U8385 ( .B1(n6621), .B2(n9811), .A(n6620), .ZN(P1_U3474) );
  MUX2_X1 U8386 ( .A(n6623), .B(n6622), .S(n8041), .Z(n6628) );
  INV_X1 U8387 ( .A(n6624), .ZN(n6625) );
  AOI22_X1 U8388 ( .A1(n6627), .A2(n6626), .B1(n6644), .B2(n6625), .ZN(n9886)
         );
  XNOR2_X1 U8389 ( .A(n6628), .B(n6647), .ZN(n9885) );
  NOR2_X1 U8390 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  AOI21_X1 U8391 ( .B1(n6647), .B2(n6628), .A(n9884), .ZN(n9910) );
  INV_X1 U8392 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9972) );
  MUX2_X1 U8393 ( .A(n6648), .B(n9972), .S(n8041), .Z(n6629) );
  NAND2_X1 U8394 ( .A1(n6629), .A2(n6649), .ZN(n6630) );
  OAI21_X1 U8395 ( .B1(n6649), .B2(n6629), .A(n6630), .ZN(n9909) );
  NOR2_X1 U8396 ( .A1(n9910), .A2(n9909), .ZN(n9908) );
  INV_X1 U8397 ( .A(n6630), .ZN(n6631) );
  NOR2_X1 U8398 ( .A1(n9908), .A2(n6631), .ZN(n6633) );
  MUX2_X1 U8399 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8041), .Z(n7004) );
  XNOR2_X1 U8400 ( .A(n7004), .B(n4505), .ZN(n6632) );
  NOR2_X1 U8401 ( .A1(n6633), .A2(n6632), .ZN(n7005) );
  AOI21_X1 U8402 ( .B1(n6633), .B2(n6632), .A(n7005), .ZN(n6654) );
  NAND2_X1 U8403 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7028) );
  OAI21_X1 U8404 ( .B1(n9906), .B2(n4505), .A(n7028), .ZN(n6642) );
  NAND2_X1 U8405 ( .A1(n6634), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6635) );
  NAND2_X1 U8406 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  OR2_X1 U8407 ( .A1(n6637), .A2(n9876), .ZN(n6638) );
  NAND2_X1 U8408 ( .A1(n6637), .A2(n9876), .ZN(n9898) );
  XNOR2_X1 U8409 ( .A(n6649), .B(n9972), .ZN(n9899) );
  NOR2_X1 U8410 ( .A1(n6639), .A2(n5151), .ZN(n7014) );
  AOI21_X1 U8411 ( .B1(n5151), .B2(n6639), .A(n7014), .ZN(n6640) );
  NOR2_X1 U8412 ( .A1(n6640), .A2(n8000), .ZN(n6641) );
  AOI211_X1 U8413 ( .C1(n9897), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n6642), .B(
        n6641), .ZN(n6653) );
  INV_X1 U8414 ( .A(n6645), .ZN(n6646) );
  XNOR2_X1 U8415 ( .A(n6649), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n9915) );
  NOR2_X1 U8416 ( .A1(n6650), .A2(n5156), .ZN(n6999) );
  AOI21_X1 U8417 ( .B1(n5156), .B2(n6650), .A(n6999), .ZN(n6651) );
  OR2_X1 U8418 ( .A1(n6651), .A2(n9891), .ZN(n6652) );
  OAI211_X1 U8419 ( .C1(n6654), .C2(n9911), .A(n6653), .B(n6652), .ZN(P2_U3191) );
  INV_X1 U8420 ( .A(n6969), .ZN(n6971) );
  NOR2_X1 U8421 ( .A1(n4425), .A2(n6655), .ZN(n6657) );
  OAI22_X1 U8422 ( .A1(n6971), .A2(n6658), .B1(n6657), .B2(n6656), .ZN(n6659)
         );
  NAND2_X1 U8423 ( .A1(n6659), .A2(n8816), .ZN(n6665) );
  INV_X1 U8424 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6660) );
  OAI22_X1 U8425 ( .A1(n6661), .A2(n8822), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6660), .ZN(n6662) );
  AOI21_X1 U8426 ( .B1(n6663), .B2(n8825), .A(n6662), .ZN(n6664) );
  OAI211_X1 U8427 ( .C1(n6666), .C2(n8828), .A(n6665), .B(n6664), .ZN(P1_U3239) );
  XNOR2_X1 U8428 ( .A(n7887), .B(n6667), .ZN(n7435) );
  XOR2_X1 U8429 ( .A(n6668), .B(n7435), .Z(n9939) );
  INV_X1 U8430 ( .A(n6670), .ZN(n6669) );
  NAND2_X1 U8431 ( .A1(n5662), .A2(n6669), .ZN(n6673) );
  NAND2_X1 U8432 ( .A1(n6671), .A2(n6670), .ZN(n6672) );
  AND2_X1 U8433 ( .A1(n6673), .A2(n6672), .ZN(n6674) );
  NAND2_X1 U8434 ( .A1(n6675), .A2(n6674), .ZN(n6682) );
  NAND2_X1 U8435 ( .A1(n6676), .A2(n7266), .ZN(n6714) );
  OR2_X1 U8436 ( .A1(n8269), .A2(n6714), .ZN(n8068) );
  XNOR2_X1 U8437 ( .A(n6677), .B(n7435), .ZN(n6680) );
  OAI22_X1 U8438 ( .A1(n6678), .A2(n8276), .B1(n6811), .B2(n8278), .ZN(n6679)
         );
  AOI21_X1 U8439 ( .B1(n6680), .B2(n8214), .A(n6679), .ZN(n6681) );
  OAI21_X1 U8440 ( .B1(n9939), .B2(n7134), .A(n6681), .ZN(n9941) );
  NAND2_X1 U8441 ( .A1(n9941), .A2(n8282), .ZN(n6685) );
  OAI22_X1 U8442 ( .A1(n8230), .A2(n9937), .B1(n6698), .B2(n8279), .ZN(n6683)
         );
  AOI21_X1 U8443 ( .B1(n8269), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6683), .ZN(
        n6684) );
  OAI211_X1 U8444 ( .C1(n9939), .C2(n8068), .A(n6685), .B(n6684), .ZN(P2_U3228) );
  INV_X1 U8445 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6691) );
  INV_X1 U8446 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6688) );
  OAI21_X1 U8447 ( .B1(n6688), .B2(n6687), .A(n6686), .ZN(n6784) );
  XNOR2_X1 U8448 ( .A(n6789), .B(n6784), .ZN(n6689) );
  NAND2_X1 U8449 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n6689), .ZN(n6785) );
  OAI211_X1 U8450 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n6689), .A(n9779), .B(
        n6785), .ZN(n6690) );
  NAND2_X1 U8451 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8821) );
  OAI211_X1 U8452 ( .C1(n9788), .C2(n6691), .A(n6690), .B(n8821), .ZN(n6696)
         );
  INV_X1 U8453 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6694) );
  AOI21_X1 U8454 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7548), .A(n6692), .ZN(
        n6790) );
  XOR2_X1 U8455 ( .A(n6790), .B(n7560), .Z(n6693) );
  NOR2_X1 U8456 ( .A1(n6694), .A2(n6693), .ZN(n6791) );
  AOI211_X1 U8457 ( .C1(n6694), .C2(n6693), .A(n6791), .B(n9241), .ZN(n6695)
         );
  AOI211_X1 U8458 ( .C1(n9781), .C2(n7560), .A(n6696), .B(n6695), .ZN(n6697)
         );
  INV_X1 U8459 ( .A(n6697), .ZN(P1_U3258) );
  INV_X1 U8460 ( .A(n6698), .ZN(n6709) );
  NAND2_X1 U8461 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9874) );
  INV_X1 U8462 ( .A(n9874), .ZN(n6699) );
  AOI21_X1 U8463 ( .B1(n7796), .B2(n7886), .A(n6699), .ZN(n6701) );
  NAND2_X1 U8464 ( .A1(n7857), .A2(n7888), .ZN(n6700) );
  OAI211_X1 U8465 ( .C1(n7853), .C2(n9937), .A(n6701), .B(n6700), .ZN(n6708)
         );
  INV_X1 U8466 ( .A(n6703), .ZN(n6705) );
  NAND3_X1 U8467 ( .A1(n6442), .A2(n6705), .A3(n6704), .ZN(n6706) );
  AOI21_X1 U8468 ( .B1(n6702), .B2(n6706), .A(n7861), .ZN(n6707) );
  AOI211_X1 U8469 ( .C1(n6709), .C2(n7850), .A(n6708), .B(n6707), .ZN(n6710)
         );
  INV_X1 U8470 ( .A(n6710), .ZN(P2_U3167) );
  INV_X1 U8471 ( .A(n6711), .ZN(n8039) );
  OAI222_X1 U8472 ( .A1(n7236), .A2(n6713), .B1(n7151), .B2(n6712), .C1(
        P2_U3151), .C2(n8039), .ZN(P2_U3277) );
  AND2_X1 U8473 ( .A1(n7134), .A2(n6714), .ZN(n6715) );
  INV_X1 U8474 ( .A(n6716), .ZN(n6718) );
  INV_X1 U8475 ( .A(n4359), .ZN(n7430) );
  INV_X1 U8476 ( .A(n7272), .ZN(n6717) );
  AOI21_X1 U8477 ( .B1(n6718), .B2(n7430), .A(n6717), .ZN(n9928) );
  XNOR2_X1 U8478 ( .A(n6719), .B(n4359), .ZN(n6720) );
  OAI22_X1 U8479 ( .A1(n8279), .A2(n6259), .B1(n9927), .B2(n8255), .ZN(n6722)
         );
  NOR2_X1 U8480 ( .A1(n9929), .A2(n6722), .ZN(n6723) );
  INV_X2 U8481 ( .A(n8269), .ZN(n8282) );
  MUX2_X1 U8482 ( .A(n6724), .B(n6723), .S(n8282), .Z(n6725) );
  OAI21_X1 U8483 ( .B1(n8287), .B2(n9928), .A(n6725), .ZN(P2_U3231) );
  INV_X1 U8484 ( .A(n7850), .ZN(n7859) );
  OAI211_X1 U8485 ( .C1(n6728), .C2(n6727), .A(n6726), .B(n7845), .ZN(n6735)
         );
  INV_X1 U8486 ( .A(n6729), .ZN(n6730) );
  AOI21_X1 U8487 ( .B1(n7796), .B2(n7885), .A(n6730), .ZN(n6732) );
  NAND2_X1 U8488 ( .A1(n7857), .A2(n7887), .ZN(n6731) );
  OAI211_X1 U8489 ( .C1(n7853), .C2(n6802), .A(n6732), .B(n6731), .ZN(n6733)
         );
  INV_X1 U8490 ( .A(n6733), .ZN(n6734) );
  OAI211_X1 U8491 ( .C1(n6766), .C2(n7859), .A(n6735), .B(n6734), .ZN(P2_U3179) );
  AOI22_X1 U8492 ( .A1(n7575), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7574), .B2(
        n9231), .ZN(n6738) );
  NAND2_X1 U8493 ( .A1(n8935), .A2(n6974), .ZN(n8933) );
  NAND2_X1 U8494 ( .A1(n8931), .A2(n8933), .ZN(n6747) );
  OAI21_X1 U8495 ( .B1(n6739), .B2(n6747), .A(n6853), .ZN(n6866) );
  INV_X1 U8496 ( .A(n6740), .ZN(n6742) );
  NAND2_X1 U8497 ( .A1(n6740), .A2(n6985), .ZN(n6839) );
  INV_X1 U8498 ( .A(n6839), .ZN(n6741) );
  AOI211_X1 U8499 ( .C1(n8935), .C2(n6742), .A(n9570), .B(n6741), .ZN(n6861)
         );
  INV_X1 U8500 ( .A(n6743), .ZN(n6744) );
  NAND2_X1 U8501 ( .A1(n6745), .A2(n6744), .ZN(n6746) );
  NAND2_X1 U8502 ( .A1(n8929), .A2(n8930), .ZN(n8926) );
  NAND2_X1 U8503 ( .A1(n6746), .A2(n8926), .ZN(n6832) );
  XNOR2_X1 U8504 ( .A(n6832), .B(n6747), .ZN(n6755) );
  NAND2_X1 U8505 ( .A1(n8867), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6753) );
  NOR2_X1 U8506 ( .A1(n6840), .A2(n4388), .ZN(n8741) );
  NAND2_X1 U8507 ( .A1(n4443), .A2(n8741), .ZN(n6752) );
  NAND2_X1 U8508 ( .A1(n8868), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6751) );
  NAND2_X1 U8509 ( .A1(n4333), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6750) );
  OAI22_X1 U8510 ( .A1(n8930), .A2(n9281), .B1(n8448), .B2(n8819), .ZN(n6982)
         );
  INV_X1 U8511 ( .A(n6982), .ZN(n6754) );
  OAI21_X1 U8512 ( .B1(n6755), .B2(n9565), .A(n6754), .ZN(n6860) );
  AOI211_X1 U8513 ( .C1(n6866), .C2(n9809), .A(n6861), .B(n6860), .ZN(n6760)
         );
  AOI22_X1 U8514 ( .A1(n8935), .A2(n9676), .B1(n9814), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n6756) );
  OAI21_X1 U8515 ( .B1(n6760), .B2(n9814), .A(n6756), .ZN(P1_U3530) );
  INV_X1 U8516 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6757) );
  OAI22_X1 U8517 ( .A1(n6985), .A2(n9722), .B1(n9725), .B2(n6757), .ZN(n6758)
         );
  INV_X1 U8518 ( .A(n6758), .ZN(n6759) );
  OAI21_X1 U8519 ( .B1(n6760), .B2(n9811), .A(n6759), .ZN(P1_U3477) );
  NAND2_X1 U8520 ( .A1(n6761), .A2(n7278), .ZN(n6762) );
  XNOR2_X1 U8521 ( .A(n6762), .B(n7439), .ZN(n6780) );
  XNOR2_X1 U8522 ( .A(n6763), .B(n7439), .ZN(n6764) );
  AOI222_X1 U8523 ( .A1(n8214), .A2(n6764), .B1(n7885), .B2(n8211), .C1(n7887), 
        .C2(n8209), .ZN(n6779) );
  MUX2_X1 U8524 ( .A(n6765), .B(n6779), .S(n8282), .Z(n6770) );
  INV_X1 U8525 ( .A(n6766), .ZN(n6767) );
  AOI22_X1 U8526 ( .A1(n8284), .A2(n6768), .B1(n8218), .B2(n6767), .ZN(n6769)
         );
  OAI211_X1 U8527 ( .C1(n8287), .C2(n6780), .A(n6770), .B(n6769), .ZN(P2_U3227) );
  INV_X1 U8528 ( .A(n6771), .ZN(n6772) );
  NOR2_X1 U8529 ( .A1(n4992), .A2(n8278), .ZN(n8361) );
  AOI21_X1 U8530 ( .B1(n6772), .B2(n8360), .A(n8361), .ZN(n6773) );
  OAI21_X1 U8531 ( .B1(n8279), .B2(n6774), .A(n6773), .ZN(n6775) );
  MUX2_X1 U8532 ( .A(n6775), .B(P2_REG2_REG_0__SCAN_IN), .S(n8269), .Z(n6776)
         );
  AOI21_X1 U8533 ( .B1(n8284), .B2(n6777), .A(n6776), .ZN(n6778) );
  INV_X1 U8534 ( .A(n6778), .ZN(P2_U3233) );
  OAI21_X1 U8535 ( .B1(n9959), .B2(n6780), .A(n6779), .ZN(n6804) );
  INV_X1 U8536 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6781) );
  OAI22_X1 U8537 ( .A1(n8357), .A2(n6802), .B1(n10192), .B2(n6781), .ZN(n6782)
         );
  AOI21_X1 U8538 ( .B1(n6804), .B2(n10192), .A(n6782), .ZN(n6783) );
  INV_X1 U8539 ( .A(n6783), .ZN(P2_U3465) );
  NAND2_X1 U8540 ( .A1(n7560), .A2(n6784), .ZN(n6786) );
  NAND2_X1 U8541 ( .A1(n6786), .A2(n6785), .ZN(n6788) );
  XNOR2_X1 U8542 ( .A(n7514), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n6787) );
  NOR2_X1 U8543 ( .A1(n6787), .A2(n6788), .ZN(n7104) );
  AOI21_X1 U8544 ( .B1(n6788), .B2(n6787), .A(n7104), .ZN(n6800) );
  NOR2_X1 U8545 ( .A1(n6790), .A2(n6789), .ZN(n6792) );
  NOR2_X1 U8546 ( .A1(n6792), .A2(n6791), .ZN(n6795) );
  NAND2_X1 U8547 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7514), .ZN(n6793) );
  OAI21_X1 U8548 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n7514), .A(n6793), .ZN(
        n6794) );
  NOR2_X1 U8549 ( .A1(n6795), .A2(n6794), .ZN(n7113) );
  AOI211_X1 U8550 ( .C1(n6795), .C2(n6794), .A(n7113), .B(n9241), .ZN(n6796)
         );
  INV_X1 U8551 ( .A(n6796), .ZN(n6799) );
  AND2_X1 U8552 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8712) );
  NOR2_X1 U8553 ( .A1(n9767), .A2(n7105), .ZN(n6797) );
  AOI211_X1 U8554 ( .C1(n9230), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n8712), .B(
        n6797), .ZN(n6798) );
  OAI211_X1 U8555 ( .C1(n6800), .C2(n7196), .A(n6799), .B(n6798), .ZN(P1_U3259) );
  INV_X1 U8556 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6801) );
  OAI22_X1 U8557 ( .A1(n6802), .A2(n8420), .B1(n9965), .B2(n6801), .ZN(n6803)
         );
  AOI21_X1 U8558 ( .B1(n6804), .B2(n9965), .A(n6803), .ZN(n6805) );
  INV_X1 U8559 ( .A(n6805), .ZN(P2_U3408) );
  OR2_X1 U8560 ( .A1(n6807), .A2(n7441), .ZN(n6808) );
  AND2_X1 U8561 ( .A1(n6806), .A2(n6808), .ZN(n6963) );
  XNOR2_X1 U8562 ( .A(n6809), .B(n7441), .ZN(n6810) );
  OAI222_X1 U8563 ( .A1(n8278), .A2(n7085), .B1(n8276), .B2(n6811), .C1(n8358), 
        .C2(n6810), .ZN(n6958) );
  AOI21_X1 U8564 ( .B1(n6963), .B2(n9933), .A(n6958), .ZN(n6816) );
  AOI22_X1 U8565 ( .A1(n5656), .A2(n6960), .B1(n10190), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n6812) );
  OAI21_X1 U8566 ( .B1(n6816), .B2(n10190), .A(n6812), .ZN(P2_U3466) );
  INV_X1 U8567 ( .A(n6960), .ZN(n6908) );
  INV_X1 U8568 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6813) );
  OAI22_X1 U8569 ( .A1(n6908), .A2(n8420), .B1(n9965), .B2(n6813), .ZN(n6814)
         );
  INV_X1 U8570 ( .A(n6814), .ZN(n6815) );
  OAI21_X1 U8571 ( .B1(n6816), .B2(n9966), .A(n6815), .ZN(P2_U3411) );
  INV_X1 U8572 ( .A(n7573), .ZN(n6818) );
  OAI222_X1 U8573 ( .A1(P2_U3151), .A2(n8046), .B1(n7151), .B2(n6818), .C1(
        n6817), .C2(n7236), .ZN(P2_U3276) );
  OAI222_X1 U8574 ( .A1(n9750), .A2(n6819), .B1(n9747), .B2(n6818), .C1(
        P1_U3086), .C2(n9035), .ZN(P1_U3336) );
  INV_X1 U8575 ( .A(n6820), .ZN(n6830) );
  NAND2_X1 U8576 ( .A1(n6822), .A2(n9790), .ZN(n6825) );
  AOI22_X1 U8577 ( .A1(n9802), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9792), .B2(
        n6823), .ZN(n6824) );
  OAI211_X1 U8578 ( .C1(n6826), .C2(n9795), .A(n6825), .B(n6824), .ZN(n6827)
         );
  AOI21_X1 U8579 ( .B1(n9799), .B2(n6828), .A(n6827), .ZN(n6829) );
  OAI21_X1 U8580 ( .B1(n6830), .B2(n9802), .A(n6829), .ZN(P1_U3290) );
  INV_X1 U8581 ( .A(n8933), .ZN(n6831) );
  OAI21_X1 U8582 ( .B1(n6832), .B2(n6831), .A(n8931), .ZN(n6837) );
  NAND2_X1 U8583 ( .A1(n6833), .A2(n8861), .ZN(n6836) );
  AOI22_X1 U8584 ( .A1(n7575), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7574), .B2(
        n6834), .ZN(n6835) );
  OR2_X1 U8585 ( .A1(n8450), .A2(n8448), .ZN(n8946) );
  NAND2_X1 U8586 ( .A1(n8450), .A2(n8448), .ZN(n8942) );
  NAND2_X1 U8587 ( .A1(n8946), .A2(n8942), .ZN(n8941) );
  XNOR2_X1 U8588 ( .A(n6837), .B(n8941), .ZN(n6838) );
  NAND2_X1 U8589 ( .A1(n6838), .A2(n9526), .ZN(n6851) );
  AOI21_X1 U8590 ( .B1(n6839), .B2(n8450), .A(n9570), .ZN(n6849) );
  OR2_X2 U8591 ( .A1(n6839), .A2(n8450), .ZN(n6894) );
  NAND2_X1 U8592 ( .A1(n8867), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6845) );
  OR2_X1 U8593 ( .A1(n6840), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6841) );
  AND2_X1 U8594 ( .A1(n6841), .A2(n6887), .ZN(n8623) );
  NAND2_X1 U8595 ( .A1(n4443), .A2(n8623), .ZN(n6844) );
  NAND2_X1 U8596 ( .A1(n8868), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U8597 ( .A1(n4333), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6842) );
  OR2_X1 U8598 ( .A1(n8461), .A2(n8819), .ZN(n6847) );
  OR2_X1 U8599 ( .A1(n6974), .A2(n9281), .ZN(n6846) );
  AND2_X1 U8600 ( .A1(n6847), .A2(n6846), .ZN(n8739) );
  INV_X1 U8601 ( .A(n8739), .ZN(n6848) );
  AOI21_X1 U8602 ( .B1(n6849), .B2(n6894), .A(n6848), .ZN(n6850) );
  NAND2_X1 U8603 ( .A1(n6851), .A2(n6850), .ZN(n9807) );
  OAI21_X1 U8604 ( .B1(n6851), .B2(n9573), .A(n9532), .ZN(n6858) );
  INV_X1 U8605 ( .A(n8450), .ZN(n9806) );
  NAND2_X1 U8606 ( .A1(n6854), .A2(n8941), .ZN(n6870) );
  OAI21_X1 U8607 ( .B1(n6854), .B2(n8941), .A(n6870), .ZN(n9810) );
  NAND2_X1 U8608 ( .A1(n9810), .A2(n9799), .ZN(n6856) );
  AOI22_X1 U8609 ( .A1(n9573), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8741), .B2(
        n9792), .ZN(n6855) );
  OAI211_X1 U8610 ( .C1(n9806), .C2(n9795), .A(n6856), .B(n6855), .ZN(n6857)
         );
  AOI21_X1 U8611 ( .B1(n9807), .B2(n6858), .A(n6857), .ZN(n6859) );
  INV_X1 U8612 ( .A(n6859), .ZN(P1_U3284) );
  INV_X1 U8613 ( .A(n6860), .ZN(n6868) );
  NAND2_X1 U8614 ( .A1(n6861), .A2(n9790), .ZN(n6864) );
  AOI22_X1 U8615 ( .A1(n9573), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6862), .B2(
        n9792), .ZN(n6863) );
  OAI211_X1 U8616 ( .C1(n6985), .C2(n9795), .A(n6864), .B(n6863), .ZN(n6865)
         );
  AOI21_X1 U8617 ( .B1(n6866), .B2(n9799), .A(n6865), .ZN(n6867) );
  OAI21_X1 U8618 ( .B1(n9573), .B2(n6868), .A(n6867), .ZN(P1_U3285) );
  INV_X1 U8619 ( .A(n8448), .ZN(n9135) );
  AOI22_X1 U8620 ( .A1(n7575), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7574), .B2(
        n6872), .ZN(n6873) );
  OR2_X1 U8621 ( .A1(n8624), .A2(n8461), .ZN(n9055) );
  OAI21_X1 U8622 ( .B1(n6875), .B2(n6886), .A(n7526), .ZN(n6914) );
  INV_X1 U8623 ( .A(n6914), .ZN(n6900) );
  NAND2_X1 U8624 ( .A1(n8946), .A2(n8931), .ZN(n6881) );
  AND2_X1 U8625 ( .A1(n8933), .A2(n8926), .ZN(n6876) );
  INV_X1 U8626 ( .A(n8927), .ZN(n6877) );
  INV_X1 U8627 ( .A(n8925), .ZN(n6880) );
  OR2_X1 U8628 ( .A1(n8929), .A2(n8930), .ZN(n8919) );
  INV_X1 U8629 ( .A(n8919), .ZN(n6879) );
  INV_X1 U8630 ( .A(n6885), .ZN(n6883) );
  INV_X1 U8631 ( .A(n9557), .ZN(n6884) );
  AOI21_X1 U8632 ( .B1(n6886), .B2(n6885), .A(n6884), .ZN(n6893) );
  NAND2_X1 U8633 ( .A1(n8867), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8634 ( .A1(n6887), .A2(n10078), .ZN(n6888) );
  AND2_X1 U8635 ( .A1(n7538), .A2(n6888), .ZN(n9572) );
  NAND2_X1 U8636 ( .A1(n4443), .A2(n9572), .ZN(n6891) );
  NAND2_X1 U8637 ( .A1(n8868), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U8638 ( .A1(n4333), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6889) );
  INV_X1 U8639 ( .A(n8689), .ZN(n9133) );
  AOI22_X1 U8640 ( .A1(n8804), .A2(n9135), .B1(n9133), .B2(n9259), .ZN(n8621)
         );
  OAI21_X1 U8641 ( .B1(n6893), .B2(n9565), .A(n8621), .ZN(n6912) );
  INV_X1 U8642 ( .A(n8624), .ZN(n6897) );
  AOI211_X1 U8643 ( .C1(n8624), .C2(n6894), .A(n9570), .B(n9567), .ZN(n6913)
         );
  NAND2_X1 U8644 ( .A1(n6913), .A2(n9790), .ZN(n6896) );
  AOI22_X1 U8645 ( .A1(n9802), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8623), .B2(
        n9792), .ZN(n6895) );
  OAI211_X1 U8646 ( .C1(n6897), .C2(n9795), .A(n6896), .B(n6895), .ZN(n6898)
         );
  AOI21_X1 U8647 ( .B1(n6912), .B2(n6473), .A(n6898), .ZN(n6899) );
  OAI21_X1 U8648 ( .B1(n6900), .B2(n9551), .A(n6899), .ZN(P1_U3283) );
  INV_X1 U8649 ( .A(n6993), .ZN(n6901) );
  AOI21_X1 U8650 ( .B1(n6903), .B2(n6902), .A(n6901), .ZN(n6911) );
  INV_X1 U8651 ( .A(n6904), .ZN(n6959) );
  NAND2_X1 U8652 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9895) );
  INV_X1 U8653 ( .A(n9895), .ZN(n6905) );
  AOI21_X1 U8654 ( .B1(n7796), .B2(n7884), .A(n6905), .ZN(n6907) );
  NAND2_X1 U8655 ( .A1(n7857), .A2(n7886), .ZN(n6906) );
  OAI211_X1 U8656 ( .C1(n7853), .C2(n6908), .A(n6907), .B(n6906), .ZN(n6909)
         );
  AOI21_X1 U8657 ( .B1(n6959), .B2(n7850), .A(n6909), .ZN(n6910) );
  OAI21_X1 U8658 ( .B1(n6911), .B2(n7861), .A(n6910), .ZN(P2_U3153) );
  AOI211_X1 U8659 ( .C1(n6914), .C2(n9809), .A(n6913), .B(n6912), .ZN(n6919)
         );
  INV_X1 U8660 ( .A(n9722), .ZN(n9732) );
  INV_X1 U8661 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6915) );
  NOR2_X1 U8662 ( .A1(n9725), .A2(n6915), .ZN(n6916) );
  AOI21_X1 U8663 ( .B1(n8624), .B2(n9732), .A(n6916), .ZN(n6917) );
  OAI21_X1 U8664 ( .B1(n6919), .B2(n9811), .A(n6917), .ZN(P1_U3483) );
  AOI22_X1 U8665 ( .A1(n8624), .A2(n9676), .B1(n9814), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n6918) );
  OAI21_X1 U8666 ( .B1(n6919), .B2(n9814), .A(n6918), .ZN(P1_U3532) );
  NAND2_X1 U8667 ( .A1(n6806), .A2(n6920), .ZN(n6921) );
  AND2_X1 U8668 ( .A1(n7295), .A2(n7304), .ZN(n7443) );
  XNOR2_X1 U8669 ( .A(n6921), .B(n7443), .ZN(n9942) );
  XOR2_X1 U8670 ( .A(n6922), .B(n7443), .Z(n6923) );
  OAI222_X1 U8671 ( .A1(n8278), .A2(n6925), .B1(n8276), .B2(n6924), .C1(n6923), 
        .C2(n8358), .ZN(n9943) );
  NAND2_X1 U8672 ( .A1(n9943), .A2(n8282), .ZN(n6928) );
  OAI22_X1 U8673 ( .A1(n8282), .A2(n6648), .B1(n6987), .B2(n8279), .ZN(n6926)
         );
  AOI21_X1 U8674 ( .B1(n8284), .B2(n9945), .A(n6926), .ZN(n6927) );
  OAI211_X1 U8675 ( .C1(n9942), .C2(n8287), .A(n6928), .B(n6927), .ZN(P2_U3225) );
  XNOR2_X1 U8676 ( .A(n6929), .B(n7431), .ZN(n9925) );
  OAI22_X1 U8677 ( .A1(n8230), .A2(n9923), .B1(n8279), .B2(n6930), .ZN(n6931)
         );
  AOI21_X1 U8678 ( .B1(n8267), .B2(n9925), .A(n6931), .ZN(n6937) );
  OAI21_X1 U8679 ( .B1(n6933), .B2(n7431), .A(n6932), .ZN(n6935) );
  AOI222_X1 U8680 ( .A1(n8214), .A2(n6935), .B1(n6934), .B2(n8209), .C1(n7890), 
        .C2(n8211), .ZN(n9922) );
  MUX2_X1 U8681 ( .A(n9922), .B(n10089), .S(n8269), .Z(n6936) );
  NAND2_X1 U8682 ( .A1(n6937), .A2(n6936), .ZN(P2_U3232) );
  INV_X1 U8683 ( .A(n7585), .ZN(n6939) );
  OAI222_X1 U8684 ( .A1(n6938), .A2(P2_U3151), .B1(n7151), .B2(n6939), .C1(
        n10075), .C2(n7236), .ZN(P2_U3275) );
  INV_X1 U8685 ( .A(n7434), .ZN(n6944) );
  XNOR2_X1 U8686 ( .A(n6940), .B(n6944), .ZN(n6941) );
  NAND2_X1 U8687 ( .A1(n6941), .A2(n8214), .ZN(n6943) );
  AOI22_X1 U8688 ( .A1(n8209), .A2(n7889), .B1(n7887), .B2(n8211), .ZN(n6942)
         );
  AND2_X1 U8689 ( .A1(n6943), .A2(n6942), .ZN(n9936) );
  NAND3_X1 U8690 ( .A1(n6945), .A2(n6944), .A3(n7284), .ZN(n6946) );
  NAND2_X1 U8691 ( .A1(n6947), .A2(n6946), .ZN(n9934) );
  AOI22_X1 U8692 ( .A1(n8284), .A2(n9931), .B1(n8218), .B2(n6948), .ZN(n6949)
         );
  OAI21_X1 U8693 ( .B1(n6348), .B2(n8282), .A(n6949), .ZN(n6950) );
  AOI21_X1 U8694 ( .B1(n8267), .B2(n9934), .A(n6950), .ZN(n6951) );
  OAI21_X1 U8695 ( .B1(n8269), .B2(n9936), .A(n6951), .ZN(P2_U3229) );
  OAI22_X1 U8696 ( .A1(n8230), .A2(n6952), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8279), .ZN(n6955) );
  MUX2_X1 U8697 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6953), .S(n8282), .Z(n6954)
         );
  AOI211_X1 U8698 ( .C1(n8267), .C2(n6956), .A(n6955), .B(n6954), .ZN(n6957)
         );
  INV_X1 U8699 ( .A(n6957), .ZN(P2_U3230) );
  INV_X1 U8700 ( .A(n6958), .ZN(n6965) );
  AOI22_X1 U8701 ( .A1(n8284), .A2(n6960), .B1(n8218), .B2(n6959), .ZN(n6961)
         );
  OAI21_X1 U8702 ( .B1(n6623), .B2(n8282), .A(n6961), .ZN(n6962) );
  AOI21_X1 U8703 ( .B1(n6963), .B2(n8267), .A(n6962), .ZN(n6964) );
  OAI21_X1 U8704 ( .B1(n6965), .B2(n8269), .A(n6964), .ZN(P2_U3226) );
  NOR2_X1 U8705 ( .A1(n6974), .A2(n8641), .ZN(n6966) );
  AOI21_X1 U8706 ( .B1(n8935), .B2(n8496), .A(n6966), .ZN(n8452) );
  INV_X1 U8707 ( .A(n6968), .ZN(n6972) );
  AOI21_X1 U8708 ( .B1(n6969), .B2(n6968), .A(n6967), .ZN(n6970) );
  NAND2_X1 U8709 ( .A1(n8935), .A2(n8646), .ZN(n6976) );
  OR2_X1 U8710 ( .A1(n6974), .A2(n8541), .ZN(n6975) );
  NAND2_X1 U8711 ( .A1(n6976), .A2(n6975), .ZN(n6977) );
  XNOR2_X1 U8712 ( .A(n6977), .B(n8644), .ZN(n8451) );
  INV_X1 U8713 ( .A(n8451), .ZN(n8454) );
  NOR2_X1 U8714 ( .A1(n8455), .A2(n8454), .ZN(n8733) );
  AOI21_X1 U8715 ( .B1(n8455), .B2(n8454), .A(n8733), .ZN(n6978) );
  NAND2_X1 U8716 ( .A1(n6978), .A2(n8452), .ZN(n8736) );
  OAI21_X1 U8717 ( .B1(n8452), .B2(n6978), .A(n8736), .ZN(n6979) );
  NAND2_X1 U8718 ( .A1(n6979), .A2(n8816), .ZN(n6984) );
  AND2_X1 U8719 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9229) );
  NOR2_X1 U8720 ( .A1(n8808), .A2(n6980), .ZN(n6981) );
  AOI211_X1 U8721 ( .C1(n8810), .C2(n6982), .A(n9229), .B(n6981), .ZN(n6983)
         );
  OAI211_X1 U8722 ( .C1(n6985), .C2(n8828), .A(n6984), .B(n6983), .ZN(P1_U3221) );
  NAND2_X1 U8723 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9920) );
  INV_X1 U8724 ( .A(n9920), .ZN(n6986) );
  AOI21_X1 U8725 ( .B1(n7796), .B2(n7883), .A(n6986), .ZN(n6991) );
  INV_X1 U8726 ( .A(n6987), .ZN(n6988) );
  NAND2_X1 U8727 ( .A1(n7850), .A2(n6988), .ZN(n6990) );
  NAND2_X1 U8728 ( .A1(n7857), .A2(n7885), .ZN(n6989) );
  NAND3_X1 U8729 ( .A1(n6991), .A2(n6990), .A3(n6989), .ZN(n6997) );
  NAND3_X1 U8730 ( .A1(n6993), .A2(n4424), .A3(n6992), .ZN(n6994) );
  AOI21_X1 U8731 ( .B1(n6995), .B2(n6994), .A(n7861), .ZN(n6996) );
  AOI211_X1 U8732 ( .C1(n9945), .C2(n7866), .A(n6997), .B(n6996), .ZN(n6998)
         );
  INV_X1 U8733 ( .A(n6998), .ZN(P2_U3161) );
  NAND2_X1 U8734 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7170), .ZN(n7001) );
  OAI21_X1 U8735 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7170), .A(n7001), .ZN(
        n7002) );
  AOI21_X1 U8736 ( .B1(n7003), .B2(n7002), .A(n7162), .ZN(n7023) );
  INV_X1 U8737 ( .A(n7004), .ZN(n7006) );
  AOI21_X1 U8738 ( .B1(n7007), .B2(n7006), .A(n7005), .ZN(n7011) );
  MUX2_X1 U8739 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8041), .Z(n7008) );
  NOR2_X1 U8740 ( .A1(n7008), .A2(n7170), .ZN(n7154) );
  AOI21_X1 U8741 ( .B1(n7170), .B2(n7008), .A(n7154), .ZN(n7009) );
  INV_X1 U8742 ( .A(n7009), .ZN(n7010) );
  NOR2_X1 U8743 ( .A1(n7011), .A2(n7010), .ZN(n7153) );
  AOI21_X1 U8744 ( .B1(n7011), .B2(n7010), .A(n7153), .ZN(n7012) );
  NOR2_X1 U8745 ( .A1(n7012), .A2(n9911), .ZN(n7021) );
  INV_X1 U8746 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7013) );
  NOR2_X1 U8747 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7013), .ZN(n7226) );
  NAND2_X1 U8748 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7170), .ZN(n7015) );
  OAI21_X1 U8749 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7170), .A(n7015), .ZN(
        n7016) );
  AOI21_X1 U8750 ( .B1(n7017), .B2(n7016), .A(n7169), .ZN(n7018) );
  NOR2_X1 U8751 ( .A1(n7018), .A2(n8000), .ZN(n7020) );
  INV_X1 U8752 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7036) );
  OAI22_X1 U8753 ( .A1(n9906), .A2(n7170), .B1(n9882), .B2(n7036), .ZN(n7019)
         );
  NOR4_X1 U8754 ( .A1(n7021), .A2(n7226), .A3(n7020), .A4(n7019), .ZN(n7022)
         );
  OAI21_X1 U8755 ( .B1(n7023), .B2(n9891), .A(n7022), .ZN(P2_U3192) );
  OAI211_X1 U8756 ( .C1(n7026), .C2(n7025), .A(n7024), .B(n7845), .ZN(n7033)
         );
  INV_X1 U8757 ( .A(n7027), .ZN(n7090) );
  NAND2_X1 U8758 ( .A1(n7857), .A2(n7884), .ZN(n7029) );
  OAI211_X1 U8759 ( .C1(n7086), .C2(n7855), .A(n7029), .B(n7028), .ZN(n7031)
         );
  INV_X1 U8760 ( .A(n7101), .ZN(n7098) );
  NOR2_X1 U8761 ( .A1(n7853), .A2(n7098), .ZN(n7030) );
  AOI211_X1 U8762 ( .C1(n7090), .C2(n7850), .A(n7031), .B(n7030), .ZN(n7032)
         );
  NAND2_X1 U8763 ( .A1(n7033), .A2(n7032), .ZN(P2_U3171) );
  INV_X1 U8764 ( .A(n7597), .ZN(n7035) );
  INV_X1 U8765 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7598) );
  OAI222_X1 U8766 ( .A1(P1_U3086), .A2(n9044), .B1(n9747), .B2(n7035), .C1(
        n7598), .C2(n9750), .ZN(P1_U3334) );
  INV_X1 U8767 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7034) );
  OAI222_X1 U8768 ( .A1(n7417), .A2(P2_U3151), .B1(n7151), .B2(n7035), .C1(
        n7034), .C2(n7236), .ZN(P2_U3274) );
  NOR2_X1 U8769 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7078) );
  NOR2_X1 U8770 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7075) );
  NOR2_X1 U8771 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7071) );
  NOR2_X1 U8772 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7068) );
  NOR2_X1 U8773 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7065) );
  NOR2_X1 U8774 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7062) );
  INV_X1 U8775 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7180) );
  AOI22_X1 U8776 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n6084), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7180), .ZN(n9996) );
  NAND2_X1 U8777 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7060) );
  INV_X1 U8778 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7211) );
  AOI22_X1 U8779 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .B1(n5920), .B2(n7211), .ZN(n9998) );
  NAND2_X1 U8780 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7058) );
  XNOR2_X1 U8781 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n7036), .ZN(n10000) );
  NOR2_X1 U8782 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7042) );
  XNOR2_X1 U8783 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10208) );
  NAND2_X1 U8784 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7040) );
  XNOR2_X1 U8785 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n10014), .ZN(n10206) );
  NAND2_X1 U8786 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7038) );
  XOR2_X1 U8787 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10204) );
  AOI21_X1 U8788 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9977) );
  NAND3_X1 U8789 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9979) );
  OAI21_X1 U8790 ( .B1(n9977), .B2(n9981), .A(n9979), .ZN(n10203) );
  NAND2_X1 U8791 ( .A1(n10204), .A2(n10203), .ZN(n7037) );
  NAND2_X1 U8792 ( .A1(n7038), .A2(n7037), .ZN(n10205) );
  NAND2_X1 U8793 ( .A1(n10206), .A2(n10205), .ZN(n7039) );
  NAND2_X1 U8794 ( .A1(n7040), .A2(n7039), .ZN(n10207) );
  NOR2_X1 U8795 ( .A1(n10208), .A2(n10207), .ZN(n7041) );
  NOR2_X1 U8796 ( .A1(n7042), .A2(n7041), .ZN(n7043) );
  NOR2_X1 U8797 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7043), .ZN(n10197) );
  AND2_X1 U8798 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7043), .ZN(n10196) );
  NOR2_X1 U8799 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10196), .ZN(n7044) );
  NOR2_X1 U8800 ( .A1(n10197), .A2(n7044), .ZN(n7045) );
  NAND2_X1 U8801 ( .A1(n7045), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7047) );
  XOR2_X1 U8802 ( .A(n7045), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10195) );
  NAND2_X1 U8803 ( .A1(n10195), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7046) );
  NAND2_X1 U8804 ( .A1(n7047), .A2(n7046), .ZN(n7048) );
  NAND2_X1 U8805 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7048), .ZN(n7050) );
  XOR2_X1 U8806 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7048), .Z(n10201) );
  NAND2_X1 U8807 ( .A1(n10201), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7049) );
  NAND2_X1 U8808 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  NAND2_X1 U8809 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7051), .ZN(n7053) );
  XOR2_X1 U8810 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7051), .Z(n10202) );
  NAND2_X1 U8811 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10202), .ZN(n7052) );
  NAND2_X1 U8812 ( .A1(n7053), .A2(n7052), .ZN(n7054) );
  NAND2_X1 U8813 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7054), .ZN(n7056) );
  INV_X1 U8814 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9771) );
  XNOR2_X1 U8815 ( .A(n9771), .B(n7054), .ZN(n10200) );
  NAND2_X1 U8816 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10200), .ZN(n7055) );
  NAND2_X1 U8817 ( .A1(n7056), .A2(n7055), .ZN(n9999) );
  NAND2_X1 U8818 ( .A1(n10000), .A2(n9999), .ZN(n7057) );
  NAND2_X1 U8819 ( .A1(n7058), .A2(n7057), .ZN(n9997) );
  NAND2_X1 U8820 ( .A1(n9998), .A2(n9997), .ZN(n7059) );
  NAND2_X1 U8821 ( .A1(n7060), .A2(n7059), .ZN(n9995) );
  INV_X1 U8822 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7063) );
  INV_X1 U8823 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7906) );
  AOI22_X1 U8824 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n7063), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n7906), .ZN(n9993) );
  NOR2_X1 U8825 ( .A1(n9994), .A2(n9993), .ZN(n7064) );
  NOR2_X1 U8826 ( .A1(n7065), .A2(n7064), .ZN(n9992) );
  INV_X1 U8827 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7066) );
  AOI22_X1 U8828 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n6242), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n7066), .ZN(n9991) );
  NOR2_X1 U8829 ( .A1(n9992), .A2(n9991), .ZN(n7067) );
  NOR2_X1 U8830 ( .A1(n7068), .A2(n7067), .ZN(n9990) );
  INV_X1 U8831 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7069) );
  AOI22_X1 U8832 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n6691), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n7069), .ZN(n9989) );
  NOR2_X1 U8833 ( .A1(n9990), .A2(n9989), .ZN(n7070) );
  NOR2_X1 U8834 ( .A1(n7071), .A2(n7070), .ZN(n9988) );
  INV_X1 U8835 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7073) );
  INV_X1 U8836 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7072) );
  AOI22_X1 U8837 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7073), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n7072), .ZN(n9987) );
  NOR2_X1 U8838 ( .A1(n9988), .A2(n9987), .ZN(n7074) );
  NOR2_X1 U8839 ( .A1(n7075), .A2(n7074), .ZN(n9986) );
  INV_X1 U8840 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9789) );
  INV_X1 U8841 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7076) );
  AOI22_X1 U8842 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9789), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n7076), .ZN(n9985) );
  NOR2_X1 U8843 ( .A1(n9986), .A2(n9985), .ZN(n7077) );
  NOR2_X1 U8844 ( .A1(n7078), .A2(n7077), .ZN(n7079) );
  AND2_X1 U8845 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7079), .ZN(n9983) );
  NOR2_X1 U8846 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n9983), .ZN(n7080) );
  NOR2_X1 U8847 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7079), .ZN(n9982) );
  NOR2_X1 U8848 ( .A1(n7080), .A2(n9982), .ZN(n7082) );
  XNOR2_X1 U8849 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7081) );
  XNOR2_X1 U8850 ( .A(n7082), .B(n7081), .ZN(ADD_1068_U4) );
  XOR2_X1 U8851 ( .A(n7445), .B(n7083), .Z(n7084) );
  OAI222_X1 U8852 ( .A1(n8278), .A2(n7086), .B1(n8276), .B2(n7085), .C1(n8358), 
        .C2(n7084), .ZN(n7095) );
  NAND2_X1 U8853 ( .A1(n7087), .A2(n7445), .ZN(n7088) );
  AND2_X1 U8854 ( .A1(n7089), .A2(n7088), .ZN(n7096) );
  NAND2_X1 U8855 ( .A1(n7096), .A2(n8267), .ZN(n7092) );
  AOI22_X1 U8856 ( .A1(n8269), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n8218), .B2(
        n7090), .ZN(n7091) );
  OAI211_X1 U8857 ( .C1(n7098), .C2(n8230), .A(n7092), .B(n7091), .ZN(n7093)
         );
  AOI21_X1 U8858 ( .B1(n7095), .B2(n8282), .A(n7093), .ZN(n7094) );
  INV_X1 U8859 ( .A(n7094), .ZN(P2_U3224) );
  AOI21_X1 U8860 ( .B1(n7096), .B2(n9933), .A(n7095), .ZN(n7103) );
  INV_X1 U8861 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7097) );
  OAI22_X1 U8862 ( .A1(n7098), .A2(n8420), .B1(n9965), .B2(n7097), .ZN(n7099)
         );
  INV_X1 U8863 ( .A(n7099), .ZN(n7100) );
  OAI21_X1 U8864 ( .B1(n7103), .B2(n9966), .A(n7100), .ZN(P2_U3417) );
  AOI22_X1 U8865 ( .A1(n5656), .A2(n7101), .B1(n10190), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7102) );
  OAI21_X1 U8866 ( .B1(n7103), .B2(n10190), .A(n7102), .ZN(P2_U3468) );
  INV_X1 U8867 ( .A(n7490), .ZN(n7126) );
  XNOR2_X1 U8868 ( .A(n7490), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n7111) );
  INV_X1 U8869 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9641) );
  XNOR2_X1 U8870 ( .A(n9780), .B(n9641), .ZN(n9777) );
  INV_X1 U8871 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7106) );
  AOI21_X1 U8872 ( .B1(n7106), .B2(n7105), .A(n7104), .ZN(n7107) );
  INV_X1 U8873 ( .A(n7107), .ZN(n9776) );
  NAND2_X1 U8874 ( .A1(n9777), .A2(n9776), .ZN(n9775) );
  OR2_X1 U8875 ( .A1(n9780), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U8876 ( .A1(n9775), .A2(n7108), .ZN(n7110) );
  INV_X1 U8877 ( .A(n7194), .ZN(n7109) );
  AOI211_X1 U8878 ( .C1(n7111), .C2(n7110), .A(n7109), .B(n7196), .ZN(n7124)
         );
  NAND2_X1 U8879 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8795) );
  INV_X1 U8880 ( .A(n8795), .ZN(n7123) );
  INV_X1 U8881 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n7112) );
  NOR2_X1 U8882 ( .A1(n9788), .A2(n7112), .ZN(n7122) );
  AOI21_X1 U8883 ( .B1(n7514), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7113), .ZN(
        n9773) );
  INV_X1 U8884 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7114) );
  XNOR2_X1 U8885 ( .A(n9780), .B(n7114), .ZN(n9774) );
  NAND2_X1 U8886 ( .A1(n9773), .A2(n9774), .ZN(n9772) );
  OR2_X1 U8887 ( .A1(n9780), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7115) );
  NAND2_X1 U8888 ( .A1(n9772), .A2(n7115), .ZN(n7120) );
  INV_X1 U8889 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7116) );
  OR2_X1 U8890 ( .A1(n7490), .A2(n7116), .ZN(n7118) );
  NAND2_X1 U8891 ( .A1(n7490), .A2(n7116), .ZN(n7117) );
  AND2_X1 U8892 ( .A1(n7118), .A2(n7117), .ZN(n7119) );
  NOR2_X1 U8893 ( .A1(n7120), .A2(n7119), .ZN(n7191) );
  AOI211_X1 U8894 ( .C1(n7120), .C2(n7119), .A(n7191), .B(n9241), .ZN(n7121)
         );
  NOR4_X1 U8895 ( .A1(n7124), .A2(n7123), .A3(n7122), .A4(n7121), .ZN(n7125)
         );
  OAI21_X1 U8896 ( .B1(n7126), .B2(n9767), .A(n7125), .ZN(P1_U3261) );
  INV_X1 U8897 ( .A(n7315), .ZN(n7127) );
  OR2_X1 U8898 ( .A1(n7300), .A2(n7127), .ZN(n7446) );
  INV_X1 U8899 ( .A(n7446), .ZN(n7128) );
  XNOR2_X1 U8900 ( .A(n7129), .B(n7128), .ZN(n9946) );
  XOR2_X1 U8901 ( .A(n7130), .B(n7446), .Z(n7131) );
  NAND2_X1 U8902 ( .A1(n7131), .A2(n8214), .ZN(n7133) );
  AOI22_X1 U8903 ( .A1(n7881), .A2(n8211), .B1(n8209), .B2(n7883), .ZN(n7132)
         );
  OAI211_X1 U8904 ( .C1(n9946), .C2(n7134), .A(n7133), .B(n7132), .ZN(n9949)
         );
  NAND2_X1 U8905 ( .A1(n9949), .A2(n8282), .ZN(n7139) );
  OAI22_X1 U8906 ( .A1(n8282), .A2(n7135), .B1(n7225), .B2(n8279), .ZN(n7136)
         );
  AOI21_X1 U8907 ( .B1(n8284), .B2(n7137), .A(n7136), .ZN(n7138) );
  OAI211_X1 U8908 ( .C1(n9946), .C2(n8068), .A(n7139), .B(n7138), .ZN(P2_U3223) );
  XNOR2_X1 U8909 ( .A(n7140), .B(n7448), .ZN(n9954) );
  NAND2_X1 U8910 ( .A1(n7142), .A2(n7141), .ZN(n7143) );
  NAND3_X1 U8911 ( .A1(n7144), .A2(n8214), .A3(n7143), .ZN(n7146) );
  AOI22_X1 U8912 ( .A1(n8209), .A2(n7882), .B1(n7880), .B2(n8211), .ZN(n7145)
         );
  NAND2_X1 U8913 ( .A1(n7146), .A2(n7145), .ZN(n9955) );
  NAND2_X1 U8914 ( .A1(n9955), .A2(n8282), .ZN(n7150) );
  OAI22_X1 U8915 ( .A1(n8282), .A2(n7147), .B1(n7822), .B2(n8279), .ZN(n7148)
         );
  AOI21_X1 U8916 ( .B1(n8284), .B2(n9957), .A(n7148), .ZN(n7149) );
  OAI211_X1 U8917 ( .C1(n8287), .C2(n9954), .A(n7150), .B(n7149), .ZN(P2_U3222) );
  INV_X1 U8918 ( .A(n7606), .ZN(n7479) );
  OAI222_X1 U8919 ( .A1(P2_U3151), .A2(n7152), .B1(n7151), .B2(n7479), .C1(
        n10083), .C2(n7236), .ZN(P2_U3273) );
  MUX2_X1 U8920 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8041), .Z(n7155) );
  NOR2_X1 U8921 ( .A1(n7155), .A2(n7212), .ZN(n7157) );
  NOR2_X1 U8922 ( .A1(n7154), .A2(n7153), .ZN(n7214) );
  AOI21_X1 U8923 ( .B1(n7155), .B2(n7212), .A(n7157), .ZN(n7156) );
  INV_X1 U8924 ( .A(n7156), .ZN(n7215) );
  NOR2_X1 U8925 ( .A1(n7214), .A2(n7215), .ZN(n7213) );
  NOR2_X1 U8926 ( .A1(n7157), .A2(n7213), .ZN(n7896) );
  INV_X1 U8927 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7158) );
  MUX2_X1 U8928 ( .A(n8281), .B(n7158), .S(n8041), .Z(n7159) );
  NOR2_X1 U8929 ( .A1(n7159), .A2(n7177), .ZN(n7894) );
  INV_X1 U8930 ( .A(n7894), .ZN(n7160) );
  NAND2_X1 U8931 ( .A1(n7159), .A2(n7177), .ZN(n7895) );
  NAND2_X1 U8932 ( .A1(n7160), .A2(n7895), .ZN(n7161) );
  XNOR2_X1 U8933 ( .A(n7896), .B(n7161), .ZN(n7183) );
  NOR2_X1 U8934 ( .A1(n7171), .A2(n7163), .ZN(n7164) );
  MUX2_X1 U8935 ( .A(n8281), .B(P2_REG2_REG_12__SCAN_IN), .S(n7177), .Z(n7165)
         );
  INV_X1 U8936 ( .A(n7165), .ZN(n7166) );
  NOR2_X1 U8937 ( .A1(n7167), .A2(n7166), .ZN(n7899) );
  AOI21_X1 U8938 ( .B1(n7167), .B2(n7166), .A(n7899), .ZN(n7168) );
  NOR2_X1 U8939 ( .A1(n7168), .A2(n9891), .ZN(n7182) );
  NOR2_X1 U8940 ( .A1(n7171), .A2(n7172), .ZN(n7173) );
  NOR2_X1 U8941 ( .A1(n7173), .A2(n7208), .ZN(n7175) );
  AOI22_X1 U8942 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7177), .B1(n7900), .B2(
        n7158), .ZN(n7174) );
  NOR2_X1 U8943 ( .A1(n7175), .A2(n7174), .ZN(n7892) );
  AOI21_X1 U8944 ( .B1(n7175), .B2(n7174), .A(n7892), .ZN(n7176) );
  OR2_X1 U8945 ( .A1(n7176), .A2(n8000), .ZN(n7179) );
  NOR2_X1 U8946 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10170), .ZN(n7738) );
  AOI21_X1 U8947 ( .B1(n9826), .B2(n7177), .A(n7738), .ZN(n7178) );
  OAI211_X1 U8948 ( .C1(n7180), .C2(n9882), .A(n7179), .B(n7178), .ZN(n7181)
         );
  AOI211_X1 U8949 ( .C1(n7183), .C2(n9867), .A(n7182), .B(n7181), .ZN(n7184)
         );
  INV_X1 U8950 ( .A(n7184), .ZN(P2_U3194) );
  INV_X1 U8951 ( .A(n7618), .ZN(n7187) );
  NAND2_X1 U8952 ( .A1(n7185), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7474) );
  NAND2_X1 U8953 ( .A1(n8438), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7186) );
  OAI211_X1 U8954 ( .C1(n7187), .C2(n7151), .A(n7474), .B(n7186), .ZN(P2_U3272) );
  NAND2_X1 U8955 ( .A1(n7618), .A2(n7188), .ZN(n7189) );
  OAI211_X1 U8956 ( .C1(n7619), .C2(n9750), .A(n7189), .B(n9108), .ZN(P1_U3332) );
  AND2_X1 U8957 ( .A1(n7490), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7190) );
  OR2_X1 U8958 ( .A1(n7191), .A2(n7190), .ZN(n7192) );
  INV_X1 U8959 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9435) );
  XNOR2_X1 U8960 ( .A(n7192), .B(n9435), .ZN(n7200) );
  INV_X1 U8961 ( .A(n7200), .ZN(n7198) );
  NAND2_X1 U8962 ( .A1(n7490), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7193) );
  NAND2_X1 U8963 ( .A1(n7194), .A2(n7193), .ZN(n7195) );
  INV_X1 U8964 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9631) );
  XNOR2_X1 U8965 ( .A(n7195), .B(n9631), .ZN(n7199) );
  OAI21_X1 U8966 ( .B1(n7196), .B2(n7199), .A(n9767), .ZN(n7197) );
  AOI21_X1 U8967 ( .B1(n7198), .B2(n9785), .A(n7197), .ZN(n7202) );
  AOI22_X1 U8968 ( .A1(n7200), .A2(n9785), .B1(n9779), .B2(n7199), .ZN(n7201)
         );
  MUX2_X1 U8969 ( .A(n7202), .B(n7201), .S(n9035), .Z(n7204) );
  NOR2_X1 U8970 ( .A1(n7578), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8637) );
  INV_X1 U8971 ( .A(n8637), .ZN(n7203) );
  OAI211_X1 U8972 ( .C1(n7205), .C2(n9788), .A(n7204), .B(n7203), .ZN(P1_U3262) );
  AOI21_X1 U8973 ( .B1(n7147), .B2(n7207), .A(n7206), .ZN(n7221) );
  AOI21_X1 U8974 ( .B1(n5198), .B2(n7209), .A(n7208), .ZN(n7210) );
  NOR2_X1 U8975 ( .A1(n7210), .A2(n8000), .ZN(n7219) );
  OAI22_X1 U8976 ( .A1(n9906), .A2(n7212), .B1(n9882), .B2(n7211), .ZN(n7218)
         );
  AOI21_X1 U8977 ( .B1(n7215), .B2(n7214), .A(n7213), .ZN(n7216) );
  NAND2_X1 U8978 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7823) );
  OAI21_X1 U8979 ( .B1(n9911), .B2(n7216), .A(n7823), .ZN(n7217) );
  NOR3_X1 U8980 ( .A1(n7219), .A2(n7218), .A3(n7217), .ZN(n7220) );
  OAI21_X1 U8981 ( .B1(n7221), .B2(n9891), .A(n7220), .ZN(P2_U3193) );
  XNOR2_X1 U8982 ( .A(n7222), .B(n7882), .ZN(n7223) );
  NOR2_X1 U8983 ( .A1(n7223), .A2(n7224), .ZN(n7819) );
  AOI21_X1 U8984 ( .B1(n7224), .B2(n7223), .A(n7819), .ZN(n7233) );
  INV_X1 U8985 ( .A(n7225), .ZN(n7231) );
  NAND2_X1 U8986 ( .A1(n7857), .A2(n7883), .ZN(n7228) );
  INV_X1 U8987 ( .A(n7226), .ZN(n7227) );
  OAI211_X1 U8988 ( .C1(n8275), .C2(n7855), .A(n7228), .B(n7227), .ZN(n7230)
         );
  NOR2_X1 U8989 ( .A1(n7853), .A2(n9948), .ZN(n7229) );
  AOI211_X1 U8990 ( .C1(n7231), .C2(n7850), .A(n7230), .B(n7229), .ZN(n7232)
         );
  OAI21_X1 U8991 ( .B1(n7233), .B2(n7861), .A(n7232), .ZN(P2_U3157) );
  INV_X1 U8992 ( .A(n7629), .ZN(n7238) );
  OAI222_X1 U8993 ( .A1(n7234), .A2(P1_U3086), .B1(n9747), .B2(n7238), .C1(
        n7630), .C2(n9750), .ZN(P1_U3331) );
  INV_X1 U8994 ( .A(n7640), .ZN(n7239) );
  AOI22_X1 U8995 ( .A1(n5617), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n8438), .ZN(n7235) );
  OAI21_X1 U8996 ( .B1(n7239), .B2(n7151), .A(n7235), .ZN(P2_U3270) );
  OAI222_X1 U8997 ( .A1(P2_U3151), .A2(n5612), .B1(n7151), .B2(n7238), .C1(
        n7237), .C2(n7236), .ZN(P2_U3271) );
  OAI222_X1 U8998 ( .A1(n7240), .A2(P1_U3086), .B1(n9747), .B2(n7239), .C1(
        n7641), .C2(n9750), .ZN(P1_U3330) );
  INV_X1 U8999 ( .A(n7652), .ZN(n7476) );
  AOI22_X1 U9000 ( .A1(n7241), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8438), .ZN(n7242) );
  OAI21_X1 U9001 ( .B1(n7476), .B2(n7151), .A(n7242), .ZN(P2_U3269) );
  MUX2_X1 U9002 ( .A(n7869), .B(n7243), .S(n7386), .Z(n7373) );
  NAND2_X1 U9003 ( .A1(n8125), .A2(n7244), .ZN(n7252) );
  AND2_X1 U9004 ( .A1(n7247), .A2(n7245), .ZN(n7250) );
  MUX2_X1 U9005 ( .A(n7247), .B(n7246), .S(n7388), .Z(n7248) );
  NAND2_X1 U9006 ( .A1(n8146), .A2(n7248), .ZN(n7355) );
  INV_X1 U9007 ( .A(n7425), .ZN(n7359) );
  OAI211_X1 U9008 ( .C1(n7250), .C2(n7355), .A(n7359), .B(n7249), .ZN(n7251)
         );
  MUX2_X1 U9009 ( .A(n7252), .B(n7251), .S(n7388), .Z(n7357) );
  INV_X1 U9010 ( .A(n7253), .ZN(n7354) );
  INV_X1 U9011 ( .A(n7428), .ZN(n7254) );
  NOR2_X1 U9012 ( .A1(n7426), .A2(n7254), .ZN(n7256) );
  AND2_X1 U9013 ( .A1(n8162), .A2(n7427), .ZN(n7255) );
  MUX2_X1 U9014 ( .A(n7256), .B(n7255), .S(n7388), .Z(n7353) );
  NAND2_X1 U9015 ( .A1(n7346), .A2(n7257), .ZN(n7454) );
  AND2_X1 U9016 ( .A1(n8187), .A2(n7258), .ZN(n7456) );
  INV_X1 U9017 ( .A(n7456), .ZN(n7259) );
  MUX2_X1 U9018 ( .A(n7454), .B(n7259), .S(n7386), .Z(n7352) );
  NAND2_X1 U9019 ( .A1(n7260), .A2(n7284), .ZN(n7263) );
  NAND2_X1 U9020 ( .A1(n7276), .A2(n7261), .ZN(n7262) );
  MUX2_X1 U9021 ( .A(n7263), .B(n7262), .S(n7388), .Z(n7274) );
  AND2_X1 U9022 ( .A1(n7265), .A2(n7264), .ZN(n7267) );
  OAI211_X1 U9023 ( .C1(n7472), .C2(n7267), .A(n4359), .B(n7266), .ZN(n7271)
         );
  INV_X1 U9024 ( .A(n7267), .ZN(n7269) );
  AOI21_X1 U9025 ( .B1(n7269), .B2(n7268), .A(n7386), .ZN(n7270) );
  AOI21_X1 U9026 ( .B1(n7272), .B2(n7271), .A(n7270), .ZN(n7273) );
  OR2_X1 U9027 ( .A1(n7274), .A2(n7273), .ZN(n7275) );
  NAND2_X1 U9028 ( .A1(n7275), .A2(n7434), .ZN(n7289) );
  INV_X1 U9029 ( .A(n7276), .ZN(n7279) );
  OAI211_X1 U9030 ( .C1(n7289), .C2(n7279), .A(n7278), .B(n7277), .ZN(n7283)
         );
  AND2_X1 U9031 ( .A1(n7290), .A2(n7286), .ZN(n7282) );
  INV_X1 U9032 ( .A(n7280), .ZN(n7281) );
  AOI21_X1 U9033 ( .B1(n7283), .B2(n7282), .A(n7281), .ZN(n7294) );
  INV_X1 U9034 ( .A(n7284), .ZN(n7288) );
  NAND2_X1 U9035 ( .A1(n7888), .A2(n7285), .ZN(n7287) );
  OAI211_X1 U9036 ( .C1(n7289), .C2(n7288), .A(n7287), .B(n7286), .ZN(n7292)
         );
  AOI21_X1 U9037 ( .B1(n7292), .B2(n7291), .A(n4766), .ZN(n7293) );
  MUX2_X1 U9038 ( .A(n7294), .B(n7293), .S(n7388), .Z(n7298) );
  AND2_X1 U9039 ( .A1(n7305), .A2(n7304), .ZN(n7297) );
  AND2_X1 U9040 ( .A1(n7301), .A2(n7295), .ZN(n7296) );
  MUX2_X1 U9041 ( .A(n7297), .B(n7296), .S(n7388), .Z(n7299) );
  NAND3_X1 U9042 ( .A1(n7298), .A2(n7299), .A3(n7441), .ZN(n7312) );
  INV_X1 U9043 ( .A(n7299), .ZN(n7307) );
  INV_X1 U9044 ( .A(n7300), .ZN(n7313) );
  OAI211_X1 U9045 ( .C1(n7307), .C2(n7302), .A(n7313), .B(n7301), .ZN(n7309)
         );
  AND2_X1 U9046 ( .A1(n7304), .A2(n7303), .ZN(n7306) );
  OAI211_X1 U9047 ( .C1(n7307), .C2(n7306), .A(n7305), .B(n7315), .ZN(n7308)
         );
  MUX2_X1 U9048 ( .A(n7309), .B(n7308), .S(n7388), .Z(n7310) );
  INV_X1 U9049 ( .A(n7310), .ZN(n7311) );
  NAND2_X1 U9050 ( .A1(n7312), .A2(n7311), .ZN(n7320) );
  NAND2_X1 U9051 ( .A1(n7320), .A2(n7313), .ZN(n7314) );
  AND2_X1 U9052 ( .A1(n7316), .A2(n7315), .ZN(n7319) );
  INV_X1 U9053 ( .A(n7317), .ZN(n7318) );
  AOI21_X1 U9054 ( .B1(n7320), .B2(n7319), .A(n7318), .ZN(n7321) );
  MUX2_X1 U9055 ( .A(n7323), .B(n7322), .S(n7388), .Z(n7324) );
  NAND2_X1 U9056 ( .A1(n7325), .A2(n7324), .ZN(n7328) );
  INV_X1 U9057 ( .A(n7328), .ZN(n7330) );
  INV_X1 U9058 ( .A(n7451), .ZN(n7327) );
  INV_X1 U9059 ( .A(n8260), .ZN(n8421) );
  MUX2_X1 U9060 ( .A(n8277), .B(n8421), .S(n7388), .Z(n7326) );
  OAI21_X1 U9061 ( .B1(n7328), .B2(n7327), .A(n7326), .ZN(n7329) );
  OAI21_X1 U9062 ( .B1(n7330), .B2(n7449), .A(n7329), .ZN(n7331) );
  NAND2_X1 U9063 ( .A1(n7331), .A2(n8251), .ZN(n7335) );
  MUX2_X1 U9064 ( .A(n7333), .B(n7332), .S(n7388), .Z(n7334) );
  NAND2_X1 U9065 ( .A1(n7335), .A2(n7334), .ZN(n7336) );
  NAND2_X1 U9066 ( .A1(n7336), .A2(n8238), .ZN(n7341) );
  NAND3_X1 U9067 ( .A1(n7341), .A2(n7342), .A3(n7337), .ZN(n7339) );
  AND2_X1 U9068 ( .A1(n7344), .A2(n7388), .ZN(n7338) );
  AOI21_X1 U9069 ( .B1(n7339), .B2(n7338), .A(n8215), .ZN(n7351) );
  NAND2_X1 U9070 ( .A1(n7341), .A2(n7340), .ZN(n7343) );
  NAND2_X1 U9071 ( .A1(n7343), .A2(n7342), .ZN(n7345) );
  NAND2_X1 U9072 ( .A1(n7345), .A2(n7344), .ZN(n7348) );
  INV_X1 U9073 ( .A(n7346), .ZN(n7347) );
  AOI21_X1 U9074 ( .B1(n7348), .B2(n7456), .A(n7347), .ZN(n7349) );
  INV_X1 U9075 ( .A(n7363), .ZN(n7365) );
  MUX2_X1 U9076 ( .A(n7365), .B(n7364), .S(n7388), .Z(n7366) );
  MUX2_X1 U9077 ( .A(n7368), .B(n7367), .S(n7386), .Z(n7369) );
  NAND2_X1 U9078 ( .A1(n7370), .A2(n7369), .ZN(n7371) );
  AOI21_X1 U9079 ( .B1(n7462), .B2(n7373), .A(n7374), .ZN(n7383) );
  NAND2_X1 U9080 ( .A1(n7374), .A2(n7373), .ZN(n7384) );
  OAI211_X1 U9081 ( .C1(n7383), .C2(n7869), .A(n7386), .B(n7384), .ZN(n7392)
         );
  INV_X1 U9082 ( .A(n7375), .ZN(n7376) );
  MUX2_X1 U9083 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4338), .Z(n7393) );
  XNOR2_X1 U9084 ( .A(n7393), .B(SI_30_), .ZN(n7394) );
  NAND2_X1 U9085 ( .A1(n8862), .A2(n7401), .ZN(n7381) );
  NAND2_X1 U9086 ( .A1(n5312), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7380) );
  INV_X1 U9087 ( .A(n7868), .ZN(n7387) );
  NAND2_X1 U9088 ( .A1(n7385), .A2(n7387), .ZN(n7463) );
  NAND2_X1 U9089 ( .A1(n7463), .A2(n7382), .ZN(n7415) );
  NOR2_X1 U9090 ( .A1(n7385), .A2(n7387), .ZN(n7465) );
  OAI21_X1 U9091 ( .B1(n7387), .B2(n7386), .A(n7385), .ZN(n7390) );
  OAI21_X1 U9092 ( .B1(n7392), .B2(n7415), .A(n7391), .ZN(n7412) );
  INV_X1 U9093 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7397) );
  INV_X1 U9094 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8829) );
  MUX2_X1 U9095 ( .A(n7397), .B(n8829), .S(n4338), .Z(n7398) );
  XNOR2_X1 U9096 ( .A(n7398), .B(SI_31_), .ZN(n7399) );
  NAND2_X1 U9097 ( .A1(n8831), .A2(n7401), .ZN(n7403) );
  NAND2_X1 U9098 ( .A1(n5312), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7402) );
  INV_X1 U9099 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7408) );
  NAND2_X1 U9100 ( .A1(n7404), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7407) );
  INV_X1 U9101 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7405) );
  OR2_X1 U9102 ( .A1(n4339), .A2(n7405), .ZN(n7406) );
  OAI211_X1 U9103 ( .C1(n7408), .C2(n5020), .A(n7407), .B(n7406), .ZN(n7409)
         );
  INV_X1 U9104 ( .A(n7409), .ZN(n7410) );
  NAND2_X1 U9105 ( .A1(n7412), .A2(n7423), .ZN(n7422) );
  AOI21_X1 U9106 ( .B1(n7468), .B2(n8370), .A(n7467), .ZN(n7416) );
  INV_X1 U9107 ( .A(n7423), .ZN(n7466) );
  INV_X1 U9108 ( .A(n8125), .ZN(n7424) );
  INV_X1 U9109 ( .A(n8135), .ZN(n8131) );
  INV_X1 U9110 ( .A(n7426), .ZN(n8175) );
  INV_X1 U9111 ( .A(n8223), .ZN(n8228) );
  NOR2_X1 U9112 ( .A1(n8360), .A2(n7429), .ZN(n7438) );
  NOR2_X1 U9113 ( .A1(n7431), .A2(n7430), .ZN(n7437) );
  INV_X1 U9114 ( .A(n7432), .ZN(n7433) );
  AND2_X1 U9115 ( .A1(n7434), .A2(n7433), .ZN(n7436) );
  AND4_X1 U9116 ( .A1(n7438), .A2(n7437), .A3(n7436), .A4(n7435), .ZN(n7442)
         );
  INV_X1 U9117 ( .A(n7439), .ZN(n7440) );
  NAND4_X1 U9118 ( .A1(n7443), .A2(n7442), .A3(n7441), .A4(n7440), .ZN(n7444)
         );
  OR3_X1 U9119 ( .A1(n7446), .A2(n7445), .A3(n7444), .ZN(n7447) );
  NOR3_X1 U9120 ( .A1(n8272), .A2(n7448), .A3(n7447), .ZN(n7452) );
  INV_X1 U9121 ( .A(n7449), .ZN(n7450) );
  OR2_X1 U9122 ( .A1(n7451), .A2(n7450), .ZN(n8263) );
  NAND4_X1 U9123 ( .A1(n8238), .A2(n8251), .A3(n7452), .A4(n8263), .ZN(n7453)
         );
  NOR3_X1 U9124 ( .A1(n7454), .A2(n8228), .A3(n7453), .ZN(n7455) );
  NAND4_X1 U9125 ( .A1(n8175), .A2(n8189), .A3(n7456), .A4(n7455), .ZN(n7457)
         );
  NOR2_X1 U9126 ( .A1(n8165), .A2(n7457), .ZN(n7458) );
  NAND4_X1 U9127 ( .A1(n8127), .A2(n8131), .A3(n8146), .A4(n7458), .ZN(n7459)
         );
  OR3_X1 U9128 ( .A1(n8097), .A2(n8112), .A3(n7459), .ZN(n7460) );
  NOR2_X1 U9129 ( .A1(n7460), .A2(n8081), .ZN(n7461) );
  NAND4_X1 U9130 ( .A1(n7463), .A2(n7462), .A3(n7461), .A4(n8074), .ZN(n7464)
         );
  NAND3_X1 U9131 ( .A1(n7470), .A2(n7469), .A3(n8041), .ZN(n7471) );
  OAI211_X1 U9132 ( .C1(n7472), .C2(n7474), .A(n7471), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7473) );
  OAI21_X1 U9133 ( .B1(n7475), .B2(n7474), .A(n7473), .ZN(P2_U3296) );
  OAI222_X1 U9134 ( .A1(n7477), .A2(P1_U3086), .B1(n9747), .B2(n7476), .C1(
        n7653), .C2(n9750), .ZN(P1_U3329) );
  OAI222_X1 U9135 ( .A1(n9750), .A2(n7607), .B1(n9747), .B2(n7479), .C1(
        P1_U3086), .C2(n7478), .ZN(P1_U3333) );
  NAND2_X1 U9136 ( .A1(n8434), .A2(n8861), .ZN(n7481) );
  OR2_X1 U9137 ( .A1(n8864), .A2(n9749), .ZN(n7480) );
  INV_X1 U9138 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7683) );
  OR2_X1 U9139 ( .A1(n8864), .A2(n7689), .ZN(n7482) );
  OR2_X1 U9140 ( .A1(n7658), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n7484) );
  INV_X1 U9141 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U9142 ( .A1(n8867), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7486) );
  NAND2_X1 U9143 ( .A1(n4333), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7485) );
  OAI211_X1 U9144 ( .C1(n7487), .C2(n10158), .A(n7486), .B(n7485), .ZN(n7488)
         );
  INV_X1 U9145 ( .A(n8803), .ZN(n9116) );
  NAND2_X1 U9146 ( .A1(n7489), .A2(n8861), .ZN(n7492) );
  AOI22_X1 U9147 ( .A1(n7575), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7574), .B2(
        n7490), .ZN(n7491) );
  INV_X1 U9148 ( .A(n9634), .ZN(n9446) );
  NAND2_X1 U9149 ( .A1(n7502), .A2(n7493), .ZN(n7494) );
  NAND2_X1 U9150 ( .A1(n7579), .A2(n7494), .ZN(n8794) );
  OR2_X1 U9151 ( .A1(n8794), .A2(n7663), .ZN(n7497) );
  AOI22_X1 U9152 ( .A1(n8867), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6062), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n7496) );
  NAND2_X1 U9153 ( .A1(n4333), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U9154 ( .A1(n7498), .A2(n8861), .ZN(n7500) );
  AOI22_X1 U9155 ( .A1(n7575), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7574), .B2(
        n9780), .ZN(n7499) );
  OR2_X1 U9156 ( .A1(n7507), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7501) );
  AND2_X1 U9157 ( .A1(n7502), .A2(n7501), .ZN(n9467) );
  NAND2_X1 U9158 ( .A1(n9467), .A2(n4443), .ZN(n7505) );
  AOI22_X1 U9159 ( .A1(n8867), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n8868), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U9160 ( .A1(n4333), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7503) );
  INV_X1 U9161 ( .A(n8709), .ZN(n9126) );
  NOR2_X1 U9162 ( .A1(n7566), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7506) );
  OR2_X1 U9163 ( .A1(n7507), .A2(n7506), .ZN(n8710) );
  INV_X1 U9164 ( .A(n8710), .ZN(n9477) );
  NAND2_X1 U9165 ( .A1(n9477), .A2(n4443), .ZN(n7512) );
  NAND2_X1 U9166 ( .A1(n8867), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U9167 ( .A1(n8868), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7508) );
  AND2_X1 U9168 ( .A1(n7509), .A2(n7508), .ZN(n7511) );
  NAND2_X1 U9169 ( .A1(n4333), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U9170 ( .A1(n7513), .A2(n8861), .ZN(n7516) );
  AOI22_X1 U9171 ( .A1(n7575), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7574), .B2(
        n7514), .ZN(n7515) );
  INV_X1 U9172 ( .A(n9645), .ZN(n9479) );
  AOI22_X1 U9173 ( .A1(n7575), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7574), .B2(
        n9248), .ZN(n7518) );
  NAND2_X1 U9174 ( .A1(n8867), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7524) );
  OR2_X1 U9175 ( .A1(n7540), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7520) );
  AND2_X1 U9176 ( .A1(n7552), .A2(n7520), .ZN(n9533) );
  NAND2_X1 U9177 ( .A1(n4443), .A2(n9533), .ZN(n7523) );
  NAND2_X1 U9178 ( .A1(n8868), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7522) );
  NAND2_X1 U9179 ( .A1(n4333), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7521) );
  INV_X1 U9180 ( .A(n8690), .ZN(n9131) );
  INV_X1 U9181 ( .A(n8461), .ZN(n9134) );
  NAND2_X1 U9182 ( .A1(n6897), .A2(n8461), .ZN(n7525) );
  NAND2_X1 U9183 ( .A1(n7527), .A2(n8861), .ZN(n7530) );
  AOI22_X1 U9184 ( .A1(n7575), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7574), .B2(
        n7528), .ZN(n7529) );
  NAND2_X1 U9185 ( .A1(n9733), .A2(n8689), .ZN(n8949) );
  NAND2_X1 U9186 ( .A1(n8948), .A2(n8949), .ZN(n9558) );
  NAND2_X1 U9187 ( .A1(n7531), .A2(n8689), .ZN(n7532) );
  AOI22_X1 U9188 ( .A1(n7575), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7574), .B2(
        n7534), .ZN(n7535) );
  NAND2_X1 U9189 ( .A1(n8867), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7544) );
  AND2_X1 U9190 ( .A1(n7538), .A2(n7537), .ZN(n7539) );
  NOR2_X1 U9191 ( .A1(n7540), .A2(n7539), .ZN(n9546) );
  NAND2_X1 U9192 ( .A1(n4443), .A2(n9546), .ZN(n7543) );
  NAND2_X1 U9193 ( .A1(n8868), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7542) );
  NAND2_X1 U9194 ( .A1(n4333), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7541) );
  AND2_X1 U9195 ( .A1(n9729), .A2(n8762), .ZN(n8952) );
  INV_X1 U9196 ( .A(n8952), .ZN(n9063) );
  NAND2_X1 U9197 ( .A1(n9524), .A2(n9063), .ZN(n9540) );
  INV_X1 U9198 ( .A(n8762), .ZN(n9132) );
  NAND2_X1 U9199 ( .A1(n7545), .A2(n8762), .ZN(n7546) );
  OR2_X1 U9200 ( .A1(n8757), .A2(n8690), .ZN(n9067) );
  NAND2_X1 U9201 ( .A1(n8757), .A2(n8690), .ZN(n9064) );
  NAND2_X1 U9202 ( .A1(n7547), .A2(n8861), .ZN(n7550) );
  AOI22_X1 U9203 ( .A1(n7575), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7574), .B2(
        n7548), .ZN(n7549) );
  NAND2_X1 U9204 ( .A1(n7552), .A2(n7551), .ZN(n7553) );
  AND2_X1 U9205 ( .A1(n7564), .A2(n7553), .ZN(n9514) );
  NAND2_X1 U9206 ( .A1(n4443), .A2(n9514), .ZN(n7557) );
  NAND2_X1 U9207 ( .A1(n8867), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7556) );
  NAND2_X1 U9208 ( .A1(n8868), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U9209 ( .A1(n4333), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7554) );
  INV_X1 U9210 ( .A(n8818), .ZN(n9130) );
  NOR2_X1 U9211 ( .A1(n9657), .A2(n9130), .ZN(n7558) );
  INV_X1 U9212 ( .A(n9657), .ZN(n9517) );
  NAND2_X1 U9213 ( .A1(n7559), .A2(n8861), .ZN(n7562) );
  AOI22_X1 U9214 ( .A1(n7575), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7574), .B2(
        n7560), .ZN(n7561) );
  AND2_X1 U9215 ( .A1(n7564), .A2(n7563), .ZN(n7565) );
  NOR2_X1 U9216 ( .A1(n7566), .A2(n7565), .ZN(n9493) );
  NAND2_X1 U9217 ( .A1(n9493), .A2(n4443), .ZN(n7570) );
  NAND2_X1 U9218 ( .A1(n8867), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7569) );
  NAND2_X1 U9219 ( .A1(n8868), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7568) );
  NAND2_X1 U9220 ( .A1(n4333), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7567) );
  NAND4_X1 U9221 ( .A1(n7570), .A2(n7569), .A3(n7568), .A4(n7567), .ZN(n9129)
         );
  INV_X1 U9222 ( .A(n9129), .ZN(n8708) );
  NAND2_X1 U9223 ( .A1(n9475), .A2(n9474), .ZN(n9473) );
  INV_X1 U9224 ( .A(n8508), .ZN(n9125) );
  INV_X1 U9225 ( .A(n9430), .ZN(n7584) );
  NAND2_X1 U9226 ( .A1(n7573), .A2(n8861), .ZN(n7577) );
  AOI22_X1 U9227 ( .A1(n7575), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7574), .B2(
        n9039), .ZN(n7576) );
  NAND2_X1 U9228 ( .A1(n7579), .A2(n7578), .ZN(n7580) );
  NAND2_X1 U9229 ( .A1(n7589), .A2(n7580), .ZN(n9434) );
  AOI22_X1 U9230 ( .A1(n8867), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n6062), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n7582) );
  NAND2_X1 U9231 ( .A1(n4333), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7581) );
  OAI211_X1 U9232 ( .C1(n9434), .C2(n7663), .A(n7582), .B(n7581), .ZN(n9124)
         );
  INV_X1 U9233 ( .A(n9124), .ZN(n7675) );
  NAND2_X1 U9234 ( .A1(n7585), .A2(n8861), .ZN(n7588) );
  OR2_X1 U9235 ( .A1(n8864), .A2(n7586), .ZN(n7587) );
  AND2_X1 U9236 ( .A1(n7589), .A2(n8753), .ZN(n7590) );
  NOR2_X1 U9237 ( .A1(n7601), .A2(n7590), .ZN(n9418) );
  INV_X1 U9238 ( .A(n7591), .ZN(n7648) );
  INV_X1 U9239 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7594) );
  NAND2_X1 U9240 ( .A1(n4333), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9241 ( .A1(n8868), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7592) );
  OAI211_X1 U9242 ( .C1(n7648), .C2(n7594), .A(n7593), .B(n7592), .ZN(n7595)
         );
  AOI21_X1 U9243 ( .B1(n9418), .B2(n4443), .A(n7595), .ZN(n8669) );
  NAND2_X1 U9244 ( .A1(n9421), .A2(n8669), .ZN(n7596) );
  INV_X1 U9245 ( .A(n8669), .ZN(n9123) );
  NAND2_X1 U9246 ( .A1(n7597), .A2(n8861), .ZN(n7600) );
  OR2_X1 U9247 ( .A1(n8864), .A2(n7598), .ZN(n7599) );
  OR2_X1 U9248 ( .A1(n7601), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7602) );
  AND2_X1 U9249 ( .A1(n7602), .A2(n7611), .ZN(n9405) );
  INV_X1 U9250 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U9251 ( .A1(n4333), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7604) );
  NAND2_X1 U9252 ( .A1(n8868), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7603) );
  OAI211_X1 U9253 ( .C1(n7648), .C2(n9621), .A(n7604), .B(n7603), .ZN(n7605)
         );
  AOI21_X1 U9254 ( .B1(n9405), .B2(n4443), .A(n7605), .ZN(n8771) );
  INV_X1 U9255 ( .A(n8771), .ZN(n9122) );
  NAND2_X1 U9256 ( .A1(n7606), .A2(n8861), .ZN(n7609) );
  OR2_X1 U9257 ( .A1(n8864), .A2(n7607), .ZN(n7608) );
  NAND2_X1 U9258 ( .A1(n7611), .A2(n7610), .ZN(n7612) );
  AND2_X1 U9259 ( .A1(n7622), .A2(n7612), .ZN(n9388) );
  INV_X1 U9260 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n7615) );
  INV_X1 U9261 ( .A(n4333), .ZN(n8872) );
  NAND2_X1 U9262 ( .A1(n8867), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7614) );
  NAND2_X1 U9263 ( .A1(n8868), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7613) );
  OAI211_X1 U9264 ( .C1(n7615), .C2(n8872), .A(n7614), .B(n7613), .ZN(n7616)
         );
  AOI21_X1 U9265 ( .B1(n9388), .B2(n4443), .A(n7616), .ZN(n8668) );
  NAND2_X1 U9266 ( .A1(n4872), .A2(n8668), .ZN(n7617) );
  INV_X1 U9267 ( .A(n8668), .ZN(n9121) );
  NAND2_X1 U9268 ( .A1(n7618), .A2(n8861), .ZN(n7621) );
  OR2_X1 U9269 ( .A1(n8864), .A2(n7619), .ZN(n7620) );
  AND2_X1 U9270 ( .A1(n7622), .A2(n8615), .ZN(n7623) );
  OR2_X1 U9271 ( .A1(n7623), .A2(n7644), .ZN(n8616) );
  INV_X1 U9272 ( .A(n8616), .ZN(n9373) );
  INV_X1 U9273 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U9274 ( .A1(n4333), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U9275 ( .A1(n8868), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7624) );
  OAI211_X1 U9276 ( .C1(n7648), .C2(n10090), .A(n7625), .B(n7624), .ZN(n7626)
         );
  AOI21_X1 U9277 ( .B1(n9373), .B2(n4443), .A(n7626), .ZN(n8770) );
  INV_X1 U9278 ( .A(n4334), .ZN(n9120) );
  NAND2_X1 U9279 ( .A1(n9372), .A2(n9120), .ZN(n7628) );
  NOR2_X1 U9280 ( .A1(n9372), .A2(n9120), .ZN(n7627) );
  NAND2_X1 U9281 ( .A1(n7629), .A2(n8861), .ZN(n7632) );
  OR2_X1 U9282 ( .A1(n8864), .A2(n7630), .ZN(n7631) );
  INV_X1 U9283 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n7633) );
  XNOR2_X1 U9284 ( .A(n7644), .B(n7633), .ZN(n9359) );
  INV_X1 U9285 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U9286 ( .A1(n4333), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U9287 ( .A1(n8868), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7634) );
  OAI211_X1 U9288 ( .C1(n7648), .C2(n10060), .A(n7635), .B(n7634), .ZN(n7636)
         );
  AOI21_X1 U9289 ( .B1(n9359), .B2(n4443), .A(n7636), .ZN(n8612) );
  NAND2_X1 U9290 ( .A1(n9701), .A2(n8612), .ZN(n7637) );
  NAND2_X1 U9291 ( .A1(n9348), .A2(n7637), .ZN(n7639) );
  INV_X1 U9292 ( .A(n8612), .ZN(n9119) );
  NAND2_X1 U9293 ( .A1(n9358), .A2(n9119), .ZN(n7638) );
  OR2_X1 U9294 ( .A1(n8864), .A2(n7641), .ZN(n7642) );
  AOI21_X1 U9295 ( .B1(n7644), .B2(P1_REG3_REG_24__SCAN_IN), .A(
        P1_REG3_REG_25__SCAN_IN), .ZN(n7645) );
  INV_X1 U9296 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U9297 ( .A1(n4333), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7647) );
  NAND2_X1 U9298 ( .A1(n8868), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7646) );
  OAI211_X1 U9299 ( .C1(n7648), .C2(n9603), .A(n7647), .B(n7646), .ZN(n7649)
         );
  INV_X1 U9300 ( .A(n7649), .ZN(n7650) );
  INV_X1 U9301 ( .A(n9118), .ZN(n8559) );
  NOR2_X1 U9302 ( .A1(n9697), .A2(n8559), .ZN(n7651) );
  NAND2_X1 U9303 ( .A1(n7652), .A2(n8861), .ZN(n7655) );
  OR2_X1 U9304 ( .A1(n8864), .A2(n7653), .ZN(n7654) );
  NOR2_X1 U9305 ( .A1(n7656), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7657) );
  INV_X1 U9306 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U9307 ( .A1(n8867), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U9308 ( .A1(n8868), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7659) );
  OAI211_X1 U9309 ( .C1(n9324), .C2(n8872), .A(n7660), .B(n7659), .ZN(n7661)
         );
  INV_X1 U9310 ( .A(n7661), .ZN(n7662) );
  NOR2_X1 U9311 ( .A1(n9323), .A2(n9117), .ZN(n7664) );
  NAND2_X1 U9312 ( .A1(n9593), .A2(n8803), .ZN(n8885) );
  NAND2_X1 U9313 ( .A1(n9007), .A2(n8885), .ZN(n8858) );
  NAND2_X1 U9314 ( .A1(n8867), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7669) );
  XNOR2_X1 U9315 ( .A(P1_REG3_REG_28__SCAN_IN), .B(n7665), .ZN(n9293) );
  NAND2_X1 U9316 ( .A1(n4443), .A2(n9293), .ZN(n7668) );
  NAND2_X1 U9317 ( .A1(n8868), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U9318 ( .A1(n4333), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7666) );
  NAND2_X1 U9319 ( .A1(n9269), .A2(n9280), .ZN(n9274) );
  NAND2_X1 U9320 ( .A1(n9006), .A2(n9274), .ZN(n9275) );
  XNOR2_X1 U9321 ( .A(n9271), .B(n9275), .ZN(n9291) );
  OR2_X1 U9322 ( .A1(n9358), .A2(n8612), .ZN(n8995) );
  NAND2_X1 U9323 ( .A1(n9358), .A2(n8612), .ZN(n8987) );
  OR2_X1 U9324 ( .A1(n9404), .A2(n8771), .ZN(n8982) );
  OR2_X1 U9325 ( .A1(n9625), .A2(n8669), .ZN(n9395) );
  NAND2_X1 U9326 ( .A1(n8982), .A2(n9395), .ZN(n8910) );
  INV_X1 U9327 ( .A(n8910), .ZN(n7677) );
  NOR2_X1 U9328 ( .A1(n9558), .A2(n8945), .ZN(n7670) );
  NAND2_X1 U9329 ( .A1(n9557), .A2(n7670), .ZN(n7671) );
  INV_X1 U9330 ( .A(n9540), .ZN(n9542) );
  INV_X1 U9331 ( .A(n9524), .ZN(n7672) );
  NOR2_X1 U9332 ( .A1(n9521), .A2(n7672), .ZN(n7673) );
  NAND2_X1 U9333 ( .A1(n9657), .A2(n8818), .ZN(n8960) );
  INV_X1 U9334 ( .A(n9505), .ZN(n9507) );
  INV_X1 U9335 ( .A(n9064), .ZN(n9508) );
  NAND2_X2 U9336 ( .A1(n7674), .A2(n8956), .ZN(n9509) );
  OR2_X1 U9337 ( .A1(n9649), .A2(n8708), .ZN(n9070) );
  NAND2_X1 U9338 ( .A1(n9649), .A2(n8708), .ZN(n8965) );
  NAND2_X1 U9339 ( .A1(n9070), .A2(n8965), .ZN(n9488) );
  INV_X1 U9340 ( .A(n9488), .ZN(n9498) );
  INV_X1 U9341 ( .A(n9474), .ZN(n9482) );
  NAND2_X1 U9342 ( .A1(n9480), .A2(n9076), .ZN(n9458) );
  OR2_X1 U9343 ( .A1(n9466), .A2(n8709), .ZN(n8912) );
  NAND2_X1 U9344 ( .A1(n9466), .A2(n8709), .ZN(n8975) );
  OR2_X1 U9345 ( .A1(n9634), .A2(n8508), .ZN(n9080) );
  NAND2_X1 U9346 ( .A1(n9634), .A2(n8508), .ZN(n8976) );
  NAND2_X1 U9347 ( .A1(n9447), .A2(n8976), .ZN(n9424) );
  OR2_X1 U9348 ( .A1(n9432), .A2(n7675), .ZN(n9081) );
  NAND2_X1 U9349 ( .A1(n9432), .A2(n7675), .ZN(n8970) );
  INV_X1 U9350 ( .A(n8970), .ZN(n9089) );
  NAND2_X1 U9351 ( .A1(n9625), .A2(n8669), .ZN(n8911) );
  NAND2_X1 U9352 ( .A1(n9404), .A2(n8771), .ZN(n8981) );
  INV_X1 U9353 ( .A(n8981), .ZN(n7676) );
  OR2_X1 U9354 ( .A1(n9387), .A2(n8668), .ZN(n8879) );
  NAND2_X1 U9355 ( .A1(n9387), .A2(n8668), .ZN(n8886) );
  OR2_X1 U9356 ( .A1(n9372), .A2(n4334), .ZN(n8985) );
  NAND2_X1 U9357 ( .A1(n9372), .A2(n4334), .ZN(n8992) );
  NAND2_X1 U9358 ( .A1(n9352), .A2(n8995), .ZN(n9334) );
  NAND2_X1 U9359 ( .A1(n9339), .A2(n8559), .ZN(n8997) );
  NAND2_X1 U9360 ( .A1(n8989), .A2(n8997), .ZN(n8857) );
  NAND2_X1 U9361 ( .A1(n9334), .A2(n9333), .ZN(n9332) );
  NAND2_X1 U9362 ( .A1(n9323), .A2(n8999), .ZN(n9092) );
  INV_X1 U9363 ( .A(n8885), .ZN(n7678) );
  XNOR2_X1 U9364 ( .A(n9276), .B(n9275), .ZN(n7681) );
  OR2_X1 U9365 ( .A1(n8803), .A2(n9281), .ZN(n7680) );
  OR2_X1 U9366 ( .A1(n8837), .A2(n8819), .ZN(n7679) );
  NAND2_X1 U9367 ( .A1(n7680), .A2(n7679), .ZN(n8654) );
  NAND2_X1 U9368 ( .A1(n9495), .A2(n9513), .ZN(n9490) );
  NAND2_X1 U9369 ( .A1(n9421), .A2(n9431), .ZN(n9415) );
  INV_X1 U9370 ( .A(n9570), .ZN(n9650) );
  OAI211_X1 U9371 ( .C1(n9295), .C2(n9307), .A(n9650), .B(n9283), .ZN(n9292)
         );
  NAND2_X1 U9372 ( .A1(n9300), .A2(n9292), .ZN(n7682) );
  AOI21_X1 U9373 ( .B1(n9291), .B2(n9809), .A(n7682), .ZN(n7685) );
  MUX2_X1 U9374 ( .A(n7683), .B(n7685), .S(n9816), .Z(n7684) );
  OAI21_X1 U9375 ( .B1(n9295), .B2(n9643), .A(n7684), .ZN(P1_U3550) );
  INV_X1 U9376 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7686) );
  MUX2_X1 U9377 ( .A(n7686), .B(n7685), .S(n9813), .Z(n7687) );
  OAI21_X1 U9378 ( .B1(n9295), .B2(n9722), .A(n7687), .ZN(P1_U3518) );
  INV_X1 U9379 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8863) );
  INV_X1 U9380 ( .A(n8862), .ZN(n8431) );
  OAI222_X1 U9381 ( .A1(n9750), .A2(n8863), .B1(n9747), .B2(n8431), .C1(n5865), 
        .C2(P1_U3086), .ZN(P1_U3325) );
  INV_X1 U9382 ( .A(n7688), .ZN(n8440) );
  OAI222_X1 U9383 ( .A1(n9750), .A2(n7689), .B1(P1_U3086), .B2(n9257), .C1(
        n9747), .C2(n8440), .ZN(P1_U3328) );
  NAND2_X1 U9384 ( .A1(n7691), .A2(n7690), .ZN(n7692) );
  NAND3_X1 U9385 ( .A1(n7693), .A2(n7845), .A3(n7692), .ZN(n7697) );
  AOI22_X1 U9386 ( .A1(n7869), .A2(n7796), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7694) );
  OAI21_X1 U9387 ( .B1(n8109), .B2(n7810), .A(n7694), .ZN(n7695) );
  AOI21_X1 U9388 ( .B1(n8087), .B2(n7850), .A(n7695), .ZN(n7696) );
  OAI211_X1 U9389 ( .C1(n8377), .C2(n7853), .A(n7697), .B(n7696), .ZN(P2_U3154) );
  INV_X1 U9390 ( .A(n7698), .ZN(n8416) );
  INV_X1 U9391 ( .A(n7699), .ZN(n7704) );
  NOR3_X1 U9392 ( .A1(n7700), .A2(n7702), .A3(n7701), .ZN(n7703) );
  OAI21_X1 U9393 ( .B1(n7704), .B2(n7703), .A(n7845), .ZN(n7708) );
  NAND2_X1 U9394 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7925) );
  OAI21_X1 U9395 ( .B1(n7855), .B2(n8248), .A(n7925), .ZN(n7706) );
  NOR2_X1 U9396 ( .A1(n7859), .A2(n8249), .ZN(n7705) );
  AOI211_X1 U9397 ( .C1(n7857), .C2(n7879), .A(n7706), .B(n7705), .ZN(n7707)
         );
  OAI211_X1 U9398 ( .C1(n8416), .C2(n7853), .A(n7708), .B(n7707), .ZN(P2_U3155) );
  AOI21_X1 U9399 ( .B1(n8150), .B2(n7709), .A(n4362), .ZN(n7714) );
  AOI22_X1 U9400 ( .A1(n7872), .A2(n7796), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7710) );
  OAI21_X1 U9401 ( .B1(n8161), .B2(n7810), .A(n7710), .ZN(n7712) );
  NOR2_X1 U9402 ( .A1(n8390), .A2(n7853), .ZN(n7711) );
  AOI211_X1 U9403 ( .C1(n8137), .C2(n7850), .A(n7712), .B(n7711), .ZN(n7713)
         );
  OAI21_X1 U9404 ( .B1(n7714), .B2(n7861), .A(n7713), .ZN(P2_U3156) );
  INV_X1 U9405 ( .A(n7715), .ZN(n8403) );
  INV_X1 U9406 ( .A(n7784), .ZN(n7719) );
  NOR3_X1 U9407 ( .A1(n7835), .A2(n7717), .A3(n7716), .ZN(n7718) );
  OAI21_X1 U9408 ( .B1(n7719), .B2(n7718), .A(n7845), .ZN(n7723) );
  INV_X1 U9409 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10005) );
  NOR2_X1 U9410 ( .A1(n10005), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8048) );
  AOI21_X1 U9411 ( .B1(n7796), .B2(n7874), .A(n8048), .ZN(n7720) );
  OAI21_X1 U9412 ( .B1(n8184), .B2(n7810), .A(n7720), .ZN(n7721) );
  AOI21_X1 U9413 ( .B1(n8190), .B2(n7850), .A(n7721), .ZN(n7722) );
  OAI211_X1 U9414 ( .C1(n8403), .C2(n7853), .A(n7723), .B(n7722), .ZN(P2_U3159) );
  INV_X1 U9415 ( .A(n7724), .ZN(n8395) );
  INV_X1 U9416 ( .A(n7725), .ZN(n7729) );
  NOR3_X1 U9417 ( .A1(n7786), .A2(n7727), .A3(n7726), .ZN(n7728) );
  OAI21_X1 U9418 ( .B1(n7729), .B2(n7728), .A(n7845), .ZN(n7734) );
  NOR2_X1 U9419 ( .A1(n7810), .A2(n8185), .ZN(n7732) );
  INV_X1 U9420 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7730) );
  OAI22_X1 U9421 ( .A1(n7855), .A2(n8161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7730), .ZN(n7731) );
  AOI211_X1 U9422 ( .C1(n8166), .C2(n7850), .A(n7732), .B(n7731), .ZN(n7733)
         );
  OAI211_X1 U9423 ( .C1(n8395), .C2(n7853), .A(n7734), .B(n7733), .ZN(P2_U3163) );
  NOR2_X1 U9424 ( .A1(n7222), .A2(n7882), .ZN(n7818) );
  NOR3_X1 U9425 ( .A1(n7819), .A2(n7818), .A3(n7817), .ZN(n7816) );
  AOI21_X1 U9426 ( .B1(n7881), .B2(n7817), .A(n7816), .ZN(n7735) );
  XOR2_X1 U9427 ( .A(n7736), .B(n7735), .Z(n7742) );
  NOR2_X1 U9428 ( .A1(n7810), .A2(n8275), .ZN(n7737) );
  AOI211_X1 U9429 ( .C1(n7796), .C2(n7879), .A(n7738), .B(n7737), .ZN(n7739)
         );
  OAI21_X1 U9430 ( .B1(n7859), .B2(n8280), .A(n7739), .ZN(n7740) );
  AOI21_X1 U9431 ( .B1(n9963), .B2(n7866), .A(n7740), .ZN(n7741) );
  OAI21_X1 U9432 ( .B1(n7742), .B2(n7861), .A(n7741), .ZN(P2_U3164) );
  INV_X1 U9433 ( .A(n7743), .ZN(n8382) );
  INV_X1 U9434 ( .A(n7744), .ZN(n7775) );
  INV_X1 U9435 ( .A(n7745), .ZN(n7747) );
  NOR3_X1 U9436 ( .A1(n7775), .A2(n7747), .A3(n7746), .ZN(n7749) );
  INV_X1 U9437 ( .A(n7748), .ZN(n7843) );
  OAI21_X1 U9438 ( .B1(n7749), .B2(n7843), .A(n7845), .ZN(n7753) );
  AOI22_X1 U9439 ( .A1(n7870), .A2(n7796), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7750) );
  OAI21_X1 U9440 ( .B1(n8134), .B2(n7810), .A(n7750), .ZN(n7751) );
  AOI21_X1 U9441 ( .B1(n8111), .B2(n7850), .A(n7751), .ZN(n7752) );
  OAI211_X1 U9442 ( .C1(n8382), .C2(n7853), .A(n7753), .B(n7752), .ZN(P2_U3165) );
  INV_X1 U9443 ( .A(n8411), .ZN(n8231) );
  OAI21_X1 U9444 ( .B1(n7860), .B2(n7755), .A(n7754), .ZN(n7756) );
  INV_X1 U9445 ( .A(n7756), .ZN(n7757) );
  OAI21_X1 U9446 ( .B1(n7764), .B2(n7757), .A(n7845), .ZN(n7761) );
  NAND2_X1 U9447 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7970) );
  OAI21_X1 U9448 ( .B1(n7855), .B2(n8224), .A(n7970), .ZN(n7759) );
  NOR2_X1 U9449 ( .A1(n7859), .A2(n8232), .ZN(n7758) );
  AOI211_X1 U9450 ( .C1(n7857), .C2(n7877), .A(n7759), .B(n7758), .ZN(n7760)
         );
  OAI211_X1 U9451 ( .C1(n8231), .C2(n7853), .A(n7761), .B(n7760), .ZN(P2_U3166) );
  INV_X1 U9452 ( .A(n8336), .ZN(n8220) );
  INV_X1 U9453 ( .A(n7833), .ZN(n7766) );
  NOR3_X1 U9454 ( .A1(n7764), .A2(n7763), .A3(n7762), .ZN(n7765) );
  OAI21_X1 U9455 ( .B1(n7766), .B2(n7765), .A(n7845), .ZN(n7770) );
  NAND2_X1 U9456 ( .A1(n7857), .A2(n8210), .ZN(n7767) );
  NAND2_X1 U9457 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7998) );
  OAI211_X1 U9458 ( .C1(n8184), .C2(n7855), .A(n7767), .B(n7998), .ZN(n7768)
         );
  AOI21_X1 U9459 ( .B1(n8217), .B2(n7850), .A(n7768), .ZN(n7769) );
  OAI211_X1 U9460 ( .C1(n8220), .C2(n7853), .A(n7770), .B(n7769), .ZN(P2_U3168) );
  INV_X1 U9461 ( .A(n7771), .ZN(n8386) );
  INV_X1 U9462 ( .A(n7772), .ZN(n7774) );
  NOR3_X1 U9463 ( .A1(n4362), .A2(n7774), .A3(n7773), .ZN(n7776) );
  OAI21_X1 U9464 ( .B1(n7776), .B2(n7775), .A(n7845), .ZN(n7780) );
  AOI22_X1 U9465 ( .A1(n8120), .A2(n7796), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7777) );
  OAI21_X1 U9466 ( .B1(n7808), .B2(n7810), .A(n7777), .ZN(n7778) );
  AOI21_X1 U9467 ( .B1(n8124), .B2(n7850), .A(n7778), .ZN(n7779) );
  OAI211_X1 U9468 ( .C1(n8386), .C2(n7853), .A(n7780), .B(n7779), .ZN(P2_U3169) );
  INV_X1 U9469 ( .A(n7781), .ZN(n8399) );
  AND3_X1 U9470 ( .A1(n7784), .A2(n7783), .A3(n7782), .ZN(n7785) );
  OAI21_X1 U9471 ( .B1(n7786), .B2(n7785), .A(n7845), .ZN(n7791) );
  NOR2_X1 U9472 ( .A1(n7810), .A2(n8197), .ZN(n7789) );
  OAI22_X1 U9473 ( .A1(n7855), .A2(n8174), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7787), .ZN(n7788) );
  AOI211_X1 U9474 ( .C1(n8177), .C2(n7850), .A(n7789), .B(n7788), .ZN(n7790)
         );
  OAI211_X1 U9475 ( .C1(n8399), .C2(n7853), .A(n7791), .B(n7790), .ZN(P2_U3173) );
  AOI21_X1 U9476 ( .B1(n7793), .B2(n7792), .A(n7700), .ZN(n7800) );
  INV_X1 U9477 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7794) );
  NOR2_X1 U9478 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7794), .ZN(n7904) );
  NOR2_X1 U9479 ( .A1(n7810), .A2(n8258), .ZN(n7795) );
  AOI211_X1 U9480 ( .C1(n7796), .C2(n7878), .A(n7904), .B(n7795), .ZN(n7797)
         );
  OAI21_X1 U9481 ( .B1(n8264), .B2(n7859), .A(n7797), .ZN(n7798) );
  AOI21_X1 U9482 ( .B1(n8260), .B2(n7866), .A(n7798), .ZN(n7799) );
  OAI21_X1 U9483 ( .B1(n7800), .B2(n7861), .A(n7799), .ZN(P2_U3174) );
  INV_X1 U9484 ( .A(n8316), .ZN(n7815) );
  XNOR2_X1 U9485 ( .A(n7801), .B(n8161), .ZN(n7803) );
  OAI21_X1 U9486 ( .B1(n7804), .B2(n7803), .A(n7802), .ZN(n7805) );
  OAI21_X1 U9487 ( .B1(n4677), .B2(n7806), .A(n7805), .ZN(n7807) );
  NAND2_X1 U9488 ( .A1(n7807), .A2(n7845), .ZN(n7814) );
  NOR2_X1 U9489 ( .A1(n7855), .A2(n7808), .ZN(n7812) );
  OAI22_X1 U9490 ( .A1(n7810), .A2(n8174), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7809), .ZN(n7811) );
  AOI211_X1 U9491 ( .C1(n8144), .C2(n7850), .A(n7812), .B(n7811), .ZN(n7813)
         );
  OAI211_X1 U9492 ( .C1(n7815), .C2(n7853), .A(n7814), .B(n7813), .ZN(P2_U3175) );
  INV_X1 U9493 ( .A(n7816), .ZN(n7821) );
  OAI21_X1 U9494 ( .B1(n7819), .B2(n7818), .A(n7817), .ZN(n7820) );
  NAND3_X1 U9495 ( .A1(n7821), .A2(n7845), .A3(n7820), .ZN(n7830) );
  INV_X1 U9496 ( .A(n7822), .ZN(n7828) );
  NAND2_X1 U9497 ( .A1(n7857), .A2(n7882), .ZN(n7824) );
  OAI211_X1 U9498 ( .C1(n8258), .C2(n7855), .A(n7824), .B(n7823), .ZN(n7827)
         );
  INV_X1 U9499 ( .A(n9957), .ZN(n7825) );
  NOR2_X1 U9500 ( .A1(n7825), .A2(n7853), .ZN(n7826) );
  AOI211_X1 U9501 ( .C1(n7828), .C2(n7850), .A(n7827), .B(n7826), .ZN(n7829)
         );
  NAND2_X1 U9502 ( .A1(n7830), .A2(n7829), .ZN(P2_U3176) );
  INV_X1 U9503 ( .A(n8201), .ZN(n8407) );
  AND3_X1 U9504 ( .A1(n7833), .A2(n7832), .A3(n7831), .ZN(n7834) );
  OAI21_X1 U9505 ( .B1(n7835), .B2(n7834), .A(n7845), .ZN(n7839) );
  NAND2_X1 U9506 ( .A1(n7857), .A2(n7876), .ZN(n7836) );
  NAND2_X1 U9507 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8023) );
  OAI211_X1 U9508 ( .C1(n8197), .C2(n7855), .A(n7836), .B(n8023), .ZN(n7837)
         );
  AOI21_X1 U9509 ( .B1(n8200), .B2(n7850), .A(n7837), .ZN(n7838) );
  OAI211_X1 U9510 ( .C1(n8407), .C2(n7853), .A(n7839), .B(n7838), .ZN(P2_U3178) );
  INV_X1 U9511 ( .A(n7840), .ZN(n7842) );
  NOR3_X1 U9512 ( .A1(n7843), .A2(n7842), .A3(n7841), .ZN(n7847) );
  INV_X1 U9513 ( .A(n7844), .ZN(n7846) );
  OAI21_X1 U9514 ( .B1(n7847), .B2(n7846), .A(n7845), .ZN(n7852) );
  AOI22_X1 U9515 ( .A1(n8120), .A2(n7857), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n7848) );
  OAI21_X1 U9516 ( .B1(n8072), .B2(n7855), .A(n7848), .ZN(n7849) );
  AOI21_X1 U9517 ( .B1(n8099), .B2(n7850), .A(n7849), .ZN(n7851) );
  OAI211_X1 U9518 ( .C1(n7854), .C2(n7853), .A(n7852), .B(n7851), .ZN(P2_U3180) );
  NAND2_X1 U9519 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7951) );
  OAI21_X1 U9520 ( .B1(n7855), .B2(n8240), .A(n7951), .ZN(n7856) );
  AOI21_X1 U9521 ( .B1(n7857), .B2(n7878), .A(n7856), .ZN(n7858) );
  OAI21_X1 U9522 ( .B1(n8241), .B2(n7859), .A(n7858), .ZN(n7865) );
  AOI211_X1 U9523 ( .C1(n7863), .C2(n7862), .A(n7861), .B(n7860), .ZN(n7864)
         );
  AOI211_X1 U9524 ( .C1(n8346), .C2(n7866), .A(n7865), .B(n7864), .ZN(n7867)
         );
  INV_X1 U9525 ( .A(n7867), .ZN(P2_U3181) );
  MUX2_X1 U9526 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8057), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9527 ( .A(n7868), .B(P2_DATAO_REG_30__SCAN_IN), .S(n7871), .Z(
        P2_U3521) );
  MUX2_X1 U9528 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n7869), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9529 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8095), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9530 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n7870), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9531 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8120), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9532 ( .A(n7872), .B(P2_DATAO_REG_24__SCAN_IN), .S(n7871), .Z(
        P2_U3515) );
  MUX2_X1 U9533 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8150), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9534 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n7873), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9535 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8149), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9536 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n7874), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9537 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n7875), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9538 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8212), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9539 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n7876), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9540 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8210), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9541 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n7877), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9542 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n7878), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9543 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n7879), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9544 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n7880), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9545 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n7881), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9546 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n7882), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9547 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n7883), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9548 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n7884), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9549 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n7885), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9550 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n7886), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9551 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n7887), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U9552 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n7888), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9553 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n7889), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9554 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n7890), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U9555 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n7891), .S(P2_U3893), .Z(
        P2_U3492) );
  AOI21_X1 U9556 ( .B1(n8355), .B2(n7893), .A(n7928), .ZN(n7910) );
  AOI21_X1 U9557 ( .B1(n7896), .B2(n7895), .A(n7894), .ZN(n7898) );
  MUX2_X1 U9558 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8041), .Z(n7918) );
  XNOR2_X1 U9559 ( .A(n7918), .B(n7927), .ZN(n7897) );
  NAND2_X1 U9560 ( .A1(n7898), .A2(n7897), .ZN(n7919) );
  OAI21_X1 U9561 ( .B1(n7898), .B2(n7897), .A(n7919), .ZN(n7908) );
  AOI21_X1 U9562 ( .B1(n7901), .B2(n8265), .A(n7912), .ZN(n7902) );
  NOR2_X1 U9563 ( .A1(n9891), .A2(n7902), .ZN(n7903) );
  AOI211_X1 U9564 ( .C1(n7927), .C2(n9826), .A(n7904), .B(n7903), .ZN(n7905)
         );
  OAI21_X1 U9565 ( .B1(n7906), .B2(n9882), .A(n7905), .ZN(n7907) );
  AOI21_X1 U9566 ( .B1(n7908), .B2(n9867), .A(n7907), .ZN(n7909) );
  OAI21_X1 U9567 ( .B1(n7910), .B2(n8000), .A(n7909), .ZN(P2_U3195) );
  NOR2_X1 U9568 ( .A1(n7927), .A2(n7911), .ZN(n7913) );
  MUX2_X1 U9569 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n7914), .S(n7930), .Z(n7915)
         );
  AOI21_X1 U9570 ( .B1(n7916), .B2(n7915), .A(n7940), .ZN(n7937) );
  MUX2_X1 U9571 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8041), .Z(n7944) );
  XNOR2_X1 U9572 ( .A(n7944), .B(n7930), .ZN(n7922) );
  OR2_X1 U9573 ( .A1(n7918), .A2(n7917), .ZN(n7920) );
  NAND2_X1 U9574 ( .A1(n7920), .A2(n7919), .ZN(n7921) );
  NAND2_X1 U9575 ( .A1(n7922), .A2(n7921), .ZN(n7945) );
  OAI21_X1 U9576 ( .B1(n7922), .B2(n7921), .A(n7945), .ZN(n7923) );
  NAND2_X1 U9577 ( .A1(n9867), .A2(n7923), .ZN(n7924) );
  OAI211_X1 U9578 ( .C1(n9906), .C2(n7943), .A(n7925), .B(n7924), .ZN(n7935)
         );
  NOR2_X1 U9579 ( .A1(n7927), .A2(n7926), .ZN(n7929) );
  AOI22_X1 U9580 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7930), .B1(n7943), .B2(
        n8351), .ZN(n7931) );
  NOR2_X1 U9581 ( .A1(n7932), .A2(n7931), .ZN(n7938) );
  AOI21_X1 U9582 ( .B1(n7932), .B2(n7931), .A(n7938), .ZN(n7933) );
  NOR2_X1 U9583 ( .A1(n7933), .A2(n8000), .ZN(n7934) );
  AOI211_X1 U9584 ( .C1(n9897), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n7935), .B(
        n7934), .ZN(n7936) );
  OAI21_X1 U9585 ( .B1(n7937), .B2(n9891), .A(n7936), .ZN(P2_U3196) );
  AOI21_X1 U9586 ( .B1(n10065), .B2(n7939), .A(n7973), .ZN(n7955) );
  XNOR2_X1 U9587 ( .A(n7972), .B(n7956), .ZN(n7941) );
  AOI21_X1 U9588 ( .B1(n7941), .B2(n8242), .A(n7957), .ZN(n7942) );
  NOR2_X1 U9589 ( .A1(n9891), .A2(n7942), .ZN(n7953) );
  MUX2_X1 U9590 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8041), .Z(n7963) );
  XNOR2_X1 U9591 ( .A(n7972), .B(n7963), .ZN(n7948) );
  OR2_X1 U9592 ( .A1(n7944), .A2(n7943), .ZN(n7946) );
  NAND2_X1 U9593 ( .A1(n7946), .A2(n7945), .ZN(n7947) );
  NAND2_X1 U9594 ( .A1(n7948), .A2(n7947), .ZN(n7964) );
  OAI21_X1 U9595 ( .B1(n7948), .B2(n7947), .A(n7964), .ZN(n7949) );
  NAND2_X1 U9596 ( .A1(n9867), .A2(n7949), .ZN(n7950) );
  OAI211_X1 U9597 ( .C1(n9906), .C2(n7962), .A(n7951), .B(n7950), .ZN(n7952)
         );
  AOI211_X1 U9598 ( .C1(n9897), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n7953), .B(
        n7952), .ZN(n7954) );
  OAI21_X1 U9599 ( .B1(n7955), .B2(n8000), .A(n7954), .ZN(P2_U3197) );
  INV_X1 U9600 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7959) );
  NOR2_X1 U9601 ( .A1(n7990), .A2(n7959), .ZN(n7958) );
  AOI21_X1 U9602 ( .B1(n7959), .B2(n7990), .A(n7958), .ZN(n7960) );
  AOI21_X1 U9603 ( .B1(n7961), .B2(n7960), .A(n7987), .ZN(n7983) );
  MUX2_X1 U9604 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8041), .Z(n7991) );
  XNOR2_X1 U9605 ( .A(n7991), .B(n7976), .ZN(n7967) );
  OR2_X1 U9606 ( .A1(n7963), .A2(n7962), .ZN(n7965) );
  NAND2_X1 U9607 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  NAND2_X1 U9608 ( .A1(n7967), .A2(n7966), .ZN(n7992) );
  OAI21_X1 U9609 ( .B1(n7967), .B2(n7966), .A(n7992), .ZN(n7968) );
  NAND2_X1 U9610 ( .A1(n9867), .A2(n7968), .ZN(n7969) );
  OAI211_X1 U9611 ( .C1(n9906), .C2(n7990), .A(n7970), .B(n7969), .ZN(n7981)
         );
  NOR2_X1 U9612 ( .A1(n7972), .A2(n7971), .ZN(n7974) );
  AOI22_X1 U9613 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n7976), .B1(n7990), .B2(
        n7975), .ZN(n7977) );
  AOI21_X1 U9614 ( .B1(n7978), .B2(n7977), .A(n7984), .ZN(n7979) );
  NOR2_X1 U9615 ( .A1(n7979), .A2(n8000), .ZN(n7980) );
  AOI211_X1 U9616 ( .C1(n9897), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n7981), .B(
        n7980), .ZN(n7982) );
  OAI21_X1 U9617 ( .B1(n7983), .B2(n9891), .A(n7982), .ZN(P2_U3198) );
  XNOR2_X1 U9618 ( .A(n8008), .B(n8007), .ZN(n7985) );
  AOI21_X1 U9619 ( .B1(n7986), .B2(n7985), .A(n8009), .ZN(n8001) );
  NOR2_X1 U9620 ( .A1(n7988), .A2(n7989), .ZN(n8003) );
  MUX2_X1 U9621 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8041), .Z(n8015) );
  XNOR2_X1 U9622 ( .A(n8015), .B(n8008), .ZN(n7995) );
  OR2_X1 U9623 ( .A1(n7991), .A2(n7990), .ZN(n7993) );
  NAND2_X1 U9624 ( .A1(n7993), .A2(n7992), .ZN(n7994) );
  NAND2_X1 U9625 ( .A1(n7995), .A2(n7994), .ZN(n8013) );
  OAI21_X1 U9626 ( .B1(n7995), .B2(n7994), .A(n8013), .ZN(n7996) );
  NAND2_X1 U9627 ( .A1(n9867), .A2(n7996), .ZN(n7997) );
  OAI211_X1 U9628 ( .C1(n9906), .C2(n8014), .A(n7998), .B(n7997), .ZN(n7999)
         );
  NOR2_X1 U9629 ( .A1(n8008), .A2(n8002), .ZN(n8004) );
  NAND2_X1 U9630 ( .A1(n8039), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8030) );
  OAI21_X1 U9631 ( .B1(n8039), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8030), .ZN(
        n8005) );
  AOI21_X1 U9632 ( .B1(n8006), .B2(n8005), .A(n8032), .ZN(n8029) );
  NOR2_X1 U9633 ( .A1(n8008), .A2(n8007), .ZN(n8010) );
  NAND2_X1 U9634 ( .A1(n8039), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8034) );
  OAI21_X1 U9635 ( .B1(n8039), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8034), .ZN(
        n8011) );
  INV_X1 U9636 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8012) );
  NOR2_X1 U9637 ( .A1(n9882), .A2(n8012), .ZN(n8026) );
  OAI21_X1 U9638 ( .B1(n8015), .B2(n8014), .A(n8013), .ZN(n8018) );
  MUX2_X1 U9639 ( .A(n8016), .B(n8334), .S(n8041), .Z(n8017) );
  NOR2_X1 U9640 ( .A1(n8018), .A2(n8017), .ZN(n8037) );
  NAND2_X1 U9641 ( .A1(n8018), .A2(n8017), .ZN(n8038) );
  INV_X1 U9642 ( .A(n8038), .ZN(n8019) );
  NOR2_X1 U9643 ( .A1(n8037), .A2(n8019), .ZN(n8020) );
  AOI21_X1 U9644 ( .B1(P2_U3893), .B2(n8020), .A(n9826), .ZN(n8024) );
  INV_X1 U9645 ( .A(n8020), .ZN(n8021) );
  NAND3_X1 U9646 ( .A1(n9867), .A2(n8039), .A3(n8021), .ZN(n8022) );
  OAI211_X1 U9647 ( .C1(n8024), .C2(n8039), .A(n8023), .B(n8022), .ZN(n8025)
         );
  OAI21_X1 U9648 ( .B1(n8029), .B2(n9891), .A(n8028), .ZN(P2_U3200) );
  INV_X1 U9649 ( .A(n8030), .ZN(n8031) );
  XNOR2_X1 U9650 ( .A(n8046), .B(n8033), .ZN(n8043) );
  INV_X1 U9651 ( .A(n8034), .ZN(n8035) );
  XNOR2_X1 U9652 ( .A(n8046), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8040) );
  XNOR2_X1 U9653 ( .A(n8036), .B(n8040), .ZN(n8052) );
  AOI21_X1 U9654 ( .B1(n8039), .B2(n8038), .A(n8037), .ZN(n8045) );
  INV_X1 U9655 ( .A(n8040), .ZN(n8042) );
  MUX2_X1 U9656 ( .A(n8043), .B(n8042), .S(n8041), .Z(n8044) );
  XNOR2_X1 U9657 ( .A(n8045), .B(n8044), .ZN(n8049) );
  NOR2_X1 U9658 ( .A1(n9906), .A2(n8046), .ZN(n8047) );
  AOI211_X1 U9659 ( .C1(n8049), .C2(n9867), .A(n8048), .B(n8047), .ZN(n8050)
         );
  OAI21_X1 U9660 ( .B1(n4739), .B2(n9882), .A(n8050), .ZN(n8051) );
  AOI21_X1 U9661 ( .B1(n8052), .B2(n9901), .A(n8051), .ZN(n8053) );
  INV_X1 U9662 ( .A(n8054), .ZN(n8055) );
  NAND2_X1 U9663 ( .A1(n8055), .A2(n8218), .ZN(n8062) );
  NAND2_X1 U9664 ( .A1(n8057), .A2(n8056), .ZN(n8365) );
  AOI21_X1 U9665 ( .B1(n8062), .B2(n8365), .A(n8269), .ZN(n8059) );
  AOI21_X1 U9666 ( .B1(n8269), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8059), .ZN(
        n8058) );
  OAI21_X1 U9667 ( .B1(n8367), .B2(n8230), .A(n8058), .ZN(P2_U3202) );
  AOI21_X1 U9668 ( .B1(n8269), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8059), .ZN(
        n8060) );
  OAI21_X1 U9669 ( .B1(n8370), .B2(n8230), .A(n8060), .ZN(P2_U3203) );
  NAND2_X1 U9670 ( .A1(n8061), .A2(n8282), .ZN(n8067) );
  OAI21_X1 U9671 ( .B1(n8282), .B2(n8063), .A(n8062), .ZN(n8064) );
  AOI21_X1 U9672 ( .B1(n8065), .B2(n8284), .A(n8064), .ZN(n8066) );
  OAI211_X1 U9673 ( .C1(n8069), .C2(n8068), .A(n8067), .B(n8066), .ZN(P2_U3204) );
  XNOR2_X1 U9674 ( .A(n8070), .B(n8074), .ZN(n8071) );
  INV_X1 U9675 ( .A(n8291), .ZN(n8080) );
  XOR2_X1 U9676 ( .A(n8075), .B(n8074), .Z(n8292) );
  AOI22_X1 U9677 ( .A1(n8076), .A2(n8218), .B1(n8269), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8077) );
  OAI21_X1 U9678 ( .B1(n8373), .B2(n8230), .A(n8077), .ZN(n8078) );
  AOI21_X1 U9679 ( .B1(n8292), .B2(n8267), .A(n8078), .ZN(n8079) );
  OAI21_X1 U9680 ( .B1(n8080), .B2(n8269), .A(n8079), .ZN(P2_U3205) );
  XNOR2_X1 U9681 ( .A(n8082), .B(n8088), .ZN(n8085) );
  OAI22_X1 U9682 ( .A1(n8083), .A2(n8278), .B1(n8109), .B2(n8276), .ZN(n8084)
         );
  INV_X1 U9683 ( .A(n8297), .ZN(n8086) );
  AOI21_X1 U9684 ( .B1(n8218), .B2(n8087), .A(n8086), .ZN(n8093) );
  XNOR2_X1 U9685 ( .A(n8089), .B(n8088), .ZN(n8295) );
  OAI22_X1 U9686 ( .A1(n8377), .A2(n8230), .B1(n8090), .B2(n8282), .ZN(n8091)
         );
  AOI21_X1 U9687 ( .B1(n8295), .B2(n8267), .A(n8091), .ZN(n8092) );
  OAI21_X1 U9688 ( .B1(n8093), .B2(n8269), .A(n8092), .ZN(P2_U3206) );
  XNOR2_X1 U9689 ( .A(n8094), .B(n8097), .ZN(n8096) );
  AOI222_X1 U9690 ( .A1(n8214), .A2(n8096), .B1(n8095), .B2(n8211), .C1(n8120), 
        .C2(n8209), .ZN(n8303) );
  XNOR2_X1 U9691 ( .A(n8098), .B(n8097), .ZN(n8301) );
  NAND2_X1 U9692 ( .A1(n8300), .A2(n8284), .ZN(n8101) );
  AOI22_X1 U9693 ( .A1(n8269), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8099), .B2(
        n8218), .ZN(n8100) );
  NAND2_X1 U9694 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  AOI21_X1 U9695 ( .B1(n8301), .B2(n8267), .A(n8102), .ZN(n8103) );
  OAI21_X1 U9696 ( .B1(n8303), .B2(n8269), .A(n8103), .ZN(P2_U3207) );
  NOR2_X1 U9697 ( .A1(n8382), .A2(n8255), .ZN(n8110) );
  INV_X1 U9698 ( .A(n8104), .ZN(n8105) );
  AOI21_X1 U9699 ( .B1(n8107), .B2(n8106), .A(n8105), .ZN(n8108) );
  OAI222_X1 U9700 ( .A1(n8278), .A2(n8109), .B1(n8276), .B2(n8134), .C1(n8358), 
        .C2(n8108), .ZN(n8304) );
  AOI211_X1 U9701 ( .C1(n8218), .C2(n8111), .A(n8110), .B(n8304), .ZN(n8115)
         );
  XNOR2_X1 U9702 ( .A(n8113), .B(n8112), .ZN(n8305) );
  AOI22_X1 U9703 ( .A1(n8305), .A2(n8267), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8269), .ZN(n8114) );
  OAI21_X1 U9704 ( .B1(n8115), .B2(n8269), .A(n8114), .ZN(P2_U3208) );
  NOR2_X1 U9705 ( .A1(n8386), .A2(n8255), .ZN(n8123) );
  INV_X1 U9706 ( .A(n8116), .ZN(n8119) );
  INV_X1 U9707 ( .A(n8127), .ZN(n8118) );
  OAI211_X1 U9708 ( .C1(n8119), .C2(n8118), .A(n8214), .B(n8117), .ZN(n8122)
         );
  AOI22_X1 U9709 ( .A1(n8120), .A2(n8211), .B1(n8209), .B2(n8150), .ZN(n8121)
         );
  NAND2_X1 U9710 ( .A1(n8122), .A2(n8121), .ZN(n8308) );
  AOI211_X1 U9711 ( .C1(n8218), .C2(n8124), .A(n8123), .B(n8308), .ZN(n8130)
         );
  NAND2_X1 U9712 ( .A1(n8126), .A2(n8125), .ZN(n8128) );
  XNOR2_X1 U9713 ( .A(n8128), .B(n8127), .ZN(n8309) );
  AOI22_X1 U9714 ( .A1(n8309), .A2(n8267), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8269), .ZN(n8129) );
  OAI21_X1 U9715 ( .B1(n8130), .B2(n8269), .A(n8129), .ZN(P2_U3209) );
  XNOR2_X1 U9716 ( .A(n8132), .B(n8131), .ZN(n8133) );
  OAI222_X1 U9717 ( .A1(n8278), .A2(n8134), .B1(n8276), .B2(n8161), .C1(n8358), 
        .C2(n8133), .ZN(n8312) );
  INV_X1 U9718 ( .A(n8312), .ZN(n8141) );
  XNOR2_X1 U9719 ( .A(n8136), .B(n8135), .ZN(n8313) );
  AOI22_X1 U9720 ( .A1(n8269), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8218), .B2(
        n8137), .ZN(n8138) );
  OAI21_X1 U9721 ( .B1(n8390), .B2(n8230), .A(n8138), .ZN(n8139) );
  AOI21_X1 U9722 ( .B1(n8313), .B2(n8267), .A(n8139), .ZN(n8140) );
  OAI21_X1 U9723 ( .B1(n8141), .B2(n8269), .A(n8140), .ZN(P2_U3210) );
  OAI21_X1 U9724 ( .B1(n8143), .B2(n8146), .A(n8142), .ZN(n8319) );
  INV_X1 U9725 ( .A(n8144), .ZN(n8152) );
  NAND3_X1 U9726 ( .A1(n8159), .A2(n8146), .A3(n8145), .ZN(n8147) );
  NAND2_X1 U9727 ( .A1(n8148), .A2(n8147), .ZN(n8151) );
  AOI222_X1 U9728 ( .A1(n8214), .A2(n8151), .B1(n8150), .B2(n8211), .C1(n8149), 
        .C2(n8209), .ZN(n8318) );
  OAI21_X1 U9729 ( .B1(n8152), .B2(n8279), .A(n8318), .ZN(n8153) );
  NAND2_X1 U9730 ( .A1(n8153), .A2(n8282), .ZN(n8155) );
  AOI22_X1 U9731 ( .A1(n8316), .A2(n8284), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n8269), .ZN(n8154) );
  OAI211_X1 U9732 ( .C1(n8319), .C2(n8287), .A(n8155), .B(n8154), .ZN(P2_U3211) );
  INV_X1 U9733 ( .A(n8165), .ZN(n8157) );
  NAND3_X1 U9734 ( .A1(n8171), .A2(n8157), .A3(n8156), .ZN(n8158) );
  AND2_X1 U9735 ( .A1(n8159), .A2(n8158), .ZN(n8160) );
  OAI222_X1 U9736 ( .A1(n8278), .A2(n8161), .B1(n8276), .B2(n8185), .C1(n8358), 
        .C2(n8160), .ZN(n8320) );
  INV_X1 U9737 ( .A(n8320), .ZN(n8170) );
  NAND2_X1 U9738 ( .A1(n8163), .A2(n8162), .ZN(n8164) );
  XOR2_X1 U9739 ( .A(n8165), .B(n8164), .Z(n8321) );
  AOI22_X1 U9740 ( .A1(n8269), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8218), .B2(
        n8166), .ZN(n8167) );
  OAI21_X1 U9741 ( .B1(n8395), .B2(n8230), .A(n8167), .ZN(n8168) );
  AOI21_X1 U9742 ( .B1(n8321), .B2(n8267), .A(n8168), .ZN(n8169) );
  OAI21_X1 U9743 ( .B1(n8170), .B2(n8269), .A(n8169), .ZN(P2_U3212) );
  INV_X1 U9744 ( .A(n8171), .ZN(n8172) );
  AOI21_X1 U9745 ( .B1(n8175), .B2(n5571), .A(n8172), .ZN(n8173) );
  OAI222_X1 U9746 ( .A1(n8278), .A2(n8174), .B1(n8276), .B2(n8197), .C1(n8358), 
        .C2(n8173), .ZN(n8324) );
  INV_X1 U9747 ( .A(n8324), .ZN(n8181) );
  XNOR2_X1 U9748 ( .A(n8176), .B(n8175), .ZN(n8325) );
  AOI22_X1 U9749 ( .A1(n8269), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8218), .B2(
        n8177), .ZN(n8178) );
  OAI21_X1 U9750 ( .B1(n8399), .B2(n8230), .A(n8178), .ZN(n8179) );
  AOI21_X1 U9751 ( .B1(n8325), .B2(n8267), .A(n8179), .ZN(n8180) );
  OAI21_X1 U9752 ( .B1(n8181), .B2(n8269), .A(n8180), .ZN(P2_U3213) );
  XNOR2_X1 U9753 ( .A(n8182), .B(n8189), .ZN(n8183) );
  OAI222_X1 U9754 ( .A1(n8278), .A2(n8185), .B1(n8276), .B2(n8184), .C1(n8358), 
        .C2(n8183), .ZN(n8327) );
  INV_X1 U9755 ( .A(n8327), .ZN(n8194) );
  NAND2_X1 U9756 ( .A1(n8186), .A2(n8187), .ZN(n8188) );
  XOR2_X1 U9757 ( .A(n8189), .B(n8188), .Z(n8328) );
  AOI22_X1 U9758 ( .A1(n8269), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8218), .B2(
        n8190), .ZN(n8191) );
  OAI21_X1 U9759 ( .B1(n8403), .B2(n8230), .A(n8191), .ZN(n8192) );
  AOI21_X1 U9760 ( .B1(n8328), .B2(n8267), .A(n8192), .ZN(n8193) );
  OAI21_X1 U9761 ( .B1(n8194), .B2(n8269), .A(n8193), .ZN(P2_U3214) );
  XOR2_X1 U9762 ( .A(n8195), .B(n8198), .Z(n8196) );
  OAI222_X1 U9763 ( .A1(n8278), .A2(n8197), .B1(n8276), .B2(n8224), .C1(n8196), 
        .C2(n8358), .ZN(n8332) );
  OAI21_X1 U9764 ( .B1(n8199), .B2(n8198), .A(n8186), .ZN(n8331) );
  AOI22_X1 U9765 ( .A1(n8269), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8218), .B2(
        n8200), .ZN(n8203) );
  NAND2_X1 U9766 ( .A1(n8201), .A2(n8284), .ZN(n8202) );
  OAI211_X1 U9767 ( .C1(n8331), .C2(n8287), .A(n8203), .B(n8202), .ZN(n8204)
         );
  AOI21_X1 U9768 ( .B1(n8332), .B2(n8282), .A(n8204), .ZN(n8205) );
  INV_X1 U9769 ( .A(n8205), .ZN(P2_U3215) );
  NAND2_X1 U9770 ( .A1(n8226), .A2(n8207), .ZN(n8208) );
  XOR2_X1 U9771 ( .A(n8208), .B(n8215), .Z(n8213) );
  AOI222_X1 U9772 ( .A1(n8214), .A2(n8213), .B1(n8212), .B2(n8211), .C1(n8210), 
        .C2(n8209), .ZN(n8339) );
  XNOR2_X1 U9773 ( .A(n8216), .B(n8215), .ZN(n8337) );
  AOI22_X1 U9774 ( .A1(n8269), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8218), .B2(
        n8217), .ZN(n8219) );
  OAI21_X1 U9775 ( .B1(n8220), .B2(n8230), .A(n8219), .ZN(n8221) );
  AOI21_X1 U9776 ( .B1(n8337), .B2(n8267), .A(n8221), .ZN(n8222) );
  OAI21_X1 U9777 ( .B1(n8339), .B2(n8269), .A(n8222), .ZN(P2_U3216) );
  AOI21_X1 U9778 ( .B1(n8206), .B2(n8223), .A(n8358), .ZN(n8227) );
  OAI22_X1 U9779 ( .A1(n8248), .A2(n8276), .B1(n8224), .B2(n8278), .ZN(n8225)
         );
  AOI21_X1 U9780 ( .B1(n8227), .B2(n8226), .A(n8225), .ZN(n8342) );
  XNOR2_X1 U9781 ( .A(n8229), .B(n8228), .ZN(n8340) );
  NOR2_X1 U9782 ( .A1(n8231), .A2(n8230), .ZN(n8234) );
  OAI22_X1 U9783 ( .A1(n8282), .A2(n7959), .B1(n8232), .B2(n8279), .ZN(n8233)
         );
  AOI211_X1 U9784 ( .C1(n8340), .C2(n8267), .A(n8234), .B(n8233), .ZN(n8235)
         );
  OAI21_X1 U9785 ( .B1(n8342), .B2(n8269), .A(n8235), .ZN(P2_U3217) );
  XOR2_X1 U9786 ( .A(n8236), .B(n8238), .Z(n8348) );
  AOI21_X1 U9787 ( .B1(n8238), .B2(n8237), .A(n4422), .ZN(n8239) );
  OAI222_X1 U9788 ( .A1(n8278), .A2(n8240), .B1(n8276), .B2(n8259), .C1(n8358), 
        .C2(n8239), .ZN(n8345) );
  NAND2_X1 U9789 ( .A1(n8345), .A2(n8282), .ZN(n8245) );
  OAI22_X1 U9790 ( .A1(n8282), .A2(n8242), .B1(n8241), .B2(n8279), .ZN(n8243)
         );
  AOI21_X1 U9791 ( .B1(n8346), .B2(n8284), .A(n8243), .ZN(n8244) );
  OAI211_X1 U9792 ( .C1(n8348), .C2(n8287), .A(n8245), .B(n8244), .ZN(P2_U3218) );
  XOR2_X1 U9793 ( .A(n8251), .B(n8246), .Z(n8247) );
  OAI222_X1 U9794 ( .A1(n8278), .A2(n8248), .B1(n8276), .B2(n8277), .C1(n8247), 
        .C2(n8358), .ZN(n8349) );
  OAI22_X1 U9795 ( .A1(n8416), .A2(n8255), .B1(n8249), .B2(n8279), .ZN(n8250)
         );
  OAI21_X1 U9796 ( .B1(n8349), .B2(n8250), .A(n8282), .ZN(n8254) );
  XNOR2_X1 U9797 ( .A(n8252), .B(n8251), .ZN(n8350) );
  AOI22_X1 U9798 ( .A1(n8350), .A2(n8267), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8269), .ZN(n8253) );
  NAND2_X1 U9799 ( .A1(n8254), .A2(n8253), .ZN(P2_U3219) );
  INV_X1 U9800 ( .A(n8255), .ZN(n8261) );
  XNOR2_X1 U9801 ( .A(n8256), .B(n8263), .ZN(n8257) );
  OAI222_X1 U9802 ( .A1(n8278), .A2(n8259), .B1(n8276), .B2(n8258), .C1(n8257), 
        .C2(n8358), .ZN(n8353) );
  AOI21_X1 U9803 ( .B1(n8261), .B2(n8260), .A(n8353), .ZN(n8270) );
  XOR2_X1 U9804 ( .A(n8263), .B(n8262), .Z(n8354) );
  OAI22_X1 U9805 ( .A1(n8282), .A2(n8265), .B1(n8264), .B2(n8279), .ZN(n8266)
         );
  AOI21_X1 U9806 ( .B1(n8354), .B2(n8267), .A(n8266), .ZN(n8268) );
  OAI21_X1 U9807 ( .B1(n8270), .B2(n8269), .A(n8268), .ZN(P2_U3220) );
  OAI21_X1 U9808 ( .B1(n4421), .B2(n4792), .A(n8271), .ZN(n9960) );
  XNOR2_X1 U9809 ( .A(n8273), .B(n8272), .ZN(n8274) );
  OAI222_X1 U9810 ( .A1(n8278), .A2(n8277), .B1(n8276), .B2(n8275), .C1(n8274), 
        .C2(n8358), .ZN(n9961) );
  NAND2_X1 U9811 ( .A1(n9961), .A2(n8282), .ZN(n8286) );
  OAI22_X1 U9812 ( .A1(n8282), .A2(n8281), .B1(n8280), .B2(n8279), .ZN(n8283)
         );
  AOI21_X1 U9813 ( .B1(n9963), .B2(n8284), .A(n8283), .ZN(n8285) );
  OAI211_X1 U9814 ( .C1(n8287), .C2(n9960), .A(n8286), .B(n8285), .ZN(P2_U3221) );
  NOR2_X1 U9815 ( .A1(n8365), .A2(n10190), .ZN(n8289) );
  AOI21_X1 U9816 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10190), .A(n8289), .ZN(
        n8288) );
  OAI21_X1 U9817 ( .B1(n8367), .B2(n8357), .A(n8288), .ZN(P2_U3490) );
  AOI21_X1 U9818 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10190), .A(n8289), .ZN(
        n8290) );
  OAI21_X1 U9819 ( .B1(n8370), .B2(n8357), .A(n8290), .ZN(P2_U3489) );
  INV_X1 U9820 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8293) );
  MUX2_X1 U9821 ( .A(n8293), .B(n8371), .S(n10192), .Z(n8294) );
  OAI21_X1 U9822 ( .B1(n8373), .B2(n8357), .A(n8294), .ZN(P2_U3487) );
  INV_X1 U9823 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U9824 ( .A1(n8295), .A2(n9933), .ZN(n8296) );
  MUX2_X1 U9825 ( .A(n8298), .B(n8374), .S(n10192), .Z(n8299) );
  OAI21_X1 U9826 ( .B1(n8377), .B2(n8357), .A(n8299), .ZN(P2_U3486) );
  AOI22_X1 U9827 ( .A1(n8301), .A2(n9933), .B1(n9964), .B2(n8300), .ZN(n8302)
         );
  NAND2_X1 U9828 ( .A1(n8303), .A2(n8302), .ZN(n8378) );
  MUX2_X1 U9829 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8378), .S(n10192), .Z(
        P2_U3485) );
  INV_X1 U9830 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8306) );
  AOI21_X1 U9831 ( .B1(n9933), .B2(n8305), .A(n8304), .ZN(n8379) );
  MUX2_X1 U9832 ( .A(n8306), .B(n8379), .S(n10192), .Z(n8307) );
  OAI21_X1 U9833 ( .B1(n8382), .B2(n8357), .A(n8307), .ZN(P2_U3484) );
  INV_X1 U9834 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8310) );
  AOI21_X1 U9835 ( .B1(n8309), .B2(n9933), .A(n8308), .ZN(n8383) );
  MUX2_X1 U9836 ( .A(n8310), .B(n8383), .S(n10192), .Z(n8311) );
  OAI21_X1 U9837 ( .B1(n8386), .B2(n8357), .A(n8311), .ZN(P2_U3483) );
  INV_X1 U9838 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8314) );
  AOI21_X1 U9839 ( .B1(n9933), .B2(n8313), .A(n8312), .ZN(n8387) );
  MUX2_X1 U9840 ( .A(n8314), .B(n8387), .S(n10192), .Z(n8315) );
  OAI21_X1 U9841 ( .B1(n8390), .B2(n8357), .A(n8315), .ZN(P2_U3482) );
  NAND2_X1 U9842 ( .A1(n8316), .A2(n9964), .ZN(n8317) );
  OAI211_X1 U9843 ( .C1(n9959), .C2(n8319), .A(n8318), .B(n8317), .ZN(n8391)
         );
  MUX2_X1 U9844 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8391), .S(n10192), .Z(
        P2_U3481) );
  INV_X1 U9845 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8322) );
  AOI21_X1 U9846 ( .B1(n8321), .B2(n9933), .A(n8320), .ZN(n8392) );
  MUX2_X1 U9847 ( .A(n8322), .B(n8392), .S(n10192), .Z(n8323) );
  OAI21_X1 U9848 ( .B1(n8395), .B2(n8357), .A(n8323), .ZN(P2_U3480) );
  INV_X1 U9849 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10171) );
  AOI21_X1 U9850 ( .B1(n8325), .B2(n9933), .A(n8324), .ZN(n8396) );
  MUX2_X1 U9851 ( .A(n10171), .B(n8396), .S(n10192), .Z(n8326) );
  OAI21_X1 U9852 ( .B1(n8399), .B2(n8357), .A(n8326), .ZN(P2_U3479) );
  AOI21_X1 U9853 ( .B1(n9933), .B2(n8328), .A(n8327), .ZN(n8400) );
  MUX2_X1 U9854 ( .A(n8329), .B(n8400), .S(n10192), .Z(n8330) );
  OAI21_X1 U9855 ( .B1(n8403), .B2(n8357), .A(n8330), .ZN(P2_U3478) );
  INV_X1 U9856 ( .A(n8331), .ZN(n8333) );
  AOI21_X1 U9857 ( .B1(n8333), .B2(n9933), .A(n8332), .ZN(n8404) );
  MUX2_X1 U9858 ( .A(n8334), .B(n8404), .S(n10192), .Z(n8335) );
  OAI21_X1 U9859 ( .B1(n8407), .B2(n8357), .A(n8335), .ZN(P2_U3477) );
  AOI22_X1 U9860 ( .A1(n8337), .A2(n9933), .B1(n9964), .B2(n8336), .ZN(n8338)
         );
  NAND2_X1 U9861 ( .A1(n8339), .A2(n8338), .ZN(n8408) );
  MUX2_X1 U9862 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8408), .S(n10192), .Z(
        P2_U3476) );
  NAND2_X1 U9863 ( .A1(n8340), .A2(n9933), .ZN(n8341) );
  NAND2_X1 U9864 ( .A1(n8342), .A2(n8341), .ZN(n8409) );
  MUX2_X1 U9865 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8409), .S(n10192), .Z(n8343) );
  AOI21_X1 U9866 ( .B1(n5656), .B2(n8411), .A(n8343), .ZN(n8344) );
  INV_X1 U9867 ( .A(n8344), .ZN(P2_U3475) );
  AOI21_X1 U9868 ( .B1(n9964), .B2(n8346), .A(n8345), .ZN(n8347) );
  OAI21_X1 U9869 ( .B1(n9959), .B2(n8348), .A(n8347), .ZN(n8413) );
  MUX2_X1 U9870 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8413), .S(n10192), .Z(
        P2_U3474) );
  AOI21_X1 U9871 ( .B1(n8350), .B2(n9933), .A(n8349), .ZN(n8414) );
  MUX2_X1 U9872 ( .A(n8351), .B(n8414), .S(n10192), .Z(n8352) );
  OAI21_X1 U9873 ( .B1(n8416), .B2(n8357), .A(n8352), .ZN(P2_U3473) );
  AOI21_X1 U9874 ( .B1(n8354), .B2(n9933), .A(n8353), .ZN(n8417) );
  MUX2_X1 U9875 ( .A(n8355), .B(n8417), .S(n10192), .Z(n8356) );
  OAI21_X1 U9876 ( .B1(n8421), .B2(n8357), .A(n8356), .ZN(P2_U3472) );
  NAND2_X1 U9877 ( .A1(n9959), .A2(n8358), .ZN(n8359) );
  NAND2_X1 U9878 ( .A1(n8360), .A2(n8359), .ZN(n8363) );
  INV_X1 U9879 ( .A(n8361), .ZN(n8362) );
  OAI211_X1 U9880 ( .C1(n9947), .C2(n8364), .A(n8363), .B(n8362), .ZN(n8422)
         );
  MUX2_X1 U9881 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8422), .S(n10192), .Z(
        P2_U3459) );
  NOR2_X1 U9882 ( .A1(n8365), .A2(n9966), .ZN(n8368) );
  AOI21_X1 U9883 ( .B1(n9966), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8368), .ZN(
        n8366) );
  OAI21_X1 U9884 ( .B1(n8367), .B2(n8420), .A(n8366), .ZN(P2_U3458) );
  AOI21_X1 U9885 ( .B1(n9966), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8368), .ZN(
        n8369) );
  OAI21_X1 U9886 ( .B1(n8370), .B2(n8420), .A(n8369), .ZN(P2_U3457) );
  INV_X1 U9887 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8372) );
  INV_X1 U9888 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8375) );
  MUX2_X1 U9889 ( .A(n8375), .B(n8374), .S(n9965), .Z(n8376) );
  OAI21_X1 U9890 ( .B1(n8377), .B2(n8420), .A(n8376), .ZN(P2_U3454) );
  MUX2_X1 U9891 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8378), .S(n9965), .Z(
        P2_U3453) );
  INV_X1 U9892 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8380) );
  MUX2_X1 U9893 ( .A(n8380), .B(n8379), .S(n9965), .Z(n8381) );
  OAI21_X1 U9894 ( .B1(n8382), .B2(n8420), .A(n8381), .ZN(P2_U3452) );
  INV_X1 U9895 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8384) );
  MUX2_X1 U9896 ( .A(n8384), .B(n8383), .S(n9965), .Z(n8385) );
  OAI21_X1 U9897 ( .B1(n8386), .B2(n8420), .A(n8385), .ZN(P2_U3451) );
  INV_X1 U9898 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8388) );
  MUX2_X1 U9899 ( .A(n8388), .B(n8387), .S(n9965), .Z(n8389) );
  OAI21_X1 U9900 ( .B1(n8390), .B2(n8420), .A(n8389), .ZN(P2_U3450) );
  MUX2_X1 U9901 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8391), .S(n9965), .Z(
        P2_U3449) );
  INV_X1 U9902 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8393) );
  MUX2_X1 U9903 ( .A(n8393), .B(n8392), .S(n9965), .Z(n8394) );
  OAI21_X1 U9904 ( .B1(n8395), .B2(n8420), .A(n8394), .ZN(P2_U3448) );
  INV_X1 U9905 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8397) );
  MUX2_X1 U9906 ( .A(n8397), .B(n8396), .S(n9965), .Z(n8398) );
  OAI21_X1 U9907 ( .B1(n8399), .B2(n8420), .A(n8398), .ZN(P2_U3447) );
  INV_X1 U9908 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8401) );
  MUX2_X1 U9909 ( .A(n8401), .B(n8400), .S(n9965), .Z(n8402) );
  OAI21_X1 U9910 ( .B1(n8403), .B2(n8420), .A(n8402), .ZN(P2_U3446) );
  MUX2_X1 U9911 ( .A(n8405), .B(n8404), .S(n9965), .Z(n8406) );
  OAI21_X1 U9912 ( .B1(n8407), .B2(n8420), .A(n8406), .ZN(P2_U3444) );
  MUX2_X1 U9913 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8408), .S(n9965), .Z(
        P2_U3441) );
  MUX2_X1 U9914 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8409), .S(n9965), .Z(n8410)
         );
  AOI21_X1 U9915 ( .B1(n5643), .B2(n8411), .A(n8410), .ZN(n8412) );
  INV_X1 U9916 ( .A(n8412), .ZN(P2_U3438) );
  MUX2_X1 U9917 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8413), .S(n9965), .Z(
        P2_U3435) );
  MUX2_X1 U9918 ( .A(n10003), .B(n8414), .S(n9965), .Z(n8415) );
  OAI21_X1 U9919 ( .B1(n8416), .B2(n8420), .A(n8415), .ZN(P2_U3432) );
  INV_X1 U9920 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8418) );
  MUX2_X1 U9921 ( .A(n8418), .B(n8417), .S(n9965), .Z(n8419) );
  OAI21_X1 U9922 ( .B1(n8421), .B2(n8420), .A(n8419), .ZN(P2_U3429) );
  MUX2_X1 U9923 ( .A(n8422), .B(P2_REG0_REG_0__SCAN_IN), .S(n9966), .Z(
        P2_U3390) );
  MUX2_X1 U9924 ( .A(n8424), .B(P2_D_REG_1__SCAN_IN), .S(n8423), .Z(P2_U3377)
         );
  INV_X1 U9925 ( .A(n8831), .ZN(n9742) );
  NOR4_X1 U9926 ( .A1(n8426), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5031), .ZN(n8427) );
  AOI21_X1 U9927 ( .B1(n8438), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8427), .ZN(
        n8428) );
  OAI21_X1 U9928 ( .B1(n9742), .B2(n7151), .A(n8428), .ZN(P2_U3264) );
  AOI22_X1 U9929 ( .A1(n8429), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8438), .ZN(n8430) );
  OAI21_X1 U9930 ( .B1(n8431), .B2(n7151), .A(n8430), .ZN(P2_U3265) );
  AOI22_X1 U9931 ( .A1(n8432), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8438), .ZN(n8433) );
  OAI21_X1 U9932 ( .B1(n9743), .B2(n7151), .A(n8433), .ZN(P2_U3266) );
  INV_X1 U9933 ( .A(n8434), .ZN(n9746) );
  AOI21_X1 U9934 ( .B1(n8438), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8435), .ZN(
        n8436) );
  OAI21_X1 U9935 ( .B1(n9746), .B2(n7151), .A(n8436), .ZN(P2_U3267) );
  AOI21_X1 U9936 ( .B1(n8438), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8437), .ZN(
        n8439) );
  OAI21_X1 U9937 ( .B1(n8440), .B2(n7151), .A(n8439), .ZN(P2_U3268) );
  MUX2_X1 U9938 ( .A(n8441), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U9939 ( .A1(n8757), .A2(n8646), .ZN(n8443) );
  OR2_X1 U9940 ( .A1(n8690), .A2(n8541), .ZN(n8442) );
  NAND2_X1 U9941 ( .A1(n8443), .A2(n8442), .ZN(n8444) );
  XNOR2_X1 U9942 ( .A(n8444), .B(n8565), .ZN(n8478) );
  AOI22_X1 U9943 ( .A1(n8757), .A2(n8640), .B1(n8567), .B2(n9131), .ZN(n8476)
         );
  INV_X1 U9944 ( .A(n8476), .ZN(n8477) );
  NAND2_X1 U9945 ( .A1(n8450), .A2(n8646), .ZN(n8446) );
  OR2_X1 U9946 ( .A1(n8448), .A2(n8541), .ZN(n8445) );
  NAND2_X1 U9947 ( .A1(n8446), .A2(n8445), .ZN(n8447) );
  XNOR2_X1 U9948 ( .A(n8447), .B(n8644), .ZN(n8457) );
  NOR2_X1 U9949 ( .A1(n8448), .A2(n8641), .ZN(n8449) );
  AOI21_X1 U9950 ( .B1(n8450), .B2(n8496), .A(n8449), .ZN(n8456) );
  XNOR2_X1 U9951 ( .A(n8457), .B(n8456), .ZN(n8735) );
  INV_X1 U9952 ( .A(n8452), .ZN(n8453) );
  NAND2_X1 U9953 ( .A1(n8624), .A2(n8646), .ZN(n8459) );
  OR2_X1 U9954 ( .A1(n8461), .A2(n8541), .ZN(n8458) );
  NAND2_X1 U9955 ( .A1(n8459), .A2(n8458), .ZN(n8460) );
  XNOR2_X1 U9956 ( .A(n8460), .B(n8644), .ZN(n8679) );
  NOR2_X1 U9957 ( .A1(n8461), .A2(n8641), .ZN(n8462) );
  AOI21_X1 U9958 ( .B1(n8624), .B2(n8640), .A(n8462), .ZN(n8680) );
  NAND2_X1 U9959 ( .A1(n9733), .A2(n8646), .ZN(n8464) );
  OR2_X1 U9960 ( .A1(n8689), .A2(n8541), .ZN(n8463) );
  NAND2_X1 U9961 ( .A1(n8464), .A2(n8463), .ZN(n8465) );
  XNOR2_X1 U9962 ( .A(n8465), .B(n8644), .ZN(n8468) );
  NOR2_X1 U9963 ( .A1(n8689), .A2(n8641), .ZN(n8466) );
  AOI21_X1 U9964 ( .B1(n9733), .B2(n8496), .A(n8466), .ZN(n8467) );
  OAI21_X1 U9965 ( .B1(n8679), .B2(n8680), .A(n8682), .ZN(n8470) );
  NAND3_X1 U9966 ( .A1(n8682), .A2(n8679), .A3(n8680), .ZN(n8469) );
  NAND2_X1 U9967 ( .A1(n8468), .A2(n8467), .ZN(n8683) );
  AOI22_X1 U9968 ( .A1(n9729), .A2(n8646), .B1(n8496), .B2(n9132), .ZN(n8471)
         );
  XOR2_X1 U9969 ( .A(n8565), .B(n8471), .Z(n8473) );
  OAI22_X1 U9970 ( .A1(n7545), .A2(n8541), .B1(n8762), .B2(n8641), .ZN(n8472)
         );
  NOR2_X1 U9971 ( .A1(n8473), .A2(n8472), .ZN(n8474) );
  AOI21_X1 U9972 ( .B1(n8473), .B2(n8472), .A(n8474), .ZN(n8684) );
  INV_X1 U9973 ( .A(n8474), .ZN(n8475) );
  XNOR2_X1 U9974 ( .A(n8478), .B(n8476), .ZN(n8760) );
  AOI22_X1 U9975 ( .A1(n9657), .A2(n8646), .B1(n8496), .B2(n9130), .ZN(n8479)
         );
  XNOR2_X1 U9976 ( .A(n8479), .B(n8565), .ZN(n8480) );
  AOI22_X1 U9977 ( .A1(n9657), .A2(n8640), .B1(n8567), .B2(n9130), .ZN(n8598)
         );
  AOI22_X1 U9978 ( .A1(n9649), .A2(n8646), .B1(n8496), .B2(n9129), .ZN(n8482)
         );
  XNOR2_X1 U9979 ( .A(n8482), .B(n8565), .ZN(n8484) );
  INV_X1 U9980 ( .A(n8484), .ZN(n8483) );
  AOI22_X1 U9981 ( .A1(n9649), .A2(n8496), .B1(n8567), .B2(n9129), .ZN(n8814)
         );
  NAND2_X1 U9982 ( .A1(n9645), .A2(n8646), .ZN(n8488) );
  INV_X1 U9983 ( .A(n8820), .ZN(n9127) );
  NAND2_X1 U9984 ( .A1(n9127), .A2(n8640), .ZN(n8487) );
  NAND2_X1 U9985 ( .A1(n8488), .A2(n8487), .ZN(n8489) );
  XNOR2_X1 U9986 ( .A(n8489), .B(n8644), .ZN(n8492) );
  INV_X1 U9987 ( .A(n8492), .ZN(n8494) );
  NOR2_X1 U9988 ( .A1(n8820), .A2(n8641), .ZN(n8490) );
  AOI21_X1 U9989 ( .B1(n9645), .B2(n8496), .A(n8490), .ZN(n8491) );
  INV_X1 U9990 ( .A(n8491), .ZN(n8493) );
  AOI21_X1 U9991 ( .B1(n8494), .B2(n8493), .A(n8716), .ZN(n8706) );
  INV_X1 U9992 ( .A(n8716), .ZN(n8495) );
  NAND2_X1 U9993 ( .A1(n9466), .A2(n8646), .ZN(n8498) );
  OR2_X1 U9994 ( .A1(n8709), .A2(n8541), .ZN(n8497) );
  NAND2_X1 U9995 ( .A1(n8498), .A2(n8497), .ZN(n8499) );
  XNOR2_X1 U9996 ( .A(n8499), .B(n8644), .ZN(n8502) );
  NOR2_X1 U9997 ( .A1(n8709), .A2(n8641), .ZN(n8500) );
  AOI21_X1 U9998 ( .B1(n9466), .B2(n8640), .A(n8500), .ZN(n8501) );
  NAND2_X1 U9999 ( .A1(n8502), .A2(n8501), .ZN(n8788) );
  OR2_X1 U10000 ( .A1(n8502), .A2(n8501), .ZN(n8503) );
  AND2_X1 U10001 ( .A1(n8788), .A2(n8503), .ZN(n8715) );
  NAND2_X1 U10002 ( .A1(n8504), .A2(n8715), .ZN(n8718) );
  NAND2_X1 U10003 ( .A1(n8718), .A2(n8788), .ZN(n8513) );
  NAND2_X1 U10004 ( .A1(n9634), .A2(n8646), .ZN(n8506) );
  NAND2_X1 U10005 ( .A1(n9125), .A2(n8640), .ZN(n8505) );
  NAND2_X1 U10006 ( .A1(n8506), .A2(n8505), .ZN(n8507) );
  XNOR2_X1 U10007 ( .A(n8507), .B(n8644), .ZN(n8511) );
  NOR2_X1 U10008 ( .A1(n8508), .A2(n8641), .ZN(n8509) );
  AOI21_X1 U10009 ( .B1(n9634), .B2(n8640), .A(n8509), .ZN(n8510) );
  NAND2_X1 U10010 ( .A1(n8511), .A2(n8510), .ZN(n8629) );
  OR2_X1 U10011 ( .A1(n8511), .A2(n8510), .ZN(n8512) );
  AND2_X1 U10012 ( .A1(n8629), .A2(n8512), .ZN(n8789) );
  NAND2_X1 U10013 ( .A1(n8513), .A2(n8789), .ZN(n8628) );
  NAND2_X1 U10014 ( .A1(n9432), .A2(n8646), .ZN(n8515) );
  NAND2_X1 U10015 ( .A1(n9124), .A2(n8640), .ZN(n8514) );
  NAND2_X1 U10016 ( .A1(n8515), .A2(n8514), .ZN(n8516) );
  XNOR2_X1 U10017 ( .A(n8516), .B(n8644), .ZN(n8518) );
  AND2_X1 U10018 ( .A1(n9124), .A2(n8567), .ZN(n8517) );
  AOI21_X1 U10019 ( .B1(n9432), .B2(n8496), .A(n8517), .ZN(n8519) );
  NAND2_X1 U10020 ( .A1(n8518), .A2(n8519), .ZN(n8744) );
  INV_X1 U10021 ( .A(n8518), .ZN(n8521) );
  INV_X1 U10022 ( .A(n8519), .ZN(n8520) );
  NAND2_X1 U10023 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  AND2_X1 U10024 ( .A1(n8744), .A2(n8522), .ZN(n8630) );
  NAND2_X1 U10025 ( .A1(n9625), .A2(n8646), .ZN(n8524) );
  OR2_X1 U10026 ( .A1(n8669), .A2(n8541), .ZN(n8523) );
  NAND2_X1 U10027 ( .A1(n8524), .A2(n8523), .ZN(n8525) );
  XNOR2_X1 U10028 ( .A(n8525), .B(n8644), .ZN(n8528) );
  NOR2_X1 U10029 ( .A1(n8669), .A2(n8641), .ZN(n8526) );
  AOI21_X1 U10030 ( .B1(n9625), .B2(n8496), .A(n8526), .ZN(n8527) );
  NAND2_X1 U10031 ( .A1(n8528), .A2(n8527), .ZN(n8530) );
  OR2_X1 U10032 ( .A1(n8528), .A2(n8527), .ZN(n8529) );
  AND2_X1 U10033 ( .A1(n8530), .A2(n8529), .ZN(n8745) );
  NAND2_X1 U10034 ( .A1(n8748), .A2(n8530), .ZN(n8665) );
  OAI22_X1 U10035 ( .A1(n9712), .A2(n6166), .B1(n8771), .B2(n8641), .ZN(n8534)
         );
  NAND2_X1 U10036 ( .A1(n9404), .A2(n8646), .ZN(n8532) );
  OR2_X1 U10037 ( .A1(n8771), .A2(n8541), .ZN(n8531) );
  NAND2_X1 U10038 ( .A1(n8532), .A2(n8531), .ZN(n8533) );
  XNOR2_X1 U10039 ( .A(n8533), .B(n8565), .ZN(n8535) );
  XOR2_X1 U10040 ( .A(n8534), .B(n8535), .Z(n8666) );
  AOI22_X1 U10041 ( .A1(n9387), .A2(n8646), .B1(n8496), .B2(n9121), .ZN(n8537)
         );
  XNOR2_X1 U10042 ( .A(n8537), .B(n8565), .ZN(n8538) );
  OAI22_X1 U10043 ( .A1(n4872), .A2(n8541), .B1(n8668), .B2(n8641), .ZN(n8769)
         );
  NAND2_X1 U10044 ( .A1(n9372), .A2(n8646), .ZN(n8543) );
  OR2_X1 U10045 ( .A1(n4334), .A2(n6166), .ZN(n8542) );
  NAND2_X1 U10046 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  XNOR2_X1 U10047 ( .A(n8544), .B(n8644), .ZN(n8547) );
  NOR2_X1 U10048 ( .A1(n4334), .A2(n8641), .ZN(n8545) );
  AOI21_X1 U10049 ( .B1(n9372), .B2(n8496), .A(n8545), .ZN(n8546) );
  NAND2_X1 U10050 ( .A1(n8547), .A2(n8546), .ZN(n8728) );
  OR2_X1 U10051 ( .A1(n8547), .A2(n8546), .ZN(n8548) );
  NAND2_X1 U10052 ( .A1(n9358), .A2(n8646), .ZN(n8551) );
  OR2_X1 U10053 ( .A1(n8612), .A2(n8541), .ZN(n8550) );
  NAND2_X1 U10054 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  XNOR2_X1 U10055 ( .A(n8552), .B(n8644), .ZN(n8555) );
  NOR2_X1 U10056 ( .A1(n8612), .A2(n8641), .ZN(n8553) );
  AOI21_X1 U10057 ( .B1(n9358), .B2(n8640), .A(n8553), .ZN(n8554) );
  NAND2_X1 U10058 ( .A1(n8555), .A2(n8554), .ZN(n8558) );
  OR2_X1 U10059 ( .A1(n8555), .A2(n8554), .ZN(n8556) );
  OAI22_X1 U10060 ( .A1(n9697), .A2(n8541), .B1(n8559), .B2(n8641), .ZN(n8570)
         );
  NAND2_X1 U10061 ( .A1(n9339), .A2(n8646), .ZN(n8561) );
  NAND2_X1 U10062 ( .A1(n9118), .A2(n8640), .ZN(n8560) );
  NAND2_X1 U10063 ( .A1(n8561), .A2(n8560), .ZN(n8562) );
  XNOR2_X1 U10064 ( .A(n8562), .B(n8565), .ZN(n8569) );
  XOR2_X1 U10065 ( .A(n8570), .B(n8569), .Z(n8698) );
  NAND2_X1 U10066 ( .A1(n9323), .A2(n8646), .ZN(n8564) );
  NAND2_X1 U10067 ( .A1(n9117), .A2(n8640), .ZN(n8563) );
  NAND2_X1 U10068 ( .A1(n8564), .A2(n8563), .ZN(n8566) );
  XNOR2_X1 U10069 ( .A(n8566), .B(n8565), .ZN(n8576) );
  AND2_X1 U10070 ( .A1(n9117), .A2(n8567), .ZN(n8568) );
  AOI21_X1 U10071 ( .B1(n9323), .B2(n8496), .A(n8568), .ZN(n8574) );
  XNOR2_X1 U10072 ( .A(n8576), .B(n8574), .ZN(n8801) );
  INV_X1 U10073 ( .A(n8569), .ZN(n8572) );
  INV_X1 U10074 ( .A(n8570), .ZN(n8571) );
  NAND2_X1 U10075 ( .A1(n8572), .A2(n8571), .ZN(n8799) );
  INV_X1 U10076 ( .A(n8574), .ZN(n8575) );
  NAND2_X1 U10077 ( .A1(n8576), .A2(n8575), .ZN(n8586) );
  NAND2_X1 U10078 ( .A1(n9593), .A2(n8646), .ZN(n8578) );
  OR2_X1 U10079 ( .A1(n8803), .A2(n8541), .ZN(n8577) );
  NAND2_X1 U10080 ( .A1(n8578), .A2(n8577), .ZN(n8579) );
  XNOR2_X1 U10081 ( .A(n8579), .B(n8644), .ZN(n8582) );
  INV_X1 U10082 ( .A(n8582), .ZN(n8584) );
  NOR2_X1 U10083 ( .A1(n8803), .A2(n8641), .ZN(n8580) );
  AOI21_X1 U10084 ( .B1(n9593), .B2(n8640), .A(n8580), .ZN(n8581) );
  INV_X1 U10085 ( .A(n8581), .ZN(n8583) );
  AOI21_X1 U10086 ( .B1(n8584), .B2(n8583), .A(n8658), .ZN(n8585) );
  AOI21_X1 U10087 ( .B1(n8590), .B2(n8586), .A(n8585), .ZN(n8591) );
  INV_X1 U10088 ( .A(n8585), .ZN(n8588) );
  INV_X1 U10089 ( .A(n8586), .ZN(n8587) );
  NOR2_X1 U10090 ( .A1(n8588), .A2(n8587), .ZN(n8589) );
  OAI21_X1 U10091 ( .B1(n8591), .B2(n8653), .A(n8816), .ZN(n8595) );
  AOI22_X1 U10092 ( .A1(n9309), .A2(n8825), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8594) );
  NAND2_X1 U10093 ( .A1(n9593), .A2(n8784), .ZN(n8593) );
  OAI22_X1 U10094 ( .A1(n8999), .A2(n9281), .B1(n9280), .B2(n8819), .ZN(n9304)
         );
  NAND2_X1 U10095 ( .A1(n9304), .A2(n8810), .ZN(n8592) );
  NAND4_X1 U10096 ( .A1(n8595), .A2(n8594), .A3(n8593), .A4(n8592), .ZN(
        P1_U3214) );
  OAI21_X1 U10097 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(n8599) );
  NAND2_X1 U10098 ( .A1(n8599), .A2(n8816), .ZN(n8605) );
  OR2_X1 U10099 ( .A1(n8690), .A2(n9281), .ZN(n8601) );
  NAND2_X1 U10100 ( .A1(n9129), .A2(n9259), .ZN(n8600) );
  AND2_X1 U10101 ( .A1(n8601), .A2(n8600), .ZN(n9511) );
  OAI21_X1 U10102 ( .B1(n9511), .B2(n8822), .A(n8602), .ZN(n8603) );
  AOI21_X1 U10103 ( .B1(n9514), .B2(n8825), .A(n8603), .ZN(n8604) );
  OAI211_X1 U10104 ( .C1(n9517), .C2(n8828), .A(n8605), .B(n8604), .ZN(
        P1_U3215) );
  INV_X1 U10105 ( .A(n9372), .ZN(n9705) );
  INV_X1 U10106 ( .A(n8606), .ZN(n8608) );
  NOR3_X1 U10107 ( .A1(n4361), .A2(n8608), .A3(n8607), .ZN(n8611) );
  INV_X1 U10108 ( .A(n8609), .ZN(n8610) );
  OAI21_X1 U10109 ( .B1(n8611), .B2(n8610), .A(n8816), .ZN(n8619) );
  OR2_X1 U10110 ( .A1(n8612), .A2(n8819), .ZN(n8614) );
  OR2_X1 U10111 ( .A1(n8668), .A2(n9281), .ZN(n8613) );
  NAND2_X1 U10112 ( .A1(n8614), .A2(n8613), .ZN(n9368) );
  OAI22_X1 U10113 ( .A1(n8616), .A2(n8808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8615), .ZN(n8617) );
  AOI21_X1 U10114 ( .B1(n9368), .B2(n8810), .A(n8617), .ZN(n8618) );
  OAI211_X1 U10115 ( .C1(n9705), .C2(n8828), .A(n8619), .B(n8618), .ZN(
        P1_U3216) );
  XOR2_X1 U10116 ( .A(n8679), .B(n8677), .Z(n8681) );
  XNOR2_X1 U10117 ( .A(n8681), .B(n8680), .ZN(n8627) );
  OAI22_X1 U10118 ( .A1(n8621), .A2(n8822), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8620), .ZN(n8622) );
  AOI21_X1 U10119 ( .B1(n8623), .B2(n8825), .A(n8622), .ZN(n8626) );
  NAND2_X1 U10120 ( .A1(n8624), .A2(n8784), .ZN(n8625) );
  OAI211_X1 U10121 ( .C1(n8627), .C2(n8786), .A(n8626), .B(n8625), .ZN(
        P1_U3217) );
  INV_X1 U10122 ( .A(n8628), .ZN(n8792) );
  INV_X1 U10123 ( .A(n8629), .ZN(n8631) );
  NOR3_X1 U10124 ( .A1(n8792), .A2(n8631), .A3(n8630), .ZN(n8633) );
  INV_X1 U10125 ( .A(n8632), .ZN(n8747) );
  OAI21_X1 U10126 ( .B1(n8633), .B2(n8747), .A(n8816), .ZN(n8639) );
  OR2_X1 U10127 ( .A1(n8669), .A2(n8819), .ZN(n8635) );
  NAND2_X1 U10128 ( .A1(n9125), .A2(n8804), .ZN(n8634) );
  NAND2_X1 U10129 ( .A1(n8635), .A2(n8634), .ZN(n9426) );
  NOR2_X1 U10130 ( .A1(n8808), .A2(n9434), .ZN(n8636) );
  AOI211_X1 U10131 ( .C1(n9426), .C2(n8810), .A(n8637), .B(n8636), .ZN(n8638)
         );
  OAI211_X1 U10132 ( .C1(n9717), .C2(n8828), .A(n8639), .B(n8638), .ZN(
        P1_U3219) );
  INV_X1 U10133 ( .A(n8653), .ZN(n8652) );
  INV_X1 U10134 ( .A(n8658), .ZN(n8651) );
  NAND2_X1 U10135 ( .A1(n9269), .A2(n8640), .ZN(n8643) );
  OR2_X1 U10136 ( .A1(n9280), .A2(n8641), .ZN(n8642) );
  NAND2_X1 U10137 ( .A1(n8643), .A2(n8642), .ZN(n8645) );
  XNOR2_X1 U10138 ( .A(n8645), .B(n8644), .ZN(n8649) );
  NAND2_X1 U10139 ( .A1(n9269), .A2(n8646), .ZN(n8647) );
  OAI21_X1 U10140 ( .B1(n9280), .B2(n8541), .A(n8647), .ZN(n8648) );
  XNOR2_X1 U10141 ( .A(n8649), .B(n8648), .ZN(n8659) );
  INV_X1 U10142 ( .A(n8659), .ZN(n8650) );
  NAND4_X1 U10143 ( .A1(n8652), .A2(n8651), .A3(n8650), .A4(n8816), .ZN(n8663)
         );
  NAND3_X1 U10144 ( .A1(n8653), .A2(n8816), .A3(n8659), .ZN(n8662) );
  INV_X1 U10145 ( .A(n8654), .ZN(n8656) );
  AOI22_X1 U10146 ( .A1(n8825), .A2(n9293), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8655) );
  OAI21_X1 U10147 ( .B1(n8656), .B2(n8822), .A(n8655), .ZN(n8657) );
  AOI21_X1 U10148 ( .B1(n9269), .B2(n8784), .A(n8657), .ZN(n8661) );
  NAND3_X1 U10149 ( .A1(n8659), .A2(n8816), .A3(n8658), .ZN(n8660) );
  NAND4_X1 U10150 ( .A1(n8663), .A2(n8662), .A3(n8661), .A4(n8660), .ZN(
        P1_U3220) );
  OAI21_X1 U10151 ( .B1(n8666), .B2(n8665), .A(n8664), .ZN(n8667) );
  NAND2_X1 U10152 ( .A1(n8667), .A2(n8816), .ZN(n8676) );
  OR2_X1 U10153 ( .A1(n8668), .A2(n8819), .ZN(n8671) );
  OR2_X1 U10154 ( .A1(n8669), .A2(n9281), .ZN(n8670) );
  NAND2_X1 U10155 ( .A1(n8671), .A2(n8670), .ZN(n9400) );
  INV_X1 U10156 ( .A(n9405), .ZN(n8673) );
  INV_X1 U10157 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8672) );
  OAI22_X1 U10158 ( .A1(n8673), .A2(n8808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8672), .ZN(n8674) );
  AOI21_X1 U10159 ( .B1(n9400), .B2(n8810), .A(n8674), .ZN(n8675) );
  OAI211_X1 U10160 ( .C1(n9712), .C2(n8828), .A(n8676), .B(n8675), .ZN(
        P1_U3223) );
  INV_X1 U10161 ( .A(n8677), .ZN(n8678) );
  OAI22_X1 U10162 ( .A1(n8681), .A2(n8680), .B1(n8679), .B2(n8678), .ZN(n8780)
         );
  NAND2_X1 U10163 ( .A1(n8682), .A2(n8683), .ZN(n8779) );
  NOR2_X1 U10164 ( .A1(n8780), .A2(n8779), .ZN(n8778) );
  INV_X1 U10165 ( .A(n8683), .ZN(n8685) );
  NOR3_X1 U10166 ( .A1(n8778), .A2(n8685), .A3(n8684), .ZN(n8688) );
  INV_X1 U10167 ( .A(n8686), .ZN(n8687) );
  OAI21_X1 U10168 ( .B1(n8688), .B2(n8687), .A(n8816), .ZN(n8696) );
  OR2_X1 U10169 ( .A1(n8689), .A2(n9281), .ZN(n8692) );
  OR2_X1 U10170 ( .A1(n8690), .A2(n8819), .ZN(n8691) );
  AND2_X1 U10171 ( .A1(n8692), .A2(n8691), .ZN(n9544) );
  OAI21_X1 U10172 ( .B1(n9544), .B2(n8822), .A(n8693), .ZN(n8694) );
  AOI21_X1 U10173 ( .B1(n9546), .B2(n8825), .A(n8694), .ZN(n8695) );
  OAI211_X1 U10174 ( .C1(n7545), .C2(n8828), .A(n8696), .B(n8695), .ZN(
        P1_U3224) );
  NAND2_X1 U10175 ( .A1(n8699), .A2(n8816), .ZN(n8703) );
  NOR2_X1 U10176 ( .A1(n9340), .A2(n8808), .ZN(n8701) );
  AOI22_X1 U10177 ( .A1(n9117), .A2(n9259), .B1(n9119), .B2(n8804), .ZN(n9335)
         );
  NOR2_X1 U10178 ( .A1(n9335), .A2(n8822), .ZN(n8700) );
  AOI211_X1 U10179 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(P1_U3086), .A(n8701), 
        .B(n8700), .ZN(n8702) );
  OAI211_X1 U10180 ( .C1(n9697), .C2(n8828), .A(n8703), .B(n8702), .ZN(
        P1_U3225) );
  OAI21_X1 U10181 ( .B1(n8706), .B2(n8705), .A(n8704), .ZN(n8707) );
  NAND2_X1 U10182 ( .A1(n8707), .A2(n8816), .ZN(n8714) );
  OAI22_X1 U10183 ( .A1(n8709), .A2(n8819), .B1(n8708), .B2(n9281), .ZN(n9483)
         );
  NOR2_X1 U10184 ( .A1(n8808), .A2(n8710), .ZN(n8711) );
  AOI211_X1 U10185 ( .C1(n8810), .C2(n9483), .A(n8712), .B(n8711), .ZN(n8713)
         );
  OAI211_X1 U10186 ( .C1(n9479), .C2(n8828), .A(n8714), .B(n8713), .ZN(
        P1_U3226) );
  INV_X1 U10187 ( .A(n8704), .ZN(n8717) );
  NOR3_X1 U10188 ( .A1(n8717), .A2(n8716), .A3(n8715), .ZN(n8719) );
  INV_X1 U10189 ( .A(n8718), .ZN(n8791) );
  OAI21_X1 U10190 ( .B1(n8719), .B2(n8791), .A(n8816), .ZN(n8723) );
  NOR2_X1 U10191 ( .A1(n8820), .A2(n9281), .ZN(n8720) );
  AOI21_X1 U10192 ( .B1(n9125), .B2(n9259), .A(n8720), .ZN(n9462) );
  NAND2_X1 U10193 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9786) );
  OAI21_X1 U10194 ( .B1(n9462), .B2(n8822), .A(n9786), .ZN(n8721) );
  AOI21_X1 U10195 ( .B1(n9467), .B2(n8825), .A(n8721), .ZN(n8722) );
  OAI211_X1 U10196 ( .C1(n4875), .C2(n8828), .A(n8723), .B(n8722), .ZN(
        P1_U3228) );
  NAND2_X1 U10197 ( .A1(n9118), .A2(n9259), .ZN(n8725) );
  OR2_X1 U10198 ( .A1(n4334), .A2(n9281), .ZN(n8724) );
  AND2_X1 U10199 ( .A1(n8725), .A2(n8724), .ZN(n9353) );
  AOI22_X1 U10200 ( .A1(n9359), .A2(n8825), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8726) );
  OAI21_X1 U10201 ( .B1(n9353), .B2(n8822), .A(n8726), .ZN(n8732) );
  NAND3_X1 U10202 ( .A1(n8609), .A2(n8728), .A3(n4859), .ZN(n8729) );
  AOI21_X1 U10203 ( .B1(n8730), .B2(n8729), .A(n8786), .ZN(n8731) );
  INV_X1 U10204 ( .A(n8733), .ZN(n8734) );
  AND3_X1 U10205 ( .A1(n8736), .A2(n8735), .A3(n8734), .ZN(n8738) );
  OAI21_X1 U10206 ( .B1(n8738), .B2(n8737), .A(n8816), .ZN(n8743) );
  NAND2_X1 U10207 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9769) );
  OAI21_X1 U10208 ( .B1(n8739), .B2(n8822), .A(n9769), .ZN(n8740) );
  AOI21_X1 U10209 ( .B1(n8741), .B2(n8825), .A(n8740), .ZN(n8742) );
  OAI211_X1 U10210 ( .C1(n9806), .C2(n8828), .A(n8743), .B(n8742), .ZN(
        P1_U3231) );
  INV_X1 U10211 ( .A(n8744), .ZN(n8746) );
  NOR3_X1 U10212 ( .A1(n8747), .A2(n8746), .A3(n8745), .ZN(n8750) );
  INV_X1 U10213 ( .A(n8748), .ZN(n8749) );
  OAI21_X1 U10214 ( .B1(n8750), .B2(n8749), .A(n8816), .ZN(n8756) );
  OR2_X1 U10215 ( .A1(n8771), .A2(n8819), .ZN(n8752) );
  NAND2_X1 U10216 ( .A1(n9124), .A2(n8804), .ZN(n8751) );
  AND2_X1 U10217 ( .A1(n8752), .A2(n8751), .ZN(n9413) );
  OAI22_X1 U10218 ( .A1(n9413), .A2(n8822), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8753), .ZN(n8754) );
  AOI21_X1 U10219 ( .B1(n9418), .B2(n8825), .A(n8754), .ZN(n8755) );
  OAI211_X1 U10220 ( .C1(n9421), .C2(n8828), .A(n8756), .B(n8755), .ZN(
        P1_U3233) );
  OAI21_X1 U10221 ( .B1(n8760), .B2(n8759), .A(n8758), .ZN(n8761) );
  NAND2_X1 U10222 ( .A1(n8761), .A2(n8816), .ZN(n8767) );
  OR2_X1 U10223 ( .A1(n8818), .A2(n8819), .ZN(n8764) );
  OR2_X1 U10224 ( .A1(n8762), .A2(n9281), .ZN(n8763) );
  AND2_X1 U10225 ( .A1(n8764), .A2(n8763), .ZN(n9529) );
  NAND2_X1 U10226 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9246) );
  OAI21_X1 U10227 ( .B1(n9529), .B2(n8822), .A(n9246), .ZN(n8765) );
  AOI21_X1 U10228 ( .B1(n9533), .B2(n8825), .A(n8765), .ZN(n8766) );
  OAI211_X1 U10229 ( .C1(n4870), .C2(n8828), .A(n8767), .B(n8766), .ZN(
        P1_U3234) );
  AOI21_X1 U10230 ( .B1(n8769), .B2(n8768), .A(n4361), .ZN(n8777) );
  OR2_X1 U10231 ( .A1(n4334), .A2(n8819), .ZN(n8773) );
  OR2_X1 U10232 ( .A1(n8771), .A2(n9281), .ZN(n8772) );
  AND2_X1 U10233 ( .A1(n8773), .A2(n8772), .ZN(n9383) );
  AOI22_X1 U10234 ( .A1(n9388), .A2(n8825), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8774) );
  OAI21_X1 U10235 ( .B1(n9383), .B2(n8822), .A(n8774), .ZN(n8775) );
  AOI21_X1 U10236 ( .B1(n9387), .B2(n8784), .A(n8775), .ZN(n8776) );
  OAI21_X1 U10237 ( .B1(n8777), .B2(n8786), .A(n8776), .ZN(P1_U3235) );
  AOI21_X1 U10238 ( .B1(n8780), .B2(n8779), .A(n8778), .ZN(n8787) );
  AOI22_X1 U10239 ( .A1(n8804), .A2(n9134), .B1(n9132), .B2(n9259), .ZN(n9562)
         );
  NAND2_X1 U10240 ( .A1(n8825), .A2(n9572), .ZN(n8781) );
  OAI211_X1 U10241 ( .C1(n9562), .C2(n8822), .A(n8782), .B(n8781), .ZN(n8783)
         );
  AOI21_X1 U10242 ( .B1(n4451), .B2(n8784), .A(n8783), .ZN(n8785) );
  OAI21_X1 U10243 ( .B1(n8787), .B2(n8786), .A(n8785), .ZN(P1_U3236) );
  INV_X1 U10244 ( .A(n8788), .ZN(n8790) );
  NOR3_X1 U10245 ( .A1(n8791), .A2(n8790), .A3(n8789), .ZN(n8793) );
  OAI21_X1 U10246 ( .B1(n8793), .B2(n8792), .A(n8816), .ZN(n8798) );
  INV_X1 U10247 ( .A(n8794), .ZN(n9444) );
  AOI22_X1 U10248 ( .A1(n9124), .A2(n9259), .B1(n9126), .B2(n8804), .ZN(n9450)
         );
  OAI21_X1 U10249 ( .B1(n9450), .B2(n8822), .A(n8795), .ZN(n8796) );
  AOI21_X1 U10250 ( .B1(n9444), .B2(n8825), .A(n8796), .ZN(n8797) );
  OAI211_X1 U10251 ( .C1(n9446), .C2(n8828), .A(n8798), .B(n8797), .ZN(
        P1_U3238) );
  AND2_X1 U10252 ( .A1(n8800), .A2(n8799), .ZN(n8802) );
  OAI211_X1 U10253 ( .C1(n8802), .C2(n8801), .A(n8816), .B(n8590), .ZN(n8812)
         );
  OR2_X1 U10254 ( .A1(n8803), .A2(n8819), .ZN(n8806) );
  NAND2_X1 U10255 ( .A1(n9118), .A2(n8804), .ZN(n8805) );
  NAND2_X1 U10256 ( .A1(n8806), .A2(n8805), .ZN(n9317) );
  INV_X1 U10257 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8807) );
  OAI22_X1 U10258 ( .A1(n9325), .A2(n8808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8807), .ZN(n8809) );
  AOI21_X1 U10259 ( .B1(n9317), .B2(n8810), .A(n8809), .ZN(n8811) );
  OAI21_X1 U10260 ( .B1(n8815), .B2(n8814), .A(n8813), .ZN(n8817) );
  NAND2_X1 U10261 ( .A1(n8817), .A2(n8816), .ZN(n8827) );
  OAI22_X1 U10262 ( .A1(n8820), .A2(n8819), .B1(n8818), .B2(n9281), .ZN(n9499)
         );
  INV_X1 U10263 ( .A(n9499), .ZN(n8823) );
  OAI21_X1 U10264 ( .B1(n8823), .B2(n8822), .A(n8821), .ZN(n8824) );
  AOI21_X1 U10265 ( .B1(n9493), .B2(n8825), .A(n8824), .ZN(n8826) );
  OAI211_X1 U10266 ( .C1(n9495), .C2(n8828), .A(n8827), .B(n8826), .ZN(
        P1_U3241) );
  INV_X1 U10267 ( .A(n9021), .ZN(n9030) );
  NOR2_X1 U10268 ( .A1(n8864), .A2(n8829), .ZN(n8830) );
  INV_X1 U10269 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U10270 ( .A1(n8867), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8833) );
  NAND2_X1 U10271 ( .A1(n8868), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8832) );
  OAI211_X1 U10272 ( .C1(n8872), .C2(n8834), .A(n8833), .B(n8832), .ZN(n9114)
         );
  AND2_X1 U10273 ( .A1(n9680), .A2(n9114), .ZN(n9099) );
  INV_X1 U10274 ( .A(n9099), .ZN(n9036) );
  INV_X1 U10275 ( .A(n9680), .ZN(n8875) );
  INV_X1 U10276 ( .A(n9114), .ZN(n9260) );
  INV_X1 U10277 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9745) );
  OR2_X1 U10278 ( .A1(n8864), .A2(n9745), .ZN(n8835) );
  NOR2_X1 U10279 ( .A1(n9587), .A2(n8837), .ZN(n9015) );
  INV_X1 U10280 ( .A(n9015), .ZN(n8876) );
  INV_X1 U10281 ( .A(n9016), .ZN(n8838) );
  INV_X1 U10282 ( .A(n9272), .ZN(n9277) );
  NAND2_X1 U10283 ( .A1(n8982), .A2(n8981), .ZN(n9397) );
  XNOR2_X1 U10284 ( .A(n9625), .B(n9123), .ZN(n9411) );
  NOR2_X1 U10285 ( .A1(n8840), .A2(n8839), .ZN(n8844) );
  NOR2_X1 U10286 ( .A1(n8841), .A2(n9025), .ZN(n8843) );
  NAND4_X1 U10287 ( .A1(n8844), .A2(n8916), .A3(n8843), .A4(n8842), .ZN(n8846)
         );
  NOR2_X1 U10288 ( .A1(n8846), .A2(n8845), .ZN(n8847) );
  NAND4_X1 U10289 ( .A1(n9060), .A2(n4943), .A3(n8848), .A4(n8847), .ZN(n8849)
         );
  NOR3_X1 U10290 ( .A1(n9540), .A2(n9558), .A3(n8849), .ZN(n8850) );
  NAND2_X1 U10291 ( .A1(n9523), .A2(n8850), .ZN(n8851) );
  OR4_X1 U10292 ( .A1(n9474), .A2(n9488), .A3(n9507), .A4(n8851), .ZN(n8852)
         );
  NOR2_X1 U10293 ( .A1(n9459), .A2(n8852), .ZN(n8853) );
  NAND4_X1 U10294 ( .A1(n9411), .A2(n9429), .A3(n9449), .A4(n8853), .ZN(n8854)
         );
  NOR2_X1 U10295 ( .A1(n9397), .A2(n8854), .ZN(n8855) );
  NAND4_X1 U10296 ( .A1(n9347), .A2(n9367), .A3(n9381), .A4(n8855), .ZN(n8856)
         );
  OR3_X1 U10297 ( .A1(n9321), .A2(n8857), .A3(n8856), .ZN(n8859) );
  OR3_X1 U10298 ( .A1(n8859), .A2(n9275), .A3(n8858), .ZN(n8860) );
  NOR2_X1 U10299 ( .A1(n9277), .A2(n8860), .ZN(n8874) );
  NAND2_X1 U10300 ( .A1(n8862), .A2(n8861), .ZN(n8866) );
  OR2_X1 U10301 ( .A1(n8864), .A2(n8863), .ZN(n8865) );
  INV_X1 U10302 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U10303 ( .A1(n8867), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U10304 ( .A1(n8868), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8869) );
  OAI211_X1 U10305 ( .C1(n8872), .C2(n8871), .A(n8870), .B(n8869), .ZN(n9115)
         );
  XNOR2_X1 U10306 ( .A(n9264), .B(n9115), .ZN(n8873) );
  NAND4_X1 U10307 ( .A1(n9036), .A2(n4411), .A3(n8874), .A4(n8873), .ZN(n9023)
         );
  OR2_X1 U10308 ( .A1(n8875), .A2(n9684), .ZN(n8898) );
  INV_X1 U10309 ( .A(n9115), .ZN(n9278) );
  AOI21_X1 U10310 ( .B1(n9264), .B2(n9278), .A(n9016), .ZN(n9097) );
  NAND2_X1 U10311 ( .A1(n8876), .A2(n9006), .ZN(n8896) );
  INV_X1 U10312 ( .A(n9007), .ZN(n8878) );
  INV_X1 U10313 ( .A(n8990), .ZN(n8877) );
  OR3_X1 U10314 ( .A1(n8896), .A2(n8878), .A3(n8877), .ZN(n9090) );
  INV_X1 U10315 ( .A(n9090), .ZN(n8884) );
  NAND2_X1 U10316 ( .A1(n8985), .A2(n8879), .ZN(n8993) );
  NAND2_X1 U10317 ( .A1(n8993), .A2(n8992), .ZN(n8880) );
  NAND2_X1 U10318 ( .A1(n8880), .A2(n8995), .ZN(n8881) );
  NAND2_X1 U10319 ( .A1(n8881), .A2(n8987), .ZN(n8882) );
  NAND2_X1 U10320 ( .A1(n8989), .A2(n8882), .ZN(n8889) );
  OR2_X1 U10321 ( .A1(n8889), .A2(n8910), .ZN(n9086) );
  OAI21_X1 U10322 ( .B1(n9086), .B2(n9412), .A(n9092), .ZN(n8883) );
  NAND2_X1 U10323 ( .A1(n8884), .A2(n8883), .ZN(n8897) );
  NAND2_X1 U10324 ( .A1(n9274), .A2(n8885), .ZN(n9012) );
  NAND2_X1 U10325 ( .A1(n8992), .A2(n8886), .ZN(n8986) );
  INV_X1 U10326 ( .A(n8986), .ZN(n8891) );
  INV_X1 U10327 ( .A(n8982), .ZN(n8887) );
  AND3_X1 U10328 ( .A1(n8987), .A2(n8891), .A3(n8887), .ZN(n8888) );
  OAI21_X1 U10329 ( .B1(n8889), .B2(n8888), .A(n8997), .ZN(n8893) );
  NAND2_X1 U10330 ( .A1(n8981), .A2(n8911), .ZN(n8909) );
  INV_X1 U10331 ( .A(n8909), .ZN(n8890) );
  NAND4_X1 U10332 ( .A1(n8997), .A2(n8891), .A3(n8890), .A4(n8987), .ZN(n8892)
         );
  AND4_X1 U10333 ( .A1(n9007), .A2(n8990), .A3(n8893), .A4(n8892), .ZN(n8894)
         );
  NOR2_X1 U10334 ( .A1(n9012), .A2(n8894), .ZN(n8895) );
  OR2_X1 U10335 ( .A1(n8896), .A2(n8895), .ZN(n9093) );
  NAND4_X1 U10336 ( .A1(n8898), .A2(n9097), .A3(n8897), .A4(n9093), .ZN(n8900)
         );
  NOR2_X1 U10337 ( .A1(n9264), .A2(n9278), .ZN(n9096) );
  AOI21_X1 U10338 ( .B1(n9096), .B2(n9114), .A(n8902), .ZN(n8899) );
  NAND3_X1 U10339 ( .A1(n8900), .A2(n8899), .A3(n4411), .ZN(n8901) );
  OAI211_X1 U10340 ( .C1(n9036), .C2(n8902), .A(n9023), .B(n8901), .ZN(n9026)
         );
  INV_X1 U10341 ( .A(n9012), .ZN(n9008) );
  NOR2_X1 U10342 ( .A1(n9118), .A2(n9021), .ZN(n8904) );
  NAND2_X1 U10343 ( .A1(n9339), .A2(n8904), .ZN(n8903) );
  OAI21_X1 U10344 ( .B1(n9021), .B2(n9117), .A(n8903), .ZN(n8908) );
  NAND2_X1 U10345 ( .A1(n9118), .A2(n9021), .ZN(n9000) );
  OAI21_X1 U10346 ( .B1(n8999), .B2(n9000), .A(n9697), .ZN(n8907) );
  NAND2_X1 U10347 ( .A1(n8999), .A2(n8904), .ZN(n8905) );
  NAND2_X1 U10348 ( .A1(n9339), .A2(n8905), .ZN(n8906) );
  AOI22_X1 U10349 ( .A1(n9323), .A2(n8908), .B1(n8907), .B2(n8906), .ZN(n9005)
         );
  MUX2_X1 U10350 ( .A(n8910), .B(n8909), .S(n9021), .Z(n8984) );
  NAND2_X1 U10351 ( .A1(n8911), .A2(n8970), .ZN(n8973) );
  AND2_X1 U10352 ( .A1(n9080), .A2(n8912), .ZN(n9077) );
  AND2_X1 U10353 ( .A1(n8922), .A2(n9021), .ZN(n8914) );
  MUX2_X1 U10354 ( .A(n8914), .B(n9030), .S(n8913), .Z(n8915) );
  NAND2_X1 U10355 ( .A1(n8915), .A2(n8918), .ZN(n8917) );
  INV_X1 U10356 ( .A(n8918), .ZN(n9047) );
  AND2_X1 U10357 ( .A1(n8927), .A2(n8924), .ZN(n8921) );
  NAND4_X1 U10358 ( .A1(n8931), .A2(n9021), .A3(n8925), .A4(n8919), .ZN(n8920)
         );
  INV_X1 U10359 ( .A(n8922), .ZN(n9050) );
  AND2_X1 U10360 ( .A1(n8925), .A2(n9053), .ZN(n8928) );
  NAND4_X1 U10361 ( .A1(n8931), .A2(n8930), .A3(n9021), .A4(n8929), .ZN(n8939)
         );
  NAND4_X1 U10362 ( .A1(n8933), .A2(n8932), .A3(n9136), .A4(n9030), .ZN(n8938)
         );
  AND2_X1 U10363 ( .A1(n4758), .A2(n9030), .ZN(n8936) );
  OAI21_X1 U10364 ( .B1(n4758), .B2(n9030), .A(n8935), .ZN(n8934) );
  OAI21_X1 U10365 ( .B1(n8936), .B2(n8935), .A(n8934), .ZN(n8937) );
  NAND3_X1 U10366 ( .A1(n8939), .A2(n8938), .A3(n8937), .ZN(n8940) );
  NAND2_X1 U10367 ( .A1(n8947), .A2(n8942), .ZN(n8943) );
  NAND2_X1 U10368 ( .A1(n8949), .A2(n9556), .ZN(n9061) );
  AOI21_X1 U10369 ( .B1(n8943), .B2(n9055), .A(n9061), .ZN(n8944) );
  NAND2_X1 U10370 ( .A1(n9524), .A2(n8948), .ZN(n9065) );
  OAI21_X1 U10371 ( .B1(n8944), .B2(n9065), .A(n9063), .ZN(n8955) );
  AOI21_X1 U10372 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n8951) );
  NAND2_X1 U10373 ( .A1(n8948), .A2(n9055), .ZN(n8950) );
  OAI21_X1 U10374 ( .B1(n8951), .B2(n8950), .A(n8949), .ZN(n8953) );
  AOI21_X1 U10375 ( .B1(n8953), .B2(n9524), .A(n8952), .ZN(n8954) );
  MUX2_X1 U10376 ( .A(n8955), .B(n8954), .S(n9021), .Z(n8961) );
  NAND2_X1 U10377 ( .A1(n8961), .A2(n9067), .ZN(n8957) );
  NAND2_X1 U10378 ( .A1(n8957), .A2(n8956), .ZN(n8958) );
  NAND2_X1 U10379 ( .A1(n9076), .A2(n9129), .ZN(n8959) );
  NAND2_X1 U10380 ( .A1(n8959), .A2(n9021), .ZN(n8967) );
  NAND2_X1 U10381 ( .A1(n8967), .A2(n9495), .ZN(n8964) );
  AND2_X1 U10382 ( .A1(n8965), .A2(n8960), .ZN(n9075) );
  NAND2_X1 U10383 ( .A1(n8961), .A2(n9064), .ZN(n8962) );
  NAND3_X1 U10384 ( .A1(n8962), .A2(n9505), .A3(n9067), .ZN(n8963) );
  AND2_X1 U10385 ( .A1(n9071), .A2(n4753), .ZN(n8966) );
  AND2_X1 U10386 ( .A1(n8967), .A2(n8966), .ZN(n8968) );
  NAND2_X1 U10387 ( .A1(n8969), .A2(n9456), .ZN(n8977) );
  NAND2_X1 U10388 ( .A1(n8970), .A2(n8976), .ZN(n8971) );
  AOI21_X1 U10389 ( .B1(n9077), .B2(n8977), .A(n8971), .ZN(n8972) );
  NAND2_X1 U10390 ( .A1(n9395), .A2(n9081), .ZN(n8974) );
  NAND2_X1 U10391 ( .A1(n8974), .A2(n9021), .ZN(n8980) );
  AND2_X1 U10392 ( .A1(n8976), .A2(n8975), .ZN(n9085) );
  NAND2_X1 U10393 ( .A1(n8977), .A2(n9085), .ZN(n8978) );
  NAND4_X1 U10394 ( .A1(n8978), .A2(n9081), .A3(n9080), .A4(n9030), .ZN(n8979)
         );
  MUX2_X1 U10395 ( .A(n8982), .B(n8981), .S(n9030), .Z(n8983) );
  OAI211_X1 U10396 ( .C1(n8994), .C2(n8986), .A(n9347), .B(n8985), .ZN(n8988)
         );
  NAND2_X1 U10397 ( .A1(n8988), .A2(n8987), .ZN(n8991) );
  NAND4_X1 U10398 ( .A1(n8991), .A2(n8990), .A3(n8989), .A4(n9030), .ZN(n9004)
         );
  OAI211_X1 U10399 ( .C1(n8994), .C2(n8993), .A(n9347), .B(n8992), .ZN(n8996)
         );
  NAND2_X1 U10400 ( .A1(n8996), .A2(n8995), .ZN(n8998) );
  NAND4_X1 U10401 ( .A1(n8998), .A2(n9092), .A3(n9021), .A4(n8997), .ZN(n9003)
         );
  OAI22_X1 U10402 ( .A1(n9339), .A2(n9000), .B1(n8999), .B2(n9030), .ZN(n9001)
         );
  NAND2_X1 U10403 ( .A1(n9693), .A2(n9001), .ZN(n9002) );
  NAND4_X1 U10404 ( .A1(n9005), .A2(n9004), .A3(n9003), .A4(n9002), .ZN(n9011)
         );
  OAI21_X1 U10405 ( .B1(n9012), .B2(n9007), .A(n9006), .ZN(n9009) );
  AOI21_X1 U10406 ( .B1(n9008), .B2(n9011), .A(n9009), .ZN(n9014) );
  INV_X1 U10407 ( .A(n9009), .ZN(n9010) );
  OAI21_X1 U10408 ( .B1(n9012), .B2(n9011), .A(n9010), .ZN(n9013) );
  MUX2_X1 U10409 ( .A(n9014), .B(n9013), .S(n9030), .Z(n9018) );
  MUX2_X1 U10410 ( .A(n9016), .B(n9015), .S(n9030), .Z(n9017) );
  MUX2_X1 U10411 ( .A(n9020), .B(n9030), .S(n9264), .Z(n9019) );
  MUX2_X1 U10412 ( .A(n9021), .B(n9020), .S(n9264), .Z(n9022) );
  INV_X1 U10413 ( .A(n9023), .ZN(n9024) );
  NOR2_X1 U10414 ( .A1(n9108), .A2(n9038), .ZN(n9031) );
  OAI211_X1 U10415 ( .C1(n9030), .C2(n9044), .A(n9027), .B(n9031), .ZN(n9113)
         );
  INV_X1 U10416 ( .A(n9028), .ZN(n9029) );
  OAI21_X1 U10417 ( .B1(n9030), .B2(n4411), .A(n9029), .ZN(n9034) );
  INV_X1 U10418 ( .A(n9031), .ZN(n9032) );
  NOR3_X1 U10419 ( .A1(n9032), .A2(n9109), .A3(n9044), .ZN(n9033) );
  OAI211_X1 U10420 ( .C1(n9036), .C2(n9035), .A(n9034), .B(n9033), .ZN(n9112)
         );
  NAND2_X1 U10421 ( .A1(n9040), .A2(n9037), .ZN(n9103) );
  NAND3_X1 U10422 ( .A1(n9040), .A2(n9039), .A3(n9038), .ZN(n9102) );
  NAND2_X1 U10423 ( .A1(n9042), .A2(n9041), .ZN(n9043) );
  AOI211_X1 U10424 ( .C1(n9045), .C2(n9142), .A(n9044), .B(n9043), .ZN(n9046)
         );
  NOR3_X1 U10425 ( .A1(n9048), .A2(n9047), .A3(n9046), .ZN(n9052) );
  INV_X1 U10426 ( .A(n9049), .ZN(n9051) );
  NOR3_X1 U10427 ( .A1(n9052), .A2(n9051), .A3(n9050), .ZN(n9054) );
  OAI21_X1 U10428 ( .B1(n9054), .B2(n4428), .A(n9053), .ZN(n9059) );
  INV_X1 U10429 ( .A(n9055), .ZN(n9058) );
  INV_X1 U10430 ( .A(n9056), .ZN(n9057) );
  AOI211_X1 U10431 ( .C1(n9060), .C2(n9059), .A(n9058), .B(n9057), .ZN(n9062)
         );
  NOR2_X1 U10432 ( .A1(n9062), .A2(n9061), .ZN(n9066) );
  OAI211_X1 U10433 ( .C1(n9066), .C2(n9065), .A(n9064), .B(n9063), .ZN(n9069)
         );
  NAND3_X1 U10434 ( .A1(n9069), .A2(n9068), .A3(n9067), .ZN(n9074) );
  INV_X1 U10435 ( .A(n9070), .ZN(n9073) );
  INV_X1 U10436 ( .A(n9071), .ZN(n9072) );
  AOI211_X1 U10437 ( .C1(n9075), .C2(n9074), .A(n9073), .B(n9072), .ZN(n9079)
         );
  INV_X1 U10438 ( .A(n9076), .ZN(n9078) );
  OAI21_X1 U10439 ( .B1(n9079), .B2(n9078), .A(n9077), .ZN(n9084) );
  INV_X1 U10440 ( .A(n9080), .ZN(n9083) );
  INV_X1 U10441 ( .A(n9081), .ZN(n9082) );
  AOI211_X1 U10442 ( .C1(n9085), .C2(n9084), .A(n9083), .B(n9082), .ZN(n9088)
         );
  INV_X1 U10443 ( .A(n9086), .ZN(n9087) );
  OAI21_X1 U10444 ( .B1(n9089), .B2(n9088), .A(n9087), .ZN(n9091) );
  AOI21_X1 U10445 ( .B1(n9092), .B2(n9091), .A(n9090), .ZN(n9095) );
  INV_X1 U10446 ( .A(n9093), .ZN(n9094) );
  NOR2_X1 U10447 ( .A1(n9095), .A2(n9094), .ZN(n9098) );
  AOI21_X1 U10448 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(n9100) );
  AOI21_X1 U10449 ( .B1(n9100), .B2(n4411), .A(n9099), .ZN(n9101) );
  MUX2_X1 U10450 ( .A(n9103), .B(n9102), .S(n9101), .Z(n9111) );
  NAND3_X1 U10451 ( .A1(n9106), .A2(n9105), .A3(n9104), .ZN(n9107) );
  OAI211_X1 U10452 ( .C1(n9109), .C2(n9108), .A(n9107), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9110) );
  NAND4_X1 U10453 ( .A1(n9113), .A2(n9112), .A3(n9111), .A4(n9110), .ZN(
        P1_U3242) );
  MUX2_X1 U10454 ( .A(n9114), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9128), .Z(
        P1_U3585) );
  MUX2_X1 U10455 ( .A(n9115), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9128), .Z(
        P1_U3584) );
  INV_X1 U10456 ( .A(n9280), .ZN(n9268) );
  MUX2_X1 U10457 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9268), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10458 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9116), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10459 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9117), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9118), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10461 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9119), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10462 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9120), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10463 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9121), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9122), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10465 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9123), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10466 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9124), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10467 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9125), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10468 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9126), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10469 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9127), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10470 ( .A(n9129), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9128), .Z(
        P1_U3569) );
  MUX2_X1 U10471 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9130), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10472 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9131), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10473 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9132), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10474 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9133), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10475 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9134), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10476 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9135), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10477 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n4758), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10478 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9136), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10479 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9137), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10480 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9138), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10481 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9139), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10482 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9140), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9141), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10484 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9142), .S(P1_U3973), .Z(
        P1_U3555) );
  NAND2_X1 U10485 ( .A1(n9781), .A2(n9143), .ZN(n9156) );
  OAI211_X1 U10486 ( .C1(n9146), .C2(n9145), .A(n9785), .B(n9144), .ZN(n9155)
         );
  AOI22_X1 U10487 ( .A1(n9230), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9154) );
  MUX2_X1 U10488 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n5894), .S(n9147), .Z(n9148)
         );
  OAI21_X1 U10489 ( .B1(n9150), .B2(n9149), .A(n9148), .ZN(n9151) );
  NAND3_X1 U10490 ( .A1(n9779), .A2(n9152), .A3(n9151), .ZN(n9153) );
  NAND4_X1 U10491 ( .A1(n9156), .A2(n9155), .A3(n9154), .A4(n9153), .ZN(
        P1_U3244) );
  AND2_X1 U10492 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9159) );
  NOR2_X1 U10493 ( .A1(n9767), .A2(n9157), .ZN(n9158) );
  AOI211_X1 U10494 ( .C1(n9230), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9159), .B(
        n9158), .ZN(n9167) );
  OAI211_X1 U10495 ( .C1(n9162), .C2(n9161), .A(n9785), .B(n9160), .ZN(n9166)
         );
  OAI211_X1 U10496 ( .C1(n9164), .C2(n9163), .A(n9779), .B(n9179), .ZN(n9165)
         );
  NAND3_X1 U10497 ( .A1(n9167), .A2(n9166), .A3(n9165), .ZN(P1_U3246) );
  INV_X1 U10498 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9169) );
  OAI21_X1 U10499 ( .B1(n9788), .B2(n9169), .A(n9168), .ZN(n9170) );
  AOI21_X1 U10500 ( .B1(n9781), .B2(n9171), .A(n9170), .ZN(n9183) );
  OAI211_X1 U10501 ( .C1(n9174), .C2(n9173), .A(n9785), .B(n9172), .ZN(n9182)
         );
  INV_X1 U10502 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9176) );
  MUX2_X1 U10503 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9176), .S(n9175), .Z(n9177)
         );
  NAND3_X1 U10504 ( .A1(n9179), .A2(n9178), .A3(n9177), .ZN(n9180) );
  NAND3_X1 U10505 ( .A1(n9779), .A2(n9194), .A3(n9180), .ZN(n9181) );
  NAND4_X1 U10506 ( .A1(n9184), .A2(n9183), .A3(n9182), .A4(n9181), .ZN(
        P1_U3247) );
  INV_X1 U10507 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9186) );
  OAI21_X1 U10508 ( .B1(n9788), .B2(n9186), .A(n9185), .ZN(n9187) );
  AOI21_X1 U10509 ( .B1(n9781), .B2(n9191), .A(n9187), .ZN(n9198) );
  OAI211_X1 U10510 ( .C1(n9190), .C2(n9189), .A(n9785), .B(n9188), .ZN(n9197)
         );
  MUX2_X1 U10511 ( .A(n5903), .B(P1_REG1_REG_5__SCAN_IN), .S(n9191), .Z(n9192)
         );
  NAND3_X1 U10512 ( .A1(n9194), .A2(n9193), .A3(n9192), .ZN(n9195) );
  NAND3_X1 U10513 ( .A1(n9779), .A2(n9207), .A3(n9195), .ZN(n9196) );
  NAND3_X1 U10514 ( .A1(n9198), .A2(n9197), .A3(n9196), .ZN(P1_U3248) );
  NAND2_X1 U10515 ( .A1(n9781), .A2(n9204), .ZN(n9212) );
  OAI211_X1 U10516 ( .C1(n9201), .C2(n9200), .A(n9785), .B(n9199), .ZN(n9211)
         );
  AND2_X1 U10517 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9203) );
  AOI21_X1 U10518 ( .B1(n9230), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9203), .ZN(
        n9210) );
  MUX2_X1 U10519 ( .A(n5906), .B(P1_REG1_REG_6__SCAN_IN), .S(n9204), .Z(n9205)
         );
  NAND3_X1 U10520 ( .A1(n9207), .A2(n9206), .A3(n9205), .ZN(n9208) );
  NAND3_X1 U10521 ( .A1(n9779), .A2(n9222), .A3(n9208), .ZN(n9209) );
  NAND4_X1 U10522 ( .A1(n9212), .A2(n9211), .A3(n9210), .A4(n9209), .ZN(
        P1_U3249) );
  INV_X1 U10523 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9214) );
  OAI21_X1 U10524 ( .B1(n9788), .B2(n9214), .A(n9213), .ZN(n9215) );
  AOI21_X1 U10525 ( .B1(n9781), .B2(n9219), .A(n9215), .ZN(n9226) );
  OAI211_X1 U10526 ( .C1(n9218), .C2(n9217), .A(n9785), .B(n9216), .ZN(n9225)
         );
  MUX2_X1 U10527 ( .A(n5909), .B(P1_REG1_REG_7__SCAN_IN), .S(n9219), .Z(n9220)
         );
  NAND3_X1 U10528 ( .A1(n9222), .A2(n9221), .A3(n9220), .ZN(n9223) );
  NAND3_X1 U10529 ( .A1(n9779), .A2(n9234), .A3(n9223), .ZN(n9224) );
  NAND3_X1 U10530 ( .A1(n9226), .A2(n9225), .A3(n9224), .ZN(P1_U3250) );
  NAND2_X1 U10531 ( .A1(n9781), .A2(n9231), .ZN(n9240) );
  OAI211_X1 U10532 ( .C1(n9228), .C2(n9227), .A(n9785), .B(n9756), .ZN(n9239)
         );
  AOI21_X1 U10533 ( .B1(n9230), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9229), .ZN(
        n9238) );
  MUX2_X1 U10534 ( .A(n5912), .B(P1_REG1_REG_8__SCAN_IN), .S(n9231), .Z(n9232)
         );
  NAND3_X1 U10535 ( .A1(n9234), .A2(n9233), .A3(n9232), .ZN(n9235) );
  NAND3_X1 U10536 ( .A1(n9779), .A2(n9236), .A3(n9235), .ZN(n9237) );
  NAND4_X1 U10537 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), .ZN(
        P1_U3251) );
  AOI211_X1 U10538 ( .C1(n9244), .C2(n9243), .A(n9242), .B(n9241), .ZN(n9245)
         );
  INV_X1 U10539 ( .A(n9245), .ZN(n9254) );
  OAI21_X1 U10540 ( .B1(n9788), .B2(n7063), .A(n9246), .ZN(n9247) );
  AOI21_X1 U10541 ( .B1(n9781), .B2(n9248), .A(n9247), .ZN(n9253) );
  OAI211_X1 U10542 ( .C1(n9251), .C2(n9250), .A(n9779), .B(n9249), .ZN(n9252)
         );
  NAND3_X1 U10543 ( .A1(n9254), .A2(n9253), .A3(n9252), .ZN(P1_U3256) );
  NAND2_X1 U10544 ( .A1(n9684), .A2(n9282), .ZN(n9255) );
  XNOR2_X1 U10545 ( .A(n9680), .B(n9255), .ZN(n9578) );
  NAND2_X1 U10546 ( .A1(n9578), .A2(n9503), .ZN(n9263) );
  INV_X1 U10547 ( .A(P1_B_REG_SCAN_IN), .ZN(n9256) );
  OR2_X1 U10548 ( .A1(n9257), .A2(n9256), .ZN(n9258) );
  NAND2_X1 U10549 ( .A1(n9259), .A2(n9258), .ZN(n9279) );
  NOR2_X1 U10550 ( .A1(n9260), .A2(n9279), .ZN(n9580) );
  INV_X1 U10551 ( .A(n9580), .ZN(n9261) );
  NOR2_X1 U10552 ( .A1(n9261), .A2(n9573), .ZN(n9265) );
  AOI21_X1 U10553 ( .B1(n9573), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9265), .ZN(
        n9262) );
  OAI211_X1 U10554 ( .C1(n9680), .C2(n9795), .A(n9263), .B(n9262), .ZN(
        P1_U3263) );
  XNOR2_X1 U10555 ( .A(n9264), .B(n9282), .ZN(n9581) );
  NAND2_X1 U10556 ( .A1(n9581), .A2(n9503), .ZN(n9267) );
  AOI21_X1 U10557 ( .B1(n9573), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9265), .ZN(
        n9266) );
  OAI211_X1 U10558 ( .C1(n9684), .C2(n9795), .A(n9267), .B(n9266), .ZN(
        P1_U3264) );
  NAND2_X1 U10559 ( .A1(n9269), .A2(n9268), .ZN(n9270) );
  XNOR2_X1 U10560 ( .A(n9273), .B(n9272), .ZN(n9584) );
  INV_X1 U10561 ( .A(n9584), .ZN(n9290) );
  INV_X1 U10562 ( .A(n9587), .ZN(n9287) );
  AOI211_X1 U10563 ( .C1(n9587), .C2(n9283), .A(n9570), .B(n9282), .ZN(n9586)
         );
  NAND2_X1 U10564 ( .A1(n9586), .A2(n9790), .ZN(n9286) );
  AOI22_X1 U10565 ( .A1(n9573), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9284), .B2(
        n9792), .ZN(n9285) );
  OAI211_X1 U10566 ( .C1(n9287), .C2(n9795), .A(n9286), .B(n9285), .ZN(n9288)
         );
  AOI21_X1 U10567 ( .B1(n9585), .B2(n6473), .A(n9288), .ZN(n9289) );
  OAI21_X1 U10568 ( .B1(n9290), .B2(n9551), .A(n9289), .ZN(P1_U3356) );
  NAND2_X1 U10569 ( .A1(n9291), .A2(n9799), .ZN(n9299) );
  INV_X1 U10570 ( .A(n9292), .ZN(n9297) );
  AOI22_X1 U10571 ( .A1(n9573), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9792), .B2(
        n9293), .ZN(n9294) );
  OAI21_X1 U10572 ( .B1(n9295), .B2(n9795), .A(n9294), .ZN(n9296) );
  AOI21_X1 U10573 ( .B1(n9297), .B2(n9790), .A(n9296), .ZN(n9298) );
  OAI211_X1 U10574 ( .C1(n9300), .C2(n9802), .A(n9299), .B(n9298), .ZN(
        P1_U3265) );
  XNOR2_X1 U10575 ( .A(n9303), .B(n9302), .ZN(n9305) );
  INV_X1 U10576 ( .A(n9590), .ZN(n9313) );
  INV_X1 U10577 ( .A(n9593), .ZN(n9689) );
  INV_X1 U10578 ( .A(n9306), .ZN(n9322) );
  INV_X1 U10579 ( .A(n9307), .ZN(n9308) );
  OAI211_X1 U10580 ( .C1(n9689), .C2(n9322), .A(n9308), .B(n9650), .ZN(n9589)
         );
  NOR2_X1 U10581 ( .A1(n9589), .A2(n9532), .ZN(n9312) );
  AOI22_X1 U10582 ( .A1(n9309), .A2(n9792), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9802), .ZN(n9310) );
  OAI21_X1 U10583 ( .B1(n9689), .B2(n9795), .A(n9310), .ZN(n9311) );
  AOI211_X1 U10584 ( .C1(n9313), .C2(n6473), .A(n9312), .B(n9311), .ZN(n9314)
         );
  OAI21_X1 U10585 ( .B1(n9591), .B2(n9551), .A(n9314), .ZN(P1_U3266) );
  XNOR2_X1 U10586 ( .A(n9315), .B(n9321), .ZN(n9316) );
  NAND2_X1 U10587 ( .A1(n9316), .A2(n9526), .ZN(n9319) );
  INV_X1 U10588 ( .A(n9317), .ZN(n9318) );
  NAND2_X1 U10589 ( .A1(n9319), .A2(n9318), .ZN(n9595) );
  INV_X1 U10590 ( .A(n9595), .ZN(n9330) );
  XNOR2_X1 U10591 ( .A(n9320), .B(n9321), .ZN(n9597) );
  NAND2_X1 U10592 ( .A1(n9597), .A2(n9799), .ZN(n9329) );
  AOI211_X1 U10593 ( .C1(n9323), .C2(n9337), .A(n9570), .B(n9322), .ZN(n9596)
         );
  NOR2_X1 U10594 ( .A1(n9693), .A2(n9795), .ZN(n9327) );
  OAI22_X1 U10595 ( .A1(n9325), .A2(n9433), .B1(n9324), .B2(n6473), .ZN(n9326)
         );
  AOI211_X1 U10596 ( .C1(n9596), .C2(n9790), .A(n9327), .B(n9326), .ZN(n9328)
         );
  OAI211_X1 U10597 ( .C1(n9802), .C2(n9330), .A(n9329), .B(n9328), .ZN(
        P1_U3267) );
  XNOR2_X1 U10598 ( .A(n9331), .B(n9333), .ZN(n9602) );
  INV_X1 U10599 ( .A(n9602), .ZN(n9346) );
  OAI211_X1 U10600 ( .C1(n9334), .C2(n9333), .A(n9332), .B(n9526), .ZN(n9336)
         );
  NAND2_X1 U10601 ( .A1(n9336), .A2(n9335), .ZN(n9600) );
  INV_X1 U10602 ( .A(n9337), .ZN(n9338) );
  AOI211_X1 U10603 ( .C1(n9339), .C2(n9355), .A(n9570), .B(n9338), .ZN(n9601)
         );
  NAND2_X1 U10604 ( .A1(n9601), .A2(n9790), .ZN(n9343) );
  INV_X1 U10605 ( .A(n9340), .ZN(n9341) );
  AOI22_X1 U10606 ( .A1(n9341), .A2(n9792), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9573), .ZN(n9342) );
  OAI211_X1 U10607 ( .C1(n9697), .C2(n9795), .A(n9343), .B(n9342), .ZN(n9344)
         );
  AOI21_X1 U10608 ( .B1(n6473), .B2(n9600), .A(n9344), .ZN(n9345) );
  OAI21_X1 U10609 ( .B1(n9346), .B2(n9551), .A(n9345), .ZN(P1_U3268) );
  XNOR2_X1 U10610 ( .A(n9348), .B(n9347), .ZN(n9607) );
  INV_X1 U10611 ( .A(n9607), .ZN(n9364) );
  NAND2_X1 U10612 ( .A1(n9350), .A2(n9349), .ZN(n9351) );
  NAND3_X1 U10613 ( .A1(n9352), .A2(n9526), .A3(n9351), .ZN(n9354) );
  NAND2_X1 U10614 ( .A1(n9354), .A2(n9353), .ZN(n9605) );
  INV_X1 U10615 ( .A(n9371), .ZN(n9357) );
  INV_X1 U10616 ( .A(n9355), .ZN(n9356) );
  AOI211_X1 U10617 ( .C1(n9358), .C2(n9357), .A(n9570), .B(n9356), .ZN(n9606)
         );
  NAND2_X1 U10618 ( .A1(n9606), .A2(n9790), .ZN(n9361) );
  AOI22_X1 U10619 ( .A1(n9359), .A2(n9792), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9573), .ZN(n9360) );
  OAI211_X1 U10620 ( .C1(n9701), .C2(n9795), .A(n9361), .B(n9360), .ZN(n9362)
         );
  AOI21_X1 U10621 ( .B1(n6473), .B2(n9605), .A(n9362), .ZN(n9363) );
  OAI21_X1 U10622 ( .B1(n9364), .B2(n9551), .A(n9363), .ZN(P1_U3269) );
  XOR2_X1 U10623 ( .A(n9367), .B(n9365), .Z(n9611) );
  INV_X1 U10624 ( .A(n9611), .ZN(n9378) );
  XOR2_X1 U10625 ( .A(n9367), .B(n9366), .Z(n9370) );
  INV_X1 U10626 ( .A(n9368), .ZN(n9369) );
  OAI21_X1 U10627 ( .B1(n9370), .B2(n9565), .A(n9369), .ZN(n9609) );
  AOI211_X1 U10628 ( .C1(n9372), .C2(n9385), .A(n9570), .B(n9371), .ZN(n9610)
         );
  NAND2_X1 U10629 ( .A1(n9610), .A2(n9790), .ZN(n9375) );
  AOI22_X1 U10630 ( .A1(n9373), .A2(n9792), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9573), .ZN(n9374) );
  OAI211_X1 U10631 ( .C1(n9705), .C2(n9795), .A(n9375), .B(n9374), .ZN(n9376)
         );
  AOI21_X1 U10632 ( .B1(n6473), .B2(n9609), .A(n9376), .ZN(n9377) );
  OAI21_X1 U10633 ( .B1(n9378), .B2(n9551), .A(n9377), .ZN(P1_U3270) );
  XNOR2_X1 U10634 ( .A(n9379), .B(n9381), .ZN(n9615) );
  INV_X1 U10635 ( .A(n9615), .ZN(n9393) );
  OAI211_X1 U10636 ( .C1(n9382), .C2(n9381), .A(n9380), .B(n9526), .ZN(n9384)
         );
  NAND2_X1 U10637 ( .A1(n9384), .A2(n9383), .ZN(n9613) );
  INV_X1 U10638 ( .A(n9385), .ZN(n9386) );
  AOI211_X1 U10639 ( .C1(n9387), .C2(n9403), .A(n9570), .B(n9386), .ZN(n9614)
         );
  NAND2_X1 U10640 ( .A1(n9614), .A2(n9790), .ZN(n9390) );
  AOI22_X1 U10641 ( .A1(n9388), .A2(n9792), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9573), .ZN(n9389) );
  OAI211_X1 U10642 ( .C1(n4872), .C2(n9795), .A(n9390), .B(n9389), .ZN(n9391)
         );
  AOI21_X1 U10643 ( .B1(n6473), .B2(n9613), .A(n9391), .ZN(n9392) );
  OAI21_X1 U10644 ( .B1(n9393), .B2(n9551), .A(n9392), .ZN(P1_U3271) );
  XNOR2_X1 U10645 ( .A(n9394), .B(n9397), .ZN(n9620) );
  INV_X1 U10646 ( .A(n9620), .ZN(n9410) );
  NAND2_X1 U10647 ( .A1(n9396), .A2(n9395), .ZN(n9398) );
  XNOR2_X1 U10648 ( .A(n9398), .B(n9397), .ZN(n9399) );
  NAND2_X1 U10649 ( .A1(n9399), .A2(n9526), .ZN(n9402) );
  INV_X1 U10650 ( .A(n9400), .ZN(n9401) );
  NAND2_X1 U10651 ( .A1(n9402), .A2(n9401), .ZN(n9618) );
  AOI211_X1 U10652 ( .C1(n9404), .C2(n9415), .A(n9570), .B(n4873), .ZN(n9619)
         );
  NAND2_X1 U10653 ( .A1(n9619), .A2(n9790), .ZN(n9407) );
  AOI22_X1 U10654 ( .A1(n9405), .A2(n9792), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9573), .ZN(n9406) );
  OAI211_X1 U10655 ( .C1(n9712), .C2(n9795), .A(n9407), .B(n9406), .ZN(n9408)
         );
  AOI21_X1 U10656 ( .B1(n6473), .B2(n9618), .A(n9408), .ZN(n9409) );
  OAI21_X1 U10657 ( .B1(n9410), .B2(n9551), .A(n9409), .ZN(P1_U3272) );
  XOR2_X1 U10658 ( .A(n9411), .B(n4408), .Z(n9627) );
  XNOR2_X1 U10659 ( .A(n9412), .B(n9411), .ZN(n9414) );
  OAI21_X1 U10660 ( .B1(n9414), .B2(n9565), .A(n9413), .ZN(n9623) );
  INV_X1 U10661 ( .A(n9431), .ZN(n9417) );
  INV_X1 U10662 ( .A(n9415), .ZN(n9416) );
  AOI211_X1 U10663 ( .C1(n9625), .C2(n9417), .A(n9570), .B(n9416), .ZN(n9624)
         );
  NAND2_X1 U10664 ( .A1(n9624), .A2(n9790), .ZN(n9420) );
  AOI22_X1 U10665 ( .A1(n9418), .A2(n9792), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9573), .ZN(n9419) );
  OAI211_X1 U10666 ( .C1(n9421), .C2(n9795), .A(n9420), .B(n9419), .ZN(n9422)
         );
  AOI21_X1 U10667 ( .B1(n6473), .B2(n9623), .A(n9422), .ZN(n9423) );
  OAI21_X1 U10668 ( .B1(n9627), .B2(n9551), .A(n9423), .ZN(P1_U3273) );
  XNOR2_X1 U10669 ( .A(n9424), .B(n9429), .ZN(n9425) );
  NAND2_X1 U10670 ( .A1(n9425), .A2(n9526), .ZN(n9428) );
  INV_X1 U10671 ( .A(n9426), .ZN(n9427) );
  NAND2_X1 U10672 ( .A1(n9428), .A2(n9427), .ZN(n9628) );
  INV_X1 U10673 ( .A(n9628), .ZN(n9440) );
  XNOR2_X1 U10674 ( .A(n9430), .B(n9429), .ZN(n9630) );
  NAND2_X1 U10675 ( .A1(n9630), .A2(n9799), .ZN(n9439) );
  AOI211_X1 U10676 ( .C1(n9432), .C2(n9442), .A(n9570), .B(n9431), .ZN(n9629)
         );
  NOR2_X1 U10677 ( .A1(n9717), .A2(n9795), .ZN(n9437) );
  OAI22_X1 U10678 ( .A1(n6473), .A2(n9435), .B1(n9434), .B2(n9433), .ZN(n9436)
         );
  AOI211_X1 U10679 ( .C1(n9629), .C2(n9790), .A(n9437), .B(n9436), .ZN(n9438)
         );
  OAI211_X1 U10680 ( .C1(n9802), .C2(n9440), .A(n9439), .B(n9438), .ZN(
        P1_U3274) );
  XOR2_X1 U10681 ( .A(n9441), .B(n9449), .Z(n9637) );
  INV_X1 U10682 ( .A(n9442), .ZN(n9443) );
  AOI211_X1 U10683 ( .C1(n9634), .C2(n9464), .A(n9570), .B(n9443), .ZN(n9633)
         );
  AOI22_X1 U10684 ( .A1(n9573), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9444), .B2(
        n9792), .ZN(n9445) );
  OAI21_X1 U10685 ( .B1(n9446), .B2(n9795), .A(n9445), .ZN(n9454) );
  OAI21_X1 U10686 ( .B1(n9449), .B2(n9448), .A(n9447), .ZN(n9452) );
  INV_X1 U10687 ( .A(n9450), .ZN(n9451) );
  AOI21_X1 U10688 ( .B1(n9452), .B2(n9526), .A(n9451), .ZN(n9636) );
  NOR2_X1 U10689 ( .A1(n9636), .A2(n9802), .ZN(n9453) );
  AOI211_X1 U10690 ( .C1(n9633), .C2(n9790), .A(n9454), .B(n9453), .ZN(n9455)
         );
  OAI21_X1 U10691 ( .B1(n9637), .B2(n9551), .A(n9455), .ZN(P1_U3275) );
  XNOR2_X1 U10692 ( .A(n9457), .B(n9456), .ZN(n9640) );
  INV_X1 U10693 ( .A(n9640), .ZN(n9472) );
  NAND2_X1 U10694 ( .A1(n9459), .A2(n9458), .ZN(n9461) );
  NAND3_X1 U10695 ( .A1(n9461), .A2(n9460), .A3(n9526), .ZN(n9463) );
  NAND2_X1 U10696 ( .A1(n9463), .A2(n9462), .ZN(n9638) );
  INV_X1 U10697 ( .A(n9464), .ZN(n9465) );
  AOI211_X1 U10698 ( .C1(n9466), .C2(n9476), .A(n9570), .B(n9465), .ZN(n9639)
         );
  NAND2_X1 U10699 ( .A1(n9639), .A2(n9790), .ZN(n9469) );
  AOI22_X1 U10700 ( .A1(n9573), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9467), .B2(
        n9792), .ZN(n9468) );
  OAI211_X1 U10701 ( .C1(n4875), .C2(n9795), .A(n9469), .B(n9468), .ZN(n9470)
         );
  AOI21_X1 U10702 ( .B1(n6473), .B2(n9638), .A(n9470), .ZN(n9471) );
  OAI21_X1 U10703 ( .B1(n9472), .B2(n9551), .A(n9471), .ZN(P1_U3276) );
  OAI21_X1 U10704 ( .B1(n9475), .B2(n9474), .A(n9473), .ZN(n9648) );
  AOI211_X1 U10705 ( .C1(n9645), .C2(n9490), .A(n9570), .B(n4876), .ZN(n9644)
         );
  AOI22_X1 U10706 ( .A1(n9573), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9477), .B2(
        n9792), .ZN(n9478) );
  OAI21_X1 U10707 ( .B1(n9479), .B2(n9795), .A(n9478), .ZN(n9486) );
  OAI21_X1 U10708 ( .B1(n9482), .B2(n9481), .A(n9480), .ZN(n9484) );
  AOI21_X1 U10709 ( .B1(n9484), .B2(n9526), .A(n9483), .ZN(n9647) );
  NOR2_X1 U10710 ( .A1(n9647), .A2(n9802), .ZN(n9485) );
  AOI211_X1 U10711 ( .C1(n9644), .C2(n9790), .A(n9486), .B(n9485), .ZN(n9487)
         );
  OAI21_X1 U10712 ( .B1(n9648), .B2(n9551), .A(n9487), .ZN(P1_U3277) );
  XNOR2_X1 U10713 ( .A(n9488), .B(n9489), .ZN(n9654) );
  INV_X1 U10714 ( .A(n9513), .ZN(n9492) );
  INV_X1 U10715 ( .A(n9490), .ZN(n9491) );
  AOI21_X1 U10716 ( .B1(n9649), .B2(n9492), .A(n9491), .ZN(n9651) );
  AOI22_X1 U10717 ( .A1(n9802), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9493), .B2(
        n9792), .ZN(n9494) );
  OAI21_X1 U10718 ( .B1(n9495), .B2(n9795), .A(n9494), .ZN(n9502) );
  OAI21_X1 U10719 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9500) );
  AOI21_X1 U10720 ( .B1(n9500), .B2(n9526), .A(n9499), .ZN(n9653) );
  NOR2_X1 U10721 ( .A1(n9653), .A2(n9573), .ZN(n9501) );
  AOI211_X1 U10722 ( .C1(n9651), .C2(n9503), .A(n9502), .B(n9501), .ZN(n9504)
         );
  OAI21_X1 U10723 ( .B1(n9654), .B2(n9551), .A(n9504), .ZN(P1_U3278) );
  XNOR2_X1 U10724 ( .A(n9506), .B(n9505), .ZN(n9661) );
  OAI21_X1 U10725 ( .B1(n9527), .B2(n9508), .A(n9507), .ZN(n9510) );
  NAND3_X1 U10726 ( .A1(n9510), .A2(n9509), .A3(n9526), .ZN(n9512) );
  NAND2_X1 U10727 ( .A1(n9512), .A2(n9511), .ZN(n9656) );
  AOI211_X1 U10728 ( .C1(n9657), .C2(n9531), .A(n9570), .B(n9513), .ZN(n9655)
         );
  NAND2_X1 U10729 ( .A1(n9655), .A2(n9790), .ZN(n9516) );
  AOI22_X1 U10730 ( .A1(n9573), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9514), .B2(
        n9792), .ZN(n9515) );
  OAI211_X1 U10731 ( .C1(n9517), .C2(n9795), .A(n9516), .B(n9515), .ZN(n9518)
         );
  AOI21_X1 U10732 ( .B1(n6473), .B2(n9656), .A(n9518), .ZN(n9519) );
  OAI21_X1 U10733 ( .B1(n9661), .B2(n9551), .A(n9519), .ZN(P1_U3279) );
  OAI21_X1 U10734 ( .B1(n9522), .B2(n9521), .A(n9520), .ZN(n9665) );
  INV_X1 U10735 ( .A(n9665), .ZN(n9538) );
  AOI21_X1 U10736 ( .B1(n9525), .B2(n9524), .A(n9523), .ZN(n9528) );
  OAI21_X1 U10737 ( .B1(n9528), .B2(n9527), .A(n9526), .ZN(n9530) );
  NAND2_X1 U10738 ( .A1(n9530), .A2(n9529), .ZN(n9664) );
  OAI211_X1 U10739 ( .C1(n4870), .C2(n4871), .A(n9650), .B(n9531), .ZN(n9662)
         );
  NOR2_X1 U10740 ( .A1(n9662), .A2(n9532), .ZN(n9536) );
  AOI22_X1 U10741 ( .A1(n9573), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9533), .B2(
        n9792), .ZN(n9534) );
  OAI21_X1 U10742 ( .B1(n4870), .B2(n9795), .A(n9534), .ZN(n9535) );
  AOI211_X1 U10743 ( .C1(n9664), .C2(n6473), .A(n9536), .B(n9535), .ZN(n9537)
         );
  OAI21_X1 U10744 ( .B1(n9538), .B2(n9551), .A(n9537), .ZN(P1_U3280) );
  OAI21_X1 U10745 ( .B1(n9541), .B2(n9540), .A(n9539), .ZN(n9669) );
  INV_X1 U10746 ( .A(n9669), .ZN(n9552) );
  XNOR2_X1 U10747 ( .A(n9543), .B(n9542), .ZN(n9545) );
  OAI21_X1 U10748 ( .B1(n9545), .B2(n9565), .A(n9544), .ZN(n9667) );
  AOI211_X1 U10749 ( .C1(n9729), .C2(n9568), .A(n9570), .B(n4871), .ZN(n9668)
         );
  NAND2_X1 U10750 ( .A1(n9668), .A2(n9790), .ZN(n9548) );
  AOI22_X1 U10751 ( .A1(n9573), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9546), .B2(
        n9792), .ZN(n9547) );
  OAI211_X1 U10752 ( .C1(n7545), .C2(n9795), .A(n9548), .B(n9547), .ZN(n9549)
         );
  AOI21_X1 U10753 ( .B1(n6473), .B2(n9667), .A(n9549), .ZN(n9550) );
  OAI21_X1 U10754 ( .B1(n9552), .B2(n9551), .A(n9550), .ZN(P1_U3281) );
  INV_X1 U10755 ( .A(n9553), .ZN(n9566) );
  OAI21_X1 U10756 ( .B1(n9555), .B2(n9558), .A(n9554), .ZN(n9674) );
  NAND2_X1 U10757 ( .A1(n9557), .A2(n9556), .ZN(n9559) );
  XNOR2_X1 U10758 ( .A(n9559), .B(n9558), .ZN(n9564) );
  INV_X1 U10759 ( .A(n9560), .ZN(n9561) );
  NAND2_X1 U10760 ( .A1(n9674), .A2(n9561), .ZN(n9563) );
  OAI211_X1 U10761 ( .C1(n9565), .C2(n9564), .A(n9563), .B(n9562), .ZN(n9672)
         );
  AOI21_X1 U10762 ( .B1(n9566), .B2(n9674), .A(n9672), .ZN(n9577) );
  INV_X1 U10763 ( .A(n9567), .ZN(n9571) );
  INV_X1 U10764 ( .A(n9568), .ZN(n9569) );
  AOI211_X1 U10765 ( .C1(n4451), .C2(n9571), .A(n9570), .B(n9569), .ZN(n9673)
         );
  AOI22_X1 U10766 ( .A1(n9573), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9572), .B2(
        n9792), .ZN(n9574) );
  OAI21_X1 U10767 ( .B1(n7531), .B2(n9795), .A(n9574), .ZN(n9575) );
  AOI21_X1 U10768 ( .B1(n9673), .B2(n9790), .A(n9575), .ZN(n9576) );
  OAI21_X1 U10769 ( .B1(n9577), .B2(n9802), .A(n9576), .ZN(P1_U3282) );
  INV_X1 U10770 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9579) );
  AOI21_X1 U10771 ( .B1(n9578), .B2(n9650), .A(n9580), .ZN(n9678) );
  INV_X1 U10772 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9582) );
  AOI21_X1 U10773 ( .B1(n9581), .B2(n9650), .A(n9580), .ZN(n9681) );
  OAI21_X1 U10774 ( .B1(n9684), .B2(n9643), .A(n9583), .ZN(P1_U3552) );
  NAND2_X1 U10775 ( .A1(n9584), .A2(n9809), .ZN(n9588) );
  MUX2_X1 U10776 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9685), .S(n9816), .Z(
        P1_U3551) );
  INV_X1 U10777 ( .A(n9809), .ZN(n9660) );
  OAI211_X1 U10778 ( .C1(n9591), .C2(n9660), .A(n9590), .B(n9589), .ZN(n9686)
         );
  AOI21_X1 U10779 ( .B1(n9676), .B2(n9593), .A(n9592), .ZN(n9594) );
  INV_X1 U10780 ( .A(n9594), .ZN(P1_U3549) );
  INV_X1 U10781 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9598) );
  AOI211_X1 U10782 ( .C1(n9597), .C2(n9809), .A(n9596), .B(n9595), .ZN(n9690)
         );
  MUX2_X1 U10783 ( .A(n9598), .B(n9690), .S(n9816), .Z(n9599) );
  OAI21_X1 U10784 ( .B1(n9693), .B2(n9643), .A(n9599), .ZN(P1_U3548) );
  AOI211_X1 U10785 ( .C1(n9602), .C2(n9809), .A(n9601), .B(n9600), .ZN(n9694)
         );
  MUX2_X1 U10786 ( .A(n9603), .B(n9694), .S(n9816), .Z(n9604) );
  OAI21_X1 U10787 ( .B1(n9697), .B2(n9643), .A(n9604), .ZN(P1_U3547) );
  AOI211_X1 U10788 ( .C1(n9607), .C2(n9809), .A(n9606), .B(n9605), .ZN(n9698)
         );
  MUX2_X1 U10789 ( .A(n10060), .B(n9698), .S(n9816), .Z(n9608) );
  OAI21_X1 U10790 ( .B1(n9701), .B2(n9643), .A(n9608), .ZN(P1_U3546) );
  AOI211_X1 U10791 ( .C1(n9611), .C2(n9809), .A(n9610), .B(n9609), .ZN(n9702)
         );
  MUX2_X1 U10792 ( .A(n10090), .B(n9702), .S(n9816), .Z(n9612) );
  OAI21_X1 U10793 ( .B1(n9705), .B2(n9643), .A(n9612), .ZN(P1_U3545) );
  INV_X1 U10794 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9616) );
  AOI211_X1 U10795 ( .C1(n9615), .C2(n9809), .A(n9614), .B(n9613), .ZN(n9706)
         );
  MUX2_X1 U10796 ( .A(n9616), .B(n9706), .S(n9816), .Z(n9617) );
  OAI21_X1 U10797 ( .B1(n4872), .B2(n9643), .A(n9617), .ZN(P1_U3544) );
  AOI211_X1 U10798 ( .C1(n9620), .C2(n9809), .A(n9619), .B(n9618), .ZN(n9709)
         );
  MUX2_X1 U10799 ( .A(n9621), .B(n9709), .S(n9816), .Z(n9622) );
  OAI21_X1 U10800 ( .B1(n9712), .B2(n9643), .A(n9622), .ZN(P1_U3543) );
  AOI211_X1 U10801 ( .C1(n9658), .C2(n9625), .A(n9624), .B(n9623), .ZN(n9626)
         );
  OAI21_X1 U10802 ( .B1(n9627), .B2(n9660), .A(n9626), .ZN(n9713) );
  MUX2_X1 U10803 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9713), .S(n9816), .Z(
        P1_U3542) );
  AOI211_X1 U10804 ( .C1(n9630), .C2(n9809), .A(n9629), .B(n9628), .ZN(n9714)
         );
  MUX2_X1 U10805 ( .A(n9631), .B(n9714), .S(n9816), .Z(n9632) );
  OAI21_X1 U10806 ( .B1(n9717), .B2(n9643), .A(n9632), .ZN(P1_U3541) );
  AOI21_X1 U10807 ( .B1(n9658), .B2(n9634), .A(n9633), .ZN(n9635) );
  OAI211_X1 U10808 ( .C1(n9637), .C2(n9660), .A(n9636), .B(n9635), .ZN(n9718)
         );
  MUX2_X1 U10809 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9718), .S(n9816), .Z(
        P1_U3540) );
  AOI211_X1 U10810 ( .C1(n9640), .C2(n9809), .A(n9639), .B(n9638), .ZN(n9719)
         );
  MUX2_X1 U10811 ( .A(n9641), .B(n9719), .S(n9816), .Z(n9642) );
  OAI21_X1 U10812 ( .B1(n4875), .B2(n9643), .A(n9642), .ZN(P1_U3539) );
  AOI21_X1 U10813 ( .B1(n9658), .B2(n9645), .A(n9644), .ZN(n9646) );
  OAI211_X1 U10814 ( .C1(n9648), .C2(n9660), .A(n9647), .B(n9646), .ZN(n9723)
         );
  MUX2_X1 U10815 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9723), .S(n9816), .Z(
        P1_U3538) );
  AOI22_X1 U10816 ( .A1(n9651), .A2(n9650), .B1(n9658), .B2(n9649), .ZN(n9652)
         );
  OAI211_X1 U10817 ( .C1(n9654), .C2(n9660), .A(n9653), .B(n9652), .ZN(n9724)
         );
  MUX2_X1 U10818 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9724), .S(n9816), .Z(
        P1_U3537) );
  AOI211_X1 U10819 ( .C1(n9658), .C2(n9657), .A(n9656), .B(n9655), .ZN(n9659)
         );
  OAI21_X1 U10820 ( .B1(n9661), .B2(n9660), .A(n9659), .ZN(n9726) );
  MUX2_X1 U10821 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9726), .S(n9816), .Z(
        P1_U3536) );
  OAI21_X1 U10822 ( .B1(n4870), .B2(n9805), .A(n9662), .ZN(n9663) );
  AOI211_X1 U10823 ( .C1(n9665), .C2(n9809), .A(n9664), .B(n9663), .ZN(n9728)
         );
  NAND2_X1 U10824 ( .A1(n9814), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9666) );
  OAI21_X1 U10825 ( .B1(n9728), .B2(n9814), .A(n9666), .ZN(P1_U3535) );
  AOI211_X1 U10826 ( .C1(n9669), .C2(n9809), .A(n9668), .B(n9667), .ZN(n9731)
         );
  AOI22_X1 U10827 ( .A1(n9729), .A2(n9676), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n9814), .ZN(n9670) );
  OAI21_X1 U10828 ( .B1(n9731), .B2(n9814), .A(n9670), .ZN(P1_U3534) );
  INV_X1 U10829 ( .A(n9671), .ZN(n9675) );
  AOI211_X1 U10830 ( .C1(n9675), .C2(n9674), .A(n9673), .B(n9672), .ZN(n9735)
         );
  AOI22_X1 U10831 ( .A1(n4451), .A2(n9676), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n9814), .ZN(n9677) );
  OAI21_X1 U10832 ( .B1(n9735), .B2(n9814), .A(n9677), .ZN(P1_U3533) );
  INV_X1 U10833 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9679) );
  INV_X1 U10834 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9682) );
  OAI21_X1 U10835 ( .B1(n9684), .B2(n9722), .A(n9683), .ZN(P1_U3520) );
  MUX2_X1 U10836 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9685), .S(n9813), .Z(
        P1_U3519) );
  MUX2_X1 U10837 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9686), .S(n9725), .Z(n9687) );
  INV_X1 U10838 ( .A(n9687), .ZN(n9688) );
  OAI21_X1 U10839 ( .B1(n9689), .B2(n9722), .A(n9688), .ZN(P1_U3517) );
  INV_X1 U10840 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9691) );
  MUX2_X1 U10841 ( .A(n9691), .B(n9690), .S(n9725), .Z(n9692) );
  OAI21_X1 U10842 ( .B1(n9693), .B2(n9722), .A(n9692), .ZN(P1_U3516) );
  INV_X1 U10843 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9695) );
  MUX2_X1 U10844 ( .A(n9695), .B(n9694), .S(n9725), .Z(n9696) );
  OAI21_X1 U10845 ( .B1(n9697), .B2(n9722), .A(n9696), .ZN(P1_U3515) );
  INV_X1 U10846 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9699) );
  MUX2_X1 U10847 ( .A(n9699), .B(n9698), .S(n9813), .Z(n9700) );
  OAI21_X1 U10848 ( .B1(n9701), .B2(n9722), .A(n9700), .ZN(P1_U3514) );
  INV_X1 U10849 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9703) );
  MUX2_X1 U10850 ( .A(n9703), .B(n9702), .S(n9813), .Z(n9704) );
  OAI21_X1 U10851 ( .B1(n9705), .B2(n9722), .A(n9704), .ZN(P1_U3513) );
  INV_X1 U10852 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9707) );
  MUX2_X1 U10853 ( .A(n9707), .B(n9706), .S(n9725), .Z(n9708) );
  OAI21_X1 U10854 ( .B1(n4872), .B2(n9722), .A(n9708), .ZN(P1_U3512) );
  INV_X1 U10855 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9710) );
  MUX2_X1 U10856 ( .A(n9710), .B(n9709), .S(n9725), .Z(n9711) );
  OAI21_X1 U10857 ( .B1(n9712), .B2(n9722), .A(n9711), .ZN(P1_U3511) );
  MUX2_X1 U10858 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9713), .S(n9725), .Z(
        P1_U3510) );
  INV_X1 U10859 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9715) );
  MUX2_X1 U10860 ( .A(n9715), .B(n9714), .S(n9725), .Z(n9716) );
  OAI21_X1 U10861 ( .B1(n9717), .B2(n9722), .A(n9716), .ZN(P1_U3509) );
  MUX2_X1 U10862 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9718), .S(n9725), .Z(
        P1_U3507) );
  INV_X1 U10863 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9720) );
  MUX2_X1 U10864 ( .A(n9720), .B(n9719), .S(n9725), .Z(n9721) );
  OAI21_X1 U10865 ( .B1(n4875), .B2(n9722), .A(n9721), .ZN(P1_U3504) );
  MUX2_X1 U10866 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9723), .S(n9725), .Z(
        P1_U3501) );
  MUX2_X1 U10867 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9724), .S(n9725), .Z(
        P1_U3498) );
  MUX2_X1 U10868 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9726), .S(n9725), .Z(
        P1_U3495) );
  NAND2_X1 U10869 ( .A1(n9811), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9727) );
  OAI21_X1 U10870 ( .B1(n9728), .B2(n9811), .A(n9727), .ZN(P1_U3492) );
  AOI22_X1 U10871 ( .A1(n9729), .A2(n9732), .B1(P1_REG0_REG_12__SCAN_IN), .B2(
        n9811), .ZN(n9730) );
  OAI21_X1 U10872 ( .B1(n9731), .B2(n9811), .A(n9730), .ZN(P1_U3489) );
  AOI22_X1 U10873 ( .A1(n4451), .A2(n9732), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n9811), .ZN(n9734) );
  OAI21_X1 U10874 ( .B1(n9735), .B2(n9811), .A(n9734), .ZN(P1_U3486) );
  MUX2_X1 U10875 ( .A(n9736), .B(P1_D_REG_1__SCAN_IN), .S(n9804), .Z(P1_U3440)
         );
  MUX2_X1 U10876 ( .A(n9737), .B(P1_D_REG_0__SCAN_IN), .S(n9804), .Z(P1_U3439)
         );
  NOR4_X1 U10877 ( .A1(n5862), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9738), .A4(
        P1_U3086), .ZN(n9739) );
  AOI21_X1 U10878 ( .B1(n9740), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9739), .ZN(
        n9741) );
  OAI21_X1 U10879 ( .B1(n9742), .B2(n9747), .A(n9741), .ZN(P1_U3324) );
  OAI222_X1 U10880 ( .A1(n9750), .A2(n9745), .B1(P1_U3086), .B2(n9744), .C1(
        n9747), .C2(n9743), .ZN(P1_U3326) );
  OAI222_X1 U10881 ( .A1(n9750), .A2(n9749), .B1(P1_U3086), .B2(n9748), .C1(
        n9747), .C2(n9746), .ZN(P1_U3327) );
  INV_X1 U10882 ( .A(n9751), .ZN(n9752) );
  MUX2_X1 U10883 ( .A(n9752), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10884 ( .A(n9753), .ZN(n9758) );
  AOI21_X1 U10885 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9757) );
  OAI21_X1 U10886 ( .B1(n9758), .B2(n9757), .A(n9785), .ZN(n9765) );
  NAND2_X1 U10887 ( .A1(n9760), .A2(n9759), .ZN(n9761) );
  NAND2_X1 U10888 ( .A1(n9762), .A2(n9761), .ZN(n9763) );
  NAND2_X1 U10889 ( .A1(n9779), .A2(n9763), .ZN(n9764) );
  OAI211_X1 U10890 ( .C1(n9767), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9768)
         );
  INV_X1 U10891 ( .A(n9768), .ZN(n9770) );
  OAI211_X1 U10892 ( .C1(n9771), .C2(n9788), .A(n9770), .B(n9769), .ZN(
        P1_U3252) );
  XNOR2_X1 U10893 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10894 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U10895 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(n9784) );
  OAI21_X1 U10896 ( .B1(n9777), .B2(n9776), .A(n9775), .ZN(n9778) );
  AOI22_X1 U10897 ( .A1(n9781), .A2(n9780), .B1(n9779), .B2(n9778), .ZN(n9782)
         );
  INV_X1 U10898 ( .A(n9782), .ZN(n9783) );
  AOI21_X1 U10899 ( .B1(n9785), .B2(n9784), .A(n9783), .ZN(n9787) );
  OAI211_X1 U10900 ( .C1(n9789), .C2(n9788), .A(n9787), .B(n9786), .ZN(
        P1_U3260) );
  NAND2_X1 U10901 ( .A1(n9791), .A2(n9790), .ZN(n9794) );
  AOI22_X1 U10902 ( .A1(n9802), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9792), .ZN(n9793) );
  OAI211_X1 U10903 ( .C1(n9796), .C2(n9795), .A(n9794), .B(n9793), .ZN(n9797)
         );
  AOI21_X1 U10904 ( .B1(n9799), .B2(n9798), .A(n9797), .ZN(n9800) );
  OAI21_X1 U10905 ( .B1(n9802), .B2(n9801), .A(n9800), .ZN(P1_U3291) );
  AND2_X1 U10906 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9804), .ZN(P1_U3294) );
  AND2_X1 U10907 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9804), .ZN(P1_U3295) );
  AND2_X1 U10908 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9804), .ZN(P1_U3296) );
  AND2_X1 U10909 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9804), .ZN(P1_U3297) );
  AND2_X1 U10910 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9804), .ZN(P1_U3298) );
  AND2_X1 U10911 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9804), .ZN(P1_U3299) );
  AND2_X1 U10912 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9804), .ZN(P1_U3300) );
  AND2_X1 U10913 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9804), .ZN(P1_U3301) );
  AND2_X1 U10914 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9804), .ZN(P1_U3302) );
  AND2_X1 U10915 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9804), .ZN(P1_U3303) );
  AND2_X1 U10916 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9804), .ZN(P1_U3304) );
  AND2_X1 U10917 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9804), .ZN(P1_U3305) );
  AND2_X1 U10918 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9804), .ZN(P1_U3306) );
  AND2_X1 U10919 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9804), .ZN(P1_U3307) );
  INV_X1 U10920 ( .A(n9804), .ZN(n9803) );
  INV_X1 U10921 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10161) );
  NOR2_X1 U10922 ( .A1(n9803), .A2(n10161), .ZN(P1_U3308) );
  AND2_X1 U10923 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9804), .ZN(P1_U3309) );
  AND2_X1 U10924 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9804), .ZN(P1_U3310) );
  AND2_X1 U10925 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9804), .ZN(P1_U3311) );
  AND2_X1 U10926 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9804), .ZN(P1_U3312) );
  AND2_X1 U10927 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9804), .ZN(P1_U3313) );
  INV_X1 U10928 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U10929 ( .A1(n9803), .A2(n10061), .ZN(P1_U3314) );
  AND2_X1 U10930 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9804), .ZN(P1_U3315) );
  INV_X1 U10931 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10103) );
  NOR2_X1 U10932 ( .A1(n9803), .A2(n10103), .ZN(P1_U3316) );
  AND2_X1 U10933 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9804), .ZN(P1_U3317) );
  AND2_X1 U10934 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9804), .ZN(P1_U3318) );
  INV_X1 U10935 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10178) );
  NOR2_X1 U10936 ( .A1(n9803), .A2(n10178), .ZN(P1_U3319) );
  INV_X1 U10937 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10155) );
  NOR2_X1 U10938 ( .A1(n9803), .A2(n10155), .ZN(P1_U3320) );
  AND2_X1 U10939 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9804), .ZN(P1_U3321) );
  AND2_X1 U10940 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9804), .ZN(P1_U3322) );
  AND2_X1 U10941 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9804), .ZN(P1_U3323) );
  NOR2_X1 U10942 ( .A1(n9806), .A2(n9805), .ZN(n9808) );
  AOI211_X1 U10943 ( .C1(n9810), .C2(n9809), .A(n9808), .B(n9807), .ZN(n9815)
         );
  INV_X1 U10944 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9812) );
  AOI22_X1 U10945 ( .A1(n9813), .A2(n9815), .B1(n9812), .B2(n9811), .ZN(
        P1_U3480) );
  AOI22_X1 U10946 ( .A1(n9816), .A2(n9815), .B1(n5916), .B2(n9814), .ZN(
        P1_U3531) );
  OAI21_X1 U10947 ( .B1(n9819), .B2(n9818), .A(n9817), .ZN(n9824) );
  OAI21_X1 U10948 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(n9823) );
  AOI22_X1 U10949 ( .A1(n9916), .A2(n9824), .B1(n9901), .B2(n9823), .ZN(n9828)
         );
  NAND2_X1 U10950 ( .A1(n9826), .A2(n9825), .ZN(n9827) );
  OAI211_X1 U10951 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6259), .A(n9828), .B(
        n9827), .ZN(n9829) );
  AOI21_X1 U10952 ( .B1(n9897), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n9829), .ZN(
        n9834) );
  XOR2_X1 U10953 ( .A(n9831), .B(n9830), .Z(n9832) );
  NAND2_X1 U10954 ( .A1(n9867), .A2(n9832), .ZN(n9833) );
  NAND2_X1 U10955 ( .A1(n9834), .A2(n9833), .ZN(P2_U3184) );
  INV_X1 U10956 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9845) );
  OR2_X1 U10957 ( .A1(n9906), .A2(n9835), .ZN(n9844) );
  INV_X1 U10958 ( .A(n9836), .ZN(n9838) );
  NAND3_X1 U10959 ( .A1(n9839), .A2(n9838), .A3(n9837), .ZN(n9840) );
  NAND2_X1 U10960 ( .A1(n9841), .A2(n9840), .ZN(n9842) );
  NAND2_X1 U10961 ( .A1(n9901), .A2(n9842), .ZN(n9843) );
  OAI211_X1 U10962 ( .C1(n9845), .C2(n9882), .A(n9844), .B(n9843), .ZN(n9846)
         );
  INV_X1 U10963 ( .A(n9846), .ZN(n9857) );
  OAI211_X1 U10964 ( .C1(n9849), .C2(n9848), .A(n9847), .B(n9867), .ZN(n9855)
         );
  OAI21_X1 U10965 ( .B1(n9852), .B2(n9851), .A(n9850), .ZN(n9853) );
  NAND2_X1 U10966 ( .A1(n9916), .A2(n9853), .ZN(n9854) );
  NAND4_X1 U10967 ( .A1(n9857), .A2(n9856), .A3(n9855), .A4(n9854), .ZN(
        P2_U3186) );
  INV_X1 U10968 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9863) );
  OR2_X1 U10969 ( .A1(n9906), .A2(n9858), .ZN(n9862) );
  OAI21_X1 U10970 ( .B1(n4431), .B2(P2_REG1_REG_5__SCAN_IN), .A(n9859), .ZN(
        n9860) );
  NAND2_X1 U10971 ( .A1(n9901), .A2(n9860), .ZN(n9861) );
  OAI211_X1 U10972 ( .C1(n9863), .C2(n9882), .A(n9862), .B(n9861), .ZN(n9864)
         );
  INV_X1 U10973 ( .A(n9864), .ZN(n9875) );
  XOR2_X1 U10974 ( .A(n9866), .B(n9865), .Z(n9868) );
  NAND2_X1 U10975 ( .A1(n9868), .A2(n9867), .ZN(n9873) );
  AOI21_X1 U10976 ( .B1(n5068), .B2(n9870), .A(n9869), .ZN(n9871) );
  OR2_X1 U10977 ( .A1(n9891), .A2(n9871), .ZN(n9872) );
  NAND4_X1 U10978 ( .A1(n9875), .A2(n9874), .A3(n9873), .A4(n9872), .ZN(
        P2_U3187) );
  INV_X1 U10979 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9881) );
  OR2_X1 U10980 ( .A1(n9906), .A2(n9876), .ZN(n9880) );
  OAI21_X1 U10981 ( .B1(n9877), .B2(P2_REG1_REG_7__SCAN_IN), .A(n9900), .ZN(
        n9878) );
  NAND2_X1 U10982 ( .A1(n9901), .A2(n9878), .ZN(n9879) );
  OAI211_X1 U10983 ( .C1(n9882), .C2(n9881), .A(n9880), .B(n9879), .ZN(n9883)
         );
  INV_X1 U10984 ( .A(n9883), .ZN(n9896) );
  AOI21_X1 U10985 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9887) );
  OR2_X1 U10986 ( .A1(n9887), .A2(n9911), .ZN(n9894) );
  INV_X1 U10987 ( .A(n9888), .ZN(n9889) );
  AOI21_X1 U10988 ( .B1(n6623), .B2(n9890), .A(n9889), .ZN(n9892) );
  OR2_X1 U10989 ( .A1(n9892), .A2(n9891), .ZN(n9893) );
  NAND4_X1 U10990 ( .A1(n9896), .A2(n9895), .A3(n9894), .A4(n9893), .ZN(
        P2_U3189) );
  NAND2_X1 U10991 ( .A1(n9897), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9905) );
  AND3_X1 U10992 ( .A1(n9900), .A2(n9899), .A3(n9898), .ZN(n9902) );
  OAI21_X1 U10993 ( .B1(n9903), .B2(n9902), .A(n9901), .ZN(n9904) );
  OAI211_X1 U10994 ( .C1(n9906), .C2(n4499), .A(n9905), .B(n9904), .ZN(n9907)
         );
  INV_X1 U10995 ( .A(n9907), .ZN(n9921) );
  AOI21_X1 U10996 ( .B1(n9910), .B2(n9909), .A(n9908), .ZN(n9912) );
  OR2_X1 U10997 ( .A1(n9912), .A2(n9911), .ZN(n9919) );
  OAI21_X1 U10998 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9917) );
  NAND2_X1 U10999 ( .A1(n9917), .A2(n9916), .ZN(n9918) );
  NAND4_X1 U11000 ( .A1(n9921), .A2(n9920), .A3(n9919), .A4(n9918), .ZN(
        P2_U3190) );
  INV_X1 U11001 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9926) );
  OAI21_X1 U11002 ( .B1(n9923), .B2(n9947), .A(n9922), .ZN(n9924) );
  AOI21_X1 U11003 ( .B1(n9933), .B2(n9925), .A(n9924), .ZN(n9967) );
  AOI22_X1 U11004 ( .A1(n9966), .A2(n9926), .B1(n9967), .B2(n9965), .ZN(
        P2_U3393) );
  OAI22_X1 U11005 ( .A1(n9928), .A2(n9959), .B1(n9927), .B2(n9947), .ZN(n9930)
         );
  OR2_X1 U11006 ( .A1(n9930), .A2(n9929), .ZN(n10191) );
  MUX2_X1 U11007 ( .A(P2_REG0_REG_2__SCAN_IN), .B(n10191), .S(n9965), .Z(
        P2_U3396) );
  AND2_X1 U11008 ( .A1(n9931), .A2(n9964), .ZN(n9932) );
  AOI21_X1 U11009 ( .B1(n9934), .B2(n9933), .A(n9932), .ZN(n9935) );
  AND2_X1 U11010 ( .A1(n9936), .A2(n9935), .ZN(n9969) );
  AOI22_X1 U11011 ( .A1(n9966), .A2(n5036), .B1(n9969), .B2(n9965), .ZN(
        P2_U3402) );
  OAI22_X1 U11012 ( .A1(n9939), .A2(n9938), .B1(n9937), .B2(n9947), .ZN(n9940)
         );
  NOR2_X1 U11013 ( .A1(n9941), .A2(n9940), .ZN(n9971) );
  AOI22_X1 U11014 ( .A1(n9966), .A2(n5062), .B1(n9971), .B2(n9965), .ZN(
        P2_U3405) );
  NOR2_X1 U11015 ( .A1(n9942), .A2(n9959), .ZN(n9944) );
  AOI211_X1 U11016 ( .C1(n9964), .C2(n9945), .A(n9944), .B(n9943), .ZN(n9973)
         );
  AOI22_X1 U11017 ( .A1(n9966), .A2(n5135), .B1(n9973), .B2(n9965), .ZN(
        P2_U3414) );
  INV_X1 U11018 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9953) );
  INV_X1 U11019 ( .A(n9946), .ZN(n9951) );
  NOR2_X1 U11020 ( .A1(n9948), .A2(n9947), .ZN(n9950) );
  AOI211_X1 U11021 ( .C1(n9952), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9974)
         );
  AOI22_X1 U11022 ( .A1(n9966), .A2(n9953), .B1(n9974), .B2(n9965), .ZN(
        P2_U3420) );
  INV_X1 U11023 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9958) );
  NOR2_X1 U11024 ( .A1(n9954), .A2(n9959), .ZN(n9956) );
  AOI211_X1 U11025 ( .C1(n9964), .C2(n9957), .A(n9956), .B(n9955), .ZN(n9975)
         );
  AOI22_X1 U11026 ( .A1(n9966), .A2(n9958), .B1(n9975), .B2(n9965), .ZN(
        P2_U3423) );
  NOR2_X1 U11027 ( .A1(n9960), .A2(n9959), .ZN(n9962) );
  AOI211_X1 U11028 ( .C1(n9964), .C2(n9963), .A(n9962), .B(n9961), .ZN(n9976)
         );
  AOI22_X1 U11029 ( .A1(n9966), .A2(n5216), .B1(n9976), .B2(n9965), .ZN(
        P2_U3426) );
  AOI22_X1 U11030 ( .A1(n10192), .A2(n9967), .B1(n6299), .B2(n10190), .ZN(
        P2_U3460) );
  AOI22_X1 U11031 ( .A1(n10192), .A2(n9969), .B1(n9968), .B2(n10190), .ZN(
        P2_U3463) );
  INV_X1 U11032 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11033 ( .A1(n10192), .A2(n9971), .B1(n9970), .B2(n10190), .ZN(
        P2_U3464) );
  AOI22_X1 U11034 ( .A1(n10192), .A2(n9973), .B1(n9972), .B2(n10190), .ZN(
        P2_U3467) );
  AOI22_X1 U11035 ( .A1(n10192), .A2(n9974), .B1(n5184), .B2(n10190), .ZN(
        P2_U3469) );
  AOI22_X1 U11036 ( .A1(n10192), .A2(n9975), .B1(n5198), .B2(n10190), .ZN(
        P2_U3470) );
  AOI22_X1 U11037 ( .A1(n10192), .A2(n9976), .B1(n7158), .B2(n10190), .ZN(
        P2_U3471) );
  INV_X1 U11038 ( .A(n9977), .ZN(n9978) );
  NAND2_X1 U11039 ( .A1(n9979), .A2(n9978), .ZN(n9980) );
  XOR2_X1 U11040 ( .A(n9981), .B(n9980), .Z(ADD_1068_U5) );
  XOR2_X1 U11041 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11042 ( .A1(n9983), .A2(n9982), .ZN(n9984) );
  XOR2_X1 U11043 ( .A(n9984), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55) );
  XNOR2_X1 U11044 ( .A(n9986), .B(n9985), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11045 ( .A(n9988), .B(n9987), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11046 ( .A(n9990), .B(n9989), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11047 ( .A(n9992), .B(n9991), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11048 ( .A(n9994), .B(n9993), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11049 ( .A(n9996), .B(n9995), .ZN(ADD_1068_U61) );
  XOR2_X1 U11050 ( .A(n9998), .B(n9997), .Z(ADD_1068_U62) );
  XOR2_X1 U11051 ( .A(n10000), .B(n9999), .Z(ADD_1068_U63) );
  INV_X1 U11052 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10002) );
  OAI22_X1 U11053 ( .A1(n10003), .A2(keyinput44), .B1(n10002), .B2(keyinput41), 
        .ZN(n10001) );
  AOI221_X1 U11054 ( .B1(n10003), .B2(keyinput44), .C1(keyinput41), .C2(n10002), .A(n10001), .ZN(n10012) );
  OAI22_X1 U11055 ( .A1(n10082), .A2(keyinput53), .B1(n10005), .B2(keyinput12), 
        .ZN(n10004) );
  AOI221_X1 U11056 ( .B1(n10082), .B2(keyinput53), .C1(keyinput12), .C2(n10005), .A(n10004), .ZN(n10011) );
  OAI22_X1 U11057 ( .A1(n10007), .A2(keyinput46), .B1(n10102), .B2(keyinput38), 
        .ZN(n10006) );
  AOI221_X1 U11058 ( .B1(n10007), .B2(keyinput46), .C1(keyinput38), .C2(n10102), .A(n10006), .ZN(n10010) );
  OAI22_X1 U11059 ( .A1(n10103), .A2(keyinput4), .B1(n10061), .B2(keyinput42), 
        .ZN(n10008) );
  AOI221_X1 U11060 ( .B1(n10103), .B2(keyinput4), .C1(keyinput42), .C2(n10061), 
        .A(n10008), .ZN(n10009) );
  NAND4_X1 U11061 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10189) );
  OAI22_X1 U11062 ( .A1(n7914), .A2(keyinput11), .B1(n10014), .B2(keyinput6), 
        .ZN(n10013) );
  AOI221_X1 U11063 ( .B1(n7914), .B2(keyinput11), .C1(keyinput6), .C2(n10014), 
        .A(n10013), .ZN(n10022) );
  OAI22_X1 U11064 ( .A1(n10063), .A2(keyinput9), .B1(n7112), .B2(keyinput20), 
        .ZN(n10015) );
  AOI221_X1 U11065 ( .B1(n10063), .B2(keyinput9), .C1(keyinput20), .C2(n7112), 
        .A(n10015), .ZN(n10021) );
  XNOR2_X1 U11066 ( .A(P2_B_REG_SCAN_IN), .B(keyinput62), .ZN(n10019) );
  XNOR2_X1 U11067 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput1), .ZN(n10018) );
  XNOR2_X1 U11068 ( .A(P1_REG3_REG_11__SCAN_IN), .B(keyinput54), .ZN(n10017)
         );
  XNOR2_X1 U11069 ( .A(keyinput59), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n10016)
         );
  AND4_X1 U11070 ( .A1(n10019), .A2(n10018), .A3(n10017), .A4(n10016), .ZN(
        n10020) );
  NAND3_X1 U11071 ( .A1(n10022), .A2(n10021), .A3(n10020), .ZN(n10188) );
  AOI22_X1 U11072 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(keyinput2), .B1(
        P1_IR_REG_1__SCAN_IN), .B2(keyinput47), .ZN(n10023) );
  OAI221_X1 U11073 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(keyinput2), .C1(
        P1_IR_REG_1__SCAN_IN), .C2(keyinput47), .A(n10023), .ZN(n10030) );
  AOI22_X1 U11074 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(keyinput16), .B1(
        P2_REG2_REG_28__SCAN_IN), .B2(keyinput43), .ZN(n10024) );
  OAI221_X1 U11075 ( .B1(P1_REG0_REG_4__SCAN_IN), .B2(keyinput16), .C1(
        P2_REG2_REG_28__SCAN_IN), .C2(keyinput43), .A(n10024), .ZN(n10029) );
  AOI22_X1 U11076 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(keyinput45), .B1(
        P2_IR_REG_24__SCAN_IN), .B2(keyinput61), .ZN(n10025) );
  OAI221_X1 U11077 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(keyinput45), .C1(
        P2_IR_REG_24__SCAN_IN), .C2(keyinput61), .A(n10025), .ZN(n10028) );
  AOI22_X1 U11078 ( .A1(P1_REG0_REG_6__SCAN_IN), .A2(keyinput15), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(keyinput17), .ZN(n10026) );
  OAI221_X1 U11079 ( .B1(P1_REG0_REG_6__SCAN_IN), .B2(keyinput15), .C1(
        P1_DATAO_REG_22__SCAN_IN), .C2(keyinput17), .A(n10026), .ZN(n10027) );
  NOR4_X1 U11080 ( .A1(n10030), .A2(n10029), .A3(n10028), .A4(n10027), .ZN(
        n10058) );
  AOI22_X1 U11081 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(keyinput48), .B1(
        P2_REG1_REG_15__SCAN_IN), .B2(keyinput49), .ZN(n10031) );
  OAI221_X1 U11082 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(keyinput48), .C1(
        P2_REG1_REG_15__SCAN_IN), .C2(keyinput49), .A(n10031), .ZN(n10038) );
  AOI22_X1 U11083 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(keyinput52), .B1(
        P2_IR_REG_28__SCAN_IN), .B2(keyinput18), .ZN(n10032) );
  OAI221_X1 U11084 ( .B1(P1_DATAO_REG_3__SCAN_IN), .B2(keyinput52), .C1(
        P2_IR_REG_28__SCAN_IN), .C2(keyinput18), .A(n10032), .ZN(n10037) );
  AOI22_X1 U11085 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(keyinput32), .B1(SI_16_), 
        .B2(keyinput39), .ZN(n10033) );
  OAI221_X1 U11086 ( .B1(P1_REG3_REG_13__SCAN_IN), .B2(keyinput32), .C1(SI_16_), .C2(keyinput39), .A(n10033), .ZN(n10036) );
  AOI22_X1 U11087 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(keyinput56), .B1(
        P2_IR_REG_1__SCAN_IN), .B2(keyinput55), .ZN(n10034) );
  OAI221_X1 U11088 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(keyinput56), .C1(
        P2_IR_REG_1__SCAN_IN), .C2(keyinput55), .A(n10034), .ZN(n10035) );
  NOR4_X1 U11089 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10035), .ZN(
        n10057) );
  AOI22_X1 U11090 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(keyinput57), .B1(
        P2_IR_REG_4__SCAN_IN), .B2(keyinput35), .ZN(n10039) );
  OAI221_X1 U11091 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(keyinput57), .C1(
        P2_IR_REG_4__SCAN_IN), .C2(keyinput35), .A(n10039), .ZN(n10046) );
  AOI22_X1 U11092 ( .A1(P1_REG1_REG_23__SCAN_IN), .A2(keyinput0), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(keyinput36), .ZN(n10040) );
  OAI221_X1 U11093 ( .B1(P1_REG1_REG_23__SCAN_IN), .B2(keyinput0), .C1(
        P1_DATAO_REG_20__SCAN_IN), .C2(keyinput36), .A(n10040), .ZN(n10045) );
  AOI22_X1 U11094 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput28), .B1(
        P2_IR_REG_25__SCAN_IN), .B2(keyinput21), .ZN(n10041) );
  OAI221_X1 U11095 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput28), .C1(
        P2_IR_REG_25__SCAN_IN), .C2(keyinput21), .A(n10041), .ZN(n10044) );
  AOI22_X1 U11096 ( .A1(P2_REG1_REG_2__SCAN_IN), .A2(keyinput37), .B1(
        P2_REG1_REG_30__SCAN_IN), .B2(keyinput29), .ZN(n10042) );
  OAI221_X1 U11097 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(keyinput37), .C1(
        P2_REG1_REG_30__SCAN_IN), .C2(keyinput29), .A(n10042), .ZN(n10043) );
  NOR4_X1 U11098 ( .A1(n10046), .A2(n10045), .A3(n10044), .A4(n10043), .ZN(
        n10056) );
  AOI22_X1 U11099 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(keyinput25), .B1(
        P2_REG0_REG_5__SCAN_IN), .B2(keyinput58), .ZN(n10047) );
  OAI221_X1 U11100 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(keyinput25), .C1(
        P2_REG0_REG_5__SCAN_IN), .C2(keyinput58), .A(n10047), .ZN(n10054) );
  AOI22_X1 U11101 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(keyinput30), .B1(
        P1_REG2_REG_22__SCAN_IN), .B2(keyinput3), .ZN(n10048) );
  OAI221_X1 U11102 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(keyinput30), .C1(
        P1_REG2_REG_22__SCAN_IN), .C2(keyinput3), .A(n10048), .ZN(n10053) );
  AOI22_X1 U11103 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput31), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput8), .ZN(n10049) );
  OAI221_X1 U11104 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput31), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput8), .A(n10049), .ZN(n10052) );
  AOI22_X1 U11105 ( .A1(SI_9_), .A2(keyinput5), .B1(n10060), .B2(keyinput34), 
        .ZN(n10050) );
  OAI221_X1 U11106 ( .B1(SI_9_), .B2(keyinput5), .C1(n10060), .C2(keyinput34), 
        .A(n10050), .ZN(n10051) );
  NOR4_X1 U11107 ( .A1(n10054), .A2(n10053), .A3(n10052), .A4(n10051), .ZN(
        n10055) );
  NAND4_X1 U11108 ( .A1(n10058), .A2(n10057), .A3(n10056), .A4(n10055), .ZN(
        n10187) );
  AOI22_X1 U11109 ( .A1(n10061), .A2(keyinput106), .B1(keyinput98), .B2(n10060), .ZN(n10059) );
  OAI221_X1 U11110 ( .B1(n10061), .B2(keyinput106), .C1(n10060), .C2(
        keyinput98), .A(n10059), .ZN(n10073) );
  AOI22_X1 U11111 ( .A1(n7135), .A2(keyinput123), .B1(keyinput73), .B2(n10063), 
        .ZN(n10062) );
  OAI221_X1 U11112 ( .B1(n7135), .B2(keyinput123), .C1(n10063), .C2(keyinput73), .A(n10062), .ZN(n10072) );
  AOI22_X1 U11113 ( .A1(n10066), .A2(keyinput107), .B1(keyinput113), .B2(
        n10065), .ZN(n10064) );
  OAI221_X1 U11114 ( .B1(n10066), .B2(keyinput107), .C1(n10065), .C2(
        keyinput113), .A(n10064), .ZN(n10071) );
  XOR2_X1 U11115 ( .A(n10067), .B(keyinput101), .Z(n10069) );
  XNOR2_X1 U11116 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput95), .ZN(n10068) );
  NAND2_X1 U11117 ( .A1(n10069), .A2(n10068), .ZN(n10070) );
  NOR4_X1 U11118 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10114) );
  AOI22_X1 U11119 ( .A1(n10076), .A2(keyinput69), .B1(n10075), .B2(keyinput100), .ZN(n10074) );
  OAI221_X1 U11120 ( .B1(n10076), .B2(keyinput69), .C1(n10075), .C2(
        keyinput100), .A(n10074), .ZN(n10087) );
  AOI22_X1 U11121 ( .A1(n10178), .A2(keyinput127), .B1(keyinput118), .B2(
        n10078), .ZN(n10077) );
  OAI221_X1 U11122 ( .B1(n10178), .B2(keyinput127), .C1(n10078), .C2(
        keyinput118), .A(n10077), .ZN(n10086) );
  AOI22_X1 U11123 ( .A1(n10080), .A2(keyinput89), .B1(n10161), .B2(keyinput114), .ZN(n10079) );
  OAI221_X1 U11124 ( .B1(n10080), .B2(keyinput89), .C1(n10161), .C2(
        keyinput114), .A(n10079), .ZN(n10085) );
  AOI22_X1 U11125 ( .A1(n10083), .A2(keyinput81), .B1(n10082), .B2(keyinput117), .ZN(n10081) );
  OAI221_X1 U11126 ( .B1(n10083), .B2(keyinput81), .C1(n10082), .C2(
        keyinput117), .A(n10081), .ZN(n10084) );
  NOR4_X1 U11127 ( .A1(n10087), .A2(n10086), .A3(n10085), .A4(n10084), .ZN(
        n10113) );
  INV_X1 U11128 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U11129 ( .A1(n10090), .A2(keyinput64), .B1(n10089), .B2(keyinput83), 
        .ZN(n10088) );
  OAI221_X1 U11130 ( .B1(n10090), .B2(keyinput64), .C1(n10089), .C2(keyinput83), .A(n10088), .ZN(n10099) );
  XOR2_X1 U11131 ( .A(P2_REG0_REG_31__SCAN_IN), .B(keyinput105), .Z(n10098) );
  XNOR2_X1 U11132 ( .A(n10091), .B(keyinput126), .ZN(n10097) );
  XNOR2_X1 U11133 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput99), .ZN(n10095) );
  XNOR2_X1 U11134 ( .A(P1_REG0_REG_27__SCAN_IN), .B(keyinput124), .ZN(n10094)
         );
  XNOR2_X1 U11135 ( .A(P2_REG1_REG_20__SCAN_IN), .B(keyinput71), .ZN(n10093)
         );
  XNOR2_X1 U11136 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput91), .ZN(n10092) );
  NAND4_X1 U11137 ( .A1(n10095), .A2(n10094), .A3(n10093), .A4(n10092), .ZN(
        n10096) );
  NOR4_X1 U11138 ( .A1(n10099), .A2(n10098), .A3(n10097), .A4(n10096), .ZN(
        n10112) );
  AOI22_X1 U11139 ( .A1(n5599), .A2(keyinput85), .B1(keyinput88), .B2(n10169), 
        .ZN(n10100) );
  OAI221_X1 U11140 ( .B1(n5599), .B2(keyinput85), .C1(n10169), .C2(keyinput88), 
        .A(n10100), .ZN(n10110) );
  AOI22_X1 U11141 ( .A1(n10103), .A2(keyinput68), .B1(n10102), .B2(keyinput102), .ZN(n10101) );
  OAI221_X1 U11142 ( .B1(n10103), .B2(keyinput68), .C1(n10102), .C2(
        keyinput102), .A(n10101), .ZN(n10109) );
  XNOR2_X1 U11143 ( .A(P1_REG3_REG_13__SCAN_IN), .B(keyinput96), .ZN(n10107)
         );
  XNOR2_X1 U11144 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput104), .ZN(n10106)
         );
  XNOR2_X1 U11145 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput116), .ZN(n10105)
         );
  XNOR2_X1 U11146 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput97), .ZN(n10104) );
  NAND4_X1 U11147 ( .A1(n10107), .A2(n10106), .A3(n10105), .A4(n10104), .ZN(
        n10108) );
  NOR3_X1 U11148 ( .A1(n10110), .A2(n10109), .A3(n10108), .ZN(n10111) );
  NAND4_X1 U11149 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n10185) );
  AOI22_X1 U11150 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(keyinput66), .B1(
        P2_REG0_REG_14__SCAN_IN), .B2(keyinput108), .ZN(n10115) );
  OAI221_X1 U11151 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(keyinput66), .C1(
        P2_REG0_REG_14__SCAN_IN), .C2(keyinput108), .A(n10115), .ZN(n10122) );
  AOI22_X1 U11152 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(keyinput94), .B1(
        P1_D_REG_5__SCAN_IN), .B2(keyinput78), .ZN(n10116) );
  OAI221_X1 U11153 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(keyinput94), .C1(
        P1_D_REG_5__SCAN_IN), .C2(keyinput78), .A(n10116), .ZN(n10121) );
  AOI22_X1 U11154 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput111), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput76), .ZN(n10117) );
  OAI221_X1 U11155 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput111), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput76), .A(n10117), .ZN(n10120) );
  AOI22_X1 U11156 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(keyinput120), .B1(
        P2_IR_REG_1__SCAN_IN), .B2(keyinput119), .ZN(n10118) );
  OAI221_X1 U11157 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(keyinput120), .C1(
        P2_IR_REG_1__SCAN_IN), .C2(keyinput119), .A(n10118), .ZN(n10119) );
  NOR4_X1 U11158 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10153) );
  AOI22_X1 U11159 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput72), .B1(
        P2_IR_REG_18__SCAN_IN), .B2(keyinput65), .ZN(n10123) );
  OAI221_X1 U11160 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput72), .C1(
        P2_IR_REG_18__SCAN_IN), .C2(keyinput65), .A(n10123), .ZN(n10130) );
  AOI22_X1 U11161 ( .A1(P2_REG0_REG_5__SCAN_IN), .A2(keyinput122), .B1(
        P2_REG2_REG_14__SCAN_IN), .B2(keyinput75), .ZN(n10124) );
  OAI221_X1 U11162 ( .B1(P2_REG0_REG_5__SCAN_IN), .B2(keyinput122), .C1(
        P2_REG2_REG_14__SCAN_IN), .C2(keyinput75), .A(n10124), .ZN(n10129) );
  AOI22_X1 U11163 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput90), .B1(
        P2_REG2_REG_3__SCAN_IN), .B2(keyinput112), .ZN(n10125) );
  OAI221_X1 U11164 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput90), .C1(
        P2_REG2_REG_3__SCAN_IN), .C2(keyinput112), .A(n10125), .ZN(n10128) );
  AOI22_X1 U11165 ( .A1(P1_REG2_REG_22__SCAN_IN), .A2(keyinput67), .B1(SI_16_), 
        .B2(keyinput103), .ZN(n10126) );
  OAI221_X1 U11166 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(keyinput67), .C1(SI_16_), .C2(keyinput103), .A(n10126), .ZN(n10127) );
  NOR4_X1 U11167 ( .A1(n10130), .A2(n10129), .A3(n10128), .A4(n10127), .ZN(
        n10152) );
  AOI22_X1 U11168 ( .A1(n10132), .A2(keyinput93), .B1(keyinput84), .B2(n7112), 
        .ZN(n10131) );
  OAI221_X1 U11169 ( .B1(n10132), .B2(keyinput93), .C1(n7112), .C2(keyinput84), 
        .A(n10131), .ZN(n10141) );
  AOI22_X1 U11170 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(keyinput109), .B1(n9324), 
        .B2(keyinput121), .ZN(n10133) );
  OAI221_X1 U11171 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(keyinput109), .C1(n9324), 
        .C2(keyinput121), .A(n10133), .ZN(n10140) );
  AOI22_X1 U11172 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(keyinput80), .B1(SI_21_), 
        .B2(keyinput74), .ZN(n10134) );
  OAI221_X1 U11173 ( .B1(P1_REG0_REG_4__SCAN_IN), .B2(keyinput80), .C1(SI_21_), 
        .C2(keyinput74), .A(n10134), .ZN(n10139) );
  XOR2_X1 U11174 ( .A(n10135), .B(keyinput79), .Z(n10137) );
  XNOR2_X1 U11175 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput87), .ZN(n10136) );
  NAND2_X1 U11176 ( .A1(n10137), .A2(n10136), .ZN(n10138) );
  NOR4_X1 U11177 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10151) );
  AOI22_X1 U11178 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput86), .B1(
        P2_IR_REG_24__SCAN_IN), .B2(keyinput125), .ZN(n10142) );
  OAI221_X1 U11179 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput86), .C1(
        P2_IR_REG_24__SCAN_IN), .C2(keyinput125), .A(n10142), .ZN(n10149) );
  AOI22_X1 U11180 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput110), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput92), .ZN(n10143) );
  OAI221_X1 U11181 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput110), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput92), .A(n10143), .ZN(n10148) );
  AOI22_X1 U11182 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(keyinput70), .B1(SI_24_), 
        .B2(keyinput115), .ZN(n10144) );
  OAI221_X1 U11183 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(keyinput70), .C1(SI_24_), 
        .C2(keyinput115), .A(n10144), .ZN(n10147) );
  AOI22_X1 U11184 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(keyinput77), .B1(
        P2_IR_REG_28__SCAN_IN), .B2(keyinput82), .ZN(n10145) );
  OAI221_X1 U11185 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(keyinput77), .C1(
        P2_IR_REG_28__SCAN_IN), .C2(keyinput82), .A(n10145), .ZN(n10146) );
  NOR4_X1 U11186 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10150) );
  NAND4_X1 U11187 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10184) );
  AOI22_X1 U11188 ( .A1(n10155), .A2(keyinput14), .B1(n5378), .B2(keyinput10), 
        .ZN(n10154) );
  OAI221_X1 U11189 ( .B1(n10155), .B2(keyinput14), .C1(n5378), .C2(keyinput10), 
        .A(n10154), .ZN(n10167) );
  INV_X1 U11190 ( .A(SI_24_), .ZN(n10157) );
  AOI22_X1 U11191 ( .A1(n10158), .A2(keyinput60), .B1(n10157), .B2(keyinput51), 
        .ZN(n10156) );
  OAI221_X1 U11192 ( .B1(n10158), .B2(keyinput60), .C1(n10157), .C2(keyinput51), .A(n10156), .ZN(n10166) );
  INV_X1 U11193 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U11194 ( .A1(n10161), .A2(keyinput50), .B1(keyinput13), .B2(n10160), 
        .ZN(n10159) );
  OAI221_X1 U11195 ( .B1(n10161), .B2(keyinput50), .C1(n10160), .C2(keyinput13), .A(n10159), .ZN(n10165) );
  XNOR2_X1 U11196 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput26), .ZN(n10163) );
  XNOR2_X1 U11197 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput23), .ZN(n10162) );
  NAND2_X1 U11198 ( .A1(n10163), .A2(n10162), .ZN(n10164) );
  NOR4_X1 U11199 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10183) );
  AOI22_X1 U11200 ( .A1(n10170), .A2(keyinput22), .B1(n10169), .B2(keyinput24), 
        .ZN(n10168) );
  OAI221_X1 U11201 ( .B1(n10170), .B2(keyinput22), .C1(n10169), .C2(keyinput24), .A(n10168), .ZN(n10181) );
  XOR2_X1 U11202 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput33), .Z(n10173) );
  XNOR2_X1 U11203 ( .A(n10171), .B(keyinput7), .ZN(n10172) );
  NOR2_X1 U11204 ( .A1(n10173), .A2(n10172), .ZN(n10177) );
  XNOR2_X1 U11205 ( .A(keyinput19), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n10176) );
  XNOR2_X1 U11206 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput40), .ZN(n10175) );
  XNOR2_X1 U11207 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput27), .ZN(n10174) );
  NAND4_X1 U11208 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n10180) );
  XNOR2_X1 U11209 ( .A(n10178), .B(keyinput63), .ZN(n10179) );
  NOR3_X1 U11210 ( .A1(n10181), .A2(n10180), .A3(n10179), .ZN(n10182) );
  OAI211_X1 U11211 ( .C1(n10185), .C2(n10184), .A(n10183), .B(n10182), .ZN(
        n10186) );
  NOR4_X1 U11212 ( .A1(n10189), .A2(n10188), .A3(n10187), .A4(n10186), .ZN(
        n10194) );
  AOI22_X1 U11213 ( .A1(n10192), .A2(n10191), .B1(P2_REG1_REG_2__SCAN_IN), 
        .B2(n10190), .ZN(n10193) );
  XNOR2_X1 U11214 ( .A(n10194), .B(n10193), .ZN(P2_U3461) );
  XOR2_X1 U11215 ( .A(n10195), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1068_U50) );
  NOR2_X1 U11216 ( .A1(n10197), .A2(n10196), .ZN(n10198) );
  XOR2_X1 U11217 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10198), .Z(ADD_1068_U51) );
  INV_X1 U11218 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10199) );
  XNOR2_X1 U11219 ( .A(n10200), .B(n10199), .ZN(ADD_1068_U47) );
  XOR2_X1 U11220 ( .A(n10201), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1068_U49) );
  XOR2_X1 U11221 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10202), .Z(ADD_1068_U48) );
  XOR2_X1 U11222 ( .A(n10204), .B(n10203), .Z(ADD_1068_U54) );
  XOR2_X1 U11223 ( .A(n10206), .B(n10205), .Z(ADD_1068_U53) );
  XNOR2_X1 U11224 ( .A(n10208), .B(n10207), .ZN(ADD_1068_U52) );
  MUX2_X1 U5069 ( .A(n9682), .B(n9681), .S(n9725), .Z(n9683) );
  CLKBUF_X1 U4864 ( .A(n8770), .Z(n4334) );
  MUX2_X1 U5070 ( .A(n9582), .B(n9681), .S(n9816), .Z(n9583) );
endmodule

